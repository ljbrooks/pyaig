module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, out1);
  input [15:0] in1, in2, in5, in8, in9, in12, in13, in16, in17, in20, in21, in24, in25;
  input in3, in4, in6, in7, in10, in11, in14, in15, in18, in19, in22, in23;
  output [31:0] out1;
  wire [15:0] in1, in2, in5, in8, in9, in12, in13, in16, in17, in20, in21, in24, in25;
  wire in3, in4, in6, in7, in10, in11, in14, in15, in18, in19, in22, in23;
  wire [31:0] out1;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__139, w__140, w__141, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__157, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__171, w__172, w__173, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__665, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__680;
  wire w__681, w__682, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__697, w__698, w__699, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__714, w__715, w__716, w__717, w__718, w__719, w__720;
  wire w__721, w__722, w__723, w__724, w__725, w__726, w__727, w__728;
  wire w__729, w__730, w__731, w__732, w__733, w__734, w__735, w__736;
  wire w__737, w__738, w__739, w__740, w__741, w__742, w__743, w__744;
  wire w__745, w__746, w__747, w__748, w__749, w__750, w__751, w__752;
  wire w__753, w__754, w__755, w__756, w__757, w__758, w__759, w__760;
  wire w__761, w__762, w__763, w__764, w__765, w__766, w__767, w__768;
  wire w__769, w__770, w__771, w__772, w__773, w__774, w__775, w__776;
  wire w__777, w__778, w__779, w__780, w__781, w__782, w__783, w__784;
  wire w__785, w__786, w__787, w__788, w__789, w__790, w__791, w__792;
  wire w__793, w__794, w__795, w__796, w__797, w__798, w__799, w__800;
  wire w__801, w__802, w__803, w__804, w__805, w__806, w__807, w__808;
  wire w__809, w__810, w__811, w__812, w__813, w__814, w__815, w__816;
  wire w__817, w__818, w__819, w__820, w__821, w__822, w__823, w__824;
  wire w__825, w__826, w__827, w__828, w__829, w__830, w__831, w__832;
  wire w__833, w__834, w__835, w__836, w__837, w__838, w__839, w__840;
  wire w__841, w__842, w__843, w__844, w__845, w__846, w__847, w__848;
  wire w__849, w__850, w__851, w__852, w__853, w__854, w__855, w__856;
  wire w__857, w__858, w__859, w__860, w__861, w__862, w__863, w__864;
  wire w__865, w__866, w__867, w__868, w__869, w__870, w__871, w__872;
  wire w__873, w__874, w__875, w__876, w__877, w__878, w__879, w__880;
  wire w__881, w__882, w__883, w__884, w__885, w__886, w__887, w__888;
  wire w__889, w__890, w__891, w__892, w__893, w__894, w__895, w__896;
  wire w__897, w__898, w__899, w__900, w__901, w__902, w__903, w__904;
  wire w__905, w__906, w__907, w__908, w__909, w__910, w__911, w__912;
  wire w__913, w__914, w__915, w__916, w__917, w__918, w__919, w__920;
  wire w__921, w__922, w__923, w__924, w__925, w__926, w__927, w__928;
  wire w__929, w__930, w__931, w__932, w__933, w__934, w__935, w__936;
  wire w__937, w__938, w__939, w__940, w__941, w__942, w__943, w__944;
  wire w__945, w__946, w__947, w__948, w__949, w__950, w__951, w__952;
  wire w__953, w__954, w__955, w__956, w__957, w__958, w__959, w__960;
  wire w__961, w__962, w__963, w__964, w__965, w__966, w__967, w__968;
  wire w__969, w__970, w__971, w__972, w__973, w__974, w__975, w__976;
  wire w__977, w__978, w__979, w__980, w__981, w__982, w__983, w__984;
  wire w__985, w__986, w__987, w__988, w__989, w__990, w__991, w__992;
  wire w__993, w__994, w__995, w__996, w__997, w__998, w__999, w__1000;
  wire w__1001, w__1002, w__1003, w__1004, w__1005, w__1006, w__1007, w__1008;
  wire w__1009, w__1010, w__1011, w__1012, w__1013, w__1014, w__1015, w__1016;
  wire w__1017, w__1018, w__1019, w__1020, w__1021, w__1022, w__1023, w__1024;
  wire w__1025, w__1026, w__1027, w__1028, w__1029, w__1030, w__1031, w__1032;
  wire w__1033, w__1034, w__1035, w__1036, w__1037, w__1038, w__1039, w__1040;
  wire w__1041, w__1042, w__1043, w__1044, w__1045, w__1046, w__1047, w__1048;
  wire w__1049, w__1050, w__1051, w__1052, w__1053, w__1054, w__1055, w__1056;
  wire w__1057, w__1058, w__1059, w__1060, w__1061, w__1062, w__1063, w__1064;
  wire w__1065, w__1066, w__1067, w__1068, w__1069, w__1070, w__1071, w__1072;
  wire w__1073, w__1074, w__1075, w__1076, w__1077, w__1078, w__1079, w__1080;
  wire w__1081, w__1082, w__1083, w__1084, w__1085, w__1086, w__1087, w__1088;
  wire w__1089, w__1090, w__1091, w__1092, w__1093, w__1094, w__1095, w__1096;
  wire w__1097, w__1098, w__1099, w__1100, w__1101, w__1102, w__1103, w__1104;
  wire w__1105, w__1106, w__1107, w__1108, w__1109, w__1110, w__1111, w__1112;
  wire w__1113, w__1114, w__1115, w__1116, w__1117, w__1118, w__1119, w__1120;
  wire w__1121, w__1122, w__1123, w__1124, w__1125, w__1126, w__1127, w__1128;
  wire w__1129, w__1130, w__1131, w__1132, w__1133, w__1134, w__1135, w__1136;
  wire w__1137, w__1138, w__1139, w__1140, w__1141, w__1142, w__1143, w__1144;
  wire w__1145, w__1146, w__1147, w__1148, w__1149, w__1150, w__1151, w__1152;
  wire w__1153, w__1154, w__1155, w__1156, w__1157, w__1158, w__1159, w__1160;
  wire w__1161, w__1162, w__1163, w__1164, w__1165, w__1166, w__1167, w__1168;
  wire w__1169, w__1170, w__1171, w__1172, w__1173, w__1174, w__1175, w__1176;
  wire w__1177, w__1178, w__1179, w__1180, w__1181, w__1182, w__1183, w__1184;
  wire w__1185, w__1186, w__1187, w__1188, w__1189, w__1190, w__1191, w__1192;
  wire w__1193, w__1194, w__1195, w__1196, w__1197, w__1198, w__1199, w__1200;
  wire w__1201, w__1202, w__1203, w__1204, w__1205, w__1206, w__1207, w__1208;
  wire w__1209, w__1210, w__1211, w__1212, w__1213, w__1214, w__1215, w__1216;
  wire w__1217, w__1218, w__1219, w__1220, w__1221, w__1222, w__1223, w__1224;
  wire w__1225, w__1226, w__1227, w__1228, w__1229, w__1230, w__1231, w__1232;
  wire w__1233, w__1234, w__1235, w__1236, w__1237, w__1238, w__1239, w__1240;
  wire w__1241, w__1242, w__1243, w__1244, w__1245, w__1246, w__1247, w__1248;
  wire w__1249, w__1250, w__1251, w__1252, w__1253, w__1254, w__1255, w__1256;
  wire w__1257, w__1258, w__1259, w__1260, w__1261, w__1262, w__1263, w__1264;
  wire w__1265, w__1266, w__1267, w__1268, w__1269, w__1270, w__1271, w__1272;
  wire w__1273, w__1274, w__1275, w__1276, w__1277, w__1278, w__1279, w__1280;
  wire w__1281, w__1282, w__1283, w__1284, w__1285, w__1286, w__1287, w__1288;
  wire w__1289, w__1290, w__1291, w__1292, w__1293, w__1294, w__1295, w__1296;
  wire w__1297, w__1298, w__1299, w__1300, w__1301, w__1302, w__1303, w__1304;
  wire w__1305, w__1306, w__1307, w__1308, w__1309, w__1310, w__1311, w__1312;
  wire w__1313, w__1314, w__1315, w__1316, w__1317, w__1318, w__1319, w__1320;
  wire w__1321, w__1322, w__1323, w__1324, w__1325, w__1326, w__1327, w__1328;
  wire w__1329, w__1330, w__1331, w__1332, w__1333, w__1334, w__1335, w__1336;
  wire w__1337, w__1338, w__1339, w__1340, w__1341, w__1342, w__1343, w__1344;
  wire w__1345, w__1346, w__1347, w__1348, w__1349, w__1350, w__1351, w__1352;
  wire w__1353, w__1354, w__1355, w__1356, w__1357, w__1358, w__1359, w__1360;
  wire w__1361, w__1362, w__1363, w__1364, w__1365, w__1366, w__1367, w__1368;
  wire w__1369, w__1370, w__1371, w__1372, w__1373, w__1374, w__1375, w__1376;
  wire w__1377, w__1378, w__1379, w__1380, w__1381, w__1382, w__1383, w__1384;
  wire w__1385, w__1386, w__1387, w__1388, w__1389, w__1390, w__1391, w__1392;
  wire w__1393, w__1394, w__1395, w__1396, w__1397, w__1398, w__1399, w__1400;
  wire w__1401, w__1402, w__1403, w__1404, w__1405, w__1406, w__1407, w__1408;
  wire w__1409, w__1410, w__1411, w__1412, w__1413, w__1414, w__1415, w__1416;
  wire w__1417, w__1418, w__1419, w__1420, w__1421, w__1422, w__1423, w__1424;
  wire w__1425, w__1426, w__1427, w__1428, w__1429, w__1430, w__1431, w__1432;
  wire w__1433, w__1434, w__1435, w__1436, w__1437, w__1438, w__1439, w__1440;
  wire w__1441, w__1442, w__1443, w__1444, w__1445, w__1446, w__1447, w__1448;
  wire w__1449, w__1450, w__1451, w__1452, w__1453, w__1454, w__1455, w__1456;
  wire w__1457, w__1458, w__1459, w__1460, w__1461, w__1462, w__1463, w__1464;
  wire w__1465, w__1466, w__1467, w__1468, w__1469, w__1470, w__1471, w__1472;
  wire w__1473, w__1474, w__1475, w__1476, w__1477, w__1478, w__1479, w__1480;
  wire w__1481, w__1482, w__1483, w__1484, w__1485, w__1486, w__1487, w__1488;
  wire w__1489, w__1490, w__1491, w__1492, w__1493, w__1494, w__1495, w__1496;
  wire w__1497, w__1498, w__1499, w__1500, w__1501, w__1502, w__1503, w__1504;
  wire w__1505, w__1506, w__1507, w__1508, w__1509, w__1510, w__1511, w__1512;
  wire w__1513, w__1514, w__1515, w__1516, w__1517, w__1518, w__1519, w__1520;
  wire w__1521, w__1522, w__1523, w__1524, w__1525, w__1526, w__1527, w__1528;
  wire w__1529, w__1530, w__1531, w__1532, w__1533, w__1534, w__1535, w__1536;
  wire w__1537, w__1538, w__1539, w__1540, w__1541, w__1542, w__1543, w__1544;
  wire w__1545, w__1546, w__1547, w__1548, w__1549, w__1550, w__1551, w__1552;
  wire w__1553, w__1554, w__1555, w__1556, w__1557, w__1558, w__1559, w__1560;
  wire w__1561, w__1562, w__1563, w__1564, w__1565, w__1566, w__1567, w__1568;
  wire w__1569, w__1570, w__1571, w__1572, w__1573, w__1574, w__1575, w__1576;
  wire w__1577, w__1578, w__1579, w__1580, w__1581, w__1582, w__1583, w__1584;
  wire w__1585, w__1586, w__1587, w__1588, w__1589, w__1590, w__1591, w__1592;
  wire w__1593, w__1594, w__1595, w__1596, w__1597, w__1598, w__1599, w__1600;
  wire w__1601, w__1602, w__1603, w__1604, w__1605, w__1606, w__1607, w__1608;
  wire w__1609, w__1610, w__1611, w__1612, w__1613, w__1614, w__1615, w__1616;
  wire w__1617, w__1618, w__1619, w__1620, w__1621, w__1622, w__1623, w__1624;
  wire w__1625, w__1626, w__1627, w__1628, w__1629, w__1630, w__1631, w__1632;
  wire w__1633, w__1634, w__1635, w__1636, w__1637, w__1638, w__1639, w__1640;
  wire w__1641, w__1642, w__1643, w__1644, w__1645, w__1646, w__1647, w__1648;
  wire w__1649, w__1650, w__1651, w__1652, w__1653, w__1654, w__1655, w__1656;
  wire w__1657, w__1658, w__1659, w__1660, w__1661, w__1662, w__1663, w__1664;
  wire w__1665, w__1666, w__1667, w__1668, w__1669, w__1670, w__1671, w__1672;
  wire w__1673, w__1674, w__1675, w__1676, w__1677, w__1678, w__1679, w__1680;
  wire w__1681, w__1682, w__1683, w__1684, w__1685, w__1686, w__1687, w__1688;
  wire w__1689, w__1690, w__1691, w__1692, w__1693, w__1694, w__1695, w__1696;
  wire w__1697, w__1698, w__1699, w__1700, w__1701, w__1702, w__1703, w__1704;
  wire w__1705, w__1706, w__1707, w__1708, w__1709, w__1710, w__1711, w__1712;
  wire w__1713, w__1714, w__1715, w__1716, w__1717, w__1718, w__1719, w__1720;
  wire w__1721, w__1722, w__1723, w__1724, w__1725, w__1726, w__1727, w__1728;
  wire w__1729, w__1730, w__1731, w__1732, w__1733, w__1734, w__1735, w__1736;
  wire w__1737, w__1738, w__1739, w__1740, w__1741, w__1742, w__1743, w__1744;
  wire w__1745, w__1746, w__1747, w__1748, w__1749, w__1750, w__1751, w__1752;
  wire w__1753, w__1754, w__1755, w__1756, w__1757, w__1758, w__1759, w__1760;
  wire w__1761, w__1762, w__1763, w__1764, w__1765, w__1766, w__1767, w__1768;
  wire w__1769, w__1770, w__1771, w__1772, w__1773, w__1774, w__1775, w__1776;
  wire w__1777, w__1778, w__1779, w__1780, w__1781, w__1782, w__1783, w__1784;
  wire w__1785, w__1786, w__1787, w__1788, w__1789, w__1790, w__1791, w__1792;
  wire w__1793, w__1794, w__1795, w__1796, w__1797, w__1798, w__1799, w__1800;
  wire w__1801, w__1802, w__1803, w__1804, w__1805, w__1806, w__1807, w__1808;
  wire w__1809, w__1810, w__1811, w__1812, w__1813, w__1814, w__1815, w__1816;
  wire w__1817, w__1818, w__1819, w__1820, w__1821, w__1822, w__1823, w__1824;
  wire w__1825, w__1826, w__1827, w__1828, w__1829, w__1830, w__1831, w__1832;
  wire w__1833, w__1834, w__1835, w__1836, w__1837, w__1838, w__1839, w__1840;
  wire w__1841, w__1842, w__1843, w__1844, w__1845, w__1846, w__1847, w__1848;
  wire w__1849, w__1850, w__1851, w__1852, w__1853, w__1854, w__1855, w__1856;
  wire w__1857, w__1858, w__1859, w__1860, w__1861, w__1862, w__1863, w__1864;
  wire w__1865, w__1866, w__1867, w__1868, w__1869, w__1870, w__1871, w__1872;
  wire w__1873, w__1874, w__1875, w__1876, w__1877, w__1878, w__1879, w__1880;
  wire w__1881, w__1882, w__1883, w__1884, w__1885, w__1886, w__1887, w__1888;
  wire w__1889, w__1890, w__1891, w__1892, w__1893, w__1894, w__1895, w__1896;
  wire w__1897, w__1898, w__1899, w__1900, w__1901, w__1902, w__1903, w__1904;
  wire w__1905, w__1906, w__1907, w__1908, w__1909, w__1910, w__1911, w__1912;
  wire w__1913, w__1914, w__1915, w__1916, w__1917, w__1918, w__1919, w__1920;
  wire w__1921, w__1922, w__1923, w__1924, w__1925, w__1926, w__1927, w__1928;
  wire w__1929, w__1930, w__1931, w__1932, w__1933, w__1934, w__1935, w__1936;
  wire w__1937, w__1938, w__1939, w__1940, w__1941, w__1942, w__1943, w__1944;
  wire w__1945, w__1946, w__1947, w__1948, w__1949, w__1950, w__1951, w__1952;
  wire w__1953, w__1954, w__1955, w__1956, w__1957, w__1958, w__1959, w__1960;
  wire w__1961, w__1962, w__1963, w__1964, w__1965, w__1966, w__1967, w__1968;
  wire w__1969, w__1970, w__1971, w__1972, w__1973, w__1974, w__1975, w__1976;
  wire w__1977, w__1978, w__1979, w__1980, w__1981, w__1982, w__1983, w__1984;
  wire w__1985, w__1986, w__1987, w__1988, w__1989, w__1990, w__1991, w__1992;
  wire w__1993, w__1994, w__1995, w__1996, w__1997, w__1998, w__1999, w__2000;
  wire w__2001, w__2002, w__2003, w__2004, w__2005, w__2006, w__2007, w__2008;
  wire w__2009, w__2010, w__2011, w__2012, w__2013, w__2014, w__2015, w__2016;
  wire w__2017, w__2018, w__2019, w__2020, w__2021, w__2022, w__2023, w__2024;
  wire w__2025, w__2026, w__2027, w__2028, w__2029, w__2030, w__2031, w__2032;
  wire w__2033, w__2034, w__2035, w__2036, w__2037, w__2038, w__2039, w__2040;
  wire w__2041, w__2042, w__2043, w__2044, w__2045, w__2046, w__2047, w__2048;
  wire w__2049, w__2050, w__2051, w__2052, w__2053, w__2054, w__2055, w__2056;
  wire w__2057, w__2058, w__2059, w__2060, w__2061, w__2062, w__2063, w__2064;
  wire w__2065, w__2066, w__2067, w__2068, w__2069, w__2070, w__2071, w__2072;
  wire w__2073, w__2074, w__2075, w__2076, w__2077, w__2078, w__2079, w__2080;
  wire w__2081, w__2082, w__2083, w__2084, w__2085, w__2086, w__2087, w__2088;
  wire w__2089, w__2090, w__2091, w__2092, w__2093, w__2094, w__2095, w__2096;
  wire w__2097, w__2098, w__2099, w__2100, w__2101, w__2102, w__2103, w__2104;
  wire w__2105, w__2106, w__2107, w__2108, w__2109, w__2110, w__2111, w__2112;
  wire w__2113, w__2114, w__2115, w__2116, w__2117, w__2118, w__2119, w__2120;
  wire w__2121, w__2122, w__2123, w__2124, w__2125, w__2126, w__2127, w__2128;
  wire w__2129, w__2130, w__2131, w__2132, w__2133, w__2134, w__2135, w__2136;
  wire w__2137, w__2138, w__2139, w__2140, w__2141, w__2142, w__2143, w__2144;
  wire w__2145, w__2146, w__2147, w__2148, w__2149, w__2150, w__2151, w__2152;
  wire w__2153, w__2154, w__2155, w__2156, w__2157, w__2158, w__2159, w__2160;
  wire w__2161, w__2162, w__2163, w__2164, w__2165, w__2166, w__2167, w__2168;
  wire w__2169, w__2170, w__2171, w__2172, w__2173, w__2174, w__2175, w__2176;
  wire w__2177, w__2178, w__2179, w__2180, w__2181, w__2182, w__2183, w__2184;
  wire w__2185, w__2186, w__2187, w__2188, w__2189, w__2190, w__2191, w__2192;
  wire w__2193, w__2194, w__2195, w__2196, w__2197, w__2198, w__2199, w__2200;
  wire w__2201, w__2202, w__2203, w__2204, w__2205, w__2206, w__2207, w__2208;
  wire w__2209, w__2210, w__2211, w__2212, w__2213, w__2214, w__2215, w__2216;
  wire w__2217, w__2218, w__2219, w__2220, w__2221, w__2222, w__2223, w__2224;
  wire w__2225, w__2226, w__2227, w__2228, w__2229, w__2230, w__2231, w__2232;
  wire w__2233, w__2234, w__2235, w__2236, w__2237, w__2238, w__2239, w__2240;
  wire w__2241, w__2242, w__2243, w__2244, w__2245, w__2246, w__2247, w__2248;
  wire w__2249, w__2250, w__2251, w__2252, w__2253, w__2254, w__2255, w__2256;
  wire w__2257, w__2258, w__2259, w__2260, w__2261, w__2262, w__2263, w__2264;
  wire w__2265, w__2266, w__2267, w__2268, w__2269, w__2270, w__2271, w__2272;
  wire w__2273, w__2274, w__2275, w__2276, w__2277, w__2278, w__2279, w__2280;
  wire w__2281, w__2282, w__2283, w__2284, w__2285, w__2286, w__2287, w__2288;
  wire w__2289, w__2290, w__2291, w__2292, w__2293, w__2294, w__2295, w__2296;
  wire w__2297, w__2298, w__2299, w__2300, w__2301, w__2302, w__2303, w__2304;
  wire w__2305, w__2306, w__2307, w__2308, w__2309, w__2310, w__2311, w__2312;
  wire w__2313, w__2314, w__2315, w__2316, w__2317, w__2318, w__2319, w__2320;
  wire w__2321, w__2322, w__2323, w__2324, w__2325, w__2326, w__2327, w__2328;
  wire w__2329, w__2330, w__2331, w__2332, w__2333, w__2334, w__2335, w__2336;
  wire w__2337, w__2338, w__2339, w__2340, w__2341, w__2342, w__2343, w__2344;
  wire w__2345, w__2346, w__2347, w__2348, w__2349, w__2350, w__2351, w__2352;
  wire w__2353, w__2354, w__2355, w__2356, w__2357, w__2358, w__2359, w__2360;
  wire w__2361, w__2362, w__2363, w__2364, w__2365, w__2366, w__2367, w__2368;
  wire w__2369, w__2370, w__2371, w__2372, w__2373, w__2374, w__2375, w__2376;
  wire w__2377, w__2378, w__2379, w__2380, w__2381, w__2382, w__2383, w__2384;
  wire w__2385, w__2386, w__2387, w__2388, w__2389, w__2390, w__2391, w__2392;
  wire w__2393, w__2394, w__2395, w__2396, w__2397, w__2398, w__2399, w__2400;
  wire w__2401, w__2402, w__2403, w__2404, w__2405, w__2406, w__2407, w__2408;
  wire w__2409, w__2410, w__2411, w__2412, w__2413, w__2414, w__2415, w__2416;
  wire w__2417, w__2418, w__2419, w__2420, w__2421, w__2422, w__2423, w__2424;
  wire w__2425, w__2426, w__2427, w__2428, w__2429, w__2430, w__2431, w__2432;
  wire w__2433, w__2434, w__2435, w__2436, w__2437, w__2438, w__2439, w__2440;
  wire w__2441, w__2442, w__2443, w__2444, w__2445, w__2446, w__2447, w__2448;
  wire w__2449, w__2450, w__2451, w__2452, w__2453, w__2454, w__2455, w__2456;
  wire w__2457, w__2458, w__2459, w__2460, w__2461, w__2462, w__2463, w__2464;
  wire w__2465, w__2466, w__2467, w__2468, w__2469, w__2470, w__2471, w__2472;
  wire w__2473, w__2474, w__2475, w__2476, w__2477, w__2478, w__2479, w__2480;
  wire w__2481, w__2482, w__2483, w__2484, w__2485, w__2486, w__2487, w__2488;
  wire w__2489, w__2490, w__2491, w__2492, w__2493, w__2494, w__2495, w__2496;
  wire w__2497, w__2498, w__2499, w__2500, w__2501, w__2502, w__2503, w__2504;
  wire w__2505, w__2506, w__2507, w__2508, w__2509, w__2510, w__2511, w__2512;
  wire w__2513, w__2514, w__2515, w__2516, w__2517, w__2518, w__2519, w__2520;
  wire w__2521, w__2522, w__2523, w__2524, w__2525, w__2526, w__2527, w__2528;
  wire w__2529, w__2530, w__2531, w__2532, w__2533, w__2534, w__2535, w__2536;
  wire w__2537, w__2538, w__2539, w__2540, w__2541, w__2542, w__2543, w__2544;
  wire w__2545, w__2546, w__2547, w__2548, w__2549, w__2550, w__2551, w__2552;
  wire w__2553, w__2554, w__2555, w__2556, w__2557, w__2558, w__2559, w__2560;
  wire w__2561, w__2562, w__2563, w__2564, w__2565, w__2566, w__2567, w__2568;
  wire w__2569, w__2570, w__2571, w__2572, w__2573, w__2574, w__2575, w__2576;
  wire w__2577, w__2578, w__2579, w__2580, w__2581, w__2582, w__2583, w__2584;
  wire w__2585, w__2586, w__2587, w__2588, w__2589, w__2590, w__2591, w__2592;
  wire w__2593, w__2594, w__2595, w__2596, w__2597, w__2598, w__2599, w__2600;
  wire w__2601, w__2602, w__2603, w__2604, w__2605, w__2606, w__2607, w__2608;
  wire w__2609, w__2610, w__2611, w__2612, w__2613, w__2614, w__2615, w__2616;
  wire w__2617, w__2618, w__2619, w__2620, w__2621, w__2622, w__2623, w__2624;
  wire w__2625, w__2626, w__2627, w__2628, w__2629, w__2630, w__2631, w__2632;
  wire w__2633, w__2634, w__2635, w__2636, w__2637, w__2638, w__2639, w__2640;
  wire w__2641, w__2642, w__2643, w__2644, w__2645, w__2646, w__2647, w__2648;
  wire w__2649, w__2650, w__2651, w__2652, w__2653, w__2654, w__2655, w__2656;
  wire w__2657, w__2658, w__2659, w__2660, w__2661, w__2662, w__2663, w__2664;
  wire w__2665, w__2666, w__2667, w__2668, w__2669, w__2670, w__2671, w__2672;
  wire w__2673, w__2674, w__2675, w__2676, w__2677, w__2678, w__2679, w__2680;
  wire w__2681, w__2682, w__2683, w__2684, w__2685, w__2686, w__2687, w__2688;
  wire w__2689, w__2690, w__2691, w__2692, w__2693, w__2694, w__2695, w__2696;
  wire w__2697, w__2698, w__2699, w__2700, w__2701, w__2702, w__2703, w__2704;
  wire w__2705, w__2706, w__2707, w__2708, w__2709, w__2710, w__2711, w__2712;
  wire w__2713, w__2714, w__2715, w__2716, w__2717, w__2718, w__2719, w__2720;
  wire w__2721, w__2722, w__2723, w__2724, w__2725, w__2726, w__2727, w__2728;
  wire w__2729, w__2730, w__2731, w__2732, w__2733, w__2734, w__2735, w__2736;
  wire w__2737, w__2738, w__2739, w__2740, w__2741, w__2742, w__2743, w__2744;
  wire w__2745, w__2746, w__2747, w__2748, w__2749, w__2750, w__2751, w__2752;
  wire w__2753, w__2754, w__2755, w__2756, w__2757, w__2758, w__2759, w__2760;
  wire w__2761, w__2762, w__2763, w__2764, w__2765, w__2766, w__2767, w__2768;
  wire w__2769, w__2770, w__2771, w__2772, w__2773, w__2774, w__2775, w__2776;
  wire w__2777, w__2778, w__2779, w__2780, w__2781, w__2782, w__2783, w__2784;
  wire w__2785, w__2786, w__2787, w__2788, w__2789, w__2790, w__2791, w__2792;
  wire w__2793, w__2794, w__2795, w__2796, w__2797, w__2798, w__2799, w__2800;
  wire w__2801, w__2802, w__2803, w__2804, w__2805, w__2806, w__2807, w__2808;
  wire w__2809, w__2810, w__2811, w__2812, w__2813, w__2814, w__2815, w__2816;
  wire w__2817, w__2818, w__2819, w__2820, w__2821, w__2822, w__2823, w__2824;
  wire w__2825, w__2826, w__2827, w__2828, w__2829, w__2830, w__2831, w__2832;
  wire w__2833, w__2834, w__2835, w__2836, w__2837, w__2838, w__2839, w__2840;
  wire w__2841, w__2842, w__2843, w__2844, w__2845, w__2846, w__2847, w__2848;
  wire w__2849, w__2850, w__2851, w__2852, w__2853, w__2854, w__2855, w__2856;
  wire w__2857, w__2858, w__2859, w__2860, w__2861, w__2862, w__2863, w__2864;
  wire w__2865, w__2866, w__2867, w__2868, w__2869, w__2870, w__2871, w__2872;
  wire w__2873, w__2874, w__2875, w__2876, w__2877, w__2878, w__2879, w__2880;
  wire w__2881, w__2882, w__2883, w__2884, w__2885, w__2886, w__2887, w__2888;
  wire w__2889, w__2890, w__2891, w__2892, w__2893, w__2894, w__2895, w__2896;
  wire w__2897, w__2898, w__2899, w__2900, w__2901, w__2902, w__2903, w__2904;
  wire w__2905, w__2906, w__2907, w__2908, w__2909, w__2910, w__2911, w__2912;
  wire w__2913, w__2914, w__2915, w__2916, w__2917, w__2918, w__2919, w__2920;
  wire w__2921, w__2922, w__2923, w__2924, w__2925, w__2926, w__2927, w__2928;
  wire w__2929, w__2930, w__2931, w__2932, w__2933, w__2934, w__2935, w__2936;
  wire w__2937, w__2938, w__2939, w__2940, w__2941, w__2942, w__2943, w__2944;
  wire w__2945, w__2946, w__2947, w__2948, w__2949, w__2950, w__2951, w__2952;
  wire w__2953, w__2954, w__2955, w__2956, w__2957, w__2958, w__2959, w__2960;
  wire w__2961, w__2962, w__2963, w__2964, w__2965, w__2966, w__2967, w__2968;
  wire w__2969, w__2970, w__2971, w__2972, w__2973, w__2974, w__2975, w__2976;
  wire w__2977, w__2978, w__2979, w__2980, w__2981, w__2982, w__2983, w__2984;
  wire w__2985, w__2986, w__2987, w__2988, w__2989, w__2990, w__2991, w__2992;
  wire w__2993, w__2994, w__2995, w__2996, w__2997, w__2998, w__2999, w__3000;
  wire w__3001, w__3002, w__3003, w__3004, w__3005, w__3006, w__3007, w__3008;
  wire w__3009, w__3010, w__3011, w__3012, w__3013, w__3014, w__3015, w__3016;
  wire w__3017, w__3018, w__3019, w__3020, w__3021, w__3022, w__3023, w__3024;
  wire w__3025, w__3026, w__3027, w__3028, w__3029, w__3030, w__3031, w__3032;
  wire w__3033, w__3034, w__3035, w__3036, w__3037, w__3038, w__3039, w__3040;
  wire w__3041, w__3042, w__3043, w__3044, w__3045, w__3046, w__3047, w__3048;
  wire w__3049, w__3050, w__3051, w__3052, w__3053, w__3054, w__3055, w__3056;
  wire w__3057, w__3058, w__3059, w__3060, w__3061, w__3062, w__3063, w__3064;
  wire w__3065, w__3066, w__3067, w__3068, w__3069, w__3070, w__3071, w__3072;
  wire w__3073, w__3074, w__3075, w__3076, w__3077, w__3078, w__3079, w__3080;
  wire w__3081, w__3082, w__3083, w__3084, w__3085, w__3086, w__3087, w__3088;
  wire w__3089, w__3090, w__3091, w__3092, w__3093, w__3094, w__3095, w__3096;
  wire w__3097, w__3098, w__3099, w__3100, w__3101, w__3102, w__3103, w__3104;
  wire w__3105, w__3106, w__3107, w__3108, w__3109, w__3110, w__3111, w__3112;
  wire w__3113, w__3114, w__3115, w__3116, w__3117, w__3118, w__3119, w__3120;
  wire w__3121, w__3122, w__3123, w__3124, w__3125, w__3126, w__3127, w__3128;
  wire w__3129, w__3130, w__3131, w__3132, w__3133, w__3134, w__3135, w__3136;
  wire w__3137, w__3138, w__3139, w__3140, w__3141, w__3142, w__3143, w__3144;
  wire w__3145, w__3146, w__3147, w__3148, w__3149, w__3150, w__3151, w__3152;
  wire w__3153, w__3154, w__3155, w__3156, w__3157, w__3158, w__3159, w__3160;
  wire w__3161, w__3162, w__3163, w__3164, w__3165, w__3166, w__3167, w__3168;
  wire w__3169, w__3170, w__3171, w__3172, w__3173, w__3174, w__3175, w__3176;
  wire w__3177, w__3178, w__3179, w__3180, w__3181, w__3182, w__3183, w__3184;
  wire w__3185, w__3186, w__3187, w__3188, w__3189, w__3190, w__3191, w__3192;
  wire w__3193, w__3194, w__3195, w__3196, w__3197, w__3198, w__3199, w__3200;
  wire w__3201, w__3202, w__3203, w__3204, w__3205, w__3206, w__3207, w__3208;
  wire w__3209, w__3210, w__3211, w__3212, w__3213, w__3214, w__3215, w__3216;
  wire w__3217, w__3218, w__3219, w__3220, w__3221, w__3222, w__3223, w__3224;
  wire w__3225, w__3226, w__3227, w__3228, w__3229, w__3230, w__3231, w__3232;
  wire w__3233, w__3234, w__3235, w__3236, w__3237, w__3238, w__3239, w__3240;
  wire w__3241, w__3242, w__3243, w__3244, w__3245, w__3246, w__3247, w__3248;
  wire w__3249, w__3250, w__3251, w__3252, w__3253, w__3254, w__3255, w__3256;
  wire w__3257, w__3258, w__3259, w__3260, w__3261, w__3262, w__3263, w__3264;
  wire w__3265, w__3266, w__3267, w__3268, w__3269, w__3270, w__3271, w__3272;
  wire w__3273, w__3274, w__3275, w__3276, w__3277, w__3278, w__3279, w__3280;
  wire w__3281, w__3282, w__3283, w__3284, w__3285, w__3286, w__3287, w__3288;
  wire w__3289, w__3290, w__3291, w__3292, w__3293, w__3294, w__3295, w__3296;
  wire w__3297, w__3298, w__3299, w__3300, w__3301, w__3302, w__3303, w__3304;
  wire w__3305, w__3306, w__3307, w__3308, w__3309, w__3310, w__3311, w__3312;
  wire w__3313, w__3314, w__3315, w__3316, w__3317, w__3318, w__3319, w__3320;
  wire w__3321, w__3322, w__3323, w__3324, w__3325, w__3326, w__3327, w__3328;
  wire w__3329, w__3330, w__3331, w__3332, w__3333, w__3334, w__3335, w__3336;
  wire w__3337, w__3338, w__3339, w__3340, w__3341, w__3342, w__3343, w__3344;
  wire w__3345, w__3346, w__3347, w__3348, w__3349, w__3350, w__3351, w__3352;
  wire w__3353, w__3354, w__3355, w__3356, w__3357, w__3358, w__3359, w__3360;
  wire w__3361, w__3362, w__3363, w__3364, w__3365, w__3366, w__3367, w__3368;
  wire w__3369, w__3370, w__3371, w__3372, w__3373, w__3374, w__3375, w__3376;
  wire w__3377, w__3378, w__3379, w__3380, w__3381, w__3382, w__3383, w__3384;
  wire w__3385, w__3386, w__3387, w__3388, w__3389, w__3390, w__3391, w__3392;
  wire w__3393, w__3394, w__3395, w__3396, w__3397, w__3398, w__3399, w__3400;
  wire w__3401, w__3402, w__3403, w__3404, w__3405, w__3406, w__3407, w__3408;
  wire w__3409, w__3410, w__3411, w__3412, w__3413, w__3414, w__3415, w__3416;
  wire w__3417, w__3418, w__3419, w__3420, w__3421, w__3422, w__3423, w__3424;
  wire w__3425, w__3426, w__3427, w__3428, w__3429, w__3430, w__3431, w__3432;
  wire w__3433, w__3434, w__3435, w__3436, w__3437, w__3438, w__3439, w__3440;
  wire w__3441, w__3442, w__3443, w__3444, w__3445, w__3446, w__3447, w__3448;
  wire w__3449, w__3450, w__3451, w__3452, w__3453, w__3454, w__3455, w__3456;
  wire w__3457, w__3458, w__3459, w__3460, w__3461, w__3462, w__3463, w__3464;
  wire w__3465, w__3466, w__3467, w__3468, w__3469, w__3470, w__3471, w__3472;
  wire w__3473, w__3474, w__3475, w__3476, w__3477, w__3478, w__3479, w__3480;
  wire w__3481, w__3482, w__3483, w__3484, w__3485, w__3486, w__3487, w__3488;
  wire w__3489, w__3490, w__3491, w__3492, w__3493, w__3494, w__3495, w__3496;
  wire w__3497, w__3498, w__3499, w__3500, w__3501, w__3502, w__3503, w__3504;
  wire w__3505, w__3506, w__3507, w__3508, w__3509, w__3510, w__3511, w__3512;
  wire w__3513, w__3514, w__3515, w__3516, w__3517, w__3518, w__3519, w__3520;
  wire w__3521, w__3522, w__3523, w__3524, w__3525, w__3526, w__3527, w__3528;
  wire w__3529, w__3530, w__3531, w__3532, w__3533, w__3534, w__3535, w__3536;
  wire w__3537, w__3538, w__3539, w__3540, w__3541, w__3542, w__3543, w__3544;
  wire w__3545, w__3546, w__3547, w__3548, w__3549, w__3550, w__3551, w__3552;
  wire w__3553, w__3554, w__3555, w__3556, w__3557, w__3558, w__3559, w__3560;
  wire w__3561, w__3562, w__3563, w__3564, w__3565, w__3566, w__3567, w__3568;
  wire w__3569, w__3570, w__3571, w__3572, w__3573, w__3574, w__3575, w__3576;
  wire w__3577, w__3578, w__3579, w__3580, w__3581, w__3582, w__3583, w__3584;
  wire w__3585, w__3586, w__3587, w__3588, w__3589, w__3590, w__3591, w__3592;
  wire w__3593, w__3594, w__3595, w__3596, w__3597, w__3598, w__3599, w__3600;
  wire w__3601, w__3602, w__3603, w__3604, w__3605, w__3606, w__3607, w__3608;
  wire w__3609, w__3610, w__3611, w__3612, w__3613, w__3614, w__3615, w__3616;
  wire w__3617, w__3618, w__3619, w__3620, w__3621, w__3622, w__3623, w__3624;
  wire w__3625, w__3626, w__3627, w__3628, w__3629, w__3630, w__3631, w__3632;
  wire w__3633, w__3634, w__3635, w__3636, w__3637, w__3638, w__3639, w__3640;
  wire w__3641, w__3642, w__3643, w__3644, w__3645, w__3646, w__3647, w__3648;
  wire w__3649, w__3650, w__3651, w__3652, w__3653, w__3654, w__3655, w__3656;
  wire w__3657, w__3658, w__3659, w__3660, w__3661, w__3662, w__3663, w__3664;
  wire w__3665, w__3666, w__3667, w__3668, w__3669, w__3670, w__3671, w__3672;
  wire w__3673, w__3674, w__3675, w__3676, w__3677, w__3678, w__3679, w__3680;
  wire w__3681, w__3682, w__3683, w__3684, w__3685, w__3686, w__3687, w__3688;
  wire w__3689, w__3690, w__3691, w__3692, w__3693, w__3694, w__3695, w__3696;
  wire w__3697, w__3698, w__3699, w__3700, w__3701, w__3702, w__3703, w__3704;
  wire w__3705, w__3706, w__3707, w__3708, w__3709, w__3710, w__3711, w__3712;
  wire w__3713, w__3714, w__3715, w__3716, w__3717, w__3718, w__3719, w__3720;
  wire w__3721, w__3722, w__3723, w__3724, w__3725, w__3726, w__3727, w__3728;
  wire w__3729, w__3730, w__3731, w__3732, w__3733, w__3734, w__3735, w__3736;
  wire w__3737, w__3738, w__3739, w__3740, w__3741, w__3742, w__3743, w__3744;
  wire w__3745, w__3746, w__3747, w__3748, w__3749, w__3750, w__3751, w__3752;
  wire w__3753, w__3754, w__3755, w__3756, w__3757, w__3758, w__3759, w__3760;
  wire w__3761, w__3762, w__3763, w__3764, w__3765, w__3766, w__3767, w__3768;
  wire w__3769, w__3770, w__3771, w__3772, w__3773, w__3774, w__3775, w__3776;
  wire w__3777, w__3778, w__3779, w__3780, w__3781, w__3782, w__3783, w__3784;
  wire w__3785, w__3786, w__3787, w__3788, w__3789, w__3790, w__3791, w__3792;
  wire w__3793, w__3794, w__3795, w__3796, w__3797, w__3798, w__3799, w__3800;
  wire w__3801, w__3802, w__3803, w__3804, w__3805, w__3806, w__3807, w__3808;
  wire w__3809, w__3810, w__3811, w__3812, w__3813, w__3814, w__3815, w__3816;
  wire w__3817, w__3818, w__3819, w__3820, w__3821, w__3822, w__3823, w__3824;
  wire w__3825, w__3826, w__3827, w__3828, w__3829, w__3830, w__3831, w__3832;
  wire w__3833, w__3834, w__3835, w__3836, w__3837, w__3838, w__3839, w__3840;
  wire w__3841, w__3842, w__3843, w__3844, w__3845, w__3846, w__3847, w__3848;
  wire w__3849, w__3850, w__3851, w__3852, w__3853, w__3854, w__3855, w__3856;
  wire w__3857, w__3858, w__3859, w__3860, w__3861, w__3862, w__3863, w__3864;
  wire w__3865, w__3866, w__3867, w__3868, w__3869, w__3870, w__3871, w__3872;
  wire w__3873, w__3874, w__3875, w__3876, w__3877, w__3878, w__3879, w__3880;
  wire w__3881, w__3882, w__3883, w__3884, w__3885, w__3886, w__3887, w__3888;
  wire w__3889, w__3890, w__3891, w__3892, w__3893, w__3894, w__3895, w__3896;
  wire w__3897, w__3898, w__3899, w__3900, w__3901, w__3902, w__3903, w__3904;
  wire w__3905, w__3906, w__3907, w__3908, w__3909, w__3910, w__3911, w__3912;
  wire w__3913, w__3914, w__3915, w__3916, w__3917, w__3918, w__3919, w__3920;
  wire w__3921, w__3922, w__3923, w__3924, w__3925, w__3926, w__3927, w__3928;
  wire w__3929, w__3930, w__3931, w__3932, w__3933, w__3934, w__3935, w__3936;
  wire w__3937, w__3938, w__3939, w__3940, w__3941, w__3942, w__3943, w__3944;
  wire w__3945, w__3946, w__3947, w__3948, w__3949, w__3950, w__3951, w__3952;
  wire w__3953, w__3954, w__3955, w__3956, w__3957, w__3958, w__3959, w__3960;
  wire w__3961, w__3962, w__3963, w__3964, w__3965, w__3966, w__3967, w__3968;
  wire w__3969, w__3970, w__3971, w__3972, w__3973, w__3974, w__3975, w__3976;
  wire w__3977, w__3978, w__3979, w__3980, w__3981, w__3982, w__3983, w__3984;
  wire w__3985, w__3986, w__3987, w__3988, w__3989, w__3990, w__3991, w__3992;
  wire w__3993, w__3994, w__3995, w__3996, w__3997, w__3998, w__3999, w__4000;
  wire w__4001, w__4002, w__4003, w__4004, w__4005, w__4006, w__4007, w__4008;
  wire w__4009, w__4010, w__4011, w__4012, w__4013, w__4014, w__4015, w__4016;
  wire w__4017, w__4018, w__4019, w__4020, w__4021, w__4022, w__4023, w__4024;
  wire w__4025, w__4026, w__4027, w__4028, w__4029, w__4030, w__4031, w__4032;
  wire w__4033, w__4034, w__4035, w__4036, w__4037, w__4038, w__4039, w__4040;
  wire w__4041, w__4042, w__4043, w__4044, w__4045, w__4046, w__4047, w__4048;
  wire w__4049, w__4050, w__4051, w__4052, w__4053, w__4054, w__4055, w__4056;
  wire w__4057, w__4058, w__4059, w__4060, w__4061, w__4062, w__4063, w__4064;
  wire w__4065, w__4066, w__4067, w__4068, w__4069, w__4070, w__4071, w__4072;
  wire w__4073, w__4074, w__4075, w__4076, w__4077, w__4078, w__4079, w__4080;
  wire w__4081, w__4082, w__4083, w__4084, w__4085, w__4086, w__4087, w__4088;
  wire w__4089, w__4090, w__4091, w__4092, w__4093, w__4094, w__4095, w__4096;
  wire w__4097, w__4098, w__4099, w__4100, w__4101, w__4102, w__4103, w__4104;
  wire w__4105, w__4106, w__4107, w__4108, w__4109, w__4110, w__4111, w__4112;
  wire w__4113, w__4114, w__4115, w__4116, w__4117, w__4118, w__4119, w__4120;
  wire w__4121, w__4122, w__4123, w__4124, w__4125, w__4126, w__4127, w__4128;
  wire w__4129, w__4130, w__4131, w__4132, w__4133, w__4134, w__4135, w__4136;
  wire w__4137, w__4138, w__4139, w__4140, w__4141, w__4142, w__4143, w__4144;
  wire w__4145, w__4146, w__4147, w__4148, w__4149, w__4150, w__4151, w__4152;
  wire w__4153, w__4154, w__4155, w__4156, w__4157, w__4158, w__4159, w__4160;
  wire w__4161, w__4162, w__4163, w__4164, w__4165, w__4166, w__4167, w__4168;
  wire w__4169, w__4170, w__4171, w__4172, w__4173, w__4174, w__4175, w__4176;
  wire w__4177, w__4178, w__4179, w__4180, w__4181, w__4182, w__4183, w__4184;
  wire w__4185, w__4186, w__4187, w__4188, w__4189, w__4190, w__4191, w__4192;
  wire w__4193, w__4194, w__4195, w__4196, w__4197, w__4198, w__4199, w__4200;
  wire w__4201, w__4202, w__4203, w__4204, w__4205, w__4206, w__4207, w__4208;
  wire w__4209, w__4210, w__4211, w__4212, w__4213, w__4214, w__4215, w__4216;
  wire w__4217, w__4218, w__4219, w__4220, w__4221, w__4222, w__4223, w__4224;
  wire w__4225, w__4226, w__4227, w__4228, w__4229, w__4230, w__4231, w__4232;
  wire w__4233, w__4234, w__4235, w__4236, w__4237, w__4238, w__4239, w__4240;
  wire w__4241, w__4242, w__4243, w__4244, w__4245, w__4246, w__4247, w__4248;
  wire w__4249, w__4250, w__4251, w__4252, w__4253, w__4254, w__4255, w__4256;
  wire w__4257, w__4258, w__4259, w__4260, w__4261, w__4262, w__4263, w__4264;
  wire w__4265, w__4266, w__4267, w__4268, w__4269, w__4270, w__4271, w__4272;
  wire w__4273, w__4274, w__4275, w__4276, w__4277, w__4278, w__4279, w__4280;
  wire w__4281, w__4282, w__4283, w__4284, w__4285, w__4286, w__4287, w__4288;
  wire w__4289, w__4290, w__4291, w__4292, w__4293, w__4294, w__4295, w__4296;
  wire w__4297, w__4298, w__4299, w__4300, w__4301, w__4302, w__4303, w__4304;
  wire w__4305, w__4306, w__4307, w__4308, w__4309, w__4310, w__4311, w__4312;
  wire w__4313, w__4314, w__4315, w__4316, w__4317, w__4318, w__4319, w__4320;
  wire w__4321, w__4322, w__4323, w__4324, w__4325, w__4326, w__4327, w__4328;
  wire w__4329, w__4330, w__4331, w__4332, w__4333, w__4334, w__4335, w__4336;
  wire w__4337, w__4338, w__4339, w__4340, w__4341, w__4342, w__4343, w__4344;
  wire w__4345, w__4346, w__4347, w__4348, w__4349, w__4350, w__4351, w__4352;
  wire w__4353, w__4354, w__4355, w__4356, w__4357, w__4358, w__4359, w__4360;
  wire w__4361, w__4362, w__4363, w__4364, w__4365, w__4366, w__4367, w__4368;
  wire w__4369, w__4370, w__4371, w__4372, w__4373, w__4374, w__4375, w__4376;
  wire w__4377, w__4378, w__4379, w__4380, w__4381, w__4382, w__4383, w__4384;
  wire w__4385, w__4386, w__4387, w__4388, w__4389, w__4390, w__4391, w__4392;
  wire w__4393, w__4394, w__4395, w__4396, w__4397, w__4398, w__4399, w__4400;
  wire w__4401, w__4402, w__4403, w__4404, w__4405, w__4406, w__4407, w__4408;
  wire w__4409, w__4410, w__4411, w__4412, w__4413, w__4414, w__4415, w__4416;
  wire w__4417, w__4418, w__4419, w__4420, w__4421, w__4422, w__4423, w__4424;
  wire w__4425, w__4426, w__4427, w__4428, w__4429, w__4430, w__4431, w__4432;
  wire w__4433, w__4434, w__4435, w__4436, w__4437, w__4438, w__4439, w__4440;
  wire w__4441, w__4442, w__4443, w__4444, w__4445, w__4446, w__4447, w__4448;
  wire w__4449, w__4450, w__4451, w__4452, w__4453, w__4454, w__4455, w__4456;
  wire w__4457, w__4458, w__4459, w__4460, w__4461, w__4462, w__4463, w__4464;
  wire w__4465, w__4466, w__4467, w__4468, w__4469, w__4470, w__4471, w__4472;
  wire w__4473, w__4474, w__4475, w__4476, w__4477, w__4478, w__4479, w__4480;
  wire w__4481, w__4482, w__4483, w__4484, w__4485, w__4486, w__4487, w__4488;
  wire w__4489, w__4490, w__4491, w__4492, w__4493, w__4494, w__4495, w__4496;
  wire w__4497, w__4498, w__4499, w__4500, w__4501, w__4502, w__4503, w__4504;
  wire w__4505, w__4506, w__4507, w__4508, w__4509, w__4510, w__4511, w__4512;
  wire w__4513, w__4514, w__4515, w__4516, w__4517, w__4518, w__4519, w__4520;
  wire w__4521, w__4522, w__4523, w__4524, w__4525, w__4526, w__4527, w__4528;
  wire w__4529, w__4530, w__4531, w__4532, w__4533, w__4534, w__4535, w__4536;
  wire w__4537, w__4538, w__4539, w__4540, w__4541, w__4542, w__4543, w__4544;
  wire w__4545, w__4546, w__4547, w__4548, w__4549, w__4550, w__4551, w__4552;
  wire w__4553, w__4554, w__4555, w__4556, w__4557, w__4558, w__4559, w__4560;
  wire w__4561, w__4562, w__4563, w__4564, w__4565, w__4566, w__4567, w__4568;
  wire w__4569, w__4570, w__4571, w__4572, w__4573, w__4574, w__4575, w__4576;
  wire w__4577, w__4578, w__4579, w__4580, w__4581, w__4582, w__4583, w__4584;
  wire w__4585, w__4586, w__4587, w__4588, w__4589, w__4590, w__4591, w__4592;
  wire w__4593, w__4594, w__4595, w__4596, w__4597, w__4598, w__4599, w__4600;
  wire w__4601, w__4602, w__4603, w__4604, w__4605, w__4606, w__4607, w__4608;
  wire w__4609, w__4610, w__4611, w__4612, w__4613, w__4614, w__4615, w__4616;
  wire w__4617, w__4618, w__4619, w__4620, w__4621, w__4622, w__4623, w__4624;
  wire w__4625, w__4626, w__4627, w__4628, w__4629, w__4630, w__4631, w__4632;
  wire w__4633, w__4634, w__4635, w__4636, w__4637, w__4638, w__4639, w__4640;
  wire w__4641, w__4642, w__4643, w__4644, w__4645, w__4646, w__4647, w__4648;
  wire w__4649, w__4650, w__4651, w__4652, w__4653, w__4654, w__4655, w__4656;
  wire w__4657, w__4658, w__4659, w__4660, w__4661, w__4662, w__4663, w__4664;
  wire w__4665, w__4666, w__4667, w__4668, w__4669, w__4670, w__4671, w__4672;
  wire w__4673, w__4674, w__4675, w__4676, w__4677, w__4678, w__4679, w__4680;
  wire w__4681, w__4682, w__4683, w__4684, w__4685, w__4686, w__4687, w__4688;
  wire w__4689, w__4690, w__4691, w__4692, w__4693, w__4694, w__4695, w__4696;
  wire w__4697, w__4698, w__4699, w__4700, w__4701, w__4702, w__4703, w__4704;
  wire w__4705, w__4706, w__4707, w__4708, w__4709, w__4710, w__4711, w__4712;
  wire w__4713, w__4714, w__4715, w__4716, w__4717, w__4718, w__4719, w__4720;
  wire w__4721, w__4722, w__4723, w__4724, w__4725, w__4726, w__4727, w__4728;
  wire w__4729, w__4730, w__4731, w__4732, w__4733, w__4734, w__4735, w__4736;
  wire w__4737, w__4738, w__4739, w__4740, w__4741, w__4742, w__4743, w__4744;
  wire w__4745, w__4746, w__4747, w__4748, w__4749, w__4750, w__4751, w__4752;
  wire w__4753, w__4754, w__4755, w__4756, w__4757, w__4758, w__4759, w__4760;
  wire w__4761, w__4762, w__4763, w__4764, w__4765, w__4766, w__4767, w__4768;
  wire w__4769, w__4770, w__4771, w__4772, w__4773, w__4774, w__4775, w__4776;
  wire w__4777, w__4778, w__4779, w__4780, w__4781, w__4782, w__4783, w__4784;
  wire w__4785, w__4786, w__4787, w__4788, w__4789, w__4790, w__4791, w__4792;
  wire w__4793, w__4794, w__4795, w__4796, w__4797, w__4798, w__4799, w__4800;
  wire w__4801, w__4802, w__4803, w__4804, w__4805, w__4806, w__4807, w__4808;
  wire w__4809, w__4810, w__4811, w__4812, w__4813, w__4814, w__4815, w__4816;
  wire w__4817, w__4818, w__4819, w__4820, w__4821, w__4822, w__4823, w__4824;
  wire w__4825, w__4826, w__4827, w__4828, w__4829, w__4830, w__4831, w__4832;
  wire w__4833, w__4834, w__4835, w__4836, w__4837, w__4838, w__4839, w__4840;
  wire w__4841, w__4842, w__4843, w__4844, w__4845, w__4846, w__4847, w__4848;
  wire w__4849, w__4850, w__4851, w__4852, w__4853, w__4854, w__4855, w__4856;
  wire w__4857, w__4858, w__4859, w__4860, w__4861, w__4862, w__4863, w__4864;
  wire w__4865, w__4866, w__4867, w__4868, w__4869, w__4870, w__4871, w__4872;
  wire w__4873, w__4874, w__4875, w__4876, w__4877, w__4878, w__4879, w__4880;
  wire w__4881, w__4882, w__4883, w__4884, w__4885, w__4886, w__4887, w__4888;
  wire w__4889, w__4890, w__4891, w__4892, w__4893, w__4894, w__4895, w__4896;
  wire w__4897, w__4898, w__4899, w__4900, w__4901, w__4902, w__4903, w__4904;
  wire w__4905, w__4906, w__4907, w__4908, w__4909, w__4910, w__4911, w__4912;
  wire w__4913, w__4914, w__4915, w__4916, w__4917, w__4918, w__4919, w__4920;
  wire w__4921, w__4922, w__4923, w__4924, w__4925, w__4926, w__4927, w__4928;
  wire w__4929, w__4930, w__4931, w__4932, w__4933, w__4934, w__4935, w__4936;
  wire w__4937, w__4938, w__4939, w__4940, w__4941, w__4942, w__4943, w__4944;
  wire w__4945, w__4946, w__4947, w__4948, w__4949, w__4950, w__4951, w__4952;
  wire w__4953, w__4954, w__4955, w__4956, w__4957, w__4958, w__4959, w__4960;
  wire w__4961, w__4962, w__4963, w__4964, w__4965, w__4966, w__4967, w__4968;
  wire w__4969, w__4970, w__4971, w__4972, w__4973, w__4974, w__4975, w__4976;
  wire w__4977, w__4978, w__4979, w__4980, w__4981, w__4982, w__4983, w__4984;
  wire w__4985, w__4986, w__4987, w__4988, w__4989, w__4990, w__4991, w__4992;
  wire w__4993, w__4994, w__4995, w__4996, w__4997, w__4998, w__4999, w__5000;
  wire w__5001, w__5002, w__5003, w__5004, w__5005, w__5006, w__5007, w__5008;
  wire w__5009, w__5010, w__5011, w__5012, w__5013, w__5014, w__5015, w__5016;
  wire w__5017, w__5018, w__5019, w__5020, w__5021, w__5022, w__5023, w__5024;
  wire w__5025, w__5026, w__5027, w__5028, w__5029, w__5030, w__5031, w__5032;
  wire w__5033, w__5034, w__5035, w__5036, w__5037, w__5038, w__5039, w__5040;
  wire w__5041, w__5042, w__5043, w__5044, w__5045, w__5046, w__5047, w__5048;
  wire w__5049, w__5050, w__5051, w__5052, w__5053, w__5054, w__5055, w__5056;
  wire w__5057, w__5058, w__5059, w__5060, w__5061, w__5062, w__5063, w__5064;
  wire w__5065, w__5066, w__5067, w__5068, w__5069, w__5070, w__5071, w__5072;
  wire w__5073, w__5074, w__5075, w__5076, w__5077, w__5078, w__5079, w__5080;
  wire w__5081, w__5082, w__5083, w__5084, w__5085, w__5086, w__5087, w__5088;
  wire w__5089, w__5090, w__5091, w__5092, w__5093, w__5094, w__5095, w__5096;
  wire w__5097, w__5098, w__5099, w__5100, w__5101, w__5102, w__5103, w__5104;
  wire w__5105, w__5106, w__5107, w__5108, w__5109, w__5110, w__5111, w__5112;
  wire w__5113, w__5114, w__5115, w__5116, w__5117, w__5118, w__5119, w__5120;
  wire w__5121, w__5122, w__5123, w__5124, w__5125, w__5126, w__5127, w__5128;
  wire w__5129, w__5130, w__5131, w__5132, w__5133, w__5134, w__5135, w__5136;
  wire w__5137, w__5138, w__5139, w__5140, w__5141, w__5142, w__5143, w__5144;
  wire w__5145, w__5146, w__5147, w__5148, w__5149, w__5150, w__5151, w__5152;
  wire w__5153, w__5154, w__5155, w__5156, w__5157, w__5158, w__5159, w__5160;
  wire w__5161, w__5162, w__5163, w__5164, w__5165, w__5166, w__5167, w__5168;
  wire w__5169, w__5170, w__5171, w__5172, w__5173, w__5174, w__5175, w__5176;
  wire w__5177, w__5178, w__5179, w__5180, w__5181, w__5182, w__5183, w__5184;
  wire w__5185, w__5186, w__5187, w__5188, w__5189, w__5190, w__5191, w__5192;
  wire w__5193, w__5194, w__5195, w__5196, w__5197, w__5198, w__5199, w__5200;
  wire w__5201, w__5202, w__5203, w__5204, w__5205, w__5206, w__5207, w__5208;
  wire w__5209, w__5210, w__5211, w__5212, w__5213, w__5214, w__5215, w__5216;
  wire w__5217, w__5218, w__5219, w__5220, w__5221, w__5222, w__5223, w__5224;
  wire w__5225, w__5226, w__5227, w__5228, w__5229, w__5230, w__5231, w__5232;
  wire w__5233, w__5234, w__5235, w__5236, w__5237, w__5238, w__5239, w__5240;
  wire w__5241, w__5242, w__5243, w__5244, w__5245, w__5246, w__5247, w__5248;
  wire w__5249, w__5250, w__5251, w__5252, w__5253, w__5254, w__5255, w__5256;
  wire w__5257, w__5258, w__5259, w__5260, w__5261, w__5262, w__5263, w__5264;
  wire w__5265, w__5266, w__5267, w__5268, w__5269, w__5270, w__5271, w__5272;
  wire w__5273, w__5274, w__5275, w__5276, w__5277, w__5278, w__5279, w__5280;
  wire w__5281, w__5282, w__5283, w__5284, w__5285, w__5286, w__5287, w__5288;
  wire w__5289, w__5290, w__5291, w__5292, w__5293, w__5294, w__5295, w__5296;
  wire w__5297, w__5298, w__5299, w__5300, w__5301, w__5302, w__5303, w__5304;
  wire w__5305, w__5306, w__5307, w__5308, w__5309, w__5310, w__5311, w__5312;
  wire w__5313, w__5314, w__5315, w__5316, w__5317, w__5318, w__5319, w__5320;
  wire w__5321, w__5322, w__5323, w__5324, w__5325, w__5326, w__5327, w__5328;
  wire w__5329, w__5330, w__5331, w__5332, w__5333, w__5334, w__5335, w__5336;
  wire w__5337, w__5338, w__5339, w__5340, w__5341, w__5342, w__5343, w__5344;
  wire w__5345, w__5346, w__5347, w__5348, w__5349, w__5350, w__5351, w__5352;
  wire w__5353, w__5354, w__5355, w__5356, w__5357, w__5358, w__5359, w__5360;
  wire w__5361, w__5362, w__5363, w__5364, w__5365, w__5366, w__5367, w__5368;
  wire w__5369, w__5370, w__5371, w__5372, w__5373, w__5374, w__5375, w__5376;
  wire w__5377, w__5378, w__5379, w__5380, w__5381, w__5382, w__5383, w__5384;
  wire w__5385, w__5386, w__5387, w__5388, w__5389, w__5390, w__5391, w__5392;
  wire w__5393, w__5394, w__5395, w__5396, w__5397, w__5398, w__5399, w__5400;
  wire w__5401, w__5402, w__5403, w__5404, w__5405, w__5406, w__5407, w__5408;
  wire w__5409, w__5410, w__5411, w__5412, w__5413, w__5414, w__5415, w__5416;
  wire w__5417, w__5418, w__5419, w__5420, w__5421, w__5422, w__5423, w__5424;
  wire w__5425, w__5426, w__5427, w__5428, w__5429, w__5430, w__5431, w__5432;
  wire w__5433, w__5434, w__5435, w__5436, w__5437, w__5438, w__5439, w__5440;
  wire w__5441, w__5442, w__5443, w__5444, w__5445, w__5446, w__5447, w__5448;
  wire w__5449, w__5450, w__5451, w__5452, w__5453, w__5454, w__5455, w__5456;
  wire w__5457, w__5458, w__5459, w__5460, w__5461, w__5462, w__5463, w__5464;
  wire w__5465, w__5466, w__5467, w__5468, w__5469, w__5470, w__5471, w__5472;
  wire w__5473, w__5474, w__5475, w__5476, w__5477, w__5478, w__5479, w__5480;
  wire w__5481, w__5482, w__5483, w__5484, w__5485, w__5486, w__5487, w__5488;
  wire w__5489, w__5490, w__5491, w__5492, w__5493, w__5494, w__5495, w__5496;
  wire w__5497, w__5498, w__5499, w__5500, w__5501, w__5502, w__5503, w__5504;
  wire w__5505, w__5506, w__5507, w__5508, w__5509, w__5510, w__5511, w__5512;
  wire w__5513, w__5514, w__5515, w__5516, w__5517, w__5518, w__5519, w__5520;
  wire w__5521, w__5522, w__5523, w__5524, w__5525, w__5526, w__5527, w__5528;
  wire w__5529, w__5530, w__5531, w__5532, w__5533, w__5534, w__5535, w__5536;
  wire w__5537, w__5538, w__5539, w__5540, w__5541, w__5542, w__5543, w__5544;
  wire w__5545, w__5546, w__5547, w__5548, w__5549, w__5550, w__5551, w__5552;
  wire w__5553, w__5554, w__5555, w__5556, w__5557, w__5558, w__5559, w__5560;
  wire w__5561, w__5562, w__5563, w__5564, w__5565, w__5566, w__5567, w__5568;
  wire w__5569, w__5570, w__5571, w__5572, w__5573, w__5574, w__5575, w__5576;
  wire w__5577, w__5578, w__5579, w__5580, w__5581, w__5582, w__5583, w__5584;
  wire w__5585, w__5586, w__5587, w__5588, w__5589, w__5590, w__5591, w__5592;
  wire w__5593, w__5594, w__5595, w__5596, w__5597, w__5598, w__5599, w__5600;
  wire w__5601, w__5602, w__5603, w__5604, w__5605, w__5606, w__5607, w__5608;
  wire w__5609, w__5610, w__5611, w__5612, w__5613, w__5614, w__5615, w__5616;
  wire w__5617, w__5618, w__5619, w__5620, w__5621, w__5622, w__5623, w__5624;
  wire w__5625, w__5626, w__5627, w__5628, w__5629, w__5630, w__5631, w__5632;
  wire w__5633, w__5634, w__5635, w__5636, w__5637, w__5638, w__5639, w__5640;
  wire w__5641, w__5642, w__5643, w__5644, w__5645, w__5646, w__5647, w__5648;
  wire w__5649, w__5650, w__5651, w__5652, w__5653, w__5654, w__5655, w__5656;
  wire w__5657, w__5658, w__5659, w__5660, w__5661, w__5662, w__5663, w__5664;
  wire w__5665, w__5666, w__5667, w__5668, w__5669, w__5670, w__5671, w__5672;
  wire w__5673, w__5674, w__5675, w__5676, w__5677, w__5678, w__5679, w__5680;
  wire w__5681, w__5682, w__5683, w__5684, w__5685, w__5686, w__5687, w__5688;
  wire w__5689, w__5690, w__5691, w__5692, w__5693, w__5694, w__5695, w__5696;
  wire w__5697, w__5698, w__5699, w__5700, w__5701, w__5702, w__5703, w__5704;
  wire w__5705, w__5706, w__5707, w__5708, w__5709, w__5710, w__5711, w__5712;
  wire w__5713, w__5714, w__5715, w__5716, w__5717, w__5718, w__5719, w__5720;
  wire w__5721, w__5722, w__5723, w__5724, w__5725, w__5726, w__5727, w__5728;
  wire w__5729, w__5730, w__5731, w__5732, w__5733, w__5734, w__5735, w__5736;
  wire w__5737, w__5738, w__5739, w__5740, w__5741, w__5742, w__5743, w__5744;
  wire w__5745, w__5746, w__5747, w__5748, w__5749, w__5750, w__5751, w__5752;
  wire w__5753, w__5754, w__5755, w__5756, w__5757, w__5758, w__5759, w__5760;
  wire w__5761, w__5762, w__5763, w__5764, w__5765, w__5766, w__5767, w__5768;
  wire w__5769, w__5770, w__5771, w__5772, w__5773, w__5774, w__5775, w__5776;
  wire w__5777, w__5778, w__5779, w__5780, w__5781, w__5782, w__5783, w__5784;
  wire w__5785, w__5786, w__5787, w__5788, w__5789, w__5790, w__5791, w__5792;
  wire w__5793, w__5794, w__5795, w__5796, w__5797, w__5798, w__5799, w__5800;
  wire w__5801, w__5802, w__5803, w__5804, w__5805, w__5806, w__5807, w__5808;
  wire w__5809, w__5810, w__5811, w__5812, w__5813, w__5814, w__5815, w__5816;
  wire w__5817, w__5818, w__5819, w__5820, w__5821, w__5822, w__5823, w__5824;
  wire w__5825, w__5826, w__5827, w__5828, w__5829, w__5830, w__5831, w__5832;
  wire w__5833, w__5834, w__5835, w__5836, w__5837, w__5838, w__5839, w__5840;
  wire w__5841, w__5842, w__5843, w__5844, w__5845, w__5846, w__5847, w__5848;
  wire w__5849, w__5850, w__5851, w__5852, w__5853, w__5854, w__5855, w__5856;
  wire w__5857, w__5858, w__5859, w__5860, w__5861, w__5862, w__5863, w__5864;
  wire w__5865, w__5866, w__5867, w__5868, w__5869, w__5870, w__5871, w__5872;
  wire w__5873, w__5874, w__5875, w__5876, w__5877, w__5878, w__5879, w__5880;
  wire w__5881, w__5882, w__5883, w__5884, w__5885, w__5886, w__5887, w__5888;
  wire w__5889, w__5890, w__5891, w__5892, w__5893, w__5894, w__5895, w__5896;
  wire w__5897, w__5898, w__5899, w__5900, w__5901, w__5902, w__5903, w__5904;
  wire w__5905, w__5906, w__5907, w__5908, w__5909, w__5910, w__5911, w__5912;
  wire w__5913, w__5914, w__5915, w__5916, w__5917, w__5918, w__5919, w__5920;
  wire w__5921, w__5922, w__5923, w__5924, w__5925, w__5926, w__5927, w__5928;
  wire w__5929, w__5930, w__5931, w__5932, w__5933, w__5934, w__5935, w__5936;
  wire w__5937, w__5938, w__5939, w__5940, w__5941, w__5942, w__5943, w__5944;
  wire w__5945, w__5946, w__5947, w__5948, w__5949, w__5950, w__5951, w__5952;
  wire w__5953, w__5954, w__5955, w__5956, w__5957, w__5958, w__5959, w__5960;
  wire w__5961, w__5962, w__5963, w__5964, w__5965, w__5966, w__5967, w__5968;
  wire w__5969, w__5970, w__5971, w__5972, w__5973, w__5974, w__5975, w__5976;
  wire w__5977, w__5978, w__5979, w__5980, w__5981, w__5982, w__5983, w__5984;
  wire w__5985, w__5986, w__5987, w__5988, w__5989, w__5990, w__5991, w__5992;
  wire w__5993, w__5994, w__5995, w__5996, w__5997, w__5998, w__5999, w__6000;
  wire w__6001, w__6002, w__6003, w__6004, w__6005, w__6006, w__6007, w__6008;
  wire w__6009, w__6010, w__6011, w__6012, w__6013, w__6014, w__6015, w__6016;
  wire w__6017, w__6018, w__6019, w__6020, w__6021, w__6022, w__6023, w__6024;
  wire w__6025, w__6026, w__6027, w__6028, w__6029, w__6030, w__6031, w__6032;
  wire w__6033, w__6034, w__6035, w__6036, w__6037, w__6038, w__6039, w__6040;
  wire w__6041, w__6042, w__6043, w__6044, w__6045, w__6046, w__6047, w__6048;
  wire w__6049, w__6050, w__6051, w__6052, w__6053, w__6054, w__6055, w__6056;
  wire w__6057, w__6058, w__6059, w__6060, w__6061, w__6062, w__6063, w__6064;
  wire w__6065, w__6066, w__6067, w__6068, w__6069, w__6070, w__6071, w__6072;
  wire w__6073, w__6074, w__6075, w__6076, w__6077, w__6078, w__6079, w__6080;
  wire w__6081, w__6082, w__6083, w__6084, w__6085, w__6086, w__6087, w__6088;
  wire w__6089, w__6090, w__6091, w__6092, w__6093, w__6094, w__6095, w__6096;
  wire w__6097, w__6098, w__6099, w__6100, w__6101, w__6102, w__6103, w__6104;
  wire w__6105, w__6106, w__6107, w__6108, w__6109, w__6110, w__6111, w__6112;
  wire w__6113, w__6114, w__6115, w__6116, w__6117, w__6118, w__6119, w__6120;
  wire w__6121, w__6122, w__6123, w__6124, w__6125, w__6126, w__6127, w__6128;
  wire w__6129, w__6130, w__6131, w__6132, w__6133, w__6134, w__6135, w__6136;
  wire w__6137, w__6138, w__6139, w__6140, w__6141, w__6142, w__6143, w__6144;
  wire w__6145, w__6146, w__6147, w__6148, w__6149, w__6150, w__6151, w__6152;
  wire w__6153, w__6154, w__6155, w__6156, w__6157, w__6158, w__6159, w__6160;
  wire w__6161, w__6162, w__6163, w__6164, w__6165, w__6166, w__6167, w__6168;
  wire w__6169, w__6170, w__6171, w__6172, w__6173, w__6174, w__6175, w__6176;
  wire w__6177, w__6178, w__6179, w__6180, w__6181, w__6182, w__6183, w__6184;
  wire w__6185, w__6186, w__6187, w__6188, w__6189, w__6190, w__6191, w__6192;
  wire w__6193, w__6194, w__6195, w__6196, w__6197, w__6198, w__6199, w__6200;
  wire w__6201, w__6202, w__6203, w__6204, w__6205, w__6206, w__6207, w__6208;
  wire w__6209, w__6210, w__6211, w__6212, w__6213, w__6214, w__6215, w__6216;
  wire w__6217, w__6218, w__6219, w__6220, w__6221, w__6222, w__6223, w__6224;
  wire w__6225, w__6226, w__6227, w__6228, w__6229, w__6230, w__6231, w__6232;
  wire w__6233, w__6234, w__6235, w__6236, w__6237, w__6238, w__6239, w__6240;
  wire w__6241, w__6242, w__6243, w__6244, w__6245, w__6246, w__6247, w__6248;
  wire w__6249, w__6250, w__6251, w__6252, w__6253, w__6254, w__6255, w__6256;
  wire w__6257, w__6258, w__6259, w__6260, w__6261, w__6262, w__6263, w__6264;
  wire w__6265, w__6266, w__6267, w__6268, w__6269, w__6270, w__6271, w__6272;
  wire w__6273, w__6274, w__6275, w__6276, w__6277, w__6278, w__6279, w__6280;
  wire w__6281, w__6282, w__6283, w__6284, w__6285, w__6286, w__6287, w__6288;
  wire w__6289, w__6290, w__6291, w__6292, w__6293, w__6294, w__6295, w__6296;
  wire w__6297, w__6298, w__6299, w__6300, w__6301, w__6302, w__6303, w__6304;
  wire w__6305, w__6306, w__6307, w__6308, w__6309, w__6310, w__6311, w__6312;
  wire w__6313, w__6314, w__6315, w__6316, w__6317, w__6318, w__6319, w__6320;
  wire w__6321, w__6322, w__6323, w__6324, w__6325, w__6326, w__6327, w__6328;
  wire w__6329, w__6330, w__6331, w__6332, w__6333, w__6334, w__6335, w__6336;
  wire w__6337, w__6338, w__6339, w__6340, w__6341, w__6342, w__6343, w__6344;
  wire w__6345, w__6346, w__6347, w__6348, w__6349, w__6350, w__6351, w__6352;
  wire w__6353, w__6354, w__6355, w__6356, w__6357, w__6358, w__6359, w__6360;
  wire w__6361, w__6362, w__6363, w__6364, w__6365, w__6366, w__6367, w__6368;
  wire w__6369, w__6370, w__6371, w__6372, w__6373, w__6374, w__6375, w__6376;
  wire w__6377, w__6378, w__6379, w__6380, w__6381, w__6382, w__6383, w__6384;
  wire w__6385, w__6386, w__6387, w__6388, w__6389, w__6390, w__6391, w__6392;
  wire w__6393, w__6394, w__6395, w__6396, w__6397, w__6398, w__6399, w__6400;
  wire w__6401, w__6402, w__6403, w__6404, w__6405, w__6406, w__6407, w__6408;
  wire w__6409, w__6410, w__6411, w__6412, w__6413, w__6414, w__6415, w__6416;
  wire w__6417, w__6418, w__6419, w__6420, w__6421, w__6422, w__6423, w__6424;
  wire w__6425, w__6426, w__6427, w__6428, w__6429, w__6430, w__6431, w__6432;
  wire w__6433, w__6434, w__6435, w__6436, w__6437, w__6438, w__6439, w__6440;
  wire w__6441, w__6442, w__6443, w__6444, w__6445, w__6446, w__6447, w__6448;
  wire w__6449, w__6450, w__6451, w__6452, w__6453, w__6454, w__6455, w__6456;
  wire w__6457, w__6458, w__6459, w__6460, w__6461, w__6462, w__6463, w__6464;
  wire w__6465, w__6466, w__6467, w__6468, w__6469, w__6470, w__6471, w__6472;
  wire w__6473, w__6474, w__6475, w__6476, w__6477, w__6478, w__6479, w__6480;
  wire w__6481, w__6482, w__6483, w__6484, w__6485, w__6486, w__6487, w__6488;
  wire w__6489, w__6490, w__6491, w__6492, w__6493, w__6494, w__6495, w__6496;
  wire w__6497, w__6498, w__6499, w__6500, w__6501, w__6502, w__6503, w__6504;
  wire w__6505, w__6506, w__6507, w__6508, w__6509, w__6510, w__6511, w__6512;
  wire w__6513, w__6514, w__6515, w__6516, w__6517, w__6518, w__6519, w__6520;
  wire w__6521, w__6522, w__6523, w__6524, w__6525, w__6526, w__6527, w__6528;
  wire w__6529, w__6530, w__6531, w__6532, w__6533, w__6534, w__6535, w__6536;
  wire w__6537, w__6538, w__6539, w__6540, w__6541, w__6542, w__6543, w__6544;
  wire w__6545, w__6546, w__6547, w__6548, w__6549, w__6550, w__6551, w__6552;
  wire w__6553, w__6554, w__6555, w__6556, w__6557, w__6558, w__6559, w__6560;
  wire w__6561, w__6562, w__6563, w__6564, w__6565, w__6566, w__6567, w__6568;
  wire w__6569, w__6570, w__6571, w__6572, w__6573, w__6574, w__6575, w__6576;
  wire w__6577, w__6578, w__6579, w__6580, w__6581, w__6582, w__6583, w__6584;
  wire w__6585, w__6586, w__6587, w__6588, w__6589, w__6590, w__6591, w__6592;
  wire w__6593, w__6594, w__6595, w__6596, w__6597, w__6598, w__6599, w__6600;
  wire w__6601, w__6602, w__6603, w__6604, w__6605, w__6606, w__6607, w__6608;
  wire w__6609, w__6610, w__6611, w__6612, w__6613, w__6614, w__6615, w__6616;
  wire w__6617, w__6618, w__6619, w__6620, w__6621, w__6622, w__6623, w__6624;
  wire w__6625, w__6626, w__6627, w__6628, w__6629, w__6630, w__6631, w__6632;
  wire w__6633, w__6634, w__6635, w__6636, w__6637, w__6638, w__6639, w__6640;
  wire w__6641, w__6642, w__6643, w__6644, w__6645, w__6646, w__6647, w__6648;
  wire w__6649, w__6650, w__6651, w__6652, w__6653, w__6654, w__6655, w__6656;
  wire w__6657, w__6658, w__6659, w__6660, w__6661, w__6662, w__6663, w__6664;
  wire w__6665, w__6666, w__6667, w__6668, w__6669, w__6670, w__6671, w__6672;
  wire w__6673, w__6674, w__6675, w__6676, w__6677, w__6678, w__6679, w__6680;
  wire w__6681, w__6682, w__6683, w__6684, w__6685, w__6686, w__6687, w__6688;
  wire w__6689, w__6690, w__6691, w__6692, w__6693, w__6694, w__6695, w__6696;
  wire w__6697, w__6698, w__6699, w__6700, w__6701, w__6702, w__6703, w__6704;
  wire w__6705, w__6706, w__6707, w__6708, w__6709, w__6710, w__6711, w__6712;
  wire w__6713, w__6714, w__6715, w__6716, w__6717, w__6718, w__6719, w__6720;
  wire w__6721, w__6722, w__6723, w__6724, w__6725, w__6726, w__6727, w__6728;
  wire w__6729, w__6730, w__6731, w__6732, w__6733, w__6734, w__6735, w__6736;
  wire w__6737, w__6738, w__6739, w__6740, w__6741, w__6742, w__6743, w__6744;
  wire w__6745, w__6746, w__6747, w__6748, w__6749, w__6750, w__6751, w__6752;
  wire w__6753, w__6754, w__6755, w__6756, w__6757, w__6758, w__6759, w__6760;
  wire w__6761, w__6762, w__6763, w__6764, w__6765, w__6766, w__6767, w__6768;
  wire w__6769, w__6770, w__6771, w__6772, w__6773, w__6774, w__6775, w__6776;
  wire w__6777, w__6778, w__6779, w__6780, w__6781, w__6782, w__6783, w__6784;
  wire w__6785, w__6786, w__6787, w__6788, w__6789, w__6790, w__6791, w__6792;
  wire w__6793, w__6794, w__6795, w__6796, w__6797, w__6798, w__6799, w__6800;
  wire w__6801, w__6802, w__6803, w__6804, w__6805, w__6806, w__6807, w__6808;
  wire w__6809, w__6810, w__6811, w__6812, w__6813, w__6814, w__6815, w__6816;
  wire w__6817, w__6818, w__6819, w__6820, w__6821, w__6822, w__6823, w__6824;
  wire w__6825, w__6826, w__6827, w__6828, w__6829, w__6830, w__6831, w__6832;
  wire w__6833, w__6834, w__6835, w__6836, w__6837, w__6838, w__6839, w__6840;
  wire w__6841, w__6842, w__6843, w__6844, w__6845, w__6846, w__6847, w__6848;
  wire w__6849, w__6850, w__6851, w__6852, w__6853, w__6854, w__6855, w__6856;
  wire w__6857, w__6858, w__6859, w__6860, w__6861, w__6862, w__6863, w__6864;
  wire w__6865, w__6866, w__6867, w__6868, w__6869, w__6870, w__6871, w__6872;
  wire w__6873, w__6874, w__6875, w__6876, w__6877, w__6878, w__6879, w__6880;
  wire w__6881, w__6882, w__6883, w__6884, w__6885, w__6886, w__6887, w__6888;
  wire w__6889, w__6890, w__6891, w__6892, w__6893, w__6894, w__6895, w__6896;
  wire w__6897, w__6898, w__6899, w__6900, w__6901, w__6902, w__6903, w__6904;
  wire w__6905, w__6906, w__6907, w__6908, w__6909, w__6910, w__6911, w__6912;
  wire w__6913, w__6914, w__6915, w__6916, w__6917, w__6918, w__6919, w__6920;
  wire w__6921, w__6922, w__6923, w__6924, w__6925, w__6926, w__6927, w__6928;
  wire w__6929, w__6930, w__6931, w__6932, w__6933, w__6934, w__6935, w__6936;
  wire w__6937, w__6938, w__6939, w__6940, w__6941, w__6942, w__6943, w__6944;
  wire w__6945, w__6946, w__6947, w__6948, w__6949, w__6950, w__6951, w__6952;
  wire w__6953, w__6954, w__6955, w__6956, w__6957, w__6958, w__6959, w__6960;
  wire w__6961, w__6962, w__6963, w__6964, w__6965, w__6966, w__6967, w__6968;
  wire w__6969, w__6970, w__6971, w__6972, w__6973, w__6974, w__6975, w__6976;
  wire w__6977, w__6978, w__6979, w__6980, w__6981, w__6982, w__6983, w__6984;
  wire w__6985, w__6986, w__6987, w__6988, w__6989, w__6990, w__6991, w__6992;
  wire w__6993, w__6994, w__6995, w__6996, w__6997, w__6998, w__6999, w__7000;
  wire w__7001, w__7002, w__7003, w__7004, w__7005, w__7006, w__7007, w__7008;
  wire w__7009, w__7010, w__7011, w__7012, w__7013, w__7014, w__7015, w__7016;
  wire w__7017, w__7018, w__7019, w__7020, w__7021, w__7022, w__7023, w__7024;
  wire w__7025, w__7026, w__7027, w__7028, w__7029, w__7030, w__7031, w__7032;
  wire w__7033, w__7034, w__7035, w__7036, w__7037, w__7038, w__7039, w__7040;
  wire w__7041, w__7042, w__7043, w__7044, w__7045, w__7046, w__7047, w__7048;
  wire w__7049, w__7050, w__7051, w__7052, w__7053, w__7054, w__7055, w__7056;
  wire w__7057, w__7058, w__7059, w__7060, w__7061, w__7062, w__7063, w__7064;
  wire w__7065, w__7066, w__7067, w__7068, w__7069, w__7070, w__7071, w__7072;
  wire w__7073, w__7074, w__7075, w__7076, w__7077, w__7078, w__7079, w__7080;
  wire w__7081, w__7082, w__7083, w__7084, w__7085, w__7086, w__7087, w__7088;
  wire w__7089, w__7090, w__7091, w__7092, w__7093, w__7094, w__7095, w__7096;
  wire w__7097, w__7098, w__7099, w__7100, w__7101, w__7102, w__7103, w__7104;
  wire w__7105, w__7106, w__7107, w__7108, w__7109, w__7110, w__7111, w__7112;
  wire w__7113, w__7114, w__7115, w__7116, w__7117, w__7118, w__7119, w__7120;
  wire w__7121, w__7122, w__7123, w__7124, w__7125, w__7126, w__7127, w__7128;
  wire w__7129, w__7130, w__7131, w__7132, w__7133, w__7134, w__7135, w__7136;
  wire w__7137, w__7138, w__7139, w__7140, w__7141, w__7142, w__7143, w__7144;
  wire w__7145, w__7146, w__7147, w__7148, w__7149, w__7150, w__7151, w__7152;
  wire w__7153, w__7154, w__7155, w__7156, w__7157, w__7158, w__7159, w__7160;
  wire w__7161, w__7162, w__7163, w__7164, w__7165, w__7166, w__7167, w__7168;
  wire w__7169, w__7170, w__7171, w__7172, w__7173, w__7174, w__7175, w__7176;
  wire w__7177, w__7178, w__7179, w__7180, w__7181, w__7182, w__7183, w__7184;
  wire w__7185, w__7186, w__7187, w__7188, w__7189, w__7190, w__7191, w__7192;
  wire w__7193, w__7194, w__7195, w__7196, w__7197, w__7198, w__7199, w__7200;
  wire w__7201, w__7202, w__7203, w__7204, w__7205, w__7206, w__7207, w__7208;
  wire w__7209, w__7210, w__7211, w__7212, w__7213, w__7214, w__7215, w__7216;
  wire w__7217, w__7218, w__7219, w__7220, w__7221, w__7222, w__7223, w__7224;
  wire w__7225, w__7226, w__7227, w__7228, w__7229, w__7230, w__7231, w__7232;
  wire w__7233, w__7234, w__7235, w__7236, w__7237, w__7238, w__7239, w__7240;
  wire w__7241, w__7242, w__7243, w__7244, w__7245, w__7246, w__7247, w__7248;
  wire w__7249, w__7250, w__7251, w__7252, w__7253, w__7254, w__7255, w__7256;
  wire w__7257, w__7258, w__7259, w__7260, w__7261, w__7262, w__7263, w__7264;
  wire w__7265, w__7266, w__7267, w__7268, w__7269, w__7270, w__7271, w__7272;
  wire w__7273, w__7274, w__7275, w__7276, w__7277, w__7278, w__7279, w__7280;
  wire w__7281, w__7282, w__7283, w__7284, w__7285, w__7286, w__7287, w__7288;
  wire w__7289, w__7290, w__7291, w__7292, w__7293, w__7294, w__7295, w__7296;
  wire w__7297, w__7298, w__7299, w__7300, w__7301, w__7302, w__7303, w__7304;
  wire w__7305, w__7306, w__7307, w__7308, w__7309, w__7310, w__7311, w__7312;
  wire w__7313, w__7314, w__7315, w__7316, w__7317, w__7318, w__7319, w__7320;
  wire w__7321, w__7322, w__7323, w__7324, w__7325, w__7326, w__7327, w__7328;
  wire w__7329, w__7330, w__7331, w__7332, w__7333, w__7334, w__7335, w__7336;
  wire w__7337, w__7338, w__7339, w__7340, w__7341, w__7342, w__7343, w__7344;
  wire w__7345, w__7346, w__7347, w__7348, w__7349, w__7350, w__7351, w__7352;
  wire w__7353, w__7354, w__7355, w__7356, w__7357, w__7358, w__7359, w__7360;
  wire w__7361, w__7362, w__7363, w__7364, w__7365, w__7366, w__7367, w__7368;
  wire w__7369, w__7370, w__7371, w__7372, w__7373, w__7374, w__7375, w__7376;
  wire w__7377, w__7378, w__7379, w__7380, w__7381, w__7382, w__7383, w__7384;
  wire w__7385, w__7386, w__7387, w__7388, w__7389, w__7390, w__7391, w__7392;
  wire w__7393, w__7394, w__7395, w__7396, w__7397, w__7398, w__7399, w__7400;
  wire w__7401, w__7402, w__7403, w__7404, w__7405, w__7406, w__7407, w__7408;
  wire w__7409, w__7410, w__7411, w__7412, w__7413, w__7414, w__7415, w__7416;
  wire w__7417, w__7418, w__7419, w__7420, w__7421, w__7422, w__7423, w__7424;
  wire w__7425, w__7426, w__7427, w__7428, w__7429, w__7430, w__7431, w__7432;
  wire w__7433, w__7434, w__7435, w__7436, w__7437, w__7438, w__7439, w__7440;
  wire w__7441, w__7442, w__7443, w__7444, w__7445, w__7446, w__7447, w__7448;
  wire w__7449, w__7450, w__7451, w__7452, w__7453, w__7454, w__7455, w__7456;
  wire w__7457, w__7458, w__7459, w__7460, w__7461, w__7462, w__7463, w__7464;
  wire w__7465, w__7466, w__7467, w__7468, w__7469, w__7470, w__7471, w__7472;
  wire w__7473, w__7474, w__7475, w__7476, w__7477, w__7478, w__7479, w__7480;
  wire w__7481, w__7482, w__7483, w__7484, w__7485, w__7486, w__7487, w__7488;
  wire w__7489, w__7490, w__7491, w__7492, w__7493, w__7494, w__7495, w__7496;
  wire w__7497, w__7498, w__7499, w__7500, w__7501, w__7502, w__7503, w__7504;
  wire w__7505, w__7506, w__7507, w__7508, w__7509, w__7510, w__7511, w__7512;
  wire w__7513, w__7514, w__7515, w__7516, w__7517, w__7518, w__7519, w__7520;
  wire w__7521, w__7522, w__7523, w__7524, w__7525, w__7526, w__7527, w__7528;
  wire w__7529, w__7530, w__7531, w__7532, w__7533, w__7534, w__7535, w__7536;
  wire w__7537, w__7538, w__7539, w__7540, w__7541, w__7542, w__7543, w__7544;
  wire w__7545, w__7546, w__7547, w__7548, w__7549, w__7550, w__7551, w__7552;
  wire w__7553, w__7554, w__7555, w__7556, w__7557, w__7558, w__7559, w__7560;
  wire w__7561, w__7562, w__7563, w__7564, w__7565, w__7566, w__7567, w__7568;
  wire w__7569, w__7570, w__7571, w__7572, w__7573, w__7574, w__7575, w__7576;
  wire w__7577, w__7578, w__7579, w__7580, w__7581, w__7582, w__7583, w__7584;
  wire w__7585, w__7586, w__7587, w__7588, w__7589, w__7590, w__7591, w__7592;
  wire w__7593, w__7594, w__7595, w__7596, w__7597, w__7598, w__7599, w__7600;
  wire w__7601, w__7602, w__7603, w__7604, w__7605, w__7606, w__7607, w__7608;
  wire w__7609, w__7610, w__7611, w__7612, w__7613, w__7614, w__7615, w__7616;
  wire w__7617, w__7618, w__7619, w__7620, w__7621, w__7622, w__7623, w__7624;
  wire w__7625, w__7626, w__7627, w__7628, w__7629, w__7630, w__7631, w__7632;
  wire w__7633, w__7634, w__7635, w__7636, w__7637, w__7638, w__7639, w__7640;
  wire w__7641, w__7642, w__7643, w__7644, w__7645, w__7646, w__7647, w__7648;
  wire w__7649, w__7650, w__7651, w__7652, w__7653, w__7654, w__7655, w__7656;
  wire w__7657, w__7658, w__7659, w__7660, w__7661, w__7662, w__7663, w__7664;
  wire w__7665, w__7666, w__7667, w__7668, w__7669, w__7670, w__7671, w__7672;
  wire w__7673, w__7674, w__7675, w__7676, w__7677, w__7678, w__7679, w__7680;
  wire w__7681, w__7682, w__7683, w__7684, w__7685, w__7686, w__7687, w__7688;
  wire w__7689, w__7690, w__7691, w__7692, w__7693, w__7694, w__7695, w__7696;
  wire w__7697, w__7698, w__7699, w__7700, w__7701, w__7702, w__7703, w__7704;
  wire w__7705, w__7706, w__7707, w__7708, w__7709, w__7710, w__7711, w__7712;
  wire w__7713, w__7714, w__7715, w__7716, w__7717, w__7718, w__7719, w__7720;
  wire w__7721, w__7722, w__7723, w__7724, w__7725, w__7726, w__7727, w__7728;
  wire w__7729, w__7730, w__7731, w__7732, w__7733, w__7734, w__7735, w__7736;
  wire w__7737, w__7738, w__7739, w__7740, w__7741, w__7742, w__7743, w__7744;
  wire w__7745, w__7746, w__7747, w__7748, w__7749, w__7750, w__7751, w__7752;
  wire w__7753, w__7754, w__7755, w__7756, w__7757, w__7758, w__7759, w__7760;
  wire w__7761, w__7762, w__7763, w__7764, w__7765, w__7766, w__7767, w__7768;
  wire w__7769, w__7770, w__7771, w__7772, w__7773, w__7774, w__7775, w__7776;
  wire w__7777, w__7778, w__7779, w__7780, w__7781, w__7782, w__7783, w__7784;
  wire w__7785, w__7786, w__7787, w__7788, w__7789, w__7790, w__7791, w__7792;
  wire w__7793, w__7794, w__7795, w__7796, w__7797, w__7798, w__7799, w__7800;
  wire w__7801, w__7802, w__7803, w__7804, w__7805, w__7806, w__7807, w__7808;
  wire w__7809, w__7810, w__7811, w__7812, w__7813, w__7814, w__7815, w__7816;
  wire w__7817, w__7818, w__7819, w__7820, w__7821, w__7822, w__7823, w__7824;
  wire w__7825, w__7826, w__7827, w__7828, w__7829, w__7830, w__7831, w__7832;
  wire w__7833, w__7834, w__7835, w__7836, w__7837, w__7838, w__7839, w__7840;
  wire w__7841, w__7842, w__7843, w__7844, w__7845, w__7846, w__7847, w__7848;
  wire w__7849, w__7850, w__7851, w__7852, w__7853, w__7854, w__7855, w__7856;
  wire w__7857, w__7858, w__7859, w__7860, w__7861, w__7862, w__7863, w__7864;
  wire w__7865, w__7866, w__7867, w__7868, w__7869, w__7870, w__7871, w__7872;
  wire w__7873, w__7874, w__7875, w__7876, w__7877, w__7878, w__7879, w__7880;
  wire w__7881, w__7882, w__7883, w__7884, w__7885, w__7886, w__7887, w__7888;
  wire w__7889, w__7890, w__7891, w__7892, w__7893, w__7894, w__7895, w__7896;
  wire w__7897, w__7898, w__7899, w__7900, w__7901, w__7902, w__7903, w__7904;
  wire w__7905, w__7906, w__7907, w__7908, w__7909, w__7910, w__7911, w__7912;
  wire w__7913, w__7914, w__7915, w__7916, w__7917, w__7918, w__7919, w__7920;
  wire w__7921, w__7922, w__7923, w__7924, w__7925, w__7926, w__7927, w__7928;
  wire w__7929, w__7930, w__7931, w__7932, w__7933, w__7934, w__7935, w__7936;
  wire w__7937, w__7938, w__7939, w__7940, w__7941, w__7942, w__7943, w__7944;
  wire w__7945, w__7946, w__7947, w__7948, w__7949, w__7950, w__7951, w__7952;
  wire w__7953, w__7954, w__7955, w__7956, w__7957, w__7958, w__7959, w__7960;
  wire w__7961, w__7962, w__7963, w__7964, w__7965, w__7966, w__7967, w__7968;
  wire w__7969, w__7970, w__7971, w__7972, w__7973, w__7974, w__7975, w__7976;
  wire w__7977, w__7978, w__7979, w__7980, w__7981, w__7982, w__7983, w__7984;
  wire w__7985, w__7986, w__7987, w__7988, w__7989, w__7990, w__7991, w__7992;
  wire w__7993, w__7994, w__7995, w__7996, w__7997, w__7998, w__7999, w__8000;
  wire w__8001, w__8002, w__8003, w__8004, w__8005, w__8006, w__8007, w__8008;
  wire w__8009, w__8010, w__8011, w__8012, w__8013, w__8014, w__8015, w__8016;
  wire w__8017, w__8018, w__8019, w__8020, w__8021, w__8022, w__8023, w__8024;
  wire w__8025, w__8026, w__8027, w__8028, w__8029, w__8030, w__8031, w__8032;
  wire w__8033, w__8034, w__8035, w__8036, w__8037, w__8038, w__8039, w__8040;
  wire w__8041, w__8042, w__8043, w__8044, w__8045, w__8046, w__8047, w__8048;
  wire w__8049, w__8050, w__8051, w__8052, w__8053, w__8054, w__8055, w__8056;
  wire w__8057, w__8058, w__8059, w__8060, w__8061, w__8062, w__8063, w__8064;
  wire w__8065, w__8066, w__8067, w__8068, w__8069, w__8070, w__8071, w__8072;
  wire w__8073, w__8074, w__8075, w__8076, w__8077, w__8078, w__8079, w__8080;
  wire w__8081, w__8082, w__8083, w__8084, w__8085, w__8086, w__8087, w__8088;
  wire w__8089, w__8090, w__8091, w__8092, w__8093, w__8094, w__8095, w__8096;
  wire w__8097, w__8098, w__8099, w__8100, w__8101, w__8102, w__8103, w__8104;
  wire w__8105, w__8106, w__8107, w__8108, w__8109, w__8110, w__8111, w__8112;
  wire w__8113, w__8114, w__8115, w__8116, w__8117, w__8118, w__8119, w__8120;
  wire w__8121, w__8122, w__8123, w__8124, w__8125, w__8126, w__8127, w__8128;
  wire w__8129, w__8130, w__8131, w__8132, w__8133, w__8134, w__8135, w__8136;
  wire w__8137, w__8138, w__8139, w__8140, w__8141, w__8142, w__8143, w__8144;
  wire w__8145, w__8146, w__8147, w__8148, w__8149, w__8150, w__8151, w__8152;
  wire w__8153, w__8154, w__8155, w__8156, w__8157, w__8158, w__8159, w__8160;
  wire w__8161, w__8162, w__8163, w__8164, w__8165, w__8166, w__8167, w__8168;
  wire w__8169, w__8170, w__8171, w__8172, w__8173, w__8174, w__8175, w__8176;
  wire w__8177, w__8178, w__8179, w__8180, w__8181, w__8182, w__8183, w__8184;
  wire w__8185, w__8186, w__8187, w__8188, w__8189, w__8190, w__8191, w__8192;
  wire w__8193, w__8194, w__8195, w__8196, w__8197, w__8198, w__8199, w__8200;
  wire w__8201, w__8202, w__8203, w__8204, w__8205, w__8206, w__8207, w__8208;
  wire w__8209, w__8210, w__8211, w__8212, w__8213, w__8214, w__8215, w__8216;
  wire w__8217, w__8218, w__8219, w__8220, w__8221, w__8222, w__8223, w__8224;
  wire w__8225, w__8226, w__8227, w__8228, w__8229, w__8230, w__8231, w__8232;
  wire w__8233, w__8234, w__8235, w__8236, w__8237, w__8238, w__8239, w__8240;
  wire w__8241, w__8242, w__8243, w__8244, w__8245, w__8246, w__8247, w__8248;
  wire w__8249, w__8250, w__8251, w__8252, w__8253, w__8254, w__8255, w__8256;
  wire w__8257, w__8258, w__8259, w__8260, w__8261, w__8262, w__8263, w__8264;
  wire w__8265, w__8266, w__8267, w__8268, w__8269, w__8270, w__8271, w__8272;
  wire w__8273, w__8274, w__8275, w__8276, w__8277, w__8278, w__8279, w__8280;
  wire w__8281, w__8282, w__8283, w__8284, w__8285, w__8286, w__8287, w__8288;
  wire w__8289, w__8290, w__8291, w__8292, w__8293, w__8294, w__8295, w__8296;
  wire w__8297, w__8298, w__8299, w__8300, w__8301, w__8302, w__8303, w__8304;
  wire w__8305, w__8306, w__8307, w__8308, w__8309, w__8310, w__8311, w__8312;
  wire w__8313, w__8314, w__8315, w__8316, w__8317, w__8318, w__8319, w__8320;
  wire w__8321, w__8322, w__8323, w__8324, w__8325, w__8326, w__8327, w__8328;
  wire w__8329, w__8330, w__8331, w__8332, w__8333, w__8334, w__8335, w__8336;
  wire w__8337, w__8338, w__8339, w__8340, w__8341, w__8342, w__8343, w__8344;
  wire w__8345, w__8346, w__8347, w__8348, w__8349, w__8350, w__8351, w__8352;
  wire w__8353, w__8354, w__8355, w__8356, w__8357, w__8358, w__8359, w__8360;
  wire w__8361, w__8362, w__8363, w__8364, w__8365, w__8366, w__8367, w__8368;
  wire w__8369, w__8370, w__8371, w__8372, w__8373, w__8374, w__8375, w__8376;
  wire w__8377, w__8378, w__8379, w__8380, w__8381, w__8382, w__8383, w__8384;
  wire w__8385, w__8386, w__8387, w__8388, w__8389, w__8390, w__8391, w__8392;
  wire w__8393, w__8394, w__8395, w__8396, w__8397, w__8398, w__8399, w__8400;
  wire w__8401, w__8402, w__8403, w__8404, w__8405, w__8406, w__8407, w__8408;
  wire w__8409, w__8410, w__8411, w__8412, w__8413, w__8414, w__8415, w__8416;
  wire w__8417, w__8418, w__8419, w__8420, w__8421, w__8422, w__8423, w__8424;
  wire w__8425, w__8426, w__8427, w__8428, w__8429, w__8430, w__8431, w__8432;
  wire w__8433, w__8434, w__8435, w__8436, w__8437, w__8438, w__8439, w__8440;
  wire w__8441, w__8442, w__8443, w__8444, w__8445, w__8446, w__8447, w__8448;
  wire w__8449, w__8450, w__8451, w__8452, w__8453, w__8454, w__8455, w__8456;
  wire w__8457, w__8458, w__8459, w__8460, w__8461, w__8462, w__8463, w__8464;
  wire w__8465, w__8466, w__8467, w__8468, w__8469, w__8470, w__8471, w__8472;
  wire w__8473, w__8474, w__8475, w__8476, w__8477, w__8478, w__8479, w__8480;
  wire w__8481, w__8482, w__8483, w__8484, w__8485, w__8486, w__8487, w__8488;
  wire w__8489, w__8490, w__8491, w__8492, w__8493, w__8494, w__8495, w__8496;
  wire w__8497, w__8498, w__8499, w__8500, w__8501, w__8502, w__8503, w__8504;
  wire w__8505, w__8506, w__8507, w__8508, w__8509, w__8510, w__8511, w__8512;
  wire w__8513, w__8514, w__8515, w__8516, w__8517, w__8518, w__8519, w__8520;
  wire w__8521, w__8522, w__8523, w__8524, w__8525, w__8526, w__8527, w__8528;
  wire w__8529, w__8530, w__8531, w__8532, w__8533, w__8534, w__8535, w__8536;
  wire w__8537, w__8538, w__8539, w__8540, w__8541, w__8542, w__8543, w__8544;
  wire w__8545, w__8546, w__8547, w__8548, w__8549, w__8550, w__8551, w__8552;
  wire w__8553, w__8554, w__8555, w__8556, w__8557, w__8558, w__8559, w__8560;
  wire w__8561, w__8562, w__8563, w__8564, w__8565, w__8566, w__8567, w__8568;
  wire w__8569, w__8570, w__8571, w__8572, w__8573, w__8574, w__8575, w__8576;
  wire w__8577, w__8578, w__8579, w__8580, w__8581, w__8582, w__8583, w__8584;
  wire w__8585, w__8586, w__8587, w__8588, w__8589, w__8590, w__8591, w__8592;
  wire w__8593, w__8594, w__8595, w__8596, w__8597, w__8598, w__8599, w__8600;
  wire w__8601, w__8602, w__8603, w__8604, w__8605, w__8606, w__8607, w__8608;
  wire w__8609, w__8610, w__8611, w__8612, w__8613, w__8614, w__8615, w__8616;
  wire w__8617, w__8618, w__8619, w__8620, w__8621, w__8622, w__8623, w__8624;
  wire w__8625, w__8626, w__8627, w__8628, w__8629, w__8630, w__8631, w__8632;
  wire w__8633, w__8634, w__8635, w__8636, w__8637, w__8638, w__8639, w__8640;
  wire w__8641, w__8642, w__8643, w__8644, w__8645, w__8646, w__8647, w__8648;
  wire w__8649, w__8650, w__8651, w__8652, w__8653, w__8654, w__8655, w__8656;
  wire w__8657, w__8658, w__8659, w__8660, w__8661, w__8662, w__8663, w__8664;
  wire w__8665, w__8666, w__8667, w__8668, w__8669, w__8670, w__8671, w__8672;
  wire w__8673, w__8674, w__8675, w__8676, w__8677, w__8678, w__8679, w__8680;
  wire w__8681, w__8682, w__8683, w__8684, w__8685, w__8686, w__8687, w__8688;
  wire w__8689, w__8690, w__8691, w__8692, w__8693, w__8694, w__8695, w__8696;
  wire w__8697, w__8698, w__8699, w__8700, w__8701, w__8702, w__8703, w__8704;
  wire w__8705, w__8706, w__8707, w__8708, w__8709, w__8710, w__8711, w__8712;
  wire w__8713, w__8714, w__8715, w__8716, w__8717, w__8718, w__8719, w__8720;
  wire w__8721, w__8722, w__8723, w__8724, w__8725, w__8726, w__8727, w__8728;
  wire w__8729, w__8730, w__8731, w__8732, w__8733, w__8734, w__8735, w__8736;
  wire w__8737, w__8738, w__8739, w__8740, w__8741, w__8742, w__8743, w__8744;
  wire w__8745, w__8746, w__8747, w__8748, w__8749, w__8750, w__8751, w__8752;
  wire w__8753, w__8754, w__8755, w__8756, w__8757, w__8758, w__8759, w__8760;
  wire w__8761, w__8762, w__8763, w__8764, w__8765, w__8766, w__8767, w__8768;
  wire w__8769, w__8770, w__8771, w__8772, w__8773, w__8774, w__8775, w__8776;
  wire w__8777, w__8778, w__8779, w__8780, w__8781, w__8782, w__8783, w__8784;
  wire w__8785, w__8786, w__8787, w__8788, w__8789, w__8790, w__8791, w__8792;
  wire w__8793, w__8794, w__8795, w__8796, w__8797, w__8798, w__8799, w__8800;
  wire w__8801, w__8802, w__8803, w__8804, w__8805, w__8806, w__8807, w__8808;
  wire w__8809, w__8810, w__8811, w__8812, w__8813, w__8814, w__8815, w__8816;
  wire w__8817, w__8818, w__8819, w__8820, w__8821, w__8822, w__8823, w__8824;
  wire w__8825, w__8826, w__8827, w__8828, w__8829, w__8830, w__8831, w__8832;
  wire w__8833, w__8834, w__8835, w__8836, w__8837, w__8838, w__8839, w__8840;
  wire w__8841, w__8842, w__8843, w__8844, w__8845, w__8846, w__8847, w__8848;
  wire w__8849, w__8850, w__8851, w__8852, w__8853, w__8854, w__8855, w__8856;
  wire w__8857, w__8858, w__8859, w__8860, w__8861, w__8862, w__8863, w__8864;
  wire w__8865, w__8866, w__8867, w__8868, w__8869, w__8870, w__8871, w__8872;
  wire w__8873, w__8874, w__8875, w__8876, w__8877, w__8878, w__8879, w__8880;
  wire w__8881, w__8882, w__8883, w__8884, w__8885, w__8886, w__8887, w__8888;
  wire w__8889, w__8890, w__8891, w__8892, w__8893, w__8894, w__8895, w__8896;
  wire w__8897, w__8898, w__8899, w__8900, w__8901, w__8902, w__8903, w__8904;
  wire w__8905, w__8906, w__8907, w__8908, w__8909, w__8910, w__8911, w__8912;
  wire w__8913, w__8914, w__8915, w__8916, w__8917, w__8918, w__8919, w__8920;
  wire w__8921, w__8922, w__8923, w__8924, w__8925, w__8926, w__8927, w__8928;
  wire w__8929, w__8930, w__8931, w__8932, w__8933, w__8934, w__8935, w__8936;
  wire w__8937, w__8938, w__8939, w__8940, w__8941, w__8942, w__8943, w__8944;
  wire w__8945, w__8946, w__8947, w__8948, w__8949, w__8950, w__8951, w__8952;
  wire w__8953, w__8954, w__8955, w__8956, w__8957, w__8958, w__8959, w__8960;
  wire w__8961, w__8962, w__8963, w__8964, w__8965, w__8966, w__8967, w__8968;
  wire w__8969, w__8970, w__8971, w__8972, w__8973, w__8974, w__8975, w__8976;
  wire w__8977, w__8978, w__8979, w__8980, w__8981, w__8982, w__8983, w__8984;
  wire w__8985, w__8986, w__8987, w__8988, w__8989, w__8990, w__8991, w__8992;
  wire w__8993, w__8994, w__8995, w__8996, w__8997, w__8998, w__8999, w__9000;
  wire w__9001, w__9002, w__9003, w__9004, w__9005, w__9006, w__9007, w__9008;
  wire w__9009, w__9010, w__9011, w__9012, w__9013, w__9014, w__9015, w__9016;
  wire w__9017, w__9018, w__9019, w__9020, w__9021, w__9022, w__9023, w__9024;
  wire w__9025, w__9026, w__9027, w__9028, w__9029, w__9030, w__9031, w__9032;
  wire w__9033, w__9034, w__9035, w__9036, w__9037, w__9038, w__9039, w__9040;
  wire w__9041, w__9042, w__9043, w__9044, w__9045, w__9046, w__9047, w__9048;
  wire w__9049, w__9050, w__9051, w__9052, w__9053, w__9054, w__9055, w__9056;
  wire w__9057, w__9058, w__9059, w__9060, w__9061, w__9062, w__9063, w__9064;
  wire w__9065, w__9066, w__9067, w__9068, w__9069, w__9070, w__9071, w__9072;
  wire w__9073, w__9074, w__9075, w__9076, w__9077, w__9078, w__9079, w__9080;
  wire w__9081, w__9082, w__9083, w__9084, w__9085, w__9086, w__9087, w__9088;
  wire w__9089, w__9090, w__9091, w__9092, w__9093, w__9094, w__9095, w__9096;
  wire w__9097, w__9098, w__9099, w__9100, w__9101, w__9102, w__9103, w__9104;
  wire w__9105, w__9106, w__9107, w__9108, w__9109, w__9110, w__9111, w__9112;
  wire w__9113, w__9114, w__9115, w__9116, w__9117, w__9118, w__9119, w__9120;
  wire w__9121, w__9122, w__9123, w__9124, w__9125, w__9126, w__9127, w__9128;
  wire w__9129, w__9130, w__9131, w__9132, w__9133, w__9134, w__9135, w__9136;
  wire w__9137, w__9138, w__9139, w__9140, w__9141, w__9142, w__9143, w__9144;
  wire w__9145, w__9146, w__9147, w__9148, w__9149, w__9150, w__9151, w__9152;
  wire w__9153, w__9154, w__9155, w__9156, w__9157, w__9158, w__9159, w__9160;
  wire w__9161, w__9162, w__9163, w__9164, w__9165, w__9166, w__9167, w__9168;
  wire w__9169, w__9170, w__9171, w__9172, w__9173, w__9174, w__9175, w__9176;
  wire w__9177, w__9178, w__9179, w__9180, w__9181, w__9182, w__9183, w__9184;
  wire w__9185, w__9186, w__9187, w__9188, w__9189, w__9190, w__9191, w__9192;
  wire w__9193, w__9194, w__9195, w__9196, w__9197, w__9198, w__9199, w__9200;
  wire w__9201, w__9202, w__9203, w__9204, w__9205, w__9206, w__9207, w__9208;
  wire w__9209, w__9210, w__9211, w__9212, w__9213, w__9214, w__9215, w__9216;
  wire w__9217, w__9218, w__9219, w__9220, w__9221, w__9222, w__9223, w__9224;
  wire w__9225, w__9226, w__9227, w__9228, w__9229, w__9230, w__9231, w__9232;
  wire w__9233, w__9234, w__9235, w__9236, w__9237, w__9238, w__9239, w__9240;
  wire w__9241, w__9242, w__9243, w__9244, w__9245, w__9246, w__9247, w__9248;
  wire w__9249, w__9250, w__9251, w__9252, w__9253, w__9254, w__9255, w__9256;
  wire w__9257, w__9258, w__9259, w__9260, w__9261, w__9262, w__9263, w__9264;
  wire w__9265, w__9266, w__9267, w__9268, w__9269, w__9270, w__9271, w__9272;
  wire w__9273, w__9274, w__9275, w__9276, w__9277, w__9278, w__9279, w__9280;
  wire w__9281, w__9282, w__9283, w__9284, w__9285, w__9286, w__9287, w__9288;
  wire w__9289, w__9290, w__9291, w__9292, w__9293, w__9294, w__9295, w__9296;
  wire w__9297, w__9298, w__9299, w__9300, w__9301, w__9302, w__9303, w__9304;
  wire w__9305, w__9306, w__9307, w__9308, w__9309, w__9310, w__9311, w__9312;
  wire w__9313, w__9314, w__9315, w__9316, w__9317, w__9318, w__9319, w__9320;
  wire w__9321, w__9322, w__9323, w__9324, w__9325, w__9326, w__9327, w__9328;
  wire w__9329, w__9330, w__9331, w__9332, w__9333, w__9334, w__9335, w__9336;
  wire w__9337, w__9338, w__9339, w__9340, w__9341, w__9342, w__9343, w__9344;
  wire w__9345, w__9346, w__9347, w__9348, w__9349, w__9350, w__9351, w__9352;
  wire w__9353, w__9354, w__9355, w__9356, w__9357, w__9358, w__9359, w__9360;
  wire w__9361, w__9362, w__9363, w__9364, w__9365, w__9366, w__9367, w__9368;
  wire w__9369, w__9370, w__9371, w__9372, w__9373, w__9374, w__9375, w__9376;
  wire w__9377, w__9378, w__9379, w__9380, w__9381, w__9382, w__9383, w__9384;
  wire w__9385, w__9386, w__9387, w__9388, w__9389, w__9390, w__9391, w__9392;
  wire w__9393, w__9394, w__9395, w__9396, w__9397, w__9398, w__9399, w__9400;
  wire w__9401, w__9402, w__9403, w__9404, w__9405, w__9406, w__9407, w__9408;
  wire w__9409, w__9410, w__9411, w__9412, w__9413, w__9414, w__9415, w__9416;
  wire w__9417, w__9418, w__9419, w__9420, w__9421, w__9422, w__9423, w__9424;
  wire w__9425, w__9426, w__9427, w__9428, w__9429, w__9430, w__9431, w__9432;
  wire w__9433, w__9434, w__9435, w__9436, w__9437, w__9438, w__9439, w__9440;
  wire w__9441, w__9442, w__9443, w__9444, w__9445, w__9446, w__9447, w__9448;
  wire w__9449, w__9450, w__9451, w__9452, w__9453, w__9454, w__9455, w__9456;
  wire w__9457, w__9458, w__9459, w__9460, w__9461, w__9462, w__9463, w__9464;
  wire w__9465, w__9466, w__9467, w__9468, w__9469, w__9470, w__9471, w__9472;
  wire w__9473, w__9474, w__9475, w__9476, w__9477, w__9478, w__9479, w__9480;
  wire w__9481, w__9482, w__9483, w__9484, w__9485, w__9486, w__9487, w__9488;
  wire w__9489, w__9490, w__9491, w__9492, w__9493, w__9494, w__9495, w__9496;
  wire w__9497, w__9498, w__9499, w__9500, w__9501, w__9502, w__9503, w__9504;
  wire w__9505, w__9506, w__9507, w__9508, w__9509, w__9510, w__9511, w__9512;
  wire w__9513, w__9514, w__9515, w__9516, w__9517, w__9518, w__9519, w__9520;
  wire w__9521, w__9522, w__9523, w__9524, w__9525, w__9526, w__9527, w__9528;
  wire w__9529, w__9530, w__9531, w__9532, w__9533, w__9534, w__9535, w__9536;
  wire w__9537, w__9538, w__9539, w__9540, w__9541, w__9542, w__9543, w__9544;
  wire w__9545, w__9546, w__9547, w__9548, w__9549, w__9550, w__9551, w__9552;
  wire w__9553, w__9554, w__9555, w__9556, w__9557, w__9558, w__9559, w__9560;
  wire w__9561, w__9562, w__9563, w__9564, w__9565, w__9566, w__9567, w__9568;
  wire w__9569, w__9570, w__9571, w__9572, w__9573, w__9574, w__9575, w__9576;
  wire w__9577, w__9578, w__9579, w__9580, w__9581, w__9582, w__9583, w__9584;
  wire w__9585, w__9586, w__9587, w__9588, w__9589, w__9590, w__9591, w__9592;
  wire w__9593, w__9594, w__9595, w__9596, w__9597, w__9598, w__9599, w__9600;
  wire w__9601, w__9602, w__9603, w__9604, w__9605, w__9606, w__9607, w__9608;
  wire w__9609, w__9610, w__9611, w__9612, w__9613, w__9614, w__9615, w__9616;
  wire w__9617, w__9618, w__9619, w__9620, w__9621, w__9622, w__9623, w__9624;
  wire w__9625, w__9626, w__9627, w__9628, w__9629, w__9630, w__9631, w__9632;
  wire w__9633, w__9634, w__9635, w__9636, w__9637, w__9638, w__9639, w__9640;
  wire w__9641, w__9642, w__9643, w__9644, w__9645, w__9646, w__9647, w__9648;
  wire w__9649, w__9650, w__9651, w__9652, w__9653, w__9654, w__9655, w__9656;
  wire w__9657, w__9658, w__9659, w__9660, w__9661, w__9662, w__9663, w__9664;
  wire w__9665, w__9666, w__9667, w__9668, w__9669, w__9670, w__9671, w__9672;
  wire w__9673, w__9674, w__9675, w__9676, w__9677, w__9678, w__9679, w__9680;
  wire w__9681, w__9682, w__9683, w__9684, w__9685, w__9686, w__9687, w__9688;
  wire w__9689, w__9690, w__9691, w__9692, w__9693, w__9694, w__9695, w__9696;
  wire w__9697, w__9698, w__9699, w__9700, w__9701, w__9702, w__9703, w__9704;
  wire w__9705, w__9706, w__9707, w__9708, w__9709, w__9710, w__9711, w__9712;
  wire w__9713, w__9714, w__9715, w__9716, w__9717, w__9718, w__9719, w__9720;
  wire w__9721, w__9722, w__9723, w__9724, w__9725, w__9726, w__9727, w__9728;
  wire w__9729, w__9730, w__9731, w__9732, w__9733, w__9734, w__9735, w__9736;
  wire w__9737, w__9738, w__9739, w__9740, w__9741, w__9742, w__9743, w__9744;
  wire w__9745, w__9746, w__9747, w__9748, w__9749, w__9750, w__9751, w__9752;
  wire w__9753, w__9754, w__9755, w__9756, w__9757, w__9758, w__9759, w__9760;
  wire w__9761, w__9762, w__9763, w__9764, w__9765, w__9766, w__9767, w__9768;
  wire w__9769, w__9770, w__9771, w__9772, w__9773, w__9774, w__9775, w__9776;
  wire w__9777, w__9778, w__9779, w__9780, w__9781, w__9782, w__9783, w__9784;
  wire w__9785, w__9786, w__9787, w__9788, w__9789, w__9790, w__9791, w__9792;
  wire w__9793, w__9794, w__9795, w__9796, w__9797, w__9798, w__9799, w__9800;
  wire w__9801, w__9802, w__9803, w__9804, w__9805, w__9806, w__9807, w__9808;
  wire w__9809, w__9810, w__9811, w__9812, w__9813, w__9814, w__9815, w__9816;
  wire w__9817, w__9818, w__9819, w__9820, w__9821, w__9822, w__9823, w__9824;
  wire w__9825, w__9826, w__9827, w__9828, w__9829, w__9830, w__9831, w__9832;
  wire w__9833, w__9834, w__9835, w__9836, w__9837, w__9838, w__9839, w__9840;
  wire w__9841, w__9842, w__9843, w__9844, w__9845, w__9846, w__9847, w__9848;
  wire w__9849, w__9850, w__9851, w__9852, w__9853, w__9854, w__9855, w__9856;
  wire w__9857, w__9858, w__9859, w__9860, w__9861, w__9862, w__9863, w__9864;
  wire w__9865, w__9866, w__9867, w__9868, w__9869, w__9870, w__9871, w__9872;
  wire w__9873, w__9874, w__9875, w__9876, w__9877, w__9878, w__9879, w__9880;
  wire w__9881, w__9882, w__9883, w__9884, w__9885, w__9886, w__9887, w__9888;
  wire w__9889, w__9890, w__9891, w__9892, w__9893, w__9894, w__9895, w__9896;
  wire w__9897, w__9898, w__9899, w__9900, w__9901, w__9902, w__9903, w__9904;
  wire w__9905, w__9906, w__9907, w__9908, w__9909, w__9910, w__9911, w__9912;
  wire w__9913, w__9914, w__9915, w__9916, w__9917, w__9918, w__9919, w__9920;
  wire w__9921, w__9922, w__9923, w__9924, w__9925, w__9926, w__9927, w__9928;
  wire w__9929, w__9930, w__9931, w__9932, w__9933, w__9934, w__9935, w__9936;
  wire w__9937, w__9938, w__9939, w__9940, w__9941, w__9942, w__9943, w__9944;
  wire w__9945, w__9946, w__9947, w__9948, w__9949, w__9950, w__9951, w__9952;
  wire w__9953, w__9954, w__9955, w__9956, w__9957, w__9958, w__9959, w__9960;
  wire w__9961, w__9962, w__9963, w__9964, w__9965, w__9966, w__9967, w__9968;
  wire w__9969, w__9970, w__9971, w__9972, w__9973, w__9974, w__9975, w__9976;
  wire w__9977, w__9978, w__9979, w__9980, w__9981, w__9982, w__9983, w__9984;
  wire w__9985, w__9986, w__9987, w__9988, w__9989, w__9990, w__9991, w__9992;
  wire w__9993, w__9994, w__9995, w__9996, w__9997, w__9998, w__9999, w__10000;
  wire w__10001, w__10002, w__10003, w__10004, w__10005, w__10006, w__10007, w__10008;
  wire w__10009, w__10010, w__10011, w__10012, w__10013, w__10014, w__10015, w__10016;
  wire w__10017, w__10018, w__10019, w__10020, w__10021, w__10022, w__10023, w__10024;
  wire w__10025, w__10026, w__10027, w__10028, w__10029, w__10030, w__10031, w__10032;
  wire w__10033, w__10034, w__10035, w__10036, w__10037, w__10038, w__10039, w__10040;
  wire w__10041, w__10042, w__10043, w__10044, w__10045, w__10046, w__10047, w__10048;
  wire w__10049, w__10050, w__10051, w__10052, w__10053, w__10054, w__10055, w__10056;
  wire w__10057, w__10058, w__10059, w__10060, w__10061, w__10062, w__10063, w__10064;
  wire w__10065, w__10066, w__10067, w__10068, w__10069, w__10070, w__10071, w__10072;
  wire w__10073, w__10074, w__10075, w__10076, w__10077, w__10078, w__10079, w__10080;
  wire w__10081, w__10082, w__10083, w__10084, w__10085, w__10086, w__10087, w__10088;
  wire w__10089, w__10090, w__10091, w__10092, w__10093, w__10094, w__10095, w__10096;
  wire w__10097, w__10098, w__10099, w__10100, w__10101, w__10102, w__10103, w__10104;
  wire w__10105, w__10106, w__10107, w__10108, w__10109, w__10110, w__10111, w__10112;
  wire w__10113, w__10114, w__10115, w__10116, w__10117, w__10118, w__10119, w__10120;
  wire w__10121, w__10122, w__10123, w__10124, w__10125, w__10126, w__10127, w__10128;
  wire w__10129, w__10130, w__10131, w__10132, w__10133, w__10134, w__10135, w__10136;
  wire w__10137, w__10138, w__10139, w__10140, w__10141, w__10142, w__10143, w__10144;
  wire w__10145, w__10146, w__10147, w__10148, w__10149, w__10150, w__10151, w__10152;
  wire w__10153, w__10154, w__10155, w__10156, w__10157, w__10158, w__10159, w__10160;
  wire w__10161, w__10162, w__10163, w__10164, w__10165, w__10166, w__10167, w__10168;
  wire w__10169, w__10170, w__10171, w__10172, w__10173, w__10174, w__10175, w__10176;
  wire w__10177, w__10178, w__10179, w__10180, w__10181, w__10182, w__10183, w__10184;
  wire w__10185, w__10186, w__10187, w__10188, w__10189, w__10190, w__10191, w__10192;
  wire w__10193, w__10194, w__10195, w__10196, w__10197, w__10198, w__10199, w__10200;
  wire w__10201, w__10202, w__10203, w__10204, w__10205, w__10206, w__10207, w__10208;
  wire w__10209, w__10210, w__10211, w__10212, w__10213, w__10214, w__10215, w__10216;
  wire w__10217, w__10218, w__10219, w__10220, w__10221, w__10222, w__10223, w__10224;
  wire w__10225, w__10226, w__10227, w__10228, w__10229, w__10230, w__10231, w__10232;
  wire w__10233, w__10234, w__10235, w__10236, w__10237, w__10238, w__10239, w__10240;
  wire w__10241, w__10242, w__10243, w__10244, w__10245, w__10246, w__10247, w__10248;
  wire w__10249, w__10250, w__10251, w__10252, w__10253, w__10254, w__10255, w__10256;
  wire w__10257, w__10258, w__10259, w__10260, w__10261, w__10262, w__10263, w__10264;
  wire w__10265, w__10266, w__10267, w__10268, w__10269, w__10270, w__10271, w__10272;
  wire w__10273, w__10274, w__10275, w__10276, w__10277, w__10278, w__10279, w__10280;
  wire w__10281, w__10282, w__10283, w__10284, w__10285, w__10286, w__10287, w__10288;
  wire w__10289, w__10290, w__10291, w__10292, w__10293, w__10294, w__10295, w__10296;
  wire w__10297, w__10298, w__10299, w__10300, w__10301, w__10302, w__10303, w__10304;
  wire w__10305, w__10306, w__10307, w__10308, w__10309, w__10310, w__10311, w__10312;
  wire w__10313, w__10314, w__10315, w__10316, w__10317, w__10318, w__10319, w__10320;
  wire w__10321, w__10322, w__10323, w__10324, w__10325, w__10326, w__10327, w__10328;
  wire w__10329, w__10330, w__10331, w__10332, w__10333, w__10334, w__10335, w__10336;
  wire w__10337, w__10338, w__10339, w__10340, w__10341, w__10342, w__10343, w__10344;
  wire w__10345, w__10346, w__10347, w__10348, w__10349, w__10350, w__10351, w__10352;
  wire w__10353, w__10354, w__10355, w__10356, w__10357, w__10358, w__10359, w__10360;
  wire w__10361, w__10362, w__10363, w__10364, w__10365, w__10366, w__10367, w__10368;
  wire w__10369, w__10370, w__10371, w__10372, w__10373, w__10374, w__10375, w__10376;
  wire w__10377, w__10378, w__10379, w__10380, w__10381, w__10382, w__10383, w__10384;
  wire w__10385, w__10386, w__10387, w__10388, w__10389, w__10390, w__10391, w__10392;
  wire w__10393, w__10394, w__10395, w__10396, w__10397, w__10398, w__10399, w__10400;
  wire w__10401, w__10402, w__10403, w__10404, w__10405, w__10406, w__10407, w__10408;
  wire w__10409, w__10410, w__10411, w__10412, w__10413, w__10414, w__10415, w__10416;
  wire w__10417, w__10418, w__10419, w__10420, w__10421, w__10422, w__10423, w__10424;
  wire w__10425, w__10426, w__10427, w__10428, w__10429, w__10430, w__10431, w__10432;
  wire w__10433, w__10434, w__10435, w__10436, w__10437, w__10438, w__10439, w__10440;
  wire w__10441, w__10442, w__10443, w__10444, w__10445, w__10446, w__10447, w__10448;
  wire w__10449, w__10450, w__10451, w__10452, w__10453, w__10454, w__10455, w__10456;
  wire w__10457, w__10458, w__10459, w__10460, w__10461, w__10462, w__10463, w__10464;
  wire w__10465, w__10466, w__10467, w__10468, w__10469, w__10470, w__10471, w__10472;
  wire w__10473, w__10474, w__10475, w__10476, w__10477, w__10478, w__10479, w__10480;
  wire w__10481, w__10482, w__10483, w__10484, w__10485, w__10486, w__10487, w__10488;
  wire w__10489, w__10490, w__10491, w__10492, w__10493, w__10494, w__10495, w__10496;
  wire w__10497, w__10498, w__10499, w__10500, w__10501, w__10502, w__10503, w__10504;
  wire w__10505, w__10506, w__10507, w__10508, w__10509, w__10510, w__10511, w__10512;
  wire w__10513, w__10514, w__10515, w__10516, w__10517, w__10518, w__10519, w__10520;
  wire w__10521, w__10522, w__10523, w__10524, w__10525, w__10526, w__10527, w__10528;
  wire w__10529, w__10530, w__10531, w__10532, w__10533, w__10534, w__10535, w__10536;
  wire w__10537, w__10538, w__10539, w__10540, w__10541, w__10542, w__10543, w__10544;
  wire w__10545, w__10546, w__10547, w__10548, w__10549, w__10550, w__10551, w__10552;
  wire w__10553, w__10554, w__10555, w__10556, w__10557, w__10558, w__10559, w__10560;
  wire w__10561, w__10562, w__10563, w__10564, w__10565, w__10566, w__10567, w__10568;
  wire w__10569, w__10570, w__10571, w__10572, w__10573, w__10574, w__10575, w__10576;
  wire w__10577, w__10578, w__10579, w__10580, w__10581, w__10582, w__10583, w__10584;
  wire w__10585, w__10586, w__10587, w__10588, w__10589, w__10590, w__10591, w__10592;
  wire w__10593, w__10594, w__10595, w__10596, w__10597, w__10598, w__10599, w__10600;
  wire w__10601, w__10602, w__10603, w__10604, w__10605, w__10606, w__10607, w__10608;
  wire w__10609, w__10610, w__10611, w__10612, w__10613, w__10614, w__10615, w__10616;
  wire w__10617, w__10618, w__10619, w__10620, w__10621, w__10622, w__10623, w__10624;
  wire w__10625, w__10626, w__10627, w__10628, w__10629, w__10630, w__10631, w__10632;
  wire w__10633, w__10634, w__10635, w__10636, w__10637, w__10638, w__10639, w__10640;
  wire w__10641, w__10642, w__10643, w__10644, w__10645, w__10646, w__10647, w__10648;
  wire w__10649, w__10650, w__10651, w__10652, w__10653, w__10654, w__10655, w__10656;
  wire w__10657, w__10658, w__10659, w__10660, w__10661, w__10662, w__10663, w__10664;
  wire w__10665, w__10666, w__10667, w__10668, w__10669, w__10670, w__10671, w__10672;
  wire w__10673, w__10674, w__10675, w__10676, w__10677, w__10678, w__10679, w__10680;
  wire w__10681, w__10682, w__10683, w__10684, w__10685, w__10686, w__10687, w__10688;
  wire w__10689, w__10690, w__10691, w__10692, w__10693, w__10694, w__10695, w__10696;
  wire w__10697, w__10698, w__10699, w__10700, w__10701, w__10702, w__10703, w__10704;
  wire w__10705, w__10706, w__10707, w__10708, w__10709, w__10710, w__10711, w__10712;
  wire w__10713, w__10714, w__10715, w__10716, w__10717, w__10718, w__10719, w__10720;
  wire w__10721, w__10722, w__10723, w__10724, w__10725, w__10726, w__10727, w__10728;
  wire w__10729, w__10730, w__10731, w__10732, w__10733, w__10734, w__10735, w__10736;
  wire w__10737, w__10738, w__10739, w__10740, w__10741, w__10742, w__10743, w__10744;
  wire w__10745, w__10746, w__10747, w__10748, w__10749, w__10750, w__10751, w__10752;
  wire w__10753, w__10754, w__10755, w__10756, w__10757, w__10758, w__10759, w__10760;
  wire w__10761, w__10762, w__10763, w__10764, w__10765, w__10766, w__10767, w__10768;
  wire w__10769, w__10770, w__10771, w__10772, w__10773, w__10774, w__10775, w__10776;
  wire w__10777, w__10778, w__10779, w__10780, w__10781, w__10782, w__10783, w__10784;
  wire w__10785, w__10786, w__10787, w__10788, w__10789, w__10790, w__10791, w__10792;
  wire w__10793, w__10794, w__10795, w__10796, w__10797, w__10798, w__10799, w__10800;
  wire w__10801, w__10802, w__10803, w__10804, w__10805, w__10806, w__10807, w__10808;
  wire w__10809, w__10810, w__10811, w__10812, w__10813, w__10814, w__10815, w__10816;
  wire w__10817, w__10818, w__10819, w__10820, w__10821, w__10822, w__10823, w__10824;
  wire w__10825, w__10826, w__10827, w__10828, w__10829, w__10830, w__10831, w__10832;
  wire w__10833, w__10834, w__10835, w__10836, w__10837, w__10838, w__10839, w__10840;
  wire w__10841, w__10842, w__10843, w__10844, w__10845, w__10846, w__10847, w__10848;
  wire w__10849, w__10850, w__10851, w__10852, w__10853, w__10854, w__10855, w__10856;
  wire w__10857, w__10858, w__10859, w__10860, w__10861, w__10862, w__10863, w__10864;
  wire w__10865, w__10866, w__10867, w__10868, w__10869, w__10870, w__10871, w__10872;
  wire w__10873, w__10874, w__10875, w__10876, w__10877, w__10878, w__10879, w__10880;
  wire w__10881, w__10882, w__10883, w__10884, w__10885, w__10886, w__10887, w__10888;
  wire w__10889, w__10890, w__10891, w__10892, w__10893, w__10894, w__10895, w__10896;
  wire w__10897, w__10898, w__10899, w__10900, w__10901, w__10902, w__10903, w__10904;
  wire w__10905, w__10906, w__10907, w__10908, w__10909, w__10910, w__10911, w__10912;
  wire w__10913, w__10914, w__10915, w__10916, w__10917, w__10918, w__10919, w__10920;
  wire w__10921, w__10922, w__10923, w__10924, w__10925, w__10926, w__10927, w__10928;
  wire w__10929, w__10930, w__10931, w__10932, w__10933, w__10934, w__10935, w__10936;
  wire w__10937, w__10938, w__10939, w__10940, w__10941, w__10942, w__10943, w__10944;
  wire w__10945, w__10946, w__10947, w__10948, w__10949, w__10950, w__10951, w__10952;
  wire w__10953, w__10954, w__10955, w__10956, w__10957, w__10958, w__10959, w__10960;
  wire w__10961, w__10962, w__10963, w__10964, w__10965, w__10966, w__10967, w__10968;
  wire w__10969, w__10970, w__10971, w__10972, w__10973, w__10974, w__10975, w__10976;
  wire w__10977, w__10978, w__10979, w__10980, w__10981, w__10982, w__10983, w__10984;
  wire w__10985, w__10986, w__10987, w__10988, w__10989, w__10990, w__10991, w__10992;
  wire w__10993, w__10994, w__10995, w__10996, w__10997, w__10998, w__10999, w__11000;
  wire w__11001, w__11002, w__11003, w__11004, w__11005, w__11006, w__11007, w__11008;
  wire w__11009, w__11010, w__11011, w__11012, w__11013, w__11014, w__11015, w__11016;
  wire w__11017, w__11018, w__11019, w__11020, w__11021, w__11022, w__11023, w__11024;
  wire w__11025, w__11026, w__11027, w__11028, w__11029, w__11030, w__11031, w__11032;
  wire w__11033, w__11034, w__11035, w__11036, w__11037, w__11038, w__11039, w__11040;
  wire w__11041, w__11042, w__11043, w__11044, w__11045, w__11046, w__11047, w__11048;
  wire w__11049, w__11050, w__11051, w__11052, w__11053, w__11054, w__11055, w__11056;
  wire w__11057, w__11058, w__11059, w__11060, w__11061, w__11062, w__11063, w__11064;
  wire w__11065, w__11066, w__11067, w__11068, w__11069, w__11070, w__11071, w__11072;
  wire w__11073, w__11074, w__11075, w__11076, w__11077, w__11078, w__11079, w__11080;
  wire w__11081, w__11082, w__11083, w__11084, w__11085, w__11086, w__11087, w__11088;
  wire w__11089, w__11090, w__11091, w__11092, w__11093, w__11094, w__11095, w__11096;
  wire w__11097, w__11098, w__11099, w__11100, w__11101, w__11102, w__11103, w__11104;
  wire w__11105, w__11106, w__11107, w__11108, w__11109, w__11110, w__11111, w__11112;
  wire w__11113, w__11114, w__11115, w__11116, w__11117, w__11118, w__11119, w__11120;
  wire w__11121, w__11122, w__11123, w__11124, w__11125, w__11126, w__11127, w__11128;
  wire w__11129, w__11130, w__11131, w__11132, w__11133, w__11134, w__11135, w__11136;
  wire w__11137, w__11138, w__11139, w__11140, w__11141, w__11142, w__11143, w__11144;
  wire w__11145, w__11146, w__11147, w__11148, w__11149, w__11150, w__11151, w__11152;
  wire w__11153, w__11154, w__11155, w__11156, w__11157, w__11158, w__11159, w__11160;
  wire w__11161, w__11162, w__11163, w__11164, w__11165, w__11166, w__11167, w__11168;
  wire w__11169, w__11170, w__11171, w__11172, w__11173, w__11174, w__11175, w__11176;
  wire w__11177, w__11178, w__11179, w__11180, w__11181, w__11182, w__11183, w__11184;
  wire w__11185, w__11186, w__11187, w__11188, w__11189, w__11190, w__11191, w__11192;
  wire w__11193, w__11194, w__11195, w__11196, w__11197, w__11198, w__11199, w__11200;
  wire w__11201, w__11202, w__11203, w__11204, w__11205, w__11206, w__11207, w__11208;
  wire w__11209, w__11210, w__11211, w__11212, w__11213, w__11214, w__11215, w__11216;
  wire w__11217, w__11218, w__11219, w__11220, w__11221, w__11222, w__11223, w__11224;
  wire w__11225, w__11226, w__11227, w__11228, w__11229, w__11230, w__11231, w__11232;
  wire w__11233, w__11234, w__11235, w__11236, w__11237, w__11238, w__11239, w__11240;
  wire w__11241, w__11242, w__11243, w__11244, w__11245, w__11246, w__11247, w__11248;
  wire w__11249, w__11250, w__11251, w__11252, w__11253, w__11254, w__11255, w__11256;
  wire w__11257, w__11258, w__11259, w__11260, w__11261, w__11262, w__11263, w__11264;
  wire w__11265, w__11266, w__11267, w__11268, w__11269, w__11270, w__11271, w__11272;
  wire w__11273, w__11274, w__11275, w__11276, w__11277, w__11278, w__11279, w__11280;
  wire w__11281, w__11282, w__11283, w__11284, w__11285, w__11286, w__11287, w__11288;
  wire w__11289, w__11290, w__11291, w__11292, w__11293, w__11294, w__11295, w__11296;
  wire w__11297, w__11298, w__11299, w__11300, w__11301, w__11302, w__11303, w__11304;
  wire w__11305, w__11306, w__11307, w__11308, w__11309, w__11310, w__11311, w__11312;
  wire w__11313, w__11314, w__11315, w__11316, w__11317, w__11318, w__11319, w__11320;
  wire w__11321, w__11322, w__11323, w__11324, w__11325, w__11326, w__11327, w__11328;
  wire w__11329, w__11330, w__11331, w__11332, w__11333, w__11334, w__11335, w__11336;
  wire w__11337, w__11338, w__11339, w__11340, w__11341, w__11342, w__11343, w__11344;
  wire w__11345, w__11346, w__11347, w__11348, w__11349, w__11350, w__11351, w__11352;
  wire w__11353, w__11354, w__11355, w__11356, w__11357, w__11358, w__11359, w__11360;
  wire w__11361, w__11362, w__11363, w__11364, w__11365, w__11366, w__11367, w__11368;
  wire w__11369, w__11370, w__11371, w__11372, w__11373, w__11374, w__11375, w__11376;
  wire w__11377, w__11378, w__11379, w__11380, w__11381, w__11382, w__11383, w__11384;
  wire w__11385, w__11386, w__11387, w__11388, w__11389, w__11390, w__11391, w__11392;
  wire w__11393, w__11394, w__11395, w__11396, w__11397, w__11398, w__11399, w__11400;
  wire w__11401, w__11402, w__11403, w__11404, w__11405, w__11406, w__11407, w__11408;
  wire w__11409, w__11410, w__11411, w__11412, w__11413, w__11414, w__11415, w__11416;
  wire w__11417, w__11418, w__11419, w__11420, w__11421, w__11422, w__11423, w__11424;
  wire w__11425, w__11426, w__11427, w__11428, w__11429, w__11430, w__11431, w__11432;
  wire w__11433, w__11434, w__11435, w__11436, w__11437, w__11438, w__11439, w__11440;
  wire w__11441, w__11442, w__11443, w__11444, w__11445, w__11446, w__11447, w__11448;
  wire w__11449, w__11450, w__11451, w__11452, w__11453, w__11454, w__11455, w__11456;
  wire w__11457, w__11458, w__11459, w__11460, w__11461, w__11462, w__11463, w__11464;
  wire w__11465, w__11466, w__11467, w__11468, w__11469, w__11470, w__11471, w__11472;
  wire w__11473, w__11474, w__11475, w__11476, w__11477, w__11478, w__11479, w__11480;
  wire w__11481, w__11482, w__11483, w__11484, w__11485, w__11486, w__11487, w__11488;
  wire w__11489, w__11490, w__11491, w__11492, w__11493, w__11494, w__11495, w__11496;
  wire w__11497, w__11498, w__11499, w__11500, w__11501, w__11502, w__11503, w__11504;
  wire w__11505, w__11506, w__11507, w__11508, w__11509, w__11510, w__11511, w__11512;
  wire w__11513, w__11514, w__11515, w__11516, w__11517, w__11518, w__11519, w__11520;
  wire w__11521, w__11522, w__11523, w__11524, w__11525, w__11526, w__11527, w__11528;
  wire w__11529, w__11530, w__11531, w__11532, w__11533, w__11534, w__11535, w__11536;
  wire w__11537, w__11538, w__11539, w__11540, w__11541, w__11542, w__11543, w__11544;
  wire w__11545, w__11546, w__11547, w__11548, w__11549, w__11550, w__11551, w__11552;
  wire w__11553, w__11554, w__11555, w__11556, w__11557, w__11558, w__11559, w__11560;
  wire w__11561, w__11562, w__11563, w__11564, w__11565, w__11566, w__11567, w__11568;
  wire w__11569, w__11570, w__11571, w__11572, w__11573, w__11574, w__11575, w__11576;
  wire w__11577, w__11578, w__11579, w__11580, w__11581, w__11582, w__11583, w__11584;
  wire w__11585, w__11586, w__11587, w__11588, w__11589, w__11590, w__11591, w__11592;
  wire w__11593, w__11594, w__11595, w__11596, w__11597, w__11598, w__11599, w__11600;
  wire w__11601, w__11602, w__11603, w__11604, w__11605, w__11606, w__11607, w__11608;
  wire w__11609, w__11610, w__11611, w__11612, w__11613, w__11614, w__11615, w__11616;
  wire w__11617, w__11618, w__11619, w__11620, w__11621, w__11622, w__11623, w__11624;
  wire w__11625, w__11626, w__11627, w__11628, w__11629, w__11630, w__11631, w__11632;
  wire w__11633, w__11634, w__11635, w__11636, w__11637, w__11638, w__11639, w__11640;
  wire w__11641, w__11642, w__11643, w__11644, w__11645, w__11646, w__11647, w__11648;
  wire w__11649, w__11650, w__11651, w__11652, w__11653, w__11654, w__11655, w__11656;
  wire w__11657, w__11658, w__11659, w__11660, w__11661, w__11662, w__11663, w__11664;
  wire w__11665, w__11666, w__11667, w__11668, w__11669, w__11670, w__11671, w__11672;
  wire w__11673, w__11674, w__11675, w__11676, w__11677, w__11678, w__11679, w__11680;
  wire w__11681, w__11682, w__11683, w__11684, w__11685, w__11686, w__11687, w__11688;
  wire w__11689, w__11690, w__11691, w__11692, w__11693, w__11694, w__11695, w__11696;
  wire w__11697, w__11698, w__11699, w__11700, w__11701, w__11702, w__11703, w__11704;
  wire w__11705, w__11706, w__11707, w__11708, w__11709, w__11710, w__11711, w__11712;
  wire w__11713, w__11714, w__11715, w__11716, w__11717, w__11718, w__11719, w__11720;
  wire w__11721, w__11722, w__11723, w__11724, w__11725, w__11726, w__11727, w__11728;
  wire w__11729, w__11730, w__11731, w__11732, w__11733, w__11734, w__11735, w__11736;
  wire w__11737, w__11738, w__11739, w__11740, w__11741, w__11742, w__11743, w__11744;
  wire w__11745, w__11746, w__11747, w__11748, w__11749, w__11750, w__11751, w__11752;
  wire w__11753, w__11754, w__11755, w__11756, w__11757, w__11758, w__11759, w__11760;
  wire w__11761, w__11762, w__11763, w__11764, w__11765, w__11766, w__11767, w__11768;
  wire w__11769, w__11770, w__11771, w__11772, w__11773, w__11774, w__11775, w__11776;
  wire w__11777, w__11778, w__11779, w__11780, w__11781, w__11782, w__11783, w__11784;
  wire w__11785, w__11786, w__11787, w__11788, w__11789, w__11790, w__11791, w__11792;
  wire w__11793, w__11794, w__11795, w__11796, w__11797, w__11798, w__11799, w__11800;
  wire w__11801, w__11802, w__11803, w__11804, w__11805, w__11806, w__11807, w__11808;
  wire w__11809, w__11810, w__11811, w__11812, w__11813, w__11814, w__11815, w__11816;
  wire w__11817, w__11818, w__11819, w__11820, w__11821, w__11822, w__11823, w__11824;
  wire w__11825, w__11826, w__11827, w__11828, w__11829, w__11830, w__11831, w__11832;
  wire w__11833, w__11834, w__11835, w__11836, w__11837, w__11838, w__11839, w__11840;
  wire w__11841, w__11842, w__11843, w__11844, w__11845, w__11846, w__11847, w__11848;
  wire w__11849, w__11850, w__11851, w__11852, w__11853, w__11854, w__11855, w__11856;
  wire w__11857, w__11858, w__11859, w__11860, w__11861, w__11862, w__11863, w__11864;
  wire w__11865, w__11866, w__11867, w__11868, w__11869, w__11870, w__11871, w__11872;
  wire w__11873, w__11874, w__11875, w__11876, w__11877, w__11878, w__11879, w__11880;
  wire w__11881, w__11882, w__11883, w__11884, w__11885, w__11886, w__11887, w__11888;
  wire w__11889, w__11890, w__11891, w__11892, w__11893, w__11894, w__11895, w__11896;
  wire w__11897, w__11898, w__11899, w__11900, w__11901, w__11902, w__11903, w__11904;
  wire w__11905, w__11906, w__11907, w__11908, w__11909, w__11910, w__11911, w__11912;
  wire w__11913, w__11914, w__11915, w__11916, w__11917, w__11918, w__11919, w__11920;
  wire w__11921, w__11922, w__11923, w__11924, w__11925, w__11926, w__11927, w__11928;
  wire w__11929, w__11930, w__11931, w__11932, w__11933, w__11934, w__11935, w__11936;
  wire w__11937, w__11938, w__11939, w__11940, w__11941, w__11942, w__11943, w__11944;
  wire w__11945, w__11946, w__11947, w__11948, w__11949, w__11950, w__11951, w__11952;
  wire w__11953, w__11954, w__11955, w__11956, w__11957, w__11958, w__11959, w__11960;
  wire w__11961, w__11962, w__11963, w__11964, w__11965, w__11966, w__11967, w__11968;
  wire w__11969, w__11970, w__11971, w__11972, w__11973, w__11974, w__11975, w__11976;
  wire w__11977, w__11978, w__11979, w__11980, w__11981, w__11982, w__11983, w__11984;
  wire w__11985, w__11986, w__11987, w__11988, w__11989, w__11990, w__11991, w__11992;
  wire w__11993, w__11994, w__11995, w__11996, w__11997, w__11998, w__11999, w__12000;
  wire w__12001, w__12002, w__12003, w__12004, w__12005, w__12006, w__12007, w__12008;
  wire w__12009, w__12010, w__12011, w__12012, w__12013, w__12014, w__12015, w__12016;
  wire w__12017, w__12018, w__12019, w__12020, w__12021, w__12022, w__12023, w__12024;
  wire w__12025, w__12026, w__12027, w__12028, w__12029, w__12030, w__12031, w__12032;
  wire w__12033, w__12034, w__12035, w__12036, w__12037, w__12038, w__12039, w__12040;
  wire w__12041, w__12042, w__12043, w__12044, w__12045, w__12046, w__12047, w__12048;
  wire w__12049, w__12050, w__12051, w__12052, w__12053, w__12054, w__12055, w__12056;
  wire w__12057, w__12058, w__12059, w__12060, w__12061, w__12062, w__12063, w__12064;
  wire w__12065, w__12066, w__12067, w__12068, w__12069, w__12070, w__12071, w__12072;
  wire w__12073, w__12074, w__12075, w__12076, w__12077, w__12078, w__12079, w__12080;
  wire w__12081, w__12082, w__12083, w__12084, w__12085, w__12086, w__12087, w__12088;
  wire w__12089, w__12090, w__12091, w__12092, w__12093, w__12094, w__12095, w__12096;
  wire w__12097, w__12098, w__12099, w__12100, w__12101, w__12102, w__12103, w__12104;
  wire w__12105, w__12106, w__12107, w__12108, w__12109, w__12110, w__12111, w__12112;
  wire w__12113, w__12114, w__12115, w__12116, w__12117, w__12118, w__12119, w__12120;
  wire w__12121, w__12122, w__12123, w__12124, w__12125, w__12126, w__12127, w__12128;
  wire w__12129, w__12130, w__12131, w__12132, w__12133, w__12134, w__12135, w__12136;
  wire w__12137, w__12138, w__12139, w__12140, w__12141, w__12142, w__12143, w__12144;
  wire w__12145, w__12146, w__12147, w__12148, w__12149, w__12150, w__12151, w__12152;
  wire w__12153, w__12154, w__12155, w__12156, w__12157, w__12158, w__12159, w__12160;
  wire w__12161, w__12162, w__12163, w__12164, w__12165, w__12166, w__12167, w__12168;
  wire w__12169, w__12170, w__12171, w__12172, w__12173, w__12174, w__12175, w__12176;
  wire w__12177, w__12178, w__12179, w__12180, w__12181, w__12182, w__12183, w__12184;
  wire w__12185, w__12186, w__12187, w__12188, w__12189, w__12190, w__12191, w__12192;
  wire w__12193, w__12194, w__12195, w__12196, w__12197, w__12198, w__12199, w__12200;
  wire w__12201, w__12202, w__12203, w__12204, w__12205, w__12206, w__12207, w__12208;
  wire w__12209, w__12210, w__12211, w__12212, w__12213, w__12214, w__12215, w__12216;
  wire w__12217, w__12218, w__12219, w__12220, w__12221, w__12222, w__12223, w__12224;
  wire w__12225, w__12226, w__12227, w__12228, w__12229, w__12230, w__12231, w__12232;
  wire w__12233, w__12234, w__12235, w__12236, w__12237, w__12238, w__12239, w__12240;
  wire w__12241, w__12242, w__12243, w__12244, w__12245, w__12246, w__12247, w__12248;
  wire w__12249, w__12250, w__12251, w__12252, w__12253, w__12254, w__12255, w__12256;
  wire w__12257, w__12258, w__12259, w__12260, w__12261, w__12262, w__12263, w__12264;
  wire w__12265, w__12266, w__12267, w__12268, w__12269, w__12270, w__12271, w__12272;
  wire w__12273, w__12274, w__12275, w__12276, w__12277, w__12278, w__12279, w__12280;
  wire w__12281, w__12282, w__12283, w__12284, w__12285, w__12286, w__12287, w__12288;
  wire w__12289, w__12290, w__12291, w__12292, w__12293, w__12294, w__12295, w__12296;
  wire w__12297, w__12298, w__12299, w__12300, w__12301, w__12302, w__12303, w__12304;
  wire w__12305, w__12306, w__12307, w__12308, w__12309, w__12310, w__12311, w__12312;
  wire w__12313, w__12314, w__12315, w__12316, w__12317, w__12318, w__12319, w__12320;
  wire w__12321, w__12322, w__12323, w__12324, w__12325, w__12326, w__12327, w__12328;
  wire w__12329, w__12330, w__12331, w__12332, w__12333, w__12334, w__12335, w__12336;
  wire w__12337, w__12338, w__12339, w__12340, w__12341, w__12342, w__12343, w__12344;
  wire w__12345, w__12346, w__12347, w__12348, w__12349, w__12350, w__12351, w__12352;
  wire w__12353, w__12354, w__12355, w__12356, w__12357, w__12358, w__12359, w__12360;
  wire w__12361, w__12362, w__12363, w__12364, w__12365, w__12366, w__12367, w__12368;
  wire w__12369, w__12370, w__12371, w__12372, w__12373, w__12374, w__12375, w__12376;
  wire w__12377, w__12378, w__12379, w__12380, w__12381, w__12382, w__12383, w__12384;
  wire w__12385, w__12386, w__12387, w__12388, w__12389, w__12390, w__12391, w__12392;
  wire w__12393, w__12394, w__12395, w__12396, w__12397, w__12398, w__12399, w__12400;
  wire w__12401, w__12402, w__12403, w__12404, w__12405, w__12406, w__12407, w__12408;
  wire w__12409, w__12410, w__12411, w__12412, w__12413, w__12414, w__12415, w__12416;
  wire w__12417, w__12418, w__12419, w__12420, w__12421, w__12422, w__12423, w__12424;
  wire w__12425, w__12426, w__12427, w__12428, w__12429, w__12430, w__12431, w__12432;
  wire w__12433, w__12434, w__12435, w__12436, w__12437, w__12438, w__12439, w__12440;
  wire w__12441, w__12442, w__12443, w__12444, w__12445, w__12446, w__12447, w__12448;
  wire w__12449, w__12450, w__12451, w__12452, w__12453, w__12454, w__12455, w__12456;
  wire w__12457, w__12458, w__12459, w__12460, w__12461, w__12462, w__12463, w__12464;
  wire w__12465, w__12466, w__12467, w__12468, w__12469, w__12470, w__12471, w__12472;
  wire w__12473, w__12474, w__12475, w__12476, w__12477, w__12478, w__12479, w__12480;
  wire w__12481, w__12482, w__12483, w__12484, w__12485, w__12486, w__12487, w__12488;
  wire w__12489, w__12490, w__12491, w__12492, w__12493, w__12494, w__12495, w__12496;
  wire w__12497, w__12498, w__12499, w__12500, w__12501, w__12502, w__12503, w__12504;
  wire w__12505, w__12506, w__12507, w__12508, w__12509, w__12510, w__12511, w__12512;
  wire w__12513, w__12514, w__12515, w__12516, w__12517, w__12518, w__12519, w__12520;
  wire w__12521, w__12522, w__12523, w__12524, w__12525, w__12526, w__12527, w__12528;
  wire w__12529, w__12530, w__12531, w__12532, w__12533, w__12534, w__12535, w__12536;
  wire w__12537, w__12538, w__12539, w__12540, w__12541, w__12542, w__12543, w__12544;
  wire w__12545, w__12546, w__12547, w__12548, w__12549, w__12550, w__12551, w__12552;
  wire w__12553, w__12554, w__12555, w__12556, w__12557, w__12558, w__12559, w__12560;
  wire w__12561, w__12562, w__12563, w__12564, w__12565, w__12566, w__12567, w__12568;
  wire w__12569, w__12570, w__12571, w__12572, w__12573, w__12574, w__12575, w__12576;
  wire w__12577, w__12578, w__12579, w__12580, w__12581, w__12582, w__12583, w__12584;
  wire w__12585, w__12586, w__12587, w__12588, w__12589, w__12590, w__12591, w__12592;
  wire w__12593, w__12594, w__12595, w__12596, w__12597, w__12598, w__12599, w__12600;
  wire w__12601, w__12602, w__12603, w__12604, w__12605, w__12606, w__12607, w__12608;
  wire w__12609, w__12610, w__12611, w__12612, w__12613, w__12614, w__12615, w__12616;
  wire w__12617, w__12618, w__12619, w__12620, w__12621, w__12622, w__12623, w__12624;
  wire w__12625, w__12626, w__12627, w__12628, w__12629, w__12630, w__12631, w__12632;
  wire w__12633, w__12634, w__12635, w__12636, w__12637, w__12638, w__12639, w__12640;
  wire w__12641, w__12642, w__12643, w__12644, w__12645, w__12646, w__12647, w__12648;
  wire w__12649, w__12650, w__12651, w__12652, w__12653, w__12654, w__12655, w__12656;
  wire w__12657, w__12658, w__12659, w__12660, w__12661, w__12662, w__12663, w__12664;
  wire w__12665, w__12666, w__12667, w__12668, w__12669, w__12670, w__12671, w__12672;
  wire w__12673, w__12674, w__12675, w__12676, w__12677, w__12678, w__12679, w__12680;
  wire w__12681, w__12682, w__12683, w__12684, w__12685, w__12686, w__12687, w__12688;
  wire w__12689, w__12690, w__12691, w__12692, w__12693, w__12694, w__12695, w__12696;
  wire w__12697, w__12698, w__12699, w__12700, w__12701, w__12702, w__12703, w__12704;
  wire w__12705, w__12706, w__12707, w__12708, w__12709, w__12710, w__12711, w__12712;
  wire w__12713, w__12714, w__12715, w__12716, w__12717, w__12718, w__12719, w__12720;
  wire w__12721, w__12722, w__12723, w__12724, w__12725, w__12726, w__12727, w__12728;
  wire w__12729, w__12730, w__12731, w__12732, w__12733, w__12734, w__12735, w__12736;
  wire w__12737, w__12738, w__12739, w__12740, w__12741, w__12742, w__12743, w__12744;
  wire w__12745, w__12746, w__12747, w__12748, w__12749, w__12750, w__12751, w__12752;
  wire w__12753, w__12754, w__12755, w__12756, w__12757, w__12758, w__12759, w__12760;
  wire w__12761, w__12762, w__12763, w__12764, w__12765, w__12766, w__12767, w__12768;
  wire w__12769, w__12770, w__12771, w__12772, w__12773, w__12774, w__12775, w__12776;
  wire w__12777, w__12778, w__12779, w__12780, w__12781, w__12782, w__12783, w__12784;
  wire w__12785, w__12786, w__12787, w__12788, w__12789, w__12790, w__12791, w__12792;
  wire w__12793, w__12794, w__12795, w__12796, w__12797, w__12798, w__12799, w__12800;
  wire w__12801, w__12802, w__12803, w__12804, w__12805, w__12806, w__12807, w__12808;
  wire w__12809, w__12810, w__12811, w__12812, w__12813, w__12814, w__12815, w__12816;
  wire w__12817, w__12818, w__12819, w__12820, w__12821, w__12822, w__12823, w__12824;
  wire w__12825, w__12826, w__12827, w__12828, w__12829, w__12830, w__12831, w__12832;
  wire w__12833, w__12834, w__12835, w__12836, w__12837, w__12838, w__12839, w__12840;
  wire w__12841, w__12842, w__12843, w__12844, w__12845, w__12846, w__12847, w__12848;
  wire w__12849, w__12850, w__12851, w__12852, w__12853, w__12854, w__12855, w__12856;
  wire w__12857, w__12858, w__12859, w__12860, w__12861, w__12862, w__12863, w__12864;
  wire w__12865, w__12866, w__12867, w__12868, w__12869, w__12870, w__12871, w__12872;
  wire w__12873, w__12874, w__12875, w__12876, w__12877, w__12878, w__12879, w__12880;
  wire w__12881, w__12882, w__12883, w__12884, w__12885, w__12886, w__12887, w__12888;
  wire w__12889, w__12890, w__12891, w__12892, w__12893, w__12894, w__12895, w__12896;
  wire w__12897, w__12898, w__12899, w__12900, w__12901, w__12902, w__12903, w__12904;
  wire w__12905, w__12906, w__12907, w__12908, w__12909, w__12910, w__12911, w__12912;
  wire w__12913, w__12914, w__12915, w__12916, w__12917, w__12918, w__12919, w__12920;
  wire w__12921, w__12922, w__12923, w__12924, w__12925, w__12926, w__12927, w__12928;
  wire w__12929, w__12930, w__12931, w__12932, w__12933, w__12934, w__12935, w__12936;
  wire w__12937, w__12938, w__12939, w__12940, w__12941, w__12942, w__12943, w__12944;
  wire w__12945, w__12946, w__12947, w__12948, w__12949, w__12950, w__12951, w__12952;
  wire w__12953, w__12954, w__12955, w__12956, w__12957, w__12958, w__12959, w__12960;
  wire w__12961, w__12962, w__12963, w__12964, w__12965, w__12966, w__12967, w__12968;
  wire w__12969, w__12970, w__12971, w__12972, w__12973, w__12974, w__12975, w__12976;
  wire w__12977, w__12978, w__12979, w__12980, w__12981, w__12982, w__12983, w__12984;
  wire w__12985, w__12986, w__12987, w__12988, w__12989, w__12990, w__12991, w__12992;
  wire w__12993, w__12994, w__12995, w__12996, w__12997, w__12998, w__12999, w__13000;
  wire w__13001, w__13002, w__13003, w__13004, w__13005, w__13006, w__13007, w__13008;
  wire w__13009, w__13010, w__13011, w__13012, w__13013, w__13014, w__13015, w__13016;
  wire w__13017, w__13018, w__13019, w__13020, w__13021, w__13022, w__13023, w__13024;
  wire w__13025, w__13026, w__13027, w__13028, w__13029, w__13030, w__13031, w__13032;
  wire w__13033, w__13034, w__13035, w__13036, w__13037, w__13038, w__13039, w__13040;
  wire w__13041, w__13042, w__13043, w__13044, w__13045, w__13046, w__13047, w__13048;
  wire w__13049, w__13050, w__13051, w__13052, w__13053, w__13054, w__13055, w__13056;
  wire w__13057, w__13058, w__13059, w__13060, w__13061, w__13062, w__13063, w__13064;
  wire w__13065, w__13066, w__13067, w__13068, w__13069, w__13070, w__13071, w__13072;
  wire w__13073, w__13074, w__13075, w__13076, w__13077, w__13078, w__13079, w__13080;
  wire w__13081, w__13082, w__13083, w__13084, w__13085, w__13086, w__13087, w__13088;
  wire w__13089, w__13090, w__13091, w__13092, w__13093, w__13094, w__13095, w__13096;
  wire w__13097, w__13098, w__13099, w__13100, w__13101, w__13102, w__13103, w__13104;
  wire w__13105, w__13106, w__13107, w__13108, w__13109, w__13110, w__13111, w__13112;
  wire w__13113, w__13114, w__13115, w__13116, w__13117, w__13118, w__13119, w__13120;
  wire w__13121, w__13122, w__13123, w__13124, w__13125, w__13126, w__13127, w__13128;
  wire w__13129, w__13130, w__13131, w__13132, w__13133, w__13134, w__13135, w__13136;
  wire w__13137, w__13138, w__13139, w__13140, w__13141, w__13142, w__13143, w__13144;
  wire w__13145, w__13146, w__13147, w__13148, w__13149, w__13150, w__13151, w__13152;
  wire w__13153, w__13154, w__13155, w__13156, w__13157, w__13158, w__13159, w__13160;
  wire w__13161, w__13162, w__13163, w__13164, w__13165, w__13166, w__13167, w__13168;
  wire w__13169, w__13170, w__13171, w__13172, w__13173, w__13174, w__13175, w__13176;
  wire w__13177, w__13178, w__13179, w__13180, w__13181, w__13182, w__13183, w__13184;
  wire w__13185, w__13186, w__13187, w__13188, w__13189, w__13190, w__13191, w__13192;
  wire w__13193, w__13194, w__13195, w__13196, w__13197, w__13198, w__13199, w__13200;
  wire w__13201, w__13202, w__13203, w__13204, w__13205, w__13206, w__13207, w__13208;
  wire w__13209, w__13210, w__13211, w__13212, w__13213, w__13214, w__13215, w__13216;
  wire w__13217, w__13218, w__13219, w__13220, w__13221, w__13222, w__13223, w__13224;
  wire w__13225, w__13226, w__13227, w__13228, w__13229, w__13230, w__13231, w__13232;
  wire w__13233, w__13234, w__13235, w__13236, w__13237, w__13238, w__13239, w__13240;
  wire w__13241, w__13242, w__13243, w__13244, w__13245, w__13246, w__13247, w__13248;
  wire w__13249, w__13250, w__13251, w__13252, w__13253, w__13254, w__13255, w__13256;
  wire w__13257, w__13258, w__13259, w__13260, w__13261, w__13262, w__13263, w__13264;
  wire w__13265, w__13266, w__13267, w__13268, w__13269, w__13270, w__13271, w__13272;
  wire w__13273, w__13274, w__13275, w__13276, w__13277, w__13278, w__13279, w__13280;
  wire w__13281, w__13282, w__13283, w__13284, w__13285, w__13286, w__13287, w__13288;
  wire w__13289, w__13290, w__13291, w__13292, w__13293, w__13294, w__13295, w__13296;
  wire w__13297, w__13298, w__13299, w__13300, w__13301, w__13302, w__13303, w__13304;
  wire w__13305, w__13306, w__13307, w__13308, w__13309, w__13310, w__13311, w__13312;
  wire w__13313, w__13314, w__13315, w__13316, w__13317, w__13318, w__13319, w__13320;
  wire w__13321, w__13322, w__13323, w__13324, w__13325, w__13326, w__13327, w__13328;
  wire w__13329, w__13330, w__13331, w__13332, w__13333, w__13334, w__13335, w__13336;
  wire w__13337, w__13338, w__13339, w__13340, w__13341, w__13342, w__13343, w__13344;
  wire w__13345, w__13346, w__13347, w__13348, w__13349, w__13350, w__13351, w__13352;
  wire w__13353, w__13354, w__13355, w__13356, w__13357, w__13358, w__13359, w__13360;
  wire w__13361, w__13362, w__13363, w__13364, w__13365, w__13366, w__13367, w__13368;
  wire w__13369, w__13370, w__13371, w__13372, w__13373, w__13374, w__13375, w__13376;
  wire w__13377, w__13378, w__13379, w__13380, w__13381, w__13382, w__13383, w__13384;
  wire w__13385, w__13386, w__13387, w__13388, w__13389, w__13390, w__13391, w__13392;
  wire w__13393, w__13394, w__13395, w__13396, w__13397, w__13398, w__13399, w__13400;
  wire w__13401, w__13402, w__13403, w__13404, w__13405, w__13406, w__13407, w__13408;
  wire w__13409, w__13410, w__13411, w__13412, w__13413, w__13414, w__13415, w__13416;
  wire w__13417, w__13418, w__13419, w__13420, w__13421, w__13422, w__13423, w__13424;
  wire w__13425, w__13426, w__13427, w__13428, w__13429, w__13430, w__13431, w__13432;
  wire w__13433, w__13434, w__13435, w__13436, w__13437, w__13438, w__13439, w__13440;
  wire w__13441, w__13442, w__13443, w__13444, w__13445, w__13446, w__13447, w__13448;
  wire w__13449, w__13450, w__13451, w__13452, w__13453, w__13454, w__13455, w__13456;
  wire w__13457, w__13458, w__13459, w__13460, w__13461, w__13462, w__13463, w__13464;
  wire w__13465, w__13466, w__13467, w__13468, w__13469, w__13470, w__13471, w__13472;
  wire w__13473, w__13474, w__13475, w__13476, w__13477, w__13478, w__13479, w__13480;
  wire w__13481, w__13482, w__13483, w__13484, w__13485, w__13486, w__13487, w__13488;
  wire w__13489, w__13490, w__13491, w__13492, w__13493, w__13494, w__13495, w__13496;
  wire w__13497, w__13498, w__13499, w__13500, w__13501, w__13502, w__13503, w__13504;
  wire w__13505, w__13506, w__13507, w__13508, w__13509, w__13510, w__13511, w__13512;
  wire w__13513, w__13514, w__13515, w__13516, w__13517, w__13518, w__13519, w__13520;
  wire w__13521, w__13522, w__13523, w__13524, w__13525, w__13526, w__13527, w__13528;
  wire w__13529, w__13530, w__13531, w__13532, w__13533, w__13534, w__13535, w__13536;
  wire w__13537, w__13538, w__13539, w__13540, w__13541, w__13542, w__13543, w__13544;
  wire w__13545, w__13546, w__13547, w__13548, w__13549, w__13550, w__13551, w__13552;
  wire w__13553, w__13554, w__13555, w__13556, w__13557, w__13558, w__13559, w__13560;
  wire w__13561, w__13562, w__13563, w__13564, w__13565, w__13566, w__13567, w__13568;
  wire w__13569, w__13570, w__13571, w__13572, w__13573, w__13574, w__13575, w__13576;
  wire w__13577, w__13578, w__13579, w__13580, w__13581, w__13582, w__13583, w__13584;
  wire w__13585, w__13586, w__13587, w__13588, w__13589, w__13590, w__13591, w__13592;
  wire w__13593, w__13594, w__13595, w__13596, w__13597, w__13598, w__13599, w__13600;
  wire w__13601, w__13602, w__13603, w__13604, w__13605, w__13606, w__13607, w__13608;
  wire w__13609, w__13610, w__13611, w__13612, w__13613, w__13614, w__13615, w__13616;
  wire w__13617, w__13618, w__13619, w__13620, w__13621, w__13622, w__13623, w__13624;
  wire w__13625, w__13626, w__13627, w__13628, w__13629, w__13630, w__13631, w__13632;
  wire w__13633, w__13634, w__13635, w__13636, w__13637, w__13638, w__13639, w__13640;
  wire w__13641, w__13642, w__13643, w__13644, w__13645, w__13646, w__13647, w__13648;
  wire w__13649, w__13650, w__13651, w__13652, w__13653, w__13654, w__13655, w__13656;
  wire w__13657, w__13658, w__13659, w__13660, w__13661, w__13662, w__13663, w__13664;
  wire w__13665, w__13666, w__13667, w__13668, w__13669, w__13670, w__13671, w__13672;
  wire w__13673, w__13674, w__13675, w__13676, w__13677, w__13678, w__13679, w__13680;
  wire w__13681, w__13682, w__13683, w__13684, w__13685, w__13686, w__13687, w__13688;
  wire w__13689, w__13690, w__13691, w__13692, w__13693, w__13694, w__13695, w__13696;
  wire w__13697, w__13698, w__13699, w__13700, w__13701, w__13702, w__13703, w__13704;
  wire w__13705, w__13706, w__13707, w__13708, w__13709, w__13710, w__13711, w__13712;
  wire w__13713, w__13714, w__13715, w__13716, w__13717, w__13718, w__13719, w__13720;
  wire w__13721, w__13722, w__13723, w__13724, w__13725, w__13726, w__13727, w__13728;
  wire w__13729, w__13730, w__13731, w__13732, w__13733, w__13734, w__13735, w__13736;
  wire w__13737, w__13738, w__13739, w__13740, w__13741, w__13742, w__13743, w__13744;
  wire w__13745, w__13746, w__13747, w__13748, w__13749, w__13750, w__13751, w__13752;
  wire w__13753, w__13754, w__13755, w__13756, w__13757, w__13758, w__13759, w__13760;
  wire w__13761, w__13762, w__13763, w__13764, w__13765, w__13766, w__13767, w__13768;
  wire w__13769, w__13770, w__13771, w__13772, w__13773, w__13774, w__13775, w__13776;
  wire w__13777, w__13778, w__13779, w__13780, w__13781, w__13782, w__13783, w__13784;
  wire w__13785, w__13786, w__13787, w__13788, w__13789, w__13790, w__13791, w__13792;
  wire w__13793, w__13794, w__13795, w__13796, w__13797, w__13798, w__13799, w__13800;
  wire w__13801, w__13802, w__13803, w__13804, w__13805, w__13806, w__13807, w__13808;
  wire w__13809, w__13810, w__13811, w__13812, w__13813, w__13814, w__13815, w__13816;
  wire w__13817, w__13818, w__13819, w__13820, w__13821, w__13822, w__13823, w__13824;
  wire w__13825, w__13826, w__13827, w__13828, w__13829, w__13830, w__13831, w__13832;
  wire w__13833, w__13834, w__13835, w__13836, w__13837, w__13838, w__13839, w__13840;
  wire w__13841, w__13842, w__13843, w__13844, w__13845, w__13846, w__13847, w__13848;
  wire w__13849, w__13850, w__13851, w__13852, w__13853, w__13854, w__13855, w__13856;
  wire w__13857, w__13858, w__13859, w__13860, w__13861, w__13862, w__13863, w__13864;
  wire w__13865, w__13866, w__13867, w__13868, w__13869, w__13870, w__13871, w__13872;
  wire w__13873, w__13874, w__13875, w__13876, w__13877, w__13878, w__13879, w__13880;
  wire w__13881, w__13882, w__13883, w__13884, w__13885, w__13886, w__13887, w__13888;
  wire w__13889, w__13890, w__13891, w__13892, w__13893, w__13894, w__13895, w__13896;
  wire w__13897, w__13898, w__13899, w__13900, w__13901, w__13902, w__13903, w__13904;
  wire w__13905, w__13906, w__13907, w__13908, w__13909, w__13910, w__13911, w__13912;
  wire w__13913, w__13914, w__13915, w__13916, w__13917, w__13918, w__13919, w__13920;
  wire w__13921, w__13922, w__13923, w__13924, w__13925, w__13926, w__13927, w__13928;
  wire w__13929, w__13930, w__13931, w__13932, w__13933, w__13934, w__13935, w__13936;
  wire w__13937, w__13938, w__13939, w__13940, w__13941, w__13942, w__13943, w__13944;
  wire w__13945, w__13946, w__13947, w__13948, w__13949, w__13950, w__13951, w__13952;
  wire w__13953, w__13954, w__13955, w__13956, w__13957, w__13958, w__13959, w__13960;
  wire w__13961, w__13962, w__13963, w__13964, w__13965, w__13966, w__13967, w__13968;
  wire w__13969, w__13970, w__13971, w__13972, w__13973, w__13974, w__13975, w__13976;
  wire w__13977, w__13978, w__13979, w__13980, w__13981, w__13982, w__13983, w__13984;
  wire w__13985, w__13986, w__13987, w__13988, w__13989, w__13990, w__13991, w__13992;
  wire w__13993, w__13994, w__13995, w__13996, w__13997, w__13998, w__13999, w__14000;
  wire w__14001, w__14002, w__14003, w__14004, w__14005, w__14006, w__14007, w__14008;
  wire w__14009, w__14010, w__14011, w__14012, w__14013, w__14014, w__14015, w__14016;
  wire w__14017, w__14018, w__14019, w__14020, w__14021, w__14022, w__14023, w__14024;
  wire w__14025, w__14026, w__14027, w__14028, w__14029, w__14030, w__14031, w__14032;
  wire w__14033, w__14034, w__14035, w__14036, w__14037, w__14038, w__14039, w__14040;
  wire w__14041, w__14042, w__14043, w__14044, w__14045, w__14046, w__14047, w__14048;
  wire w__14049, w__14050, w__14051, w__14052, w__14053, w__14054, w__14055, w__14056;
  wire w__14057, w__14058, w__14059, w__14060, w__14061, w__14062, w__14063, w__14064;
  wire w__14065, w__14066, w__14067, w__14068, w__14069, w__14070, w__14071, w__14072;
  wire w__14073, w__14074, w__14075, w__14076, w__14077, w__14078, w__14079, w__14080;
  wire w__14081, w__14082, w__14083, w__14084, w__14085, w__14086, w__14087, w__14088;
  wire w__14089, w__14090, w__14091, w__14092, w__14093, w__14094, w__14095, w__14096;
  wire w__14097, w__14098, w__14099, w__14100, w__14101, w__14102, w__14103, w__14104;
  wire w__14105, w__14106, w__14107, w__14108, w__14109, w__14110, w__14111, w__14112;
  wire w__14113, w__14114, w__14115, w__14116, w__14117, w__14118, w__14119, w__14120;
  wire w__14121, w__14122, w__14123, w__14124, w__14125, w__14126, w__14127, w__14128;
  wire w__14129, w__14130, w__14131, w__14132, w__14133, w__14134, w__14135, w__14136;
  wire w__14137, w__14138, w__14139, w__14140, w__14141, w__14142, w__14143, w__14144;
  wire w__14145, w__14146, w__14147, w__14148, w__14149, w__14150, w__14151, w__14152;
  wire w__14153, w__14154, w__14155, w__14156, w__14157, w__14158, w__14159, w__14160;
  wire w__14161, w__14162, w__14163, w__14164, w__14165, w__14166, w__14167, w__14168;
  wire w__14169, w__14170, w__14171, w__14172, w__14173, w__14174, w__14175, w__14176;
  wire w__14177, w__14178, w__14179, w__14180, w__14181, w__14182, w__14183, w__14184;
  wire w__14185, w__14186, w__14187, w__14188, w__14189, w__14190, w__14191, w__14192;
  wire w__14193, w__14194, w__14195, w__14196, w__14197, w__14198, w__14199, w__14200;
  wire w__14201, w__14202, w__14203, w__14204, w__14205, w__14206, w__14207, w__14208;
  wire w__14209, w__14210, w__14211, w__14212, w__14213, w__14214, w__14215, w__14216;
  wire w__14217, w__14218, w__14219, w__14220, w__14221, w__14222, w__14223, w__14224;
  wire w__14225, w__14226, w__14227, w__14228, w__14229, w__14230, w__14231, w__14232;
  wire w__14233, w__14234, w__14235, w__14236, w__14237, w__14238, w__14239, w__14240;
  wire w__14241, w__14242, w__14243, w__14244, w__14245, w__14246, w__14247, w__14248;
  wire w__14249, w__14250, w__14251, w__14252, w__14253, w__14254, w__14255, w__14256;
  wire w__14257, w__14258, w__14259, w__14260, w__14261, w__14262, w__14263, w__14264;
  wire w__14265, w__14266, w__14267, w__14268, w__14269, w__14270, w__14271, w__14272;
  wire w__14273, w__14274, w__14275, w__14276, w__14277, w__14278, w__14279, w__14280;
  wire w__14281, w__14282, w__14283, w__14284, w__14285, w__14286, w__14287, w__14288;
  wire w__14289, w__14290, w__14291, w__14292, w__14293, w__14294, w__14295, w__14296;
  wire w__14297, w__14298, w__14299, w__14300, w__14301, w__14302, w__14303, w__14304;
  wire w__14305, w__14306, w__14307, w__14308, w__14309, w__14310, w__14311, w__14312;
  wire w__14313, w__14314, w__14315, w__14316, w__14317, w__14318, w__14319, w__14320;
  wire w__14321, w__14322, w__14323, w__14324, w__14325, w__14326, w__14327, w__14328;
  wire w__14329, w__14330, w__14331, w__14332, w__14333, w__14334, w__14335, w__14336;
  wire w__14337, w__14338, w__14339;
  buf g__1(w__13188 ,w__13057);
  buf g__2(w__13187 ,w__13058);
  buf g__3(w__13186 ,w__13056);
  buf g__4(w__13185 ,w__13055);
  buf g__5(w__13184 ,w__13053);
  buf g__6(w__13183 ,w__13054);
  buf g__7(w__13182 ,w__13052);
  buf g__8(w__13181 ,w__13051);
  buf g__9(w__13148 ,w__13050);
  buf g__10(w__13147 ,w__13049);
  buf g__11(w__13146 ,w__13048);
  buf g__12(w__13145 ,w__13047);
  buf g__13(w__13144 ,w__13030);
  buf g__14(w__13143 ,w__13045);
  buf g__15(w__13142 ,w__13044);
  buf g__16(w__13141 ,w__13043);
  buf g__17(w__13140 ,w__13042);
  buf g__18(w__13139 ,w__13041);
  buf g__19(w__13138 ,w__13040);
  buf g__20(w__13137 ,w__13039);
  buf g__21(w__13136 ,w__13038);
  buf g__22(w__13135 ,w__13037);
  buf g__23(w__13134 ,w__13036);
  buf g__24(w__13133 ,w__13035);
  buf g__25(w__13132 ,w__13034);
  buf g__26(w__13131 ,w__13033);
  buf g__27(w__13130 ,w__13032);
  buf g__28(w__13129 ,w__13031);
  buf g__29(w__13128 ,w__13046);
  buf g__30(w__13127 ,w__13061);
  buf g__31(w__13126 ,w__13060);
  buf g__32(w__13125 ,w__13059);
  and g__33(w__13008 ,w__13181 ,w__13063);
  and g__34(w__13028 ,w__13129 ,w__13084);
  and g__35(w__13026 ,w__13131 ,w__13069);
  and g__36(w__13022 ,w__13135 ,w__13073);
  and g__37(w__13014 ,w__13143 ,w__13067);
  and g__38(w__12998 ,w__13127 ,w__13079);
  and g__39(w__13013 ,w__13128 ,w__13075);
  and g__40(w__13021 ,w__13136 ,w__13067);
  and g__41(w__13012 ,w__13145 ,w__13075);
  and g__42(w__13011 ,w__13146 ,w__13079);
  and g__43(w__13025 ,w__13132 ,w__13073);
  and g__44(w__13020 ,w__13137 ,w__13078);
  and g__45(w__13010 ,w__13147 ,w__13081);
  and g__46(w__13009 ,w__13148 ,w__13072);
  and g__47(w__13019 ,w__13138 ,w__13070);
  and g__48(w__13029 ,w__13144 ,w__13082);
  and g__49(w__13124 ,w__13126 ,w__13070);
  and g__50(w__13027 ,w__13130 ,w__13064);
  and g__51(w__13024 ,w__13133 ,w__13116);
  and g__52(w__13018 ,w__13139 ,w__13081);
  and g__53(w__13006 ,w__13184 ,w__13066);
  and g__54(w__13005 ,w__13183 ,w__13116);
  and g__55(w__13017 ,w__13140 ,w__13076);
  and g__56(w__13123 ,w__13185 ,w__13072);
  and g__57(w__13122 ,w__13186 ,w__13076);
  and g__58(w__13023 ,w__13134 ,w__13078);
  and g__59(w__13016 ,w__13141 ,w__13069);
  and g__60(w__13121 ,w__13188 ,w__13082);
  and g__61(w__13001 ,w__13187 ,w__13066);
  and g__62(w__13015 ,w__13142 ,w__13064);
  and g__63(w__13000 ,w__13125 ,w__13084);
  and g__64(w__13007 ,w__13182 ,w__13063);
  not g__65(w__13120 ,in22);
  not g__66(w__13119 ,in22);
  not g__67(w__13118 ,in22);
  not g__68(w__13117 ,in22);
  buf g__69(w__13004 ,w__13123);
  buf g__70(w__12999 ,w__13124);
  buf g__71(w__13003 ,w__13122);
  buf g__72(w__13002 ,w__13121);
  not g__73(w__13116 ,w__13083);
  not g__74(w__13084 ,w__13083);
  not g__75(w__13083 ,w__13120);
  not g__76(w__13082 ,w__13080);
  not g__77(w__13081 ,w__13080);
  not g__78(w__13080 ,w__13119);
  not g__79(w__13079 ,w__13077);
  not g__80(w__13078 ,w__13077);
  not g__81(w__13077 ,w__13119);
  not g__82(w__13076 ,w__13074);
  not g__83(w__13075 ,w__13074);
  not g__84(w__13074 ,w__13118);
  not g__85(w__13073 ,w__13071);
  not g__86(w__13072 ,w__13071);
  not g__87(w__13071 ,w__13118);
  not g__88(w__13070 ,w__13068);
  not g__89(w__13069 ,w__13068);
  not g__90(w__13068 ,w__13117);
  not g__91(w__13067 ,w__13065);
  not g__92(w__13066 ,w__13065);
  not g__93(w__13065 ,w__13117);
  not g__94(w__13064 ,w__13062);
  not g__95(w__13063 ,w__13062);
  not g__96(w__13062 ,w__13120);
  buf g__97(w__13328 ,w__13101);
  buf g__98(w__13327 ,w__13115);
  buf g__99(w__13326 ,w__13114);
  buf g__100(w__13325 ,w__13113);
  buf g__101(w__13324 ,w__13112);
  buf g__102(w__13323 ,w__13111);
  buf g__103(w__13322 ,w__13110);
  buf g__104(w__13321 ,w__13109);
  buf g__105(w__13320 ,w__13108);
  buf g__106(w__13319 ,w__13107);
  buf g__107(w__13318 ,w__13106);
  buf g__108(w__13317 ,w__13105);
  buf g__109(w__13316 ,w__13104);
  buf g__110(w__13315 ,w__13103);
  buf g__111(w__13314 ,w__13102);
  buf g__112(w__13313 ,w__13085);
  buf g__113(w__13312 ,w__13100);
  buf g__114(w__13311 ,w__13099);
  buf g__115(w__13310 ,w__13098);
  buf g__116(w__13309 ,w__13097);
  buf g__117(w__13276 ,w__13096);
  buf g__118(w__13275 ,w__13095);
  buf g__119(w__13274 ,w__13094);
  buf g__120(w__13273 ,w__13093);
  buf g__121(w__13272 ,w__13092);
  buf g__122(w__13271 ,w__13091);
  buf g__123(w__13270 ,w__13089);
  buf g__124(w__13269 ,w__13088);
  buf g__125(w__13268 ,w__13087);
  buf g__126(w__13267 ,w__13090);
  buf g__127(w__13266 ,w__13086);
  and g__128(w__12976 ,w__13318 ,w__13190);
  and g__129(w__13265 ,w__13266 ,w__13211);
  and g__130(w__13264 ,w__13269 ,w__13208);
  and g__131(w__13263 ,w__13272 ,w__13200);
  and g__132(w__13262 ,w__13312 ,w__13206);
  and g__133(w__12981 ,w__13328 ,w__13202);
  and g__134(w__13261 ,w__13273 ,w__13206);
  and g__135(w__12980 ,w__13314 ,w__13202);
  and g__136(w__13260 ,w__13315 ,w__13194);
  and g__137(w__12993 ,w__13270 ,w__13200);
  and g__138(w__13259 ,w__13274 ,w__13193);
  and g__139(w__12978 ,w__13316 ,w__13196);
  and g__140(w__12977 ,w__13317 ,w__13199);
  and g__141(w__13258 ,w__13275 ,w__13209);
  and g__142(w__12997 ,w__13313 ,w__13197);
  and g__143(w__13257 ,w__13327 ,w__13209);
  and g__144(w__12995 ,w__13268 ,w__13191);
  and g__145(w__12992 ,w__13267 ,w__13212);
  and g__146(w__13256 ,w__13276 ,w__13196);
  and g__147(w__12974 ,w__13320 ,w__13205);
  and g__148(w__12973 ,w__13321 ,w__13212);
  and g__149(w__13255 ,w__13309 ,w__13203);
  and g__150(w__13254 ,w__13322 ,w__13199);
  and g__151(w__13253 ,w__13323 ,w__13203);
  and g__152(w__13252 ,w__13271 ,w__13193);
  and g__153(w__13251 ,w__13310 ,w__13208);
  and g__154(w__13250 ,w__13324 ,w__13197);
  and g__155(w__12969 ,w__13325 ,w__13205);
  and g__156(w__13249 ,w__13311 ,w__13191);
  and g__157(w__13248 ,w__13326 ,w__13211);
  and g__158(w__12975 ,w__13319 ,w__13190);
  not g__159(w__13247 ,in22);
  not g__160(w__13246 ,in22);
  not g__161(w__13245 ,in22);
  not g__162(w__13244 ,in22);
  buf g__163(w__12989 ,w__13261);
  buf g__164(w__12994 ,w__13264);
  buf g__165(w__12990 ,w__13263);
  buf g__166(w__12986 ,w__13256);
  buf g__167(w__12984 ,w__13251);
  buf g__168(w__12991 ,w__13252);
  buf g__169(w__12987 ,w__13258);
  buf g__170(w__12983 ,w__13249);
  buf g__171(w__12985 ,w__13255);
  buf g__172(w__12982 ,w__13262);
  buf g__173(w__12996 ,w__13265);
  buf g__174(w__12979 ,w__13260);
  buf g__175(w__12988 ,w__13259);
  buf g__176(w__12968 ,w__13248);
  buf g__177(w__12967 ,w__13257);
  buf g__178(w__12972 ,w__13254);
  buf g__179(w__12970 ,w__13250);
  buf g__180(w__12971 ,w__13253);
  not g__181(w__13212 ,w__13210);
  not g__182(w__13211 ,w__13210);
  not g__183(w__13210 ,w__13247);
  not g__184(w__13209 ,w__13207);
  not g__185(w__13208 ,w__13207);
  not g__186(w__13207 ,w__13244);
  not g__187(w__13206 ,w__13204);
  not g__188(w__13205 ,w__13204);
  not g__189(w__13204 ,w__13244);
  not g__190(w__13203 ,w__13201);
  not g__191(w__13202 ,w__13201);
  not g__192(w__13201 ,w__13245);
  not g__193(w__13200 ,w__13198);
  not g__194(w__13199 ,w__13198);
  not g__195(w__13198 ,w__13245);
  not g__196(w__13197 ,w__13195);
  not g__197(w__13196 ,w__13195);
  not g__198(w__13195 ,w__13246);
  not g__199(w__13194 ,w__13192);
  not g__200(w__13193 ,w__13192);
  not g__201(w__13192 ,w__13246);
  not g__202(w__13191 ,w__13189);
  not g__203(w__13190 ,w__13189);
  not g__204(w__13189 ,w__13247);
  buf g__205(w__13459 ,w__13170);
  buf g__206(w__13458 ,w__13172);
  buf g__207(w__13457 ,w__13174);
  buf g__208(w__13456 ,w__13165);
  buf g__209(w__13455 ,w__13180);
  buf g__210(w__13454 ,w__13178);
  buf g__211(w__13453 ,w__13179);
  buf g__212(w__13452 ,w__13177);
  buf g__213(w__13451 ,w__13176);
  buf g__214(w__13450 ,w__13175);
  buf g__215(w__13449 ,w__13173);
  buf g__216(w__13448 ,w__13171);
  buf g__217(w__13447 ,w__13169);
  buf g__218(w__13446 ,w__13168);
  buf g__219(w__13445 ,w__13167);
  buf g__220(w__13444 ,w__13166);
  buf g__221(w__13443 ,w__13149);
  buf g__222(w__13442 ,w__13164);
  buf g__223(w__13441 ,w__13163);
  buf g__224(w__13440 ,w__13162);
  buf g__225(w__13439 ,w__13161);
  buf g__226(w__13438 ,w__13160);
  buf g__227(w__13437 ,w__13159);
  buf g__228(w__13436 ,w__13158);
  buf g__229(w__13403 ,w__13157);
  buf g__230(w__13402 ,w__13156);
  buf g__231(w__13401 ,w__13155);
  buf g__232(w__13400 ,w__13154);
  buf g__233(w__13399 ,w__13153);
  buf g__234(w__13398 ,w__13152);
  buf g__235(w__13397 ,w__13151);
  buf g__236(w__13396 ,w__13150);
  and g__237(w__12945 ,w__13459 ,w__13330);
  and g__238(w__12965 ,w__13396 ,w__13382);
  and g__239(w__12963 ,w__13398 ,w__13379);
  and g__240(w__12959 ,w__13402 ,w__13371);
  and g__241(w__13395 ,w__13442 ,w__13377);
  and g__242(w__13394 ,w__13455 ,w__13334);
  and g__243(w__12950 ,w__13456 ,w__13373);
  and g__244(w__12958 ,w__13403 ,w__13377);
  and g__245(w__12949 ,w__13444 ,w__13373);
  and g__246(w__13393 ,w__13445 ,w__13334);
  and g__247(w__12962 ,w__13399 ,w__13371);
  and g__248(w__12957 ,w__13436 ,w__13333);
  and g__249(w__12947 ,w__13446 ,w__13336);
  and g__250(w__12946 ,w__13447 ,w__13339);
  and g__251(w__12956 ,w__13437 ,w__13380);
  and g__252(w__12966 ,w__13443 ,w__13337);
  and g__253(w__13392 ,w__13453 ,w__13380);
  and g__254(w__12964 ,w__13397 ,w__13331);
  and g__255(w__12961 ,w__13400 ,w__13383);
  and g__256(w__12955 ,w__13438 ,w__13336);
  and g__257(w__12943 ,w__13458 ,w__13376);
  and g__258(w__12942 ,w__13449 ,w__13383);
  and g__259(w__12954 ,w__13439 ,w__13374);
  and g__260(w__13391 ,w__13457 ,w__13339);
  and g__261(w__13390 ,w__13450 ,w__13374);
  and g__262(w__12960 ,w__13401 ,w__13333);
  and g__263(w__12953 ,w__13440 ,w__13379);
  and g__264(w__12939 ,w__13451 ,w__13337);
  and g__265(w__12938 ,w__13452 ,w__13376);
  and g__266(w__13389 ,w__13441 ,w__13331);
  and g__267(w__13388 ,w__13454 ,w__13382);
  and g__268(w__12944 ,w__13448 ,w__13330);
  not g__269(w__13387 ,in18);
  not g__270(w__13386 ,in18);
  not g__271(w__13385 ,in18);
  not g__272(w__13384 ,in18);
  buf g__273(w__12952 ,w__13389);
  buf g__274(w__12935 ,w__13394);
  buf g__275(w__12941 ,w__13391);
  buf g__276(w__12951 ,w__13395);
  buf g__277(w__12948 ,w__13393);
  buf g__278(w__12936 ,w__13392);
  buf g__279(w__12940 ,w__13390);
  buf g__280(w__12937 ,w__13388);
  not g__281(w__13383 ,w__13381);
  not g__282(w__13382 ,w__13381);
  not g__283(w__13381 ,w__13387);
  not g__284(w__13380 ,w__13378);
  not g__285(w__13379 ,w__13378);
  not g__286(w__13378 ,w__13384);
  not g__287(w__13377 ,w__13375);
  not g__288(w__13376 ,w__13375);
  not g__289(w__13375 ,w__13384);
  not g__290(w__13374 ,w__13372);
  not g__291(w__13373 ,w__13372);
  not g__292(w__13372 ,w__13385);
  not g__293(w__13371 ,w__13338);
  not g__294(w__13339 ,w__13338);
  not g__295(w__13338 ,w__13385);
  not g__296(w__13337 ,w__13335);
  not g__297(w__13336 ,w__13335);
  not g__298(w__13335 ,w__13386);
  not g__299(w__13334 ,w__13332);
  not g__300(w__13333 ,w__13332);
  not g__301(w__13332 ,w__13386);
  not g__302(w__13331 ,w__13329);
  not g__303(w__13330 ,w__13329);
  not g__304(w__13329 ,w__13387);
  buf g__305(w__13631 ,w__13234);
  buf g__306(w__13630 ,w__13235);
  buf g__307(w__13629 ,w__13237);
  buf g__308(w__13628 ,w__13239);
  buf g__309(w__13627 ,w__13238);
  buf g__310(w__13626 ,w__13241);
  buf g__311(w__13594 ,w__13240);
  buf g__312(w__13593 ,w__13229);
  buf g__313(w__13592 ,w__13243);
  buf g__314(w__13591 ,w__13242);
  buf g__315(w__13590 ,w__13236);
  buf g__316(w__13589 ,w__13233);
  buf g__317(w__13588 ,w__13232);
  buf g__318(w__13587 ,w__13231);
  buf g__319(w__13586 ,w__13230);
  buf g__320(w__13585 ,w__13213);
  buf g__321(w__13584 ,w__13228);
  buf g__322(w__13583 ,w__13227);
  buf g__323(w__13582 ,w__13226);
  buf g__324(w__13581 ,w__13225);
  buf g__325(w__13580 ,w__13224);
  buf g__326(w__13579 ,w__13223);
  buf g__327(w__13578 ,w__13222);
  buf g__328(w__13577 ,w__13221);
  buf g__329(w__13576 ,w__13220);
  buf g__330(w__13575 ,w__13219);
  buf g__331(w__13574 ,w__13218);
  buf g__332(w__13573 ,w__13217);
  buf g__333(w__13572 ,w__13216);
  buf g__334(w__13571 ,w__13215);
  buf g__335(w__13570 ,w__13214);
  and g__336(w__13569 ,w__13631 ,w__13461);
  and g__337(w__12933 ,w__13570 ,w__13513);
  and g__338(w__12931 ,w__13572 ,w__13510);
  and g__339(w__12927 ,w__13576 ,w__13502);
  and g__340(w__12919 ,w__13584 ,w__13508);
  and g__341(w__13568 ,w__13593 ,w__13504);
  and g__342(w__12926 ,w__13577 ,w__13508);
  and g__343(w__13567 ,w__13586 ,w__13504);
  and g__344(w__13566 ,w__13587 ,w__13465);
  and g__345(w__13565 ,w__13573 ,w__13502);
  and g__346(w__12925 ,w__13578 ,w__13464);
  and g__347(w__13564 ,w__13588 ,w__13467);
  and g__348(w__13531 ,w__13589 ,w__13501);
  and g__349(w__12924 ,w__13579 ,w__13511);
  and g__350(w__12934 ,w__13585 ,w__13499);
  and g__351(w__13530 ,w__13592 ,w__13511);
  and g__352(w__13529 ,w__13571 ,w__13462);
  and g__353(w__13528 ,w__13574 ,w__13514);
  and g__354(w__12923 ,w__13580 ,w__13467);
  and g__355(w__13527 ,w__13590 ,w__13507);
  and g__356(w__13526 ,w__13629 ,w__13514);
  and g__357(w__12922 ,w__13581 ,w__13505);
  and g__358(w__13525 ,w__13627 ,w__13501);
  and g__359(w__13524 ,w__13628 ,w__13505);
  and g__360(w__12928 ,w__13575 ,w__13464);
  and g__361(w__13523 ,w__13582 ,w__13510);
  and g__362(w__13522 ,w__13594 ,w__13499);
  and g__363(w__13521 ,w__13626 ,w__13507);
  and g__364(w__12920 ,w__13583 ,w__13462);
  and g__365(w__13520 ,w__13591 ,w__13513);
  and g__366(w__13519 ,w__13630 ,w__13461);
  not g__367(w__13518 ,in18);
  not g__368(w__13517 ,in18);
  not g__369(w__13516 ,in18);
  not g__370(w__13515 ,in18);
  buf g__371(w__12907 ,w__13522);
  buf g__372(w__12921 ,w__13523);
  buf g__373(w__12912 ,w__13519);
  buf g__374(w__12913 ,w__13569);
  buf g__375(w__12909 ,w__13525);
  buf g__376(w__12910 ,w__13526);
  buf g__377(w__12908 ,w__13524);
  buf g__378(w__12905 ,w__13520);
  buf g__379(w__12932 ,w__13529);
  buf g__380(w__12904 ,w__13530);
  buf g__381(w__12930 ,w__13565);
  buf g__382(w__12929 ,w__13528);
  buf g__383(w__12917 ,w__13567);
  buf g__384(w__12916 ,w__13566);
  buf g__385(w__12906 ,w__13521);
  buf g__386(w__12918 ,w__13568);
  buf g__387(w__12911 ,w__13527);
  buf g__388(w__12914 ,w__13531);
  buf g__389(w__12915 ,w__13564);
  not g__390(w__13514 ,w__13512);
  not g__391(w__13513 ,w__13512);
  not g__392(w__13512 ,w__13518);
  not g__393(w__13511 ,w__13509);
  not g__394(w__13510 ,w__13509);
  not g__395(w__13509 ,w__13515);
  not g__396(w__13508 ,w__13506);
  not g__397(w__13507 ,w__13506);
  not g__398(w__13506 ,w__13515);
  not g__399(w__13505 ,w__13503);
  not g__400(w__13504 ,w__13503);
  not g__401(w__13503 ,w__13516);
  not g__402(w__13502 ,w__13500);
  not g__403(w__13501 ,w__13500);
  not g__404(w__13500 ,w__13516);
  not g__405(w__13499 ,w__13466);
  not g__406(w__13467 ,w__13466);
  not g__407(w__13466 ,w__13517);
  not g__408(w__13465 ,w__13463);
  not g__409(w__13464 ,w__13463);
  not g__410(w__13463 ,w__13517);
  not g__411(w__13462 ,w__13460);
  not g__412(w__13461 ,w__13460);
  not g__413(w__13460 ,w__13518);
  buf g__414(w__13782 ,w__13293);
  buf g__415(w__13781 ,w__13308);
  buf g__416(w__13780 ,w__13307);
  buf g__417(w__13779 ,w__13306);
  buf g__418(w__13778 ,w__13305);
  buf g__419(w__13777 ,w__13304);
  buf g__420(w__13776 ,w__13303);
  buf g__421(w__13775 ,w__13302);
  buf g__422(w__13774 ,w__13301);
  buf g__423(w__13773 ,w__13300);
  buf g__424(w__13772 ,w__13299);
  buf g__425(w__13771 ,w__13298);
  buf g__426(w__13770 ,w__13297);
  buf g__427(w__13769 ,w__13296);
  buf g__428(w__13768 ,w__13295);
  buf g__429(w__13767 ,w__13294);
  buf g__430(w__13766 ,w__13277);
  buf g__431(w__13765 ,w__13292);
  buf g__432(w__13764 ,w__13291);
  buf g__433(w__13763 ,w__13290);
  buf g__434(w__13762 ,w__13289);
  buf g__435(w__13761 ,w__13288);
  buf g__436(w__13760 ,w__13287);
  buf g__437(w__13759 ,w__13286);
  buf g__438(w__13758 ,w__13285);
  buf g__439(w__13757 ,w__13284);
  buf g__440(w__13756 ,w__13283);
  buf g__441(w__13755 ,w__13282);
  buf g__442(w__13754 ,w__13281);
  buf g__443(w__13722 ,w__13280);
  buf g__444(w__13721 ,w__13279);
  buf g__445(w__13720 ,w__13278);
  and g__446(w__13719 ,w__13771 ,w__13633);
  and g__447(w__13718 ,w__13720 ,w__13654);
  and g__448(w__13717 ,w__13722 ,w__13639);
  and g__449(w__13716 ,w__13757 ,w__13649);
  and g__450(w__13715 ,w__13765 ,w__13637);
  and g__451(w__12872 ,w__13781 ,w__13643);
  and g__452(w__13714 ,w__13782 ,w__13651);
  and g__453(w__13713 ,w__13758 ,w__13637);
  and g__454(w__13712 ,w__13767 ,w__13651);
  and g__455(w__12885 ,w__13768 ,w__13643);
  and g__456(w__13711 ,w__13754 ,w__13649);
  and g__457(w__13710 ,w__13759 ,w__13642);
  and g__458(w__13709 ,w__13769 ,w__13645);
  and g__459(w__13708 ,w__13770 ,w__13648);
  and g__460(w__13707 ,w__13760 ,w__13640);
  and g__461(w__12903 ,w__13766 ,w__13646);
  and g__462(w__13706 ,w__13780 ,w__13640);
  and g__463(w__13705 ,w__13721 ,w__13634);
  and g__464(w__13704 ,w__13755 ,w__13655);
  and g__465(w__13703 ,w__13761 ,w__13645);
  and g__466(w__13702 ,w__13773 ,w__13636);
  and g__467(w__13701 ,w__13774 ,w__13655);
  and g__468(w__13700 ,w__13762 ,w__13652);
  and g__469(w__13699 ,w__13775 ,w__13648);
  and g__470(w__13698 ,w__13776 ,w__13652);
  and g__471(w__13697 ,w__13756 ,w__13642);
  and g__472(w__13696 ,w__13763 ,w__13639);
  and g__473(w__13695 ,w__13777 ,w__13646);
  and g__474(w__13694 ,w__13778 ,w__13636);
  and g__475(w__13693 ,w__13764 ,w__13634);
  and g__476(w__12874 ,w__13779 ,w__13654);
  and g__477(w__13692 ,w__13772 ,w__13633);
  not g__478(w__13691 ,in14);
  not g__479(w__13658 ,in14);
  not g__480(w__13657 ,in14);
  not g__481(w__13656 ,in14);
  buf g__482(w__12879 ,w__13701);
  buf g__483(w__12883 ,w__13708);
  buf g__484(w__12881 ,w__13692);
  buf g__485(w__12899 ,w__13711);
  buf g__486(w__12882 ,w__13719);
  buf g__487(w__12886 ,w__13712);
  buf g__488(w__12880 ,w__13702);
  buf g__489(w__12878 ,w__13699);
  buf g__490(w__12877 ,w__13698);
  buf g__491(w__12887 ,w__13714);
  buf g__492(w__12875 ,w__13694);
  buf g__493(w__12876 ,w__13695);
  buf g__494(w__12893 ,w__13707);
  buf g__495(w__12898 ,w__13704);
  buf g__496(w__12900 ,w__13717);
  buf g__497(w__12896 ,w__13716);
  buf g__498(w__12884 ,w__13709);
  buf g__499(w__12901 ,w__13705);
  buf g__500(w__12897 ,w__13697);
  buf g__501(w__12888 ,w__13715);
  buf g__502(w__12902 ,w__13718);
  buf g__503(w__12890 ,w__13696);
  buf g__504(w__12892 ,w__13703);
  buf g__505(w__12894 ,w__13710);
  buf g__506(w__12889 ,w__13693);
  buf g__507(w__12873 ,w__13706);
  buf g__508(w__12891 ,w__13700);
  buf g__509(w__12895 ,w__13713);
  not g__510(w__13655 ,w__13653);
  not g__511(w__13654 ,w__13653);
  not g__512(w__13653 ,w__13691);
  not g__513(w__13652 ,w__13650);
  not g__514(w__13651 ,w__13650);
  not g__515(w__13650 ,w__13657);
  not g__516(w__13649 ,w__13647);
  not g__517(w__13648 ,w__13647);
  not g__518(w__13647 ,w__13657);
  not g__519(w__13646 ,w__13644);
  not g__520(w__13645 ,w__13644);
  not g__521(w__13644 ,w__13658);
  not g__522(w__13643 ,w__13641);
  not g__523(w__13642 ,w__13641);
  not g__524(w__13641 ,w__13658);
  not g__525(w__13640 ,w__13638);
  not g__526(w__13639 ,w__13638);
  not g__527(w__13638 ,w__13656);
  not g__528(w__13637 ,w__13635);
  not g__529(w__13636 ,w__13635);
  not g__530(w__13635 ,w__13656);
  not g__531(w__13634 ,w__13632);
  not g__532(w__13633 ,w__13632);
  not g__533(w__13632 ,w__13691);
  buf g__534(w__13865 ,w__13341);
  buf g__535(w__13864 ,w__13356);
  buf g__536(w__13863 ,w__13370);
  buf g__537(w__13862 ,w__13369);
  buf g__538(w__13861 ,w__13368);
  buf g__539(w__13860 ,w__13367);
  buf g__540(w__13859 ,w__13366);
  buf g__541(w__13858 ,w__13365);
  buf g__542(w__13857 ,w__13364);
  buf g__543(w__13856 ,w__13363);
  buf g__544(w__13855 ,w__13362);
  buf g__545(w__13854 ,w__13361);
  buf g__546(w__13853 ,w__13360);
  buf g__547(w__13852 ,w__13359);
  buf g__548(w__13851 ,w__13358);
  buf g__549(w__13850 ,w__13357);
  buf g__550(w__13849 ,w__13340);
  buf g__551(w__13848 ,w__13355);
  buf g__552(w__13847 ,w__13354);
  buf g__553(w__13846 ,w__13353);
  buf g__554(w__13845 ,w__13352);
  buf g__555(w__13844 ,w__13351);
  buf g__556(w__13843 ,w__13350);
  buf g__557(w__13842 ,w__13349);
  buf g__558(w__13841 ,w__13348);
  buf g__559(w__13840 ,w__13347);
  buf g__560(w__13839 ,w__13346);
  buf g__561(w__13838 ,w__13345);
  buf g__562(w__13837 ,w__13344);
  buf g__563(w__13836 ,w__13343);
  buf g__564(w__13835 ,w__13342);
  and g__565(w__13834 ,w__13854 ,w__13784);
  and g__566(w__13833 ,w__13865 ,w__13805);
  and g__567(w__13832 ,w__13836 ,w__13802);
  and g__568(w__13831 ,w__13840 ,w__13794);
  and g__569(w__13830 ,w__13848 ,w__13800);
  and g__570(w__13829 ,w__13864 ,w__13796);
  and g__571(w__13828 ,w__13841 ,w__13800);
  and g__572(w__13827 ,w__13850 ,w__13796);
  and g__573(w__13826 ,w__13851 ,w__13788);
  and g__574(w__12867 ,w__13837 ,w__13794);
  and g__575(w__13825 ,w__13842 ,w__13787);
  and g__576(w__13824 ,w__13852 ,w__13790);
  and g__577(w__13823 ,w__13853 ,w__13793);
  and g__578(w__13822 ,w__13843 ,w__13803);
  and g__579(w__12871 ,w__13849 ,w__13791);
  and g__580(w__13821 ,w__13863 ,w__13803);
  and g__581(w__12869 ,w__13835 ,w__13785);
  and g__582(w__12866 ,w__13838 ,w__13806);
  and g__583(w__13820 ,w__13844 ,w__13790);
  and g__584(w__13819 ,w__13856 ,w__13799);
  and g__585(w__13818 ,w__13857 ,w__13806);
  and g__586(w__13817 ,w__13845 ,w__13797);
  and g__587(w__12846 ,w__13858 ,w__13793);
  and g__588(w__12845 ,w__13859 ,w__13797);
  and g__589(w__13816 ,w__13839 ,w__13787);
  and g__590(w__13815 ,w__13846 ,w__13802);
  and g__591(w__13814 ,w__13860 ,w__13791);
  and g__592(w__13813 ,w__13861 ,w__13799);
  and g__593(w__13812 ,w__13847 ,w__13785);
  and g__594(w__12842 ,w__13862 ,w__13805);
  and g__595(w__13811 ,w__13855 ,w__13784);
  not g__596(w__13810 ,in14);
  not g__597(w__13809 ,in14);
  not g__598(w__13808 ,in14);
  not g__599(w__13807 ,in14);
  buf g__600(w__12858 ,w__13815);
  buf g__601(w__12859 ,w__13817);
  buf g__602(w__12847 ,w__13818);
  buf g__603(w__12850 ,w__13834);
  buf g__604(w__12844 ,w__13814);
  buf g__605(w__12849 ,w__13811);
  buf g__606(w__12865 ,w__13816);
  buf g__607(w__12853 ,w__13826);
  buf g__608(w__12854 ,w__13827);
  buf g__609(w__12848 ,w__13819);
  buf g__610(w__12860 ,w__13820);
  buf g__611(w__12863 ,w__13828);
  buf g__612(w__12861 ,w__13822);
  buf g__613(w__12856 ,w__13830);
  buf g__614(w__12852 ,w__13824);
  buf g__615(w__12862 ,w__13825);
  buf g__616(w__12870 ,w__13833);
  buf g__617(w__12855 ,w__13829);
  buf g__618(w__12841 ,w__13821);
  buf g__619(w__12868 ,w__13832);
  buf g__620(w__12857 ,w__13812);
  buf g__621(w__12864 ,w__13831);
  buf g__622(w__12851 ,w__13823);
  buf g__623(w__12843 ,w__13813);
  not g__624(w__13806 ,w__13804);
  not g__625(w__13805 ,w__13804);
  not g__626(w__13804 ,w__13810);
  not g__627(w__13803 ,w__13801);
  not g__628(w__13802 ,w__13801);
  not g__629(w__13801 ,w__13807);
  not g__630(w__13800 ,w__13798);
  not g__631(w__13799 ,w__13798);
  not g__632(w__13798 ,w__13807);
  not g__633(w__13797 ,w__13795);
  not g__634(w__13796 ,w__13795);
  not g__635(w__13795 ,w__13808);
  not g__636(w__13794 ,w__13792);
  not g__637(w__13793 ,w__13792);
  not g__638(w__13792 ,w__13808);
  not g__639(w__13791 ,w__13789);
  not g__640(w__13790 ,w__13789);
  not g__641(w__13789 ,w__13809);
  not g__642(w__13788 ,w__13786);
  not g__643(w__13787 ,w__13786);
  not g__644(w__13786 ,w__13809);
  not g__645(w__13785 ,w__13783);
  not g__646(w__13784 ,w__13783);
  not g__647(w__13783 ,w__13810);
  buf g__648(w__13954 ,w__13420);
  buf g__649(w__13953 ,w__13435);
  buf g__650(w__13952 ,w__13434);
  buf g__651(w__13951 ,w__13433);
  buf g__652(w__13950 ,w__13432);
  buf g__653(w__13949 ,w__13431);
  buf g__654(w__13948 ,w__13430);
  buf g__655(w__13947 ,w__13429);
  buf g__656(w__13946 ,w__13428);
  buf g__657(w__13945 ,w__13427);
  buf g__658(w__13944 ,w__13426);
  buf g__659(w__13943 ,w__13425);
  buf g__660(w__13942 ,w__13424);
  buf g__661(w__13941 ,w__13423);
  buf g__662(w__13940 ,w__13422);
  buf g__663(w__13939 ,w__13421);
  buf g__664(w__13938 ,w__13404);
  buf g__665(w__13937 ,w__13419);
  buf g__666(w__13936 ,w__13418);
  buf g__667(w__13935 ,w__13417);
  buf g__668(w__13934 ,w__13416);
  buf g__669(w__13933 ,w__13415);
  buf g__670(w__13932 ,w__13414);
  buf g__671(w__13931 ,w__13413);
  buf g__672(w__13930 ,w__13412);
  buf g__673(w__13929 ,w__13411);
  buf g__674(w__13928 ,w__13410);
  buf g__675(w__13927 ,w__13409);
  buf g__676(w__13926 ,w__13408);
  buf g__677(w__13925 ,w__13407);
  buf g__678(w__13924 ,w__13406);
  buf g__679(w__13923 ,w__13405);
  and g__680(w__13922 ,w__13943 ,w__13867);
  and g__681(w__13921 ,w__13923 ,w__13888);
  and g__682(w__13920 ,w__13925 ,w__13879);
  and g__683(w__13919 ,w__13929 ,w__13871);
  and g__684(w__13918 ,w__13937 ,w__13877);
  and g__685(w__13917 ,w__13953 ,w__13883);
  and g__686(w__13916 ,w__13954 ,w__13873);
  and g__687(w__13915 ,w__13930 ,w__13877);
  and g__688(w__13914 ,w__13939 ,w__13873);
  and g__689(w__13913 ,w__13940 ,w__13883);
  and g__690(w__13912 ,w__13926 ,w__13871);
  and g__691(w__13911 ,w__13931 ,w__13882);
  and g__692(w__13910 ,w__13941 ,w__13885);
  and g__693(w__13909 ,w__13942 ,w__13870);
  and g__694(w__13908 ,w__13932 ,w__13880);
  and g__695(w__12840 ,w__13938 ,w__13886);
  and g__696(w__13907 ,w__13952 ,w__13880);
  and g__697(w__13906 ,w__13924 ,w__13868);
  and g__698(w__13905 ,w__13927 ,w__13889);
  and g__699(w__13904 ,w__13933 ,w__13885);
  and g__700(w__13903 ,w__13945 ,w__13876);
  and g__701(w__13902 ,w__13946 ,w__13889);
  and g__702(w__13901 ,w__13934 ,w__13874);
  and g__703(w__12815 ,w__13947 ,w__13870);
  and g__704(w__12814 ,w__13948 ,w__13874);
  and g__705(w__13900 ,w__13928 ,w__13882);
  and g__706(w__13899 ,w__13935 ,w__13879);
  and g__707(w__13898 ,w__13949 ,w__13886);
  and g__708(w__13897 ,w__13950 ,w__13876);
  and g__709(w__13896 ,w__13936 ,w__13868);
  and g__710(w__13895 ,w__13951 ,w__13888);
  and g__711(w__13894 ,w__13944 ,w__13867);
  not g__712(w__13893 ,in10);
  not g__713(w__13892 ,in10);
  not g__714(w__13891 ,in10);
  not g__715(w__13890 ,in10);
  buf g__716(w__12813 ,w__13898);
  buf g__717(w__12809 ,w__13917);
  buf g__718(w__12830 ,w__13908);
  buf g__719(w__12826 ,w__13896);
  buf g__720(w__12812 ,w__13897);
  buf g__721(w__12831 ,w__13911);
  buf g__722(w__12810 ,w__13907);
  buf g__723(w__12834 ,w__13900);
  buf g__724(w__12828 ,w__13901);
  buf g__725(w__12816 ,w__13902);
  buf g__726(w__12817 ,w__13903);
  buf g__727(w__12829 ,w__13904);
  buf g__728(w__12835 ,w__13905);
  buf g__729(w__12838 ,w__13906);
  buf g__730(w__12832 ,w__13915);
  buf g__731(w__12824 ,w__13916);
  buf g__732(w__12820 ,w__13909);
  buf g__733(w__12821 ,w__13910);
  buf g__734(w__12827 ,w__13899);
  buf g__735(w__12836 ,w__13912);
  buf g__736(w__12822 ,w__13913);
  buf g__737(w__12823 ,w__13914);
  buf g__738(w__12839 ,w__13921);
  buf g__739(w__12818 ,w__13894);
  buf g__740(w__12837 ,w__13920);
  buf g__741(w__12825 ,w__13918);
  buf g__742(w__12833 ,w__13919);
  buf g__743(w__12819 ,w__13922);
  buf g__744(w__12811 ,w__13895);
  not g__745(w__13889 ,w__13887);
  not g__746(w__13888 ,w__13887);
  not g__747(w__13887 ,w__13893);
  not g__748(w__13886 ,w__13884);
  not g__749(w__13885 ,w__13884);
  not g__750(w__13884 ,w__13892);
  not g__751(w__13883 ,w__13881);
  not g__752(w__13882 ,w__13881);
  not g__753(w__13881 ,w__13892);
  not g__754(w__13880 ,w__13878);
  not g__755(w__13879 ,w__13878);
  not g__756(w__13878 ,w__13890);
  not g__757(w__13877 ,w__13875);
  not g__758(w__13876 ,w__13875);
  not g__759(w__13875 ,w__13890);
  not g__760(w__13874 ,w__13872);
  not g__761(w__13873 ,w__13872);
  not g__762(w__13872 ,w__13891);
  not g__763(w__13871 ,w__13869);
  not g__764(w__13870 ,w__13869);
  not g__765(w__13869 ,w__13891);
  not g__766(w__13868 ,w__13866);
  not g__767(w__13867 ,w__13866);
  not g__768(w__13866 ,w__13893);
  buf g__769(w__14033 ,w__13484);
  buf g__770(w__14032 ,w__13498);
  buf g__771(w__14031 ,w__13497);
  buf g__772(w__14030 ,w__13496);
  buf g__773(w__14029 ,w__13495);
  buf g__774(w__14028 ,w__13494);
  buf g__775(w__14027 ,w__13493);
  buf g__776(w__14026 ,w__13492);
  buf g__777(w__14025 ,w__13491);
  buf g__778(w__14024 ,w__13490);
  buf g__779(w__14023 ,w__13489);
  buf g__780(w__14022 ,w__13488);
  buf g__781(w__14021 ,w__13487);
  buf g__782(w__14020 ,w__13486);
  buf g__783(w__14019 ,w__13485);
  buf g__784(w__14018 ,w__13468);
  buf g__785(w__14017 ,w__13483);
  buf g__786(w__14016 ,w__13482);
  buf g__787(w__14015 ,w__13481);
  buf g__788(w__14014 ,w__13480);
  buf g__789(w__14013 ,w__13479);
  buf g__790(w__14012 ,w__13478);
  buf g__791(w__14011 ,w__13477);
  buf g__792(w__14010 ,w__13476);
  buf g__793(w__14009 ,w__13475);
  buf g__794(w__14008 ,w__13474);
  buf g__795(w__14007 ,w__13473);
  buf g__796(w__14006 ,w__13472);
  buf g__797(w__14005 ,w__13471);
  buf g__798(w__14004 ,w__13470);
  buf g__799(w__14003 ,w__13469);
  and g__800(w__14002 ,w__14023 ,w__13956);
  and g__801(w__12807 ,w__14003 ,w__13977);
  and g__802(w__12805 ,w__14005 ,w__13974);
  and g__803(w__12801 ,w__14009 ,w__13966);
  and g__804(w__14001 ,w__14017 ,w__13972);
  and g__805(w__14000 ,w__14033 ,w__13968);
  and g__806(w__13999 ,w__14010 ,w__13972);
  and g__807(w__13998 ,w__14019 ,w__13968);
  and g__808(w__13997 ,w__14020 ,w__13960);
  and g__809(w__13996 ,w__14006 ,w__13966);
  and g__810(w__13995 ,w__14011 ,w__13959);
  and g__811(w__13994 ,w__14021 ,w__13962);
  and g__812(w__13993 ,w__14022 ,w__13965);
  and g__813(w__13992 ,w__14012 ,w__13975);
  and g__814(w__12808 ,w__14018 ,w__13963);
  and g__815(w__13991 ,w__14032 ,w__13975);
  and g__816(w__13990 ,w__14004 ,w__13957);
  and g__817(w__13989 ,w__14007 ,w__13978);
  and g__818(w__12797 ,w__14013 ,w__13962);
  and g__819(w__13988 ,w__14025 ,w__13971);
  and g__820(w__13987 ,w__14026 ,w__13978);
  and g__821(w__12796 ,w__14014 ,w__13969);
  and g__822(w__12783 ,w__14027 ,w__13965);
  and g__823(w__12782 ,w__14028 ,w__13969);
  and g__824(w__12802 ,w__14008 ,w__13959);
  and g__825(w__12795 ,w__14015 ,w__13974);
  and g__826(w__12781 ,w__14029 ,w__13963);
  and g__827(w__13986 ,w__14030 ,w__13971);
  and g__828(w__13985 ,w__14016 ,w__13957);
  and g__829(w__13984 ,w__14031 ,w__13977);
  and g__830(w__13983 ,w__14024 ,w__13956);
  not g__831(w__13982 ,in10);
  not g__832(w__13981 ,in10);
  not g__833(w__13980 ,in10);
  not g__834(w__13979 ,in10);
  buf g__835(w__12786 ,w__13983);
  buf g__836(w__12780 ,w__13986);
  buf g__837(w__12779 ,w__13984);
  buf g__838(w__12794 ,w__13985);
  buf g__839(w__12799 ,w__13995);
  buf g__840(w__12784 ,w__13987);
  buf g__841(w__12785 ,w__13988);
  buf g__842(w__12803 ,w__13989);
  buf g__843(w__12806 ,w__13990);
  buf g__844(w__12790 ,w__13997);
  buf g__845(w__12778 ,w__13991);
  buf g__846(w__12791 ,w__13998);
  buf g__847(w__12793 ,w__14001);
  buf g__848(w__12800 ,w__13999);
  buf g__849(w__12804 ,w__13996);
  buf g__850(w__12792 ,w__14000);
  buf g__851(w__12788 ,w__13993);
  buf g__852(w__12787 ,w__14002);
  buf g__853(w__12798 ,w__13992);
  buf g__854(w__12789 ,w__13994);
  not g__855(w__13978 ,w__13976);
  not g__856(w__13977 ,w__13976);
  not g__857(w__13976 ,w__13982);
  not g__858(w__13975 ,w__13973);
  not g__859(w__13974 ,w__13973);
  not g__860(w__13973 ,w__13979);
  not g__861(w__13972 ,w__13970);
  not g__862(w__13971 ,w__13970);
  not g__863(w__13970 ,w__13979);
  not g__864(w__13969 ,w__13967);
  not g__865(w__13968 ,w__13967);
  not g__866(w__13967 ,w__13980);
  not g__867(w__13966 ,w__13964);
  not g__868(w__13965 ,w__13964);
  not g__869(w__13964 ,w__13980);
  not g__870(w__13963 ,w__13961);
  not g__871(w__13962 ,w__13961);
  not g__872(w__13961 ,w__13981);
  not g__873(w__13960 ,w__13958);
  not g__874(w__13959 ,w__13958);
  not g__875(w__13958 ,w__13981);
  not g__876(w__13957 ,w__13955);
  not g__877(w__13956 ,w__13955);
  not g__878(w__13955 ,w__13982);
  buf g__879(w__14113 ,w__13548);
  buf g__880(w__14112 ,w__13563);
  buf g__881(w__14111 ,w__13562);
  buf g__882(w__14110 ,w__13561);
  buf g__883(w__14109 ,w__13560);
  buf g__884(w__14108 ,w__13559);
  buf g__885(w__14107 ,w__13558);
  buf g__886(w__14106 ,w__13557);
  buf g__887(w__14105 ,w__13556);
  buf g__888(w__14104 ,w__13555);
  buf g__889(w__14103 ,w__13554);
  buf g__890(w__14102 ,w__13553);
  buf g__891(w__14101 ,w__13552);
  buf g__892(w__14100 ,w__13551);
  buf g__893(w__14099 ,w__13550);
  buf g__894(w__14098 ,w__13549);
  buf g__895(w__14097 ,w__13532);
  buf g__896(w__14096 ,w__13547);
  buf g__897(w__14095 ,w__13546);
  buf g__898(w__14094 ,w__13545);
  buf g__899(w__14093 ,w__13544);
  buf g__900(w__14092 ,w__13543);
  buf g__901(w__14091 ,w__13542);
  buf g__902(w__14090 ,w__13541);
  buf g__903(w__14089 ,w__13540);
  buf g__904(w__14088 ,w__13539);
  buf g__905(w__14087 ,w__13538);
  buf g__906(w__14086 ,w__13537);
  buf g__907(w__14085 ,w__13534);
  buf g__908(w__14084 ,w__13533);
  buf g__909(w__14083 ,w__13536);
  buf g__910(w__14082 ,w__13535);
  and g__911(w__14081 ,w__14102 ,w__14035);
  and g__912(w__14080 ,w__14084 ,w__14056);
  and g__913(w__12774 ,w__14082 ,w__14053);
  and g__914(w__12770 ,w__14088 ,w__14045);
  and g__915(w__14079 ,w__14096 ,w__14051);
  and g__916(w__14078 ,w__14112 ,w__14039);
  and g__917(w__14077 ,w__14113 ,w__14047);
  and g__918(w__14076 ,w__14089 ,w__14051);
  and g__919(w__14075 ,w__14098 ,w__14047);
  and g__920(w__14074 ,w__14099 ,w__14039);
  and g__921(w__12773 ,w__14083 ,w__14045);
  and g__922(w__14073 ,w__14090 ,w__14038);
  and g__923(w__14072 ,w__14100 ,w__14041);
  and g__924(w__14071 ,w__14101 ,w__14044);
  and g__925(w__14070 ,w__14091 ,w__14054);
  and g__926(w__12777 ,w__14097 ,w__14042);
  and g__927(w__12747 ,w__14111 ,w__14054);
  and g__928(w__12775 ,w__14085 ,w__14036);
  and g__929(w__12772 ,w__14086 ,w__14057);
  and g__930(w__12766 ,w__14092 ,w__14041);
  and g__931(w__14069 ,w__14104 ,w__14050);
  and g__932(w__14068 ,w__14105 ,w__14057);
  and g__933(w__12765 ,w__14093 ,w__14048);
  and g__934(w__14067 ,w__14106 ,w__14044);
  and g__935(w__14066 ,w__14107 ,w__14048);
  and g__936(w__12771 ,w__14087 ,w__14038);
  and g__937(w__12764 ,w__14094 ,w__14053);
  and g__938(w__12750 ,w__14108 ,w__14042);
  and g__939(w__14065 ,w__14109 ,w__14050);
  and g__940(w__14064 ,w__14095 ,w__14036);
  and g__941(w__14063 ,w__14110 ,w__14056);
  and g__942(w__14062 ,w__14103 ,w__14035);
  not g__943(w__14061 ,in3);
  not g__944(w__14060 ,in3);
  not g__945(w__14059 ,in3);
  not g__946(w__14058 ,in3);
  buf g__947(w__12760 ,w__14075);
  buf g__948(w__12759 ,w__14074);
  buf g__949(w__12753 ,w__14068);
  buf g__950(w__12769 ,w__14076);
  buf g__951(w__12752 ,w__14067);
  buf g__952(w__12761 ,w__14077);
  buf g__953(w__12748 ,w__14063);
  buf g__954(w__12756 ,w__14081);
  buf g__955(w__12754 ,w__14069);
  buf g__956(w__12751 ,w__14066);
  buf g__957(w__12767 ,w__14070);
  buf g__958(w__12758 ,w__14072);
  buf g__959(w__12749 ,w__14065);
  buf g__960(w__12768 ,w__14073);
  buf g__961(w__12763 ,w__14064);
  buf g__962(w__12762 ,w__14079);
  buf g__963(w__12755 ,w__14062);
  buf g__964(w__12757 ,w__14071);
  buf g__965(w__12776 ,w__14080);
  buf g__966(w__12746 ,w__14078);
  not g__967(w__14057 ,w__14055);
  not g__968(w__14056 ,w__14055);
  not g__969(w__14055 ,w__14061);
  not g__970(w__14054 ,w__14052);
  not g__971(w__14053 ,w__14052);
  not g__972(w__14052 ,w__14058);
  not g__973(w__14051 ,w__14049);
  not g__974(w__14050 ,w__14049);
  not g__975(w__14049 ,w__14058);
  not g__976(w__14048 ,w__14046);
  not g__977(w__14047 ,w__14046);
  not g__978(w__14046 ,w__14059);
  not g__979(w__14045 ,w__14043);
  not g__980(w__14044 ,w__14043);
  not g__981(w__14043 ,w__14059);
  not g__982(w__14042 ,w__14040);
  not g__983(w__14041 ,w__14040);
  not g__984(w__14040 ,w__14060);
  not g__985(w__14039 ,w__14037);
  not g__986(w__14038 ,w__14037);
  not g__987(w__14037 ,w__14060);
  not g__988(w__14036 ,w__14034);
  not g__989(w__14035 ,w__14034);
  not g__990(w__14034 ,w__14061);
  buf g__991(w__14193 ,w__13596);
  buf g__992(w__14192 ,w__13611);
  buf g__993(w__14191 ,w__13625);
  buf g__994(w__14190 ,w__13624);
  buf g__995(w__14189 ,w__13623);
  buf g__996(w__14188 ,w__13622);
  buf g__997(w__14187 ,w__13621);
  buf g__998(w__14186 ,w__13620);
  buf g__999(w__14185 ,w__13619);
  buf g__1000(w__14184 ,w__13618);
  buf g__1001(w__14183 ,w__13617);
  buf g__1002(w__14182 ,w__13616);
  buf g__1003(w__14181 ,w__13615);
  buf g__1004(w__14180 ,w__13614);
  buf g__1005(w__14179 ,w__13613);
  buf g__1006(w__14178 ,w__13612);
  buf g__1007(w__14177 ,w__13595);
  buf g__1008(w__14176 ,w__13610);
  buf g__1009(w__14175 ,w__13609);
  buf g__1010(w__14174 ,w__13608);
  buf g__1011(w__14173 ,w__13607);
  buf g__1012(w__14172 ,w__13606);
  buf g__1013(w__14171 ,w__13605);
  buf g__1014(w__14170 ,w__13604);
  buf g__1015(w__14169 ,w__13603);
  buf g__1016(w__14168 ,w__13602);
  buf g__1017(w__14167 ,w__13601);
  buf g__1018(w__14166 ,w__13600);
  buf g__1019(w__14165 ,w__13599);
  buf g__1020(w__14164 ,w__13598);
  buf g__1021(w__14163 ,w__13597);
  and g__1022(w__14162 ,w__14182 ,w__14115);
  and g__1023(w__12744 ,w__14193 ,w__14136);
  and g__1024(w__14161 ,w__14164 ,w__14133);
  and g__1025(w__14160 ,w__14168 ,w__14125);
  and g__1026(w__12730 ,w__14176 ,w__14131);
  and g__1027(w__14159 ,w__14192 ,w__14127);
  and g__1028(w__12737 ,w__14169 ,w__14131);
  and g__1029(w__14158 ,w__14178 ,w__14127);
  and g__1030(w__12727 ,w__14179 ,w__14119);
  and g__1031(w__14157 ,w__14165 ,w__14125);
  and g__1032(w__12736 ,w__14170 ,w__14118);
  and g__1033(w__14156 ,w__14180 ,w__14121);
  and g__1034(w__14155 ,w__14181 ,w__14124);
  and g__1035(w__12735 ,w__14171 ,w__14134);
  and g__1036(w__12745 ,w__14177 ,w__14122);
  and g__1037(w__12715 ,w__14191 ,w__14134);
  and g__1038(w__14154 ,w__14163 ,w__14116);
  and g__1039(w__14153 ,w__14166 ,w__14137);
  and g__1040(w__14152 ,w__14172 ,w__14121);
  and g__1041(w__14151 ,w__14184 ,w__14130);
  and g__1042(w__14150 ,w__14185 ,w__14137);
  and g__1043(w__14149 ,w__14173 ,w__14128);
  and g__1044(w__14148 ,w__14186 ,w__14124);
  and g__1045(w__14147 ,w__14187 ,w__14128);
  and g__1046(w__14146 ,w__14167 ,w__14118);
  and g__1047(w__14145 ,w__14174 ,w__14133);
  and g__1048(w__14144 ,w__14188 ,w__14122);
  and g__1049(w__14143 ,w__14189 ,w__14130);
  and g__1050(w__12731 ,w__14175 ,w__14116);
  and g__1051(w__12716 ,w__14190 ,w__14136);
  and g__1052(w__14142 ,w__14183 ,w__14115);
  not g__1053(w__14141 ,in3);
  not g__1054(w__14140 ,in3);
  not g__1055(w__14139 ,in3);
  not g__1056(w__14138 ,in3);
  buf g__1057(w__12723 ,w__14142);
  buf g__1058(w__12740 ,w__14153);
  buf g__1059(w__12734 ,w__14152);
  buf g__1060(w__12718 ,w__14144);
  buf g__1061(w__12732 ,w__14145);
  buf g__1062(w__12739 ,w__14146);
  buf g__1063(w__12729 ,w__14159);
  buf g__1064(w__12720 ,w__14148);
  buf g__1065(w__12733 ,w__14149);
  buf g__1066(w__12721 ,w__14150);
  buf g__1067(w__12738 ,w__14160);
  buf g__1068(w__12724 ,w__14162);
  buf g__1069(w__12728 ,w__14158);
  buf g__1070(w__12743 ,w__14154);
  buf g__1071(w__12725 ,w__14155);
  buf g__1072(w__12726 ,w__14156);
  buf g__1073(w__12722 ,w__14151);
  buf g__1074(w__12741 ,w__14157);
  buf g__1075(w__12719 ,w__14147);
  buf g__1076(w__12742 ,w__14161);
  buf g__1077(w__12717 ,w__14143);
  not g__1078(w__14137 ,w__14135);
  not g__1079(w__14136 ,w__14135);
  not g__1080(w__14135 ,w__14141);
  not g__1081(w__14134 ,w__14132);
  not g__1082(w__14133 ,w__14132);
  not g__1083(w__14132 ,w__14138);
  not g__1084(w__14131 ,w__14129);
  not g__1085(w__14130 ,w__14129);
  not g__1086(w__14129 ,w__14138);
  not g__1087(w__14128 ,w__14126);
  not g__1088(w__14127 ,w__14126);
  not g__1089(w__14126 ,w__14139);
  not g__1090(w__14125 ,w__14123);
  not g__1091(w__14124 ,w__14123);
  not g__1092(w__14123 ,w__14139);
  not g__1093(w__14122 ,w__14120);
  not g__1094(w__14121 ,w__14120);
  not g__1095(w__14120 ,w__14140);
  not g__1096(w__14119 ,w__14117);
  not g__1097(w__14118 ,w__14117);
  not g__1098(w__14117 ,w__14140);
  not g__1099(w__14116 ,w__14114);
  not g__1100(w__14115 ,w__14114);
  not g__1101(w__14114 ,w__14141);
  buf g__1102(w__14276 ,w__13675);
  buf g__1103(w__14275 ,w__13689);
  buf g__1104(w__14274 ,w__13688);
  buf g__1105(w__14273 ,w__13687);
  buf g__1106(w__14272 ,w__13685);
  buf g__1107(w__14271 ,w__13684);
  buf g__1108(w__14270 ,w__13683);
  buf g__1109(w__14269 ,w__13681);
  buf g__1110(w__14268 ,w__13680);
  buf g__1111(w__14267 ,w__13679);
  buf g__1112(w__14266 ,w__13678);
  buf g__1113(w__14265 ,w__13677);
  buf g__1114(w__14264 ,w__13676);
  buf g__1115(w__14263 ,w__13659);
  buf g__1116(w__14262 ,w__13673);
  buf g__1117(w__14261 ,w__13672);
  buf g__1118(w__14260 ,w__13671);
  buf g__1119(w__14259 ,w__13669);
  buf g__1120(w__14258 ,w__13668);
  buf g__1121(w__14257 ,w__13667);
  buf g__1122(w__14256 ,w__13666);
  buf g__1123(w__14255 ,w__13665);
  buf g__1124(w__14254 ,w__13664);
  buf g__1125(w__14253 ,w__13663);
  buf g__1126(w__14252 ,w__13662);
  buf g__1127(w__14251 ,w__13661);
  buf g__1128(w__14250 ,w__13660);
  buf g__1129(w__14249 ,w__13670);
  buf g__1130(w__14248 ,w__13674);
  buf g__1131(w__14247 ,w__13682);
  buf g__1132(w__14246 ,w__13686);
  buf g__1133(w__14245 ,w__13690);
  and g__1134(w__14244 ,w__14268 ,w__14195);
  and g__1135(w__14243 ,w__14250 ,w__14216);
  and g__1136(w__14242 ,w__14252 ,w__14213);
  and g__1137(w__14241 ,w__14256 ,w__14205);
  and g__1138(w__12699 ,w__14248 ,w__14211);
  and g__1139(w__14240 ,w__14245 ,w__14199);
  and g__1140(w__14239 ,w__14276 ,w__14207);
  and g__1141(w__12706 ,w__14257 ,w__14211);
  and g__1142(w__14238 ,w__14264 ,w__14207);
  and g__1143(w__14237 ,w__14265 ,w__14199);
  and g__1144(w__14236 ,w__14253 ,w__14205);
  and g__1145(w__12705 ,w__14258 ,w__14198);
  and g__1146(w__14235 ,w__14266 ,w__14201);
  and g__1147(w__14234 ,w__14267 ,w__14204);
  and g__1148(w__12704 ,w__14259 ,w__14214);
  and g__1149(w__12714 ,w__14263 ,w__14202);
  and g__1150(w__14233 ,w__14275 ,w__14214);
  and g__1151(w__14232 ,w__14251 ,w__14196);
  and g__1152(w__14231 ,w__14254 ,w__14217);
  and g__1153(w__14230 ,w__14249 ,w__14201);
  and g__1154(w__14229 ,w__14247 ,w__14210);
  and g__1155(w__14228 ,w__14270 ,w__14217);
  and g__1156(w__14227 ,w__14260 ,w__14208);
  and g__1157(w__12689 ,w__14271 ,w__14204);
  and g__1158(w__12688 ,w__14272 ,w__14208);
  and g__1159(w__14226 ,w__14255 ,w__14198);
  and g__1160(w__14225 ,w__14261 ,w__14213);
  and g__1161(w__12687 ,w__14246 ,w__14202);
  and g__1162(w__14224 ,w__14273 ,w__14210);
  and g__1163(w__12700 ,w__14262 ,w__14196);
  and g__1164(w__14223 ,w__14274 ,w__14216);
  and g__1165(w__14222 ,w__14269 ,w__14195);
  not g__1166(w__14221 ,in6);
  not g__1167(w__14220 ,in6);
  not g__1168(w__14219 ,in6);
  not g__1169(w__14218 ,in6);
  buf g__1170(w__12710 ,w__14236);
  buf g__1171(w__12690 ,w__14228);
  buf g__1172(w__12702 ,w__14227);
  buf g__1173(w__12701 ,w__14225);
  buf g__1174(w__12697 ,w__14238);
  buf g__1175(w__12683 ,w__14240);
  buf g__1176(w__12707 ,w__14241);
  buf g__1177(w__12696 ,w__14237);
  buf g__1178(w__12691 ,w__14229);
  buf g__1179(w__12703 ,w__14230);
  buf g__1180(w__12709 ,w__14231);
  buf g__1181(w__12698 ,w__14239);
  buf g__1182(w__12712 ,w__14232);
  buf g__1183(w__12694 ,w__14234);
  buf g__1184(w__12713 ,w__14243);
  buf g__1185(w__12684 ,w__14233);
  buf g__1186(w__12693 ,w__14244);
  buf g__1187(w__12711 ,w__14242);
  buf g__1188(w__12695 ,w__14235);
  buf g__1189(w__12685 ,w__14223);
  buf g__1190(w__12692 ,w__14222);
  buf g__1191(w__12708 ,w__14226);
  buf g__1192(w__12686 ,w__14224);
  not g__1193(w__14217 ,w__14215);
  not g__1194(w__14216 ,w__14215);
  not g__1195(w__14215 ,w__14221);
  not g__1196(w__14214 ,w__14212);
  not g__1197(w__14213 ,w__14212);
  not g__1198(w__14212 ,w__14218);
  not g__1199(w__14211 ,w__14209);
  not g__1200(w__14210 ,w__14209);
  not g__1201(w__14209 ,w__14218);
  not g__1202(w__14208 ,w__14206);
  not g__1203(w__14207 ,w__14206);
  not g__1204(w__14206 ,w__14219);
  not g__1205(w__14205 ,w__14203);
  not g__1206(w__14204 ,w__14203);
  not g__1207(w__14203 ,w__14219);
  not g__1208(w__14202 ,w__14200);
  not g__1209(w__14201 ,w__14200);
  not g__1210(w__14200 ,w__14220);
  not g__1211(w__14199 ,w__14197);
  not g__1212(w__14198 ,w__14197);
  not g__1213(w__14197 ,w__14220);
  not g__1214(w__14196 ,w__14194);
  not g__1215(w__14195 ,w__14194);
  not g__1216(w__14194 ,w__14221);
  buf g__1217(w__14339 ,w__13731);
  buf g__1218(w__14338 ,w__13739);
  buf g__1219(w__14337 ,w__13753);
  buf g__1220(w__14336 ,w__13752);
  buf g__1221(w__14335 ,w__13751);
  buf g__1222(w__14334 ,w__13750);
  buf g__1223(w__14333 ,w__13749);
  buf g__1224(w__14332 ,w__13748);
  buf g__1225(w__14331 ,w__13747);
  buf g__1226(w__14330 ,w__13746);
  buf g__1227(w__14329 ,w__13745);
  buf g__1228(w__14328 ,w__13744);
  buf g__1229(w__14327 ,w__13743);
  buf g__1230(w__14326 ,w__13742);
  buf g__1231(w__14325 ,w__13741);
  buf g__1232(w__14324 ,w__13740);
  buf g__1233(w__14323 ,w__13723);
  buf g__1234(w__14322 ,w__13738);
  buf g__1235(w__14321 ,w__13737);
  buf g__1236(w__14320 ,w__13736);
  buf g__1237(w__14319 ,w__13735);
  buf g__1238(w__14318 ,w__13734);
  buf g__1239(w__14317 ,w__13733);
  buf g__1240(w__14316 ,w__13732);
  buf g__1241(w__14315 ,w__13730);
  buf g__1242(w__14314 ,w__13729);
  buf g__1243(w__14313 ,w__13728);
  buf g__1244(w__14312 ,w__13727);
  buf g__1245(w__14311 ,w__13726);
  buf g__1246(w__14310 ,w__13725);
  buf g__1247(w__14309 ,w__13724);
  and g__1248(w__12661 ,w__14328 ,w__14278);
  and g__1249(w__12681 ,w__14309 ,w__14299);
  and g__1250(w__12679 ,w__14311 ,w__14284);
  and g__1251(w__12675 ,w__14315 ,w__14288);
  and g__1252(w__12667 ,w__14322 ,w__14282);
  and g__1253(w__12666 ,w__14338 ,w__14290);
  and g__1254(w__12674 ,w__14339 ,w__14282);
  and g__1255(w__12665 ,w__14324 ,w__14290);
  and g__1256(w__12664 ,w__14325 ,w__14294);
  and g__1257(w__12678 ,w__14312 ,w__14288);
  and g__1258(w__12673 ,w__14316 ,w__14293);
  and g__1259(w__12663 ,w__14326 ,w__14296);
  and g__1260(w__12662 ,w__14327 ,w__14287);
  and g__1261(w__12672 ,w__14317 ,w__14285);
  and g__1262(w__12682 ,w__14323 ,w__14297);
  and g__1263(w__12652 ,w__14337 ,w__14285);
  and g__1264(w__12680 ,w__14310 ,w__14279);
  and g__1265(w__12677 ,w__14313 ,w__14300);
  and g__1266(w__12671 ,w__14318 ,w__14296);
  and g__1267(w__12659 ,w__14330 ,w__14281);
  and g__1268(w__12658 ,w__14331 ,w__14300);
  and g__1269(w__12670 ,w__14319 ,w__14291);
  and g__1270(w__14308 ,w__14332 ,w__14287);
  and g__1271(w__14307 ,w__14333 ,w__14291);
  and g__1272(w__12676 ,w__14314 ,w__14293);
  and g__1273(w__12669 ,w__14320 ,w__14284);
  and g__1274(w__14306 ,w__14334 ,w__14297);
  and g__1275(w__12654 ,w__14335 ,w__14281);
  and g__1276(w__12668 ,w__14321 ,w__14279);
  and g__1277(w__14305 ,w__14336 ,w__14299);
  and g__1278(w__12660 ,w__14329 ,w__14278);
  not g__1279(w__14304 ,in6);
  not g__1280(w__14303 ,in6);
  not g__1281(w__14302 ,in6);
  not g__1282(w__14301 ,in6);
  buf g__1283(w__12656 ,w__14307);
  buf g__1284(w__12657 ,w__14308);
  buf g__1285(w__12653 ,w__14305);
  buf g__1286(w__12655 ,w__14306);
  not g__1287(w__14300 ,w__14298);
  not g__1288(w__14299 ,w__14298);
  not g__1289(w__14298 ,w__14304);
  not g__1290(w__14297 ,w__14295);
  not g__1291(w__14296 ,w__14295);
  not g__1292(w__14295 ,w__14303);
  not g__1293(w__14294 ,w__14292);
  not g__1294(w__14293 ,w__14292);
  not g__1295(w__14292 ,w__14303);
  not g__1296(w__14291 ,w__14289);
  not g__1297(w__14290 ,w__14289);
  not g__1298(w__14289 ,w__14302);
  not g__1299(w__14288 ,w__14286);
  not g__1300(w__14287 ,w__14286);
  not g__1301(w__14286 ,w__14302);
  not g__1302(w__14285 ,w__14283);
  not g__1303(w__14284 ,w__14283);
  not g__1304(w__14283 ,w__14301);
  not g__1305(w__14282 ,w__14280);
  not g__1306(w__14281 ,w__14280);
  not g__1307(w__14280 ,w__14301);
  not g__1308(w__14279 ,w__14277);
  not g__1309(w__14278 ,w__14277);
  not g__1310(w__14277 ,w__14304);
  xnor g__1311(out1[31] ,w__2397 ,w__2341);
  nor g__1312(w__2397 ,w__2396 ,w__2280);
  xnor g__1313(out1[30] ,w__2395 ,w__2340);
  and g__1314(w__2396 ,w__2286 ,w__2395);
  or g__1315(w__2395 ,w__2278 ,w__2394);
  xnor g__1316(out1[29] ,w__2393 ,w__2339);
  nor g__1317(w__2394 ,w__2287 ,w__2393);
  and g__1318(w__2393 ,w__2392 ,w__2289);
  or g__1319(w__2392 ,w__2318 ,w__2391);
  and g__1320(w__2391 ,w__2296 ,w__2390);
  xnor g__1321(out1[27] ,w__2389 ,w__2337);
  or g__1322(w__2390 ,w__2282 ,w__2389);
  and g__1323(w__2389 ,w__2388 ,w__2291);
  or g__1324(w__2388 ,w__2304 ,w__2387);
  and g__1325(w__2387 ,w__2279 ,w__2386);
  xnor g__1326(out1[25] ,w__2385 ,w__2335);
  or g__1327(w__2386 ,w__2385 ,w__2281);
  and g__1328(w__2385 ,w__2384 ,w__2292);
  or g__1329(w__2384 ,w__2319 ,w__2383);
  and g__1330(w__2383 ,w__2316 ,w__2382);
  xnor g__1331(out1[23] ,w__2381 ,w__2334);
  or g__1332(w__2382 ,w__2381 ,w__2293);
  and g__1333(w__2381 ,w__2285 ,w__2380);
  or g__1334(w__2380 ,w__2283 ,w__2379);
  and g__1335(w__2379 ,w__2310 ,w__2378);
  xnor g__1336(out1[21] ,w__2377 ,w__2331);
  or g__1337(w__2378 ,w__2377 ,w__2294);
  and g__1338(w__2377 ,w__2306 ,w__2376);
  or g__1339(w__2376 ,w__2302 ,w__2375);
  and g__1340(w__2375 ,w__2301 ,w__2374);
  xnor g__1341(out1[19] ,w__2373 ,w__2329);
  or g__1342(w__2374 ,w__2373 ,w__2295);
  and g__1343(w__2373 ,w__2251 ,w__2372);
  xnor g__1344(out1[18] ,w__2370 ,w__2273);
  or g__1345(w__2372 ,w__2245 ,w__2371);
  not g__1346(w__2371 ,w__2370);
  or g__1347(w__2370 ,w__2246 ,w__2369);
  xnor g__1348(out1[17] ,w__2368 ,w__2277);
  and g__1349(w__2369 ,w__2368 ,w__2252);
  or g__1350(w__2368 ,w__2288 ,w__2367);
  xnor g__1351(out1[16] ,w__2366 ,w__2342);
  nor g__1352(w__2367 ,w__2366 ,w__2284);
  and g__1353(w__2366 ,w__2365 ,w__2248);
  or g__1354(w__2365 ,w__2242 ,w__2364);
  and g__1355(w__2364 ,w__2317 ,w__2363);
  or g__1356(w__2363 ,w__2362 ,w__2300);
  and g__1357(w__2362 ,w__2315 ,w__2361);
  or g__1358(w__2361 ,w__2314 ,w__2360);
  and g__1359(w__2360 ,w__2359 ,w__2297);
  or g__1360(w__2359 ,w__2313 ,w__2358);
  and g__1361(w__2358 ,w__2312 ,w__2357);
  or g__1362(w__2357 ,w__2356 ,w__2298);
  and g__1363(w__2356 ,w__2311 ,w__2355);
  or g__1364(w__2355 ,w__2309 ,w__2354);
  and g__1365(w__2354 ,w__2353 ,w__2299);
  or g__1366(w__2353 ,w__2308 ,w__2352);
  and g__1367(w__2352 ,w__2351 ,w__2290);
  or g__1368(w__2351 ,w__2307 ,w__2350);
  and g__1369(w__2350 ,w__2305 ,w__2349);
  xnor g__1370(out1[7] ,w__2348 ,w__2328);
  or g__1371(w__2349 ,w__2303 ,w__2348);
  and g__1372(w__2348 ,w__2347 ,w__2249);
  or g__1373(w__2347 ,w__2247 ,w__2346);
  and g__1374(w__2346 ,w__2244 ,w__2345);
  or g__1375(w__2345 ,w__2243 ,w__2344);
  and g__1376(w__2344 ,w__2163 ,w__2343);
  xnor g__1377(out1[4] ,w__2320 ,w__2209);
  or g__1378(w__2343 ,w__2162 ,w__2320);
  xnor g__1379(w__2342 ,w__2263 ,w__2215);
  xnor g__1380(w__2341 ,w__2160 ,w__2210);
  xnor g__1381(w__2340 ,w__2156 ,w__2232);
  xnor g__1382(w__2339 ,w__2159 ,w__2236);
  xnor g__1383(w__2338 ,w__2208 ,w__2231);
  xnor g__1384(w__2337 ,w__2206 ,w__2226);
  xnor g__1385(w__2336 ,w__2168 ,w__2221);
  xnor g__1386(w__2335 ,w__2127 ,w__2239);
  xnor g__1387(w__2334 ,w__2197 ,w__2233);
  xnor g__1388(w__2333 ,w__2155 ,w__2235);
  xnor g__1389(w__2332 ,w__2260 ,w__2256);
  xnor g__1390(w__2331 ,w__2201 ,w__2227);
  xnor g__1391(w__2330 ,w__2196 ,w__2224);
  xnor g__1392(w__2329 ,w__2157 ,w__2222);
  xnor g__1393(w__2328 ,w__2194 ,w__2241);
  xnor g__1394(w__2327 ,w__2262 ,w__2258);
  xnor g__1395(w__2326 ,w__2200 ,w__2229);
  xnor g__1396(w__2325 ,w__2254 ,w__2266);
  xnor g__1397(w__2324 ,w__2272 ,w__2214);
  xnor g__1398(w__2323 ,w__2204 ,w__2212);
  xnor g__1399(w__2322 ,w__2270 ,w__2219);
  xnor g__1400(w__2321 ,w__2268 ,w__2217);
  nor g__1401(w__2319 ,w__2155 ,w__2235);
  nor g__1402(w__2318 ,w__2208 ,w__2231);
  or g__1403(w__2317 ,w__2261 ,w__2257);
  or g__1404(w__2316 ,w__2198 ,w__2233);
  or g__1405(w__2315 ,w__2259 ,w__2255);
  nor g__1406(w__2314 ,w__2260 ,w__2256);
  nor g__1407(w__2313 ,w__2254 ,w__2266);
  or g__1408(w__2312 ,w__2271 ,w__2213);
  or g__1409(w__2311 ,w__2203 ,w__2211);
  or g__1410(w__2310 ,w__2202 ,w__2227);
  nor g__1411(w__2309 ,w__2204 ,w__2212);
  nor g__1412(w__2308 ,w__2270 ,w__2219);
  nor g__1413(w__2307 ,w__2268 ,w__2217);
  or g__1414(w__2306 ,w__2195 ,w__2223);
  or g__1415(w__2305 ,w__2194 ,w__2240);
  nor g__1416(w__2304 ,w__2168 ,w__2221);
  nor g__1417(w__2303 ,w__2193 ,w__2241);
  nor g__1418(w__2302 ,w__2196 ,w__2224);
  or g__1419(w__2301 ,w__2158 ,w__2222);
  nor g__1420(w__2300 ,w__2262 ,w__2258);
  or g__1421(w__2299 ,w__2269 ,w__2218);
  nor g__1422(w__2298 ,w__2272 ,w__2214);
  or g__1423(w__2297 ,w__2253 ,w__2265);
  and g__1424(w__2320 ,w__2123 ,w__2250);
  or g__1425(w__2296 ,w__2206 ,w__2225);
  and g__1426(w__2295 ,w__2158 ,w__2222);
  and g__1427(w__2294 ,w__2202 ,w__2227);
  and g__1428(w__2293 ,w__2198 ,w__2233);
  or g__1429(w__2292 ,w__2154 ,w__2234);
  or g__1430(w__2291 ,w__2167 ,w__2220);
  or g__1431(w__2290 ,w__2267 ,w__2216);
  or g__1432(w__2289 ,w__2207 ,w__2230);
  nor g__1433(w__2288 ,w__2264 ,w__2215);
  and g__1434(w__2287 ,w__2159 ,w__2237);
  or g__1435(w__2286 ,w__2156 ,w__2232);
  or g__1436(w__2285 ,w__2199 ,w__2228);
  and g__1437(w__2284 ,w__2264 ,w__2215);
  nor g__1438(w__2283 ,w__2200 ,w__2229);
  nor g__1439(w__2282 ,w__2205 ,w__2226);
  nor g__1440(w__2281 ,w__2126 ,w__2239);
  and g__1441(w__2280 ,w__2156 ,w__2232);
  or g__1442(w__2279 ,w__2127 ,w__2238);
  nor g__1443(w__2278 ,w__2159 ,w__2237);
  xnor g__1444(out1[3] ,w__2183 ,w__2161);
  xnor g__1445(w__2277 ,w__2180 ,w__2175);
  xnor g__1446(w__2276 ,w__2166 ,w__2174);
  xnor g__1447(w__2275 ,w__2179 ,w__2172);
  xnor g__1448(w__2274 ,w__2192 ,w__2177);
  xnor g__1449(w__2273 ,w__2182 ,w__2170);
  not g__1450(w__2271 ,w__2272);
  not g__1451(w__2269 ,w__2270);
  not g__1452(w__2267 ,w__2268);
  not g__1453(w__2265 ,w__2266);
  not g__1454(w__2264 ,w__2263);
  not g__1455(w__2261 ,w__2262);
  not g__1456(w__2259 ,w__2260);
  not g__1457(w__2257 ,w__2258);
  not g__1458(w__2255 ,w__2256);
  not g__1459(w__2253 ,w__2254);
  or g__1460(w__2252 ,w__2180 ,w__2175);
  or g__1461(w__2251 ,w__2181 ,w__2169);
  or g__1462(w__2250 ,w__2184 ,w__2121);
  or g__1463(w__2249 ,w__2165 ,w__2173);
  or g__1464(w__2248 ,w__2191 ,w__2176);
  nor g__1465(w__2247 ,w__2166 ,w__2174);
  and g__1466(w__2246 ,w__2180 ,w__2175);
  nor g__1467(w__2245 ,w__2182 ,w__2170);
  or g__1468(w__2244 ,w__2178 ,w__2171);
  nor g__1469(w__2243 ,w__2179 ,w__2172);
  nor g__1470(w__2242 ,w__2192 ,w__2177);
  or g__1471(w__2272 ,w__2142 ,w__2190);
  or g__1472(w__2270 ,w__2137 ,w__2187);
  or g__1473(w__2268 ,w__2135 ,w__2189);
  xnor g__1474(w__2266 ,w__2058 ,w__2099);
  or g__1475(w__2263 ,w__2119 ,w__2164);
  or g__1476(w__2262 ,w__2151 ,w__2188);
  or g__1477(w__2260 ,w__2147 ,w__2186);
  xnor g__1478(w__2258 ,w__2006 ,w__2101);
  xnor g__1479(w__2256 ,w__2062 ,w__2100);
  or g__1480(w__2254 ,w__2145 ,w__2185);
  not g__1481(w__2240 ,w__2241);
  not g__1482(w__2239 ,w__2238);
  not g__1483(w__2237 ,w__2236);
  not g__1484(w__2235 ,w__2234);
  not g__1485(w__2231 ,w__2230);
  not g__1486(w__2229 ,w__2228);
  not g__1487(w__2226 ,w__2225);
  not g__1488(w__2224 ,w__2223);
  not g__1489(w__2221 ,w__2220);
  not g__1490(w__2218 ,w__2219);
  not g__1491(w__2216 ,w__2217);
  not g__1492(w__2213 ,w__2214);
  not g__1493(w__2211 ,w__2212);
  xor g__1494(out1[2] ,w__2035 ,w__2116);
  xnor g__1495(w__2210 ,w__1955 ,w__2103);
  xnor g__1496(w__2209 ,w__2094 ,w__2125);
  xnor g__1497(w__2241 ,w__2060 ,w__2104);
  xnor g__1498(w__2238 ,w__1990 ,w__2115);
  xnor g__1499(w__2236 ,w__1977 ,w__2114);
  xnor g__1500(w__2234 ,w__1960 ,w__2113);
  xnor g__1501(w__2233 ,w__1979 ,w__2112);
  xnor g__1502(w__2232 ,w__2034 ,w__2110);
  xnor g__1503(w__2230 ,w__1964 ,w__2111);
  xnor g__1504(w__2228 ,w__1983 ,w__2109);
  xnor g__1505(w__2227 ,w__1986 ,w__2108);
  xnor g__1506(w__2225 ,w__1984 ,w__2107);
  xnor g__1507(w__2223 ,w__1985 ,w__2106);
  xnor g__1508(w__2222 ,w__1982 ,w__2117);
  xnor g__1509(w__2220 ,w__1988 ,w__2102);
  xnor g__1510(w__2219 ,w__2067 ,w__2096);
  xnor g__1511(w__2217 ,w__2061 ,w__2095);
  xnor g__1512(w__2215 ,w__2016 ,w__2105);
  xnor g__1513(w__2214 ,w__2064 ,w__2098);
  xnor g__1514(w__2212 ,w__2063 ,w__2097);
  not g__1515(w__2207 ,w__2208);
  not g__1516(w__2206 ,w__2205);
  not g__1517(w__2203 ,w__2204);
  not g__1518(w__2202 ,w__2201);
  not g__1519(w__2200 ,w__2199);
  not g__1520(w__2198 ,w__2197);
  not g__1521(w__2195 ,w__2196);
  not g__1522(w__2194 ,w__2193);
  not g__1523(w__2191 ,w__2192);
  nor g__1524(w__2190 ,w__2038 ,w__2141);
  nor g__1525(w__2189 ,w__2042 ,w__2133);
  nor g__1526(w__2188 ,w__2039 ,w__2148);
  nor g__1527(w__2187 ,w__2041 ,w__2136);
  nor g__1528(w__2186 ,w__2036 ,w__2146);
  nor g__1529(w__2185 ,w__2037 ,w__2143);
  or g__1530(w__2208 ,w__2088 ,w__2150);
  or g__1531(w__2205 ,w__2082 ,w__2153);
  or g__1532(w__2204 ,w__2081 ,w__2138);
  or g__1533(w__2201 ,w__2092 ,w__2139);
  and g__1534(w__2199 ,w__2084 ,w__2144);
  or g__1535(w__2197 ,w__2086 ,w__2149);
  or g__1536(w__2196 ,w__2050 ,w__2134);
  or g__1537(w__2193 ,w__2022 ,w__2132);
  or g__1538(w__2192 ,w__2091 ,w__2152);
  not g__1539(w__2184 ,w__2183);
  not g__1540(w__2181 ,w__2182);
  not g__1541(w__2179 ,w__2178);
  not g__1542(w__2176 ,w__2177);
  not g__1543(w__2174 ,w__2173);
  not g__1544(w__2172 ,w__2171);
  not g__1545(w__2170 ,w__2169);
  not g__1546(w__2167 ,w__2168);
  not g__1547(w__2165 ,w__2166);
  nor g__1548(w__2164 ,w__1967 ,w__2140);
  or g__1549(w__2163 ,w__2093 ,w__2125);
  nor g__1550(w__2162 ,w__2094 ,w__2124);
  xnor g__1551(w__2161 ,w__2059 ,w__1909);
  nor g__1552(w__2160 ,w__2056 ,w__2120);
  or g__1553(w__2183 ,w__2069 ,w__2122);
  or g__1554(w__2182 ,w__2068 ,w__2128);
  or g__1555(w__2180 ,w__2052 ,w__2118);
  and g__1556(w__2178 ,w__2071 ,w__2130);
  xnor g__1557(w__2177 ,w__2065 ,w__2047);
  xnor g__1558(w__2175 ,w__2011 ,w__2043);
  xnor g__1559(w__2173 ,w__2066 ,w__2045);
  xnor g__1560(w__2171 ,w__2003 ,w__2044);
  xnor g__1561(w__2169 ,w__1989 ,w__2046);
  or g__1562(w__2168 ,w__2075 ,w__2129);
  or g__1563(w__2166 ,w__2074 ,w__2131);
  not g__1564(w__2158 ,w__2157);
  not g__1565(w__2154 ,w__2155);
  and g__1566(w__2153 ,w__1988 ,w__2076);
  nor g__1567(w__2152 ,w__2040 ,w__2089);
  and g__1568(w__2151 ,w__1831 ,w__2062);
  and g__1569(w__2150 ,w__1984 ,w__2083);
  and g__1570(w__2149 ,w__1983 ,w__2085);
  nor g__1571(w__2148 ,w__1831 ,w__2062);
  and g__1572(w__2147 ,w__1824 ,w__2058);
  nor g__1573(w__2146 ,w__1824 ,w__2058);
  and g__1574(w__2145 ,w__1821 ,w__2064);
  or g__1575(w__2144 ,w__1987 ,w__2080);
  nor g__1576(w__2143 ,w__1821 ,w__2064);
  and g__1577(w__2142 ,w__1818 ,w__2063);
  nor g__1578(w__2141 ,w__1818 ,w__2063);
  nor g__1579(w__2140 ,w__1789 ,w__2065);
  and g__1580(w__2139 ,w__1985 ,w__2077);
  and g__1581(w__2138 ,w__2078 ,w__2067);
  and g__1582(w__2137 ,w__1810 ,w__2061);
  nor g__1583(w__2136 ,w__1810 ,w__2061);
  and g__1584(w__2135 ,w__1807 ,w__2060);
  and g__1585(w__2134 ,w__1982 ,w__2049);
  nor g__1586(w__2133 ,w__1807 ,w__2060);
  nor g__1587(w__2132 ,w__2023 ,w__2066);
  nor g__1588(w__2131 ,w__1981 ,w__2072);
  or g__1589(w__2130 ,w__1870 ,w__2070);
  and g__1590(w__2129 ,w__1990 ,w__2054);
  nor g__1591(w__2128 ,w__1965 ,w__2053);
  and g__1592(w__2159 ,w__2032 ,w__2090);
  or g__1593(w__2157 ,w__2024 ,w__2073);
  or g__1594(w__2156 ,w__2028 ,w__2057);
  or g__1595(w__2155 ,w__2031 ,w__2087);
  not g__1596(w__2127 ,w__2126);
  not g__1597(w__2125 ,w__2124);
  or g__1598(w__2123 ,w__1909 ,w__2059);
  and g__1599(w__2122 ,w__2035 ,w__2048);
  and g__1600(w__2121 ,w__1909 ,w__2059);
  and g__1601(w__2120 ,w__2055 ,w__2018);
  and g__1602(w__2119 ,w__1789 ,w__2065);
  and g__1603(w__2118 ,w__2016 ,w__2051);
  xnor g__1604(w__2117 ,w__1786 ,w__2008);
  xnor g__1605(w__2116 ,w__1797 ,w__1997);
  xnor g__1606(w__2115 ,w__1803 ,w__2005);
  xnor g__1607(w__2114 ,w__1865 ,w__2019);
  xnor g__1608(w__2113 ,w__1780 ,w__2021);
  xnor g__1609(w__2112 ,w__1788 ,w__2017);
  xnor g__1610(w__2111 ,w__1794 ,w__2020);
  xnor g__1611(w__2110 ,w__1815 ,w__2018);
  xnor g__1612(w__2109 ,w__1826 ,w__2015);
  xnor g__1613(w__2108 ,w__1908 ,w__2013);
  xnor g__1614(w__2107 ,w__1830 ,w__2000);
  xnor g__1615(w__2106 ,w__1812 ,w__2010);
  xnor g__1616(w__2105 ,w__1792 ,w__1995);
  xor g__1617(w__2104 ,w__1807 ,w__2042);
  xnor g__1618(w__2103 ,w__1690 ,w__1991);
  xnor g__1619(w__2102 ,w__1911 ,w__2002);
  xor g__1620(w__2101 ,w__1779 ,w__2040);
  xor g__1621(w__2100 ,w__1831 ,w__2039);
  xor g__1622(w__2099 ,w__1824 ,w__2036);
  xor g__1623(w__2098 ,w__1821 ,w__2037);
  xor g__1624(w__2097 ,w__1818 ,w__2038);
  xnor g__1625(w__2096 ,w__1814 ,w__2033);
  xor g__1626(w__2095 ,w__1810 ,w__2041);
  or g__1627(w__2126 ,w__1992 ,w__2079);
  xnor g__1628(w__2124 ,w__1998 ,w__1948);
  not g__1629(w__2093 ,w__2094);
  nor g__1630(w__2092 ,w__1811 ,w__2010);
  and g__1631(w__2091 ,w__1779 ,w__2006);
  or g__1632(w__2090 ,w__2029 ,w__2020);
  nor g__1633(w__2089 ,w__1779 ,w__2006);
  nor g__1634(w__2088 ,w__1829 ,w__2000);
  and g__1635(w__2087 ,w__2027 ,w__2017);
  nor g__1636(w__2086 ,w__1825 ,w__2015);
  or g__1637(w__2085 ,w__1826 ,w__2014);
  or g__1638(w__2084 ,w__1907 ,w__2013);
  or g__1639(w__2083 ,w__1830 ,w__1999);
  nor g__1640(w__2082 ,w__1910 ,w__2002);
  and g__1641(w__2081 ,w__1814 ,w__2033);
  nor g__1642(w__2080 ,w__1908 ,w__2012);
  and g__1643(w__2079 ,w__2030 ,w__2021);
  or g__1644(w__2078 ,w__1814 ,w__2033);
  or g__1645(w__2077 ,w__1812 ,w__2009);
  or g__1646(w__2076 ,w__1911 ,w__2001);
  nor g__1647(w__2075 ,w__1802 ,w__2005);
  nor g__1648(w__2074 ,w__1801 ,w__2003);
  and g__1649(w__2073 ,w__1989 ,w__2025);
  and g__1650(w__2072 ,w__1801 ,w__2003);
  or g__1651(w__2071 ,w__1782 ,w__1998);
  and g__1652(w__2070 ,w__1782 ,w__1998);
  nor g__1653(w__2069 ,w__1796 ,w__1997);
  and g__1654(w__2068 ,w__1798 ,w__2011);
  or g__1655(w__2094 ,w__1914 ,w__2026);
  and g__1656(w__2057 ,w__1993 ,w__2019);
  and g__1657(w__2056 ,w__1815 ,w__2034);
  or g__1658(w__2055 ,w__1815 ,w__2034);
  or g__1659(w__2054 ,w__1803 ,w__2004);
  nor g__1660(w__2053 ,w__1798 ,w__2011);
  nor g__1661(w__2052 ,w__1791 ,w__1995);
  or g__1662(w__2051 ,w__1792 ,w__1994);
  nor g__1663(w__2050 ,w__1786 ,w__2007);
  or g__1664(w__2049 ,w__1785 ,w__2008);
  or g__1665(w__2048 ,w__1797 ,w__1996);
  xnor g__1666(out1[1] ,w__1722 ,w__1953);
  xor g__1667(w__2047 ,w__1789 ,w__1967);
  xnor g__1668(w__2046 ,w__1800 ,w__1962);
  xnor g__1669(w__2045 ,w__1804 ,w__1980);
  xnor g__1670(w__2044 ,w__1981 ,w__1801);
  xor g__1671(w__2043 ,w__1798 ,w__1965);
  xnor g__1672(w__2067 ,w__1745 ,w__1952);
  xnor g__1673(w__2066 ,w__1768 ,w__1950);
  xnor g__1674(w__2065 ,w__1724 ,w__1957);
  xnor g__1675(w__2064 ,w__1747 ,w__1945);
  xnor g__1676(w__2063 ,w__1761 ,w__1949);
  xnor g__1677(w__2062 ,w__1833 ,w__1947);
  xnor g__1678(w__2061 ,w__1754 ,w__1954);
  xnor g__1679(w__2060 ,w__1864 ,w__1956);
  xnor g__1680(w__2059 ,w__1966 ,w__1951);
  xnor g__1681(w__2058 ,w__1756 ,w__1946);
  or g__1682(w__2032 ,w__1793 ,w__1963);
  nor g__1683(w__2031 ,w__1788 ,w__1978);
  or g__1684(w__2030 ,w__1781 ,w__1960);
  nor g__1685(w__2029 ,w__1794 ,w__1964);
  and g__1686(w__2028 ,w__1865 ,w__1977);
  or g__1687(w__2027 ,w__1787 ,w__1979);
  and g__1688(w__2026 ,w__1913 ,w__1966);
  or g__1689(w__2025 ,w__1800 ,w__1961);
  nor g__1690(w__2024 ,w__1799 ,w__1962);
  nor g__1691(w__2023 ,w__1804 ,w__1980);
  and g__1692(w__2022 ,w__1804 ,w__1980);
  and g__1693(w__2042 ,w__1921 ,w__1976);
  and g__1694(w__2041 ,w__1925 ,w__1969);
  and g__1695(w__2040 ,w__1942 ,w__1968);
  and g__1696(w__2039 ,w__1938 ,w__1975);
  and g__1697(w__2038 ,w__1930 ,w__1972);
  and g__1698(w__2037 ,w__1933 ,w__1973);
  and g__1699(w__2036 ,w__1936 ,w__1974);
  or g__1700(w__2035 ,w__1905 ,w__1959);
  or g__1701(w__2034 ,w__1844 ,w__1971);
  or g__1702(w__2033 ,w__1927 ,w__1970);
  not g__1703(w__2015 ,w__2014);
  not g__1704(w__2013 ,w__2012);
  not g__1705(w__2010 ,w__2009);
  not g__1706(w__2008 ,w__2007);
  not g__1707(w__2005 ,w__2004);
  not g__1708(w__2002 ,w__2001);
  not g__1709(w__2000 ,w__1999);
  not g__1710(w__1996 ,w__1997);
  not g__1711(w__1994 ,w__1995);
  or g__1712(w__1993 ,w__1865 ,w__1977);
  and g__1713(w__1992 ,w__1781 ,w__1960);
  xnor g__1714(w__1991 ,w__1896 ,w__1879);
  xnor g__1715(w__2021 ,w__1868 ,w__1892);
  xnor g__1716(w__2020 ,w__1766 ,w__1893);
  xnor g__1717(w__2019 ,w__1912 ,w__1889);
  xnor g__1718(w__2018 ,w__1876 ,w__1883);
  xnor g__1719(w__2017 ,w__1723 ,w__1894);
  or g__1720(w__2016 ,w__1902 ,w__1958);
  xnor g__1721(w__2014 ,w__1866 ,w__1888);
  xnor g__1722(w__2012 ,w__1878 ,w__1887);
  xnor g__1723(w__2011 ,w__1869 ,w__1891);
  xnor g__1724(w__2009 ,w__1873 ,w__1885);
  xnor g__1725(w__2007 ,w__1875 ,w__1884);
  xnor g__1726(w__2006 ,w__1749 ,w__1880);
  xnor g__1727(w__2004 ,w__1877 ,w__1881);
  xnor g__1728(w__2003 ,w__1713 ,w__1882);
  xnor g__1729(w__2001 ,w__1872 ,w__1886);
  xnor g__1730(w__1999 ,w__1874 ,w__1890);
  xnor g__1731(w__1998 ,w__1704 ,w__1898);
  xnor g__1732(w__1997 ,w__1721 ,w__1897);
  xnor g__1733(w__1995 ,w__1725 ,w__1895);
  not g__1734(w__1987 ,w__1986);
  not g__1735(w__1978 ,w__1979);
  or g__1736(w__1976 ,w__1769 ,w__1920);
  or g__1737(w__1975 ,w__1759 ,w__1937);
  or g__1738(w__1974 ,w__1760 ,w__1935);
  or g__1739(w__1973 ,w__1762 ,w__1931);
  or g__1740(w__1972 ,w__1764 ,w__1944);
  and g__1741(w__1971 ,w__1843 ,w__1912);
  nor g__1742(w__1970 ,w__1684 ,w__1926);
  or g__1743(w__1969 ,w__1767 ,w__1922);
  or g__1744(w__1968 ,w__1867 ,w__1939);
  or g__1745(w__1990 ,w__1848 ,w__1906);
  or g__1746(w__1989 ,w__1850 ,w__1915);
  or g__1747(w__1988 ,w__1842 ,w__1924);
  or g__1748(w__1986 ,w__1847 ,w__1929);
  or g__1749(w__1985 ,w__1841 ,w__1923);
  or g__1750(w__1984 ,w__1853 ,w__1932);
  or g__1751(w__1983 ,w__1852 ,w__1934);
  or g__1752(w__1982 ,w__1731 ,w__1919);
  and g__1753(w__1981 ,w__1845 ,w__1916);
  or g__1754(w__1980 ,w__1839 ,w__1918);
  or g__1755(w__1979 ,w__1858 ,w__1940);
  or g__1756(w__1977 ,w__1834 ,w__1917);
  not g__1757(w__1963 ,w__1964);
  not g__1758(w__1962 ,w__1961);
  and g__1759(w__1959 ,w__1722 ,w__1904);
  and g__1760(w__1958 ,w__1724 ,w__1900);
  xnor g__1761(w__1957 ,w__1708 ,w__1790);
  xor g__1762(w__1956 ,w__1767 ,w__1809);
  or g__1763(w__1955 ,w__1837 ,w__1903);
  xor g__1764(w__1954 ,w__1684 ,w__1813);
  xnor g__1765(w__1953 ,w__1494 ,w__1795);
  xor g__1766(w__1952 ,w__1764 ,w__1817);
  xnor g__1767(w__1951 ,w__1697 ,w__1784);
  xnor g__1768(w__1950 ,w__1758 ,w__1806);
  xnor g__1769(w__1949 ,w__1753 ,w__1820);
  xor g__1770(w__1948 ,w__1782 ,w__1870);
  xor g__1771(w__1947 ,w__1867 ,w__1743);
  xor g__1772(w__1946 ,w__1759 ,w__1828);
  xor g__1773(w__1945 ,w__1760 ,w__1823);
  and g__1774(w__1967 ,w__1773 ,w__1928);
  or g__1775(w__1966 ,w__1836 ,w__1899);
  and g__1776(w__1965 ,w__1862 ,w__1943);
  or g__1777(w__1964 ,w__1774 ,w__1941);
  xnor g__1778(w__1961 ,w__1871 ,w__1771);
  or g__1779(w__1960 ,w__1775 ,w__1901);
  nor g__1780(w__1944 ,w__1745 ,w__1817);
  or g__1781(w__1943 ,w__1726 ,w__1778);
  or g__1782(w__1942 ,w__1742 ,w__1832);
  and g__1783(w__1941 ,w__1861 ,w__1874);
  and g__1784(w__1940 ,w__1856 ,w__1866);
  nor g__1785(w__1939 ,w__1743 ,w__1833);
  or g__1786(w__1938 ,w__1755 ,w__1827);
  nor g__1787(w__1937 ,w__1756 ,w__1828);
  or g__1788(w__1936 ,w__1746 ,w__1822);
  nor g__1789(w__1935 ,w__1747 ,w__1823);
  and g__1790(w__1934 ,w__1851 ,w__1878);
  or g__1791(w__1933 ,w__1752 ,w__1819);
  and g__1792(w__1932 ,w__1849 ,w__1872);
  nor g__1793(w__1931 ,w__1753 ,w__1820);
  or g__1794(w__1930 ,w__1744 ,w__1816);
  nor g__1795(w__1929 ,w__1846 ,w__1873);
  or g__1796(w__1928 ,w__1765 ,w__1857);
  and g__1797(w__1927 ,w__1754 ,w__1813);
  nor g__1798(w__1926 ,w__1754 ,w__1813);
  or g__1799(w__1925 ,w__1863 ,w__1808);
  nor g__1800(w__1924 ,w__1838 ,w__1877);
  and g__1801(w__1923 ,w__1875 ,w__1835);
  nor g__1802(w__1922 ,w__1864 ,w__1809);
  or g__1803(w__1921 ,w__1758 ,w__1805);
  nor g__1804(w__1920 ,w__1757 ,w__1806);
  and g__1805(w__1919 ,w__1733 ,w__1871);
  nor g__1806(w__1918 ,w__1763 ,w__1840);
  and g__1807(w__1917 ,w__1766 ,w__1776);
  or g__1808(w__1916 ,w__1770 ,w__1854);
  and g__1809(w__1915 ,w__1869 ,w__1855);
  nor g__1810(w__1914 ,w__1696 ,w__1784);
  or g__1811(w__1913 ,w__1697 ,w__1783);
  not g__1812(w__1910 ,w__1911);
  not g__1813(w__1907 ,w__1908);
  and g__1814(w__1906 ,w__1859 ,w__1868);
  and g__1815(w__1905 ,w__1494 ,w__1795);
  or g__1816(w__1904 ,w__1494 ,w__1795);
  and g__1817(w__1903 ,w__1876 ,w__1777);
  and g__1818(w__1902 ,w__1708 ,w__1790);
  and g__1819(w__1901 ,w__1723 ,w__1860);
  or g__1820(w__1900 ,w__1708 ,w__1790);
  xnor g__1821(out1[0] ,w__847 ,w__1693);
  and g__1822(w__1899 ,w__1721 ,w__1772);
  xor g__1823(w__1898 ,w__1486 ,w__1770);
  xnor g__1824(w__1897 ,w__1484 ,w__1702);
  xnor g__1825(w__1896 ,w__1454 ,w__1692);
  xnor g__1826(w__1895 ,w__1750 ,w__1705);
  xnor g__1827(w__1894 ,w__1628 ,w__1707);
  xnor g__1828(w__1893 ,w__1677 ,w__1699);
  xnor g__1829(w__1892 ,w__1672 ,w__1710);
  xnor g__1830(w__1891 ,w__1673 ,w__1712);
  xnor g__1831(w__1890 ,w__1627 ,w__1709);
  xnor g__1832(w__1889 ,w__1678 ,w__1720);
  xnor g__1833(w__1888 ,w__1671 ,w__1700);
  xnor g__1834(w__1887 ,w__1681 ,w__1719);
  xnor g__1835(w__1886 ,w__1675 ,w__1718);
  xnor g__1836(w__1885 ,w__1679 ,w__1717);
  xnor g__1837(w__1884 ,w__1573 ,w__1716);
  xnor g__1838(w__1883 ,w__1674 ,w__1711);
  xnor g__1839(w__1882 ,w__1491 ,w__1763);
  xnor g__1840(w__1881 ,w__1682 ,w__1714);
  xor g__1841(w__1880 ,w__1765 ,w__1706);
  xnor g__1842(w__1879 ,w__1610 ,w__1687);
  xnor g__1843(w__1912 ,w__1501 ,w__1688);
  xnor g__1844(w__1911 ,w__1496 ,w__1691);
  xnor g__1845(w__1909 ,w__1482 ,w__1686);
  xnor g__1846(w__1908 ,w__1469 ,w__1689);
  not g__1847(w__1863 ,w__1864);
  or g__1848(w__1862 ,w__1751 ,w__1705);
  or g__1849(w__1861 ,w__1627 ,w__1709);
  or g__1850(w__1860 ,w__1628 ,w__1707);
  or g__1851(w__1859 ,w__1672 ,w__1710);
  and g__1852(w__1858 ,w__1671 ,w__1700);
  nor g__1853(w__1857 ,w__2 ,w__1749);
  or g__1854(w__1856 ,w__1671 ,w__1700);
  or g__1855(w__1855 ,w__1673 ,w__1712);
  nor g__1856(w__1854 ,w__1486 ,w__1703);
  and g__1857(w__1853 ,w__1675 ,w__1718);
  and g__1858(w__1852 ,w__1681 ,w__1719);
  or g__1859(w__1851 ,w__1681 ,w__1719);
  and g__1860(w__1850 ,w__1673 ,w__1712);
  or g__1861(w__1849 ,w__1675 ,w__1718);
  and g__1862(w__1848 ,w__1672 ,w__1710);
  nor g__1863(w__1847 ,w__1680 ,w__1717);
  and g__1864(w__1846 ,w__1680 ,w__1717);
  or g__1865(w__1845 ,w__1485 ,w__1704);
  and g__1866(w__1844 ,w__1678 ,w__1720);
  or g__1867(w__1843 ,w__1678 ,w__1720);
  nor g__1868(w__1842 ,w__1683 ,w__1714);
  nor g__1869(w__1841 ,w__1572 ,w__1716);
  nor g__1870(w__1840 ,w__1491 ,w__1713);
  and g__1871(w__1839 ,w__1491 ,w__1713);
  and g__1872(w__1838 ,w__1683 ,w__1714);
  and g__1873(w__1837 ,w__1674 ,w__1711);
  nor g__1874(w__1836 ,w__1483 ,w__1702);
  or g__1875(w__1835 ,w__1573 ,w__1715);
  nor g__1876(w__1834 ,w__1676 ,w__1699);
  or g__1877(w__1878 ,w__1652 ,w__1734);
  and g__1878(w__1877 ,w__1631 ,w__1729);
  or g__1879(w__1876 ,w__1658 ,w__1736);
  or g__1880(w__1875 ,w__1535 ,w__1727);
  or g__1881(w__1874 ,w__1668 ,w__1740);
  and g__1882(w__1873 ,w__1643 ,w__1730);
  or g__1883(w__1872 ,w__1648 ,w__1732);
  or g__1884(w__1871 ,w__1638 ,w__1735);
  and g__1885(w__1870 ,w__1613 ,w__1694);
  or g__1886(w__1869 ,w__1625 ,w__1695);
  or g__1887(w__1868 ,w__1649 ,w__1741);
  and g__1888(w__1867 ,w__1662 ,w__1738);
  or g__1889(w__1866 ,w__1663 ,w__1737);
  or g__1890(w__1865 ,w__1655 ,w__1739);
  or g__1891(w__1864 ,w__1636 ,w__1728);
  not g__1892(w__1832 ,w__1833);
  not g__1893(w__1829 ,w__1830);
  not g__1894(w__1827 ,w__1828);
  not g__1895(w__1825 ,w__1826);
  not g__1896(w__1822 ,w__1823);
  not g__1897(w__1819 ,w__1820);
  not g__1898(w__1816 ,w__1817);
  not g__1899(w__1811 ,w__1812);
  not g__1900(w__1808 ,w__1809);
  not g__1901(w__1805 ,w__1806);
  not g__1902(w__1802 ,w__1803);
  not g__1903(w__1799 ,w__1800);
  not g__1904(w__1796 ,w__1797);
  not g__1905(w__1793 ,w__1794);
  not g__1906(w__1791 ,w__1792);
  not g__1907(w__1788 ,w__1787);
  not g__1908(w__1786 ,w__1785);
  not g__1909(w__1783 ,w__1784);
  not g__1910(w__1781 ,w__1780);
  and g__1911(w__1778 ,w__1751 ,w__1705);
  or g__1912(w__1777 ,w__1674 ,w__1711);
  or g__1913(w__1776 ,w__1677 ,w__1698);
  and g__1914(w__1775 ,w__1628 ,w__1707);
  and g__1915(w__1774 ,w__1627 ,w__1709);
  or g__1916(w__1773 ,w__10 ,w__1748);
  or g__1917(w__1772 ,w__1484 ,w__1701);
  xnor g__1918(w__1771 ,w__1487 ,w__1629);
  xnor g__1919(w__1833 ,w__1306 ,w__1603);
  xnor g__1920(w__1831 ,w__1507 ,w__1602);
  xnor g__1921(w__1830 ,w__1505 ,w__1601);
  xnor g__1922(w__1828 ,w__1473 ,w__1600);
  xnor g__1923(w__1826 ,w__1508 ,w__1599);
  xnor g__1924(w__1824 ,w__1360 ,w__1598);
  xnor g__1925(w__1823 ,w__1504 ,w__1597);
  xnor g__1926(w__1821 ,w__1356 ,w__1596);
  xnor g__1927(w__1820 ,w__1286 ,w__1595);
  xnor g__1928(w__1818 ,w__1503 ,w__1594);
  xnor g__1929(w__1817 ,w__1498 ,w__1593);
  xnor g__1930(w__1815 ,w__1510 ,w__1587);
  xnor g__1931(w__1814 ,w__1351 ,w__1592);
  xnor g__1932(w__1813 ,w__1497 ,w__1591);
  xnor g__1933(w__1812 ,w__1480 ,w__1590);
  xnor g__1934(w__1810 ,w__1344 ,w__1589);
  xnor g__1935(w__1809 ,w__1279 ,w__1588);
  xnor g__1936(w__1807 ,w__1509 ,w__1586);
  xnor g__1937(w__1806 ,w__1495 ,w__1585);
  xnor g__1938(w__1804 ,w__1338 ,w__1584);
  xnor g__1939(w__1803 ,w__1477 ,w__1583);
  xor g__1940(w__1801 ,w__1574 ,w__1582);
  xnor g__1941(w__1800 ,w__1685 ,w__1579);
  xnor g__1942(w__1798 ,w__1490 ,w__1581);
  xnor g__1943(w__1797 ,w__1364 ,w__1580);
  xnor g__1944(w__1795 ,w__1329 ,w__1578);
  xnor g__1945(w__1794 ,w__1489 ,w__1577);
  xnor g__1946(w__1792 ,w__1488 ,w__1611);
  xnor g__1947(w__1790 ,w__1502 ,w__1608);
  xnor g__1948(w__1789 ,w__1328 ,w__1612);
  xnor g__1949(w__1787 ,w__1479 ,w__1605);
  xnor g__1950(w__1785 ,w__1471 ,w__1607);
  xnor g__1951(w__1784 ,w__1296 ,w__1609);
  xnor g__1952(w__1782 ,w__1321 ,w__1606);
  xnor g__1953(w__1780 ,w__1493 ,w__1);
  xnor g__1954(w__1779 ,w__1500 ,w__1604);
  not g__1955(w__1769 ,w__1768);
  not g__1956(w__1762 ,w__1761);
  not g__1957(w__1758 ,w__1757);
  not g__1958(w__1755 ,w__1756);
  not g__1959(w__1752 ,w__1753);
  not g__1960(w__1751 ,w__1750);
  not g__1961(w__1748 ,w__1749);
  not g__1962(w__1746 ,w__1747);
  not g__1963(w__1744 ,w__1745);
  not g__1964(w__1742 ,w__1743);
  nor g__1965(w__1741 ,w__1370 ,w__1619);
  nor g__1966(w__1740 ,w__1506 ,w__1664);
  nor g__1967(w__1739 ,w__1435 ,w__1632);
  or g__1968(w__1738 ,w__1298 ,w__1661);
  nor g__1969(w__1737 ,w__1439 ,w__1660);
  and g__1970(w__1736 ,w__1501 ,w__1666);
  nor g__1971(w__1735 ,w__1437 ,w__1657);
  nor g__1972(w__1734 ,w__1434 ,w__1650);
  or g__1973(w__1733 ,w__1487 ,w__1629);
  nor g__1974(w__1732 ,w__1425 ,w__1642);
  and g__1975(w__1731 ,w__1487 ,w__1629);
  or g__1976(w__1730 ,w__1426 ,w__1640);
  or g__1977(w__1729 ,w__1423 ,w__1646);
  nor g__1978(w__1728 ,w__1429 ,w__1635);
  and g__1979(w__1727 ,w__1533 ,w__1685);
  and g__1980(w__1770 ,w__1521 ,w__1626);
  or g__1981(w__1768 ,w__1528 ,w__1633);
  and g__1982(w__1767 ,w__1534 ,w__1634);
  or g__1983(w__1766 ,w__1524 ,w__1616);
  and g__1984(w__1765 ,w__1567 ,w__1667);
  and g__1985(w__1764 ,w__1542 ,w__1641);
  and g__1986(w__1763 ,w__1525 ,w__1653);
  or g__1987(w__1761 ,w__1548 ,w__1645);
  and g__1988(w__1760 ,w__1553 ,w__1651);
  and g__1989(w__1759 ,w__1559 ,w__1656);
  or g__1990(w__1757 ,w__1530 ,w__1630);
  or g__1991(w__1756 ,w__1561 ,w__1659);
  or g__1992(w__1754 ,w__1540 ,w__1639);
  or g__1993(w__1753 ,w__1550 ,w__1647);
  or g__1994(w__1750 ,w__1545 ,w__1621);
  or g__1995(w__1749 ,w__1539 ,w__1669);
  or g__1996(w__1747 ,w__1556 ,w__1654);
  or g__1997(w__1745 ,w__1544 ,w__1670);
  or g__1998(w__1743 ,w__1563 ,w__1665);
  not g__1999(w__1726 ,w__1725);
  not g__2000(w__1716 ,w__1715);
  not g__2001(w__1703 ,w__1704);
  not g__2002(w__1701 ,w__1702);
  not g__2003(w__1699 ,w__1698);
  not g__2004(w__1696 ,w__1697);
  nor g__2005(w__1695 ,w__1369 ,w__1637);
  or g__2006(w__1694 ,w__1576 ,w__1624);
  xnor g__2007(w__1693 ,w__813 ,w__1499);
  xnor g__2008(w__1692 ,w__1207 ,w__1457);
  xor g__2009(w__1691 ,w__1506 ,w__1414);
  or g__2010(w__1690 ,w__1516 ,w__1618);
  xor g__2011(w__1689 ,w__1439 ,w__1476);
  xnor g__2012(w__1688 ,w__1406 ,w__1478);
  xnor g__2013(w__1687 ,w__1311 ,w__1445);
  xnor g__2014(w__1686 ,w__1575 ,w__1475);
  or g__2015(w__1725 ,w__1526 ,w__1617);
  or g__2016(w__1724 ,w__1527 ,w__1614);
  or g__2017(w__1723 ,w__1564 ,w__1644);
  or g__2018(w__1722 ,w__1079 ,w__1620);
  or g__2019(w__1721 ,w__1512 ,w__1622);
  xnor g__2020(w__1720 ,w__1433 ,w__1453);
  xnor g__2021(w__1719 ,w__1305 ,w__1455);
  xnor g__2022(w__1718 ,w__1235 ,w__1460);
  xnor g__2023(w__1717 ,w__1222 ,w__1452);
  xnor g__2024(w__1715 ,w__1226 ,w__1450);
  xnor g__2025(w__1714 ,w__1428 ,w__1449);
  xnor g__2026(w__1713 ,w__1334 ,w__1448);
  xnor g__2027(w__1712 ,w__1303 ,w__1442);
  xnor g__2028(w__1711 ,w__1293 ,w__1447);
  xnor g__2029(w__1710 ,w__1294 ,w__1446);
  xnor g__2030(w__1709 ,w__1373 ,w__1444);
  or g__2031(w__1708 ,w__1467 ,w__1615);
  xnor g__2032(w__1707 ,w__1424 ,w__1441);
  xnor g__2033(w__1706 ,w__1324 ,w__1443);
  xnor g__2034(w__1705 ,w__1374 ,w__1458);
  xnor g__2035(w__1704 ,w__1084 ,w__1440);
  xnor g__2036(w__1702 ,w__972 ,w__1459);
  xnor g__2037(w__1700 ,w__1236 ,w__1456);
  xnor g__2038(w__1698 ,w__1309 ,w__1451);
  or g__2039(w__1697 ,w__1514 ,w__1623);
  not g__2040(w__1683 ,w__1682);
  not g__2041(w__1680 ,w__1679);
  not g__2042(w__1676 ,w__1677);
  and g__2043(w__1670 ,w__1543 ,w__1497);
  and g__2044(w__1669 ,w__1569 ,w__1507);
  and g__2045(w__1668 ,w__1414 ,w__1496);
  or g__2046(w__1667 ,w__1307 ,w__1565);
  or g__2047(w__1666 ,w__1406 ,w__1478);
  nor g__2048(w__1665 ,w__1304 ,w__1562);
  nor g__2049(w__1664 ,w__1414 ,w__1496);
  and g__2050(w__1663 ,w__1476 ,w__1469);
  or g__2051(w__1662 ,w__1359 ,w__1472);
  nor g__2052(w__1661 ,w__1358 ,w__1473);
  nor g__2053(w__1660 ,w__1476 ,w__1469);
  and g__2054(w__1659 ,w__1560 ,w__1504);
  and g__2055(w__1658 ,w__1406 ,w__1478);
  nor g__2056(w__1657 ,w__1332 ,w__1490);
  or g__2057(w__1656 ,w__1436 ,w__1558);
  and g__2058(w__1655 ,w__1348 ,w__1489);
  and g__2059(w__1654 ,w__1555 ,w__1503);
  or g__2060(w__1653 ,w__1438 ,w__1522);
  and g__2061(w__1652 ,w__1352 ,w__1480);
  or g__2062(w__1651 ,w__1295 ,w__1551);
  nor g__2063(w__1650 ,w__1352 ,w__1480);
  and g__2064(w__1649 ,w__1361 ,w__1479);
  and g__2065(w__1648 ,w__1350 ,w__1477);
  nor g__2066(w__1647 ,w__1430 ,w__1549);
  nor g__2067(w__1646 ,w__1335 ,w__1493);
  and g__2068(w__1645 ,w__1547 ,w__1498);
  and g__2069(w__1644 ,w__1508 ,w__1570);
  or g__2070(w__1643 ,w__1346 ,w__1470);
  nor g__2071(w__1642 ,w__1350 ,w__1477);
  or g__2072(w__1641 ,w__1301 ,w__1541);
  nor g__2073(w__1640 ,w__1345 ,w__1471);
  and g__2074(w__1639 ,w__1571 ,w__1509);
  and g__2075(w__1638 ,w__1332 ,w__1490);
  nor g__2076(w__1637 ,w__1331 ,w__1488);
  and g__2077(w__1636 ,w__1340 ,w__1495);
  nor g__2078(w__1635 ,w__1340 ,w__1495);
  or g__2079(w__1634 ,w__1427 ,w__1532);
  and g__2080(w__1633 ,w__1574 ,w__1568);
  nor g__2081(w__1632 ,w__1348 ,w__1489);
  or g__2082(w__1631 ,w__9 ,w__1492);
  nor g__2083(w__1630 ,w__1302 ,w__1529);
  or g__2084(w__1685 ,w__1378 ,w__1531);
  and g__2085(w__1684 ,w__1385 ,w__1537);
  or g__2086(w__1682 ,w__1383 ,w__1536);
  or g__2087(w__1681 ,w__1396 ,w__1557);
  or g__2088(w__1679 ,w__1402 ,w__1546);
  or g__2089(w__1678 ,w__1394 ,w__1552);
  or g__2090(w__1677 ,w__1380 ,w__1466);
  or g__2091(w__1675 ,w__1397 ,w__1554);
  or g__2092(w__1674 ,w__1398 ,w__1520);
  or g__2093(w__1673 ,w__1388 ,w__1519);
  or g__2094(w__1672 ,w__1391 ,w__1515);
  or g__2095(w__1671 ,w__1389 ,w__1566);
  or g__2096(w__1626 ,w__1297 ,w__1518);
  and g__2097(w__1625 ,w__1331 ,w__1488);
  nor g__2098(w__1624 ,w__1482 ,w__1474);
  nor g__2099(w__1623 ,w__1376 ,w__1513);
  nor g__2100(w__1622 ,w__1372 ,w__1511);
  nor g__2101(w__1621 ,w__1368 ,w__1517);
  and g__2102(w__1620 ,w__1057 ,w__1499);
  nor g__2103(w__1619 ,w__1361 ,w__1479);
  and g__2104(w__1618 ,w__1510 ,w__1523);
  and g__2105(w__1617 ,w__1463 ,w__1502);
  and g__2106(w__1616 ,w__1505 ,w__1462);
  nor g__2107(w__1615 ,w__1291 ,w__1464);
  and g__2108(w__1614 ,w__1500 ,w__1468);
  or g__2109(w__1613 ,w__1481 ,w__1475);
  xnor g__2110(w__1612 ,w__1215 ,w__1367);
  xor g__2111(w__1611 ,w__1369 ,w__1331);
  or g__2112(w__1610 ,w__1314 ,w__1538);
  xnor g__2113(w__1609 ,w__1416 ,w__1366);
  xnor g__2114(w__1608 ,w__1217 ,w__1325);
  xnor g__2115(w__1607 ,w__1426 ,w__1346);
  xnor g__2116(w__1606 ,w__1438 ,w__1418);
  xor g__2117(w__1605 ,w__1370 ,w__1361);
  xnor g__2118(w__1604 ,w__1318 ,w__1323);
  xnor g__2119(w__1603 ,w__1281 ,w__1404);
  xnor g__2120(w__1602 ,w__1363 ,w__1362);
  xnor g__2121(w__1601 ,w__1413 ,w__1327);
  xnor g__2122(w__1600 ,w__1359 ,w__1298);
  xnor g__2123(w__1599 ,w__1319 ,w__1322);
  xor g__2124(w__1598 ,w__1304 ,w__1405);
  xnor g__2125(w__1597 ,w__1357 ,w__1407);
  xor g__2126(w__1596 ,w__1436 ,w__1283);
  xor g__2127(w__1595 ,w__1295 ,w__1409);
  xnor g__2128(w__1594 ,w__1354 ,w__1353);
  xnor g__2129(w__1593 ,w__1349 ,w__1410);
  xor g__2130(w__1592 ,w__1430 ,w__1284);
  xnor g__2131(w__1591 ,w__1347 ,w__1411);
  xor g__2132(w__1590 ,w__1352 ,w__1434);
  xor g__2133(w__1589 ,w__1301 ,w__1422);
  xnor g__2134(w__1588 ,w__1290 ,w__1431);
  xnor g__2135(w__1587 ,w__1420 ,w__1336);
  xnor g__2136(w__1586 ,w__1342 ,w__1341);
  xor g__2137(w__1585 ,w__1340 ,w__1429);
  xor g__2138(w__1584 ,w__1427 ,w__1277);
  xor g__2139(w__1583 ,w__1425 ,w__1350);
  xnor g__2140(w__1582 ,w__1412 ,w__1333);
  xor g__2141(w__1581 ,w__1437 ,w__1332);
  xnor g__2142(w__1580 ,w__1375 ,w__1330);
  xnor g__2143(w__1579 ,w__1419 ,w__1339);
  xnor g__2144(w__1578 ,w__1371 ,w__1326);
  xor g__2145(w__1577 ,w__1435 ,w__1348);
  xnor g__2146(w__1629 ,w__1308 ,w__1310);
  or g__2147(w__1628 ,w__1313 ,w__1465);
  or g__2148(w__1627 ,w__1312 ,w__1461);
  not g__2149(w__1576 ,w__1575);
  not g__2150(w__1572 ,w__1573);
  or g__2151(w__1571 ,w__1342 ,w__1341);
  or g__2152(w__1570 ,w__1319 ,w__1322);
  or g__2153(w__1569 ,w__1363 ,w__1362);
  or g__2154(w__1568 ,w__1412 ,w__1333);
  or g__2155(w__1567 ,w__1280 ,w__1403);
  and g__2156(w__1566 ,w__1305 ,w__1399);
  nor g__2157(w__1565 ,w__1281 ,w__1404);
  and g__2158(w__1564 ,w__1319 ,w__1322);
  and g__2159(w__1563 ,w__1405 ,w__1360);
  nor g__2160(w__1562 ,w__1405 ,w__1360);
  and g__2161(w__1561 ,w__1357 ,w__1407);
  or g__2162(w__1560 ,w__1357 ,w__1407);
  or g__2163(w__1559 ,w__1282 ,w__1355);
  nor g__2164(w__1558 ,w__1283 ,w__1356);
  nor g__2165(w__1557 ,w__1292 ,w__1393);
  and g__2166(w__1556 ,w__1354 ,w__1353);
  or g__2167(w__1555 ,w__1354 ,w__1353);
  and g__2168(w__1554 ,w__1395 ,w__1428);
  or g__2169(w__1553 ,w__1285 ,w__1408);
  and g__2170(w__1552 ,w__1309 ,w__1392);
  nor g__2171(w__1551 ,w__1286 ,w__1409);
  and g__2172(w__1550 ,w__1284 ,w__1351);
  nor g__2173(w__1549 ,w__1284 ,w__1351);
  and g__2174(w__1548 ,w__1349 ,w__1410);
  or g__2175(w__1547 ,w__1349 ,w__1410);
  nor g__2176(w__1546 ,w__1299 ,w__1386);
  and g__2177(w__1545 ,w__1215 ,w__1328);
  and g__2178(w__1544 ,w__1347 ,w__1411);
  or g__2179(w__1543 ,w__1347 ,w__1411);
  or g__2180(w__1542 ,w__1421 ,w__1343);
  nor g__2181(w__1541 ,w__1422 ,w__1344);
  and g__2182(w__1540 ,w__1342 ,w__1341);
  and g__2183(w__1539 ,w__1363 ,w__1362);
  and g__2184(w__1538 ,w__1293 ,w__1316);
  or g__2185(w__1537 ,w__1382 ,w__1432);
  and g__2186(w__1536 ,w__1294 ,w__1379);
  and g__2187(w__1535 ,w__1419 ,w__1339);
  or g__2188(w__1534 ,w__1276 ,w__1337);
  or g__2189(w__1533 ,w__1419 ,w__1339);
  nor g__2190(w__1532 ,w__1277 ,w__1338);
  and g__2191(w__1531 ,w__1303 ,w__1377);
  and g__2192(w__1530 ,w__1168 ,w__1334);
  nor g__2193(w__1529 ,w__1168 ,w__1334);
  and g__2194(w__1528 ,w__1412 ,w__1333);
  and g__2195(w__1527 ,w__1318 ,w__1323);
  and g__2196(w__1526 ,w__1217 ,w__1325);
  or g__2197(w__1525 ,w__1320 ,w__1417);
  and g__2198(w__1524 ,w__1413 ,w__1327);
  or g__2199(w__1523 ,w__1420 ,w__1336);
  nor g__2200(w__1522 ,w__1321 ,w__1418);
  or g__2201(w__1521 ,w__1415 ,w__1366);
  and g__2202(w__1520 ,w__1387 ,w__1433);
  and g__2203(w__1519 ,w__1400 ,w__1374);
  nor g__2204(w__1518 ,w__1416 ,w__1365);
  nor g__2205(w__1517 ,w__1215 ,w__1328);
  and g__2206(w__1516 ,w__1420 ,w__1336);
  and g__2207(w__1515 ,w__1401 ,w__1424);
  and g__2208(w__1514 ,w__1330 ,w__1364);
  nor g__2209(w__1513 ,w__1330 ,w__1364);
  and g__2210(w__1512 ,w__1326 ,w__1329);
  nor g__2211(w__1511 ,w__1326 ,w__1329);
  or g__2212(w__1574 ,w__1241 ,w__1384);
  or g__2213(w__1573 ,w__1238 ,w__1381);
  not g__2214(w__1492 ,w__1493);
  not g__2215(w__1485 ,w__1486);
  not g__2216(w__1483 ,w__1484);
  not g__2217(w__1482 ,w__1481);
  not g__2218(w__1474 ,w__1475);
  not g__2219(w__1472 ,w__1473);
  not g__2220(w__1470 ,w__1471);
  or g__2221(w__1468 ,w__1318 ,w__1323);
  and g__2222(w__1467 ,w__1216 ,w__1324);
  and g__2223(w__1466 ,w__1373 ,w__1390);
  and g__2224(w__1465 ,w__1236 ,w__1315);
  nor g__2225(w__1464 ,w__1216 ,w__1324);
  or g__2226(w__1463 ,w__1217 ,w__1325);
  or g__2227(w__1462 ,w__1413 ,w__1327);
  and g__2228(w__1461 ,w__1235 ,w__1317);
  xnor g__2229(w__1460 ,w__967 ,w__1221);
  xnor g__2230(w__1458 ,w__1288 ,w__1230);
  xnor g__2231(w__1457 ,w__615 ,w__1202);
  xnor g__2232(w__1456 ,w__976 ,w__1225);
  xnor g__2233(w__1455 ,w__968 ,w__1220);
  xnor g__2234(w__1454 ,w__897 ,w__1204);
  xnor g__2235(w__1453 ,w__1163 ,w__1219);
  xnor g__2236(w__1452 ,w__973 ,w__1292);
  xnor g__2237(w__1451 ,w__1165 ,w__1232);
  xnor g__2238(w__1450 ,w__1299 ,w__1164);
  xnor g__2239(w__1449 ,w__982 ,w__1224);
  xor g__2240(w__1448 ,w__1302 ,w__1168);
  xnor g__2241(w__1447 ,w__1081 ,w__1218);
  xnor g__2242(w__1446 ,w__970 ,w__1228);
  xnor g__2243(w__1445 ,w__895 ,w__1188);
  xnor g__2244(w__1444 ,w__1167 ,w__1231);
  xor g__2245(w__1443 ,w__1291 ,w__1216);
  xnor g__2246(w__1442 ,w__1166 ,w__1233);
  xnor g__2247(w__1441 ,w__835 ,w__1234);
  xnor g__2248(w__1440 ,w__856 ,w__1300);
  xnor g__2249(w__1510 ,w__657 ,w__1189);
  xnor g__2250(w__1509 ,w__821 ,w__1187);
  xnor g__2251(w__1508 ,w__882 ,w__1184);
  xnor g__2252(w__1507 ,w__875 ,w__1182);
  xor g__2253(w__1506 ,w__766 ,w__1180);
  xnor g__2254(w__1505 ,w__871 ,w__1203);
  xnor g__2255(w__1504 ,w__983 ,w__1175);
  xnor g__2256(w__1503 ,w__791 ,w__1174);
  xnor g__2257(w__1502 ,w__877 ,w__1205);
  xnor g__2258(w__1501 ,w__828 ,w__1183);
  xnor g__2259(w__1500 ,w__887 ,w__1206);
  xnor g__2260(w__1498 ,w__797 ,w__1171);
  xnor g__2261(w__1497 ,w__808 ,w__1170);
  xnor g__2262(w__1496 ,w__888 ,w__1181);
  xnor g__2263(w__1495 ,w__842 ,w__1191);
  xnor g__2264(w__1494 ,w__824 ,w__1200);
  xnor g__2265(w__1493 ,w__735 ,w__1193);
  xnor g__2266(w__1491 ,w__980 ,w__1194);
  xnor g__2267(w__1490 ,w__864 ,w__1198);
  xnor g__2268(w__1489 ,w__719 ,w__1192);
  xnor g__2269(w__1488 ,w__845 ,w__1196);
  xnor g__2270(w__1487 ,w__833 ,w__1186);
  xnor g__2271(w__1486 ,w__848 ,w__1195);
  xnor g__2272(w__1484 ,w__874 ,w__1199);
  xnor g__2273(w__1481 ,w__841 ,w__1185);
  xnor g__2274(w__1480 ,w__978 ,w__1173);
  xnor g__2275(w__1479 ,w__1002 ,w__1197);
  xnor g__2276(w__1478 ,w__738 ,w__1176);
  xnor g__2277(w__1477 ,w__993 ,w__1172);
  xnor g__2278(w__1476 ,w__643 ,w__1179);
  xnor g__2279(w__1475 ,w__831 ,w__1190);
  xnor g__2280(w__1473 ,w__990 ,w__1178);
  xnor g__2281(w__1471 ,w__799 ,w__1169);
  xnor g__2282(w__1469 ,w__878 ,w__1177);
  not g__2283(w__1432 ,w__1431);
  not g__2284(w__1421 ,w__1422);
  not g__2285(w__1417 ,w__1418);
  not g__2286(w__1415 ,w__1416);
  not g__2287(w__1408 ,w__1409);
  not g__2288(w__1403 ,w__1404);
  nor g__2289(w__1402 ,w__1164 ,w__1227);
  or g__2290(w__1401 ,w__835 ,w__1234);
  or g__2291(w__1400 ,w__1288 ,w__1229);
  or g__2292(w__1399 ,w__968 ,w__1220);
  and g__2293(w__1398 ,w__1163 ,w__1219);
  nor g__2294(w__1397 ,w__982 ,w__1223);
  and g__2295(w__1396 ,w__973 ,w__1222);
  or g__2296(w__1395 ,w__981 ,w__1224);
  and g__2297(w__1394 ,w__1165 ,w__1232);
  nor g__2298(w__1393 ,w__973 ,w__1222);
  or g__2299(w__1392 ,w__1165 ,w__1232);
  and g__2300(w__1391 ,w__835 ,w__1234);
  or g__2301(w__1390 ,w__1167 ,w__1231);
  and g__2302(w__1389 ,w__968 ,w__1220);
  nor g__2303(w__1388 ,w__1287 ,w__1230);
  or g__2304(w__1387 ,w__1163 ,w__1219);
  and g__2305(w__1386 ,w__1164 ,w__1227);
  or g__2306(w__1385 ,w__1289 ,w__1278);
  and g__2307(w__1384 ,w__1300 ,w__1256);
  and g__2308(w__1383 ,w__970 ,w__1228);
  nor g__2309(w__1382 ,w__1290 ,w__1279);
  and g__2310(w__1381 ,w__1308 ,w__1209);
  and g__2311(w__1380 ,w__1167 ,w__1231);
  or g__2312(w__1379 ,w__970 ,w__1228);
  and g__2313(w__1378 ,w__1166 ,w__1233);
  or g__2314(w__1377 ,w__1166 ,w__1233);
  and g__2315(w__1439 ,w__1146 ,w__1266);
  and g__2316(w__1438 ,w__1108 ,w__1261);
  and g__2317(w__1437 ,w__1070 ,w__1259);
  and g__2318(w__1436 ,w__1138 ,w__1263);
  and g__2319(w__1435 ,w__1142 ,w__1245);
  and g__2320(w__1434 ,w__1129 ,w__1253);
  or g__2321(w__1433 ,w__1130 ,w__1254);
  or g__2322(w__1431 ,w__1102 ,w__1237);
  and g__2323(w__1430 ,w__1122 ,w__1250);
  and g__2324(w__1429 ,w__1099 ,w__1239);
  or g__2325(w__1428 ,w__1134 ,w__1255);
  and g__2326(w__1427 ,w__1093 ,w__1252);
  and g__2327(w__1426 ,w__1059 ,w__1242);
  and g__2328(w__1425 ,w__1118 ,w__1247);
  or g__2329(w__1424 ,w__1071 ,w__1271);
  and g__2330(w__1423 ,w__1088 ,w__1251);
  or g__2331(w__1422 ,w__1111 ,w__1244);
  or g__2332(w__1420 ,w__1089 ,w__1243);
  or g__2333(w__1419 ,w__1098 ,w__1240);
  or g__2334(w__1418 ,w__1061 ,w__1257);
  or g__2335(w__1416 ,w__1105 ,w__1264);
  or g__2336(w__1414 ,w__1124 ,w__1272);
  or g__2337(w__1413 ,w__1162 ,w__1262);
  or g__2338(w__1412 ,w__1092 ,w__1248);
  or g__2339(w__1411 ,w__1115 ,w__1246);
  or g__2340(w__1410 ,w__1119 ,w__1249);
  or g__2341(w__1409 ,w__1132 ,w__1258);
  or g__2342(w__1407 ,w__1143 ,w__1265);
  or g__2343(w__1406 ,w__1150 ,w__1268);
  or g__2344(w__1405 ,w__1153 ,w__1270);
  or g__2345(w__1404 ,w__1160 ,w__1274);
  not g__2346(w__1376 ,w__1375);
  not g__2347(w__1372 ,w__1371);
  not g__2348(w__1368 ,w__1367);
  not g__2349(w__1365 ,w__1366);
  not g__2350(w__1359 ,w__1358);
  not g__2351(w__1355 ,w__1356);
  not g__2352(w__1346 ,w__1345);
  not g__2353(w__1343 ,w__1344);
  not g__2354(w__1337 ,w__1338);
  not g__2355(w__1321 ,w__1320);
  or g__2356(w__1317 ,w__967 ,w__1221);
  or g__2357(w__1316 ,w__1081 ,w__1218);
  or g__2358(w__1315 ,w__976 ,w__1225);
  and g__2359(w__1314 ,w__1081 ,w__1218);
  and g__2360(w__1313 ,w__976 ,w__1225);
  and g__2361(w__1312 ,w__967 ,w__1221);
  or g__2362(w__1311 ,w__1048 ,w__1210);
  xnor g__2363(w__1310 ,w__839 ,w__1082);
  or g__2364(w__1375 ,w__1062 ,w__1275);
  or g__2365(w__1374 ,w__1073 ,w__1267);
  or g__2366(w__1373 ,w__1080 ,w__1260);
  and g__2367(w__1370 ,w__1140 ,w__1213);
  and g__2368(w__1369 ,w__1065 ,w__1273);
  or g__2369(w__1367 ,w__1058 ,w__1212);
  xnor g__2370(w__1366 ,w__750 ,w__1039);
  or g__2371(w__1364 ,w__1077 ,w__1269);
  xnor g__2372(w__1363 ,w__640 ,w__1038);
  xnor g__2373(w__1362 ,w__859 ,w__1037);
  xnor g__2374(w__1361 ,w__858 ,w__1028);
  xnor g__2375(w__1360 ,w__994 ,w__1036);
  xnor g__2376(w__1358 ,w__762 ,w__1035);
  xnor g__2377(w__1357 ,w__754 ,w__1034);
  xnor g__2378(w__1356 ,w__998 ,w__1033);
  xnor g__2379(w__1354 ,w__747 ,w__1032);
  xnor g__2380(w__1353 ,w__969 ,w__1031);
  xnor g__2381(w__1352 ,w__745 ,w__1030);
  xnor g__2382(w__1351 ,w__880 ,w__1029);
  xnor g__2383(w__1350 ,w__634 ,w__1027);
  xnor g__2384(w__1349 ,w__764 ,w__1006);
  xnor g__2385(w__1348 ,w__846 ,w__1023);
  xnor g__2386(w__1347 ,w__711 ,w__1025);
  xnor g__2387(w__1345 ,w__660 ,w__1024);
  xnor g__2388(w__1344 ,w__812 ,w__1005);
  xnor g__2389(w__1342 ,w__716 ,w__1022);
  xnor g__2390(w__1341 ,w__819 ,w__1009);
  xnor g__2391(w__1340 ,w__663 ,w__1020);
  xnor g__2392(w__1339 ,w__684 ,w__1018);
  xnor g__2393(w__1338 ,w__867 ,w__1019);
  xnor g__2394(w__1336 ,w__889 ,w__1013);
  xnor g__2395(w__1335 ,w__818 ,w__1017);
  xnor g__2396(w__1334 ,w__641 ,w__1016);
  xnor g__2397(w__1333 ,w__854 ,w__1021);
  xnor g__2398(w__1332 ,w__860 ,w__1007);
  xnor g__2399(w__1331 ,w__682 ,w__1004);
  xnor g__2400(w__1330 ,w__673 ,w__1015);
  xnor g__2401(w__1329 ,w__820 ,w__1008);
  xnor g__2402(w__1328 ,w__823 ,w__1014);
  xnor g__2403(w__1327 ,w__876 ,w__1010);
  xnor g__2404(w__1325 ,w__748 ,w__1026);
  xnor g__2405(w__1324 ,w__742 ,w__1012);
  xnor g__2406(w__1323 ,w__862 ,w__1040);
  xnor g__2407(w__1322 ,w__826 ,w__1041);
  xnor g__2408(w__1320 ,w__683 ,w__1011);
  or g__2409(w__1319 ,w__1045 ,w__1214);
  or g__2410(w__1318 ,w__1047 ,w__1211);
  not g__2411(w__1307 ,w__1306);
  not g__2412(w__1297 ,w__1296);
  not g__2413(w__1289 ,w__1290);
  not g__2414(w__1287 ,w__1288);
  not g__2415(w__1285 ,w__1286);
  not g__2416(w__1282 ,w__1283);
  not g__2417(w__1280 ,w__1281);
  not g__2418(w__1278 ,w__1279);
  not g__2419(w__1276 ,w__1277);
  nor g__2420(w__1275 ,w__680 ,w__1156);
  nor g__2421(w__1274 ,w__996 ,w__1158);
  or g__2422(w__1273 ,w__761 ,w__1155);
  and g__2423(w__1272 ,w__993 ,w__1154);
  nor g__2424(w__1271 ,w__678 ,w__1064);
  nor g__2425(w__1270 ,w__997 ,w__1151);
  nor g__2426(w__1269 ,w__879 ,w__1063);
  nor g__2427(w__1268 ,w__676 ,w__1148);
  and g__2428(w__1267 ,w__877 ,w__1068);
  or g__2429(w__1266 ,w__1001 ,w__1144);
  nor g__2430(w__1265 ,w__690 ,w__1141);
  and g__2431(w__1264 ,w__874 ,w__1076);
  or g__2432(w__1263 ,w__891 ,w__1137);
  and g__2433(w__1262 ,w__888 ,w__1067);
  or g__2434(w__1261 ,w__992 ,w__1078);
  and g__2435(w__1260 ,w__766 ,w__1136);
  or g__2436(w__1259 ,w__873 ,w__1046);
  nor g__2437(w__1258 ,w__893 ,w__1131);
  and g__2438(w__1257 ,w__868 ,w__1042);
  or g__2439(w__1256 ,w__856 ,w__1083);
  nor g__2440(w__1255 ,w__890 ,w__1125);
  nor g__2441(w__1254 ,w__886 ,w__1127);
  or g__2442(w__1253 ,w__892 ,w__1072);
  or g__2443(w__1252 ,w__881 ,w__1091);
  or g__2444(w__1251 ,w__1003 ,w__1120);
  or g__2445(w__1250 ,w__885 ,w__1121);
  nor g__2446(w__1249 ,w__759 ,w__1117);
  nor g__2447(w__1248 ,w__884 ,w__1107);
  or g__2448(w__1247 ,w__757 ,w__1112);
  nor g__2449(w__1246 ,w__758 ,w__1113);
  or g__2450(w__1245 ,w__872 ,w__1090);
  nor g__2451(w__1244 ,w__995 ,w__1060);
  nor g__2452(w__1243 ,w__767 ,w__1087);
  or g__2453(w__1242 ,w__1000 ,w__1109);
  nor g__2454(w__1241 ,w__855 ,w__1084);
  and g__2455(w__1240 ,w__864 ,w__1094);
  or g__2456(w__1239 ,w__672 ,w__1097);
  and g__2457(w__1238 ,w__839 ,w__1082);
  nor g__2458(w__1237 ,w__863 ,w__1101);
  or g__2459(w__1309 ,w__938 ,w__1114);
  or g__2460(w__1308 ,w__954 ,w__1100);
  or g__2461(w__1306 ,w__961 ,w__1157);
  or g__2462(w__1305 ,w__958 ,w__1152);
  and g__2463(w__1304 ,w__957 ,w__1149);
  or g__2464(w__1303 ,w__913 ,w__1085);
  and g__2465(w__1302 ,w__966 ,w__1086);
  and g__2466(w__1301 ,w__928 ,w__1110);
  or g__2467(w__1300 ,w__911 ,w__1104);
  and g__2468(w__1299 ,w__931 ,w__1116);
  and g__2469(w__1298 ,w__953 ,w__1145);
  or g__2470(w__1296 ,w__907 ,w__1074);
  and g__2471(w__1295 ,w__940 ,w__1128);
  or g__2472(w__1294 ,w__965 ,w__1096);
  or g__2473(w__1293 ,w__903 ,w__1126);
  and g__2474(w__1292 ,w__944 ,w__1135);
  and g__2475(w__1291 ,w__947 ,w__1056);
  or g__2476(w__1290 ,w__909 ,w__1106);
  or g__2477(w__1288 ,w__908 ,w__1075);
  or g__2478(w__1286 ,w__943 ,w__1133);
  or g__2479(w__1284 ,w__936 ,w__1123);
  or g__2480(w__1283 ,w__949 ,w__1139);
  or g__2481(w__1281 ,w__964 ,w__1161);
  or g__2482(w__1279 ,w__922 ,w__1103);
  or g__2483(w__1277 ,w__917 ,w__1095);
  not g__2484(w__1229 ,w__1230);
  not g__2485(w__1227 ,w__1226);
  not g__2486(w__1223 ,w__1224);
  and g__2487(w__1214 ,w__878 ,w__1043);
  or g__2488(w__1213 ,w__883 ,w__1055);
  and g__2489(w__1212 ,w__887 ,w__1049);
  and g__2490(w__1211 ,w__875 ,w__1044);
  nor g__2491(w__1210 ,w__870 ,w__1051);
  or g__2492(w__1209 ,w__839 ,w__1082);
  nor g__2493(w__1208 ,w__866 ,w__1147);
  or g__2494(w__1207 ,w__950 ,w__1052);
  xnor g__2495(w__1206 ,w__814 ,w__827);
  xnor g__2496(w__1205 ,w__829 ,w__843);
  xnor g__2497(w__1204 ,w__616 ,w__778);
  xnor g__2498(w__1203 ,w__752 ,w__811);
  xnor g__2499(w__1202 ,w__619 ,w__779);
  xnor g__2500(w__1201 ,w__865 ,w__12809);
  xor g__2501(w__1200 ,w__879 ,w__825);
  xnor g__2502(w__1199 ,w__630 ,w__849);
  xnor g__2503(w__1198 ,w__636 ,w__857);
  xnor g__2504(w__1197 ,w__668 ,w__804);
  xor g__2505(w__1196 ,w__873 ,w__793);
  xor g__2506(w__1195 ,w__884 ,w__838);
  xor g__2507(w__1194 ,w__881 ,w__806);
  xor g__2508(w__1193 ,w__890 ,w__795);
  xor g__2509(w__1192 ,w__886 ,w__815);
  xor g__2510(w__1191 ,w__863 ,w__816);
  xnor g__2511(w__1190 ,w__868 ,w__789);
  xnor g__2512(w__1189 ,w__805 ,w__869);
  xnor g__2513(w__1188 ,w__126 ,w__780);
  xor g__2514(w__1187 ,w__995 ,w__985);
  xor g__2515(w__1186 ,w__1000 ,w__837);
  xnor g__2516(w__1185 ,w__638 ,w__992);
  xnor g__2517(w__1184 ,w__723 ,w__852);
  xor g__2518(w__1183 ,w__767 ,w__987);
  xnor g__2519(w__1182 ,w__800 ,w__850);
  xnor g__2520(w__1181 ,w__628 ,w__834);
  xnor g__2521(w__1180 ,w__746 ,w__986);
  xnor g__2522(w__1179 ,w__633 ,w__861);
  xor g__2523(w__1178 ,w__996 ,w__991);
  xnor g__2524(w__1177 ,w__629 ,w__796);
  xnor g__2525(w__1176 ,w__717 ,w__894);
  xor g__2526(w__1175 ,w__997 ,w__984);
  xor g__2527(w__1174 ,w__891 ,w__786);
  xor g__2528(w__1173 ,w__1001 ,w__975);
  xnor g__2529(w__1172 ,w__988 ,w__989);
  xor g__2530(w__1171 ,w__893 ,w__794);
  xor g__2531(w__1170 ,w__885 ,w__809);
  xor g__2532(w__1169 ,w__892 ,w__802);
  or g__2533(w__1236 ,w__910 ,w__1050);
  or g__2534(w__1235 ,w__924 ,w__1159);
  xnor g__2535(w__1234 ,w__237 ,w__772);
  xnor g__2536(w__1233 ,w__239 ,w__771);
  xnor g__2537(w__1232 ,w__356 ,w__773);
  xnor g__2538(w__1231 ,w__241 ,w__777);
  xnor g__2539(w__1230 ,w__756 ,w__770);
  xnor g__2540(w__1228 ,w__354 ,w__785);
  xnor g__2541(w__1226 ,w__350 ,w__775);
  xnor g__2542(w__1225 ,w__353 ,w__783);
  xnor g__2543(w__1224 ,w__349 ,w__782);
  xnor g__2544(w__1222 ,w__234 ,w__784);
  xnor g__2545(w__1221 ,w__240 ,w__781);
  xnor g__2546(w__1220 ,w__236 ,w__896);
  xnor g__2547(w__1219 ,w__357 ,w__776);
  xnor g__2548(w__1218 ,w__235 ,w__774);
  or g__2549(w__1217 ,w__900 ,w__1054);
  or g__2550(w__1216 ,w__935 ,w__1053);
  or g__2551(w__1215 ,w__945 ,w__1066);
  and g__2552(w__1162 ,w__628 ,w__834);
  and g__2553(w__1161 ,w__762 ,w__963);
  and g__2554(w__1160 ,w__991 ,w__990);
  nor g__2555(w__1159 ,w__691 ,w__960);
  nor g__2556(w__1158 ,w__991 ,w__990);
  and g__2557(w__1157 ,w__959 ,w__994);
  nor g__2558(w__1156 ,w__714 ,w__820);
  nor g__2559(w__1155 ,w__662 ,w__823);
  or g__2560(w__1154 ,w__988 ,w__989);
  and g__2561(w__1153 ,w__984 ,w__983);
  nor g__2562(w__1152 ,w__769 ,w__956);
  nor g__2563(w__1151 ,w__984 ,w__983);
  and g__2564(w__1150 ,w__666 ,w__846);
  or g__2565(w__1149 ,w__768 ,w__955);
  nor g__2566(w__1148 ,w__666 ,w__846);
  or g__2567(w__1146 ,w__977 ,w__974);
  or g__2568(w__1145 ,w__952 ,w__999);
  nor g__2569(w__1144 ,w__978 ,w__975);
  and g__2570(w__1143 ,w__755 ,w__969);
  or g__2571(w__1142 ,w__751 ,w__810);
  nor g__2572(w__1141 ,w__755 ,w__969);
  or g__2573(w__1140 ,w__722 ,w__851);
  nor g__2574(w__1139 ,w__763 ,w__948);
  or g__2575(w__1138 ,w__6 ,w__790);
  nor g__2576(w__1137 ,w__4 ,w__791);
  or g__2577(w__1136 ,w__746 ,w__986);
  or g__2578(w__1135 ,w__760 ,w__942);
  and g__2579(w__1134 ,w__735 ,w__795);
  and g__2580(w__1133 ,w__941 ,w__880);
  and g__2581(w__1132 ,w__794 ,w__797);
  nor g__2582(w__1131 ,w__794 ,w__797);
  and g__2583(w__1130 ,w__719 ,w__815);
  or g__2584(w__1129 ,w__798 ,w__801);
  or g__2585(w__1128 ,w__765 ,w__937);
  nor g__2586(w__1127 ,w__719 ,w__815);
  and g__2587(w__1126 ,w__951 ,w__894);
  nor g__2588(w__1125 ,w__735 ,w__795);
  and g__2589(w__1124 ,w__988 ,w__989);
  nor g__2590(w__1123 ,w__681 ,w__934);
  or g__2591(w__1122 ,w__8 ,w__807);
  nor g__2592(w__1121 ,w__5 ,w__808);
  nor g__2593(w__1120 ,w__668 ,w__804);
  and g__2594(w__1119 ,w__647 ,w__812);
  or g__2595(w__1118 ,w__725 ,w__817);
  nor g__2596(w__1117 ,w__647 ,w__812);
  or g__2597(w__1116 ,w__685 ,w__930);
  and g__2598(w__1115 ,w__718 ,w__819);
  and g__2599(w__1114 ,w__929 ,w__876);
  nor g__2600(w__1113 ,w__718 ,w__819);
  nor g__2601(w__1112 ,w__724 ,w__818);
  and g__2602(w__1111 ,w__985 ,w__821);
  or g__2603(w__1110 ,w__677 ,w__926);
  nor g__2604(w__1109 ,w__833 ,w__837);
  or g__2605(w__1108 ,w__637 ,w__840);
  nor g__2606(w__1107 ,w__838 ,w__848);
  nor g__2607(w__1106 ,w__689 ,w__923);
  and g__2608(w__1105 ,w__630 ,w__849);
  and g__2609(w__1104 ,w__679 ,w__962);
  and g__2610(w__1103 ,w__921 ,w__867);
  and g__2611(w__1102 ,w__816 ,w__842);
  nor g__2612(w__1101 ,w__816 ,w__842);
  and g__2613(w__1100 ,w__918 ,w__860);
  or g__2614(w__1099 ,w__653 ,w__853);
  and g__2615(w__1098 ,w__636 ,w__857);
  nor g__2616(w__1097 ,w__652 ,w__854);
  and g__2617(w__1096 ,w__916 ,w__858);
  nor g__2618(w__1095 ,w__688 ,w__915);
  or g__2619(w__1094 ,w__636 ,w__857);
  or g__2620(w__1093 ,w__7 ,w__979);
  and g__2621(w__1092 ,w__838 ,w__848);
  nor g__2622(w__1091 ,w__3 ,w__980);
  nor g__2623(w__1090 ,w__752 ,w__811);
  and g__2624(w__1089 ,w__828 ,w__987);
  or g__2625(w__1088 ,w__667 ,w__803);
  nor g__2626(w__1087 ,w__828 ,w__987);
  or g__2627(w__1086 ,w__683 ,w__912);
  and g__2628(w__1085 ,w__682 ,w__904);
  or g__2629(w__1168 ,w__527 ,w__933);
  or g__2630(w__1167 ,w__700 ,w__901);
  or g__2631(w__1166 ,w__704 ,w__914);
  or g__2632(w__1165 ,w__706 ,w__920);
  and g__2633(w__1164 ,w__698 ,w__932);
  or g__2634(w__1163 ,w__709 ,w__939);
  not g__2635(w__1083 ,w__1084);
  and g__2636(w__1080 ,w__746 ,w__986);
  and g__2637(w__1079 ,w__847 ,w__813);
  nor g__2638(w__1078 ,w__638 ,w__841);
  and g__2639(w__1077 ,w__825 ,w__824);
  or g__2640(w__1076 ,w__630 ,w__849);
  nor g__2641(w__1075 ,w__671 ,w__906);
  and g__2642(w__1074 ,w__673 ,w__905);
  and g__2643(w__1073 ,w__829 ,w__843);
  nor g__2644(w__1072 ,w__799 ,w__802);
  and g__2645(w__1071 ,w__712 ,w__826);
  or g__2646(w__1070 ,w__844 ,w__792);
  nor g__2647(w__1069 ,w__971 ,w__787);
  or g__2648(w__1068 ,w__829 ,w__843);
  or g__2649(w__1067 ,w__628 ,w__834);
  nor g__2650(w__1066 ,w__687 ,w__927);
  or g__2651(w__1065 ,w__661 ,w__822);
  nor g__2652(w__1064 ,w__712 ,w__826);
  nor g__2653(w__1063 ,w__825 ,w__824);
  and g__2654(w__1062 ,w__714 ,w__820);
  nor g__2655(w__1061 ,w__830 ,w__789);
  nor g__2656(w__1060 ,w__985 ,w__821);
  or g__2657(w__1059 ,w__832 ,w__836);
  and g__2658(w__1058 ,w__814 ,w__827);
  or g__2659(w__1057 ,w__847 ,w__813);
  or g__2660(w__1056 ,w__675 ,w__919);
  nor g__2661(w__1055 ,w__723 ,w__852);
  and g__2662(w__1054 ,w__899 ,w__862);
  and g__2663(w__1053 ,w__925 ,w__859);
  and g__2664(w__1052 ,w__898 ,w__889);
  nor g__2665(w__1051 ,w__657 ,w__805);
  and g__2666(w__1050 ,w__946 ,w__861);
  or g__2667(w__1049 ,w__814 ,w__827);
  and g__2668(w__1048 ,w__657 ,w__805);
  and g__2669(w__1047 ,w__800 ,w__850);
  nor g__2670(w__1046 ,w__845 ,w__793);
  and g__2671(w__1045 ,w__629 ,w__796);
  or g__2672(w__1044 ,w__800 ,w__850);
  or g__2673(w__1043 ,w__629 ,w__796);
  or g__2674(w__1042 ,w__831 ,w__788);
  xor g__2675(w__1041 ,w__678 ,w__712);
  xnor g__2676(w__1040 ,w__650 ,w__649);
  xnor g__2677(w__1039 ,w__475 ,w__679);
  xnor g__2678(w__1038 ,w__674 ,w__12759);
  xnor g__2679(w__1037 ,w__644 ,w__656);
  xnor g__2680(w__1036 ,w__744 ,w__739);
  xnor g__2681(w__1035 ,w__731 ,w__12884);
  xor g__2682(w__1034 ,w__768 ,w__12883);
  xnor g__2683(w__1033 ,w__730 ,w__727);
  xor g__2684(w__1032 ,w__763 ,w__12882);
  xor g__2685(w__1031 ,w__690 ,w__755);
  xor g__2686(w__1030 ,w__769 ,w__710);
  xnor g__2687(w__1029 ,w__734 ,w__733);
  xnor g__2688(w__1028 ,w__631 ,w__651);
  xor g__2689(w__1027 ,w__691 ,w__635);
  xnor g__2690(w__1026 ,w__670 ,w__12887);
  xor g__2691(w__1025 ,w__681 ,w__12880);
  xor g__2692(w__1024 ,w__760 ,w__741);
  xor g__2693(w__1023 ,w__676 ,w__666);
  xor g__2694(w__1022 ,w__677 ,w__12879);
  xnor g__2695(w__1021 ,w__653 ,w__672);
  xor g__2696(w__1020 ,w__689 ,w__12878);
  xnor g__2697(w__1019 ,w__669 ,w__626);
  xnor g__2698(w__1018 ,w__665 ,w__721);
  xnor g__2699(w__1017 ,w__757 ,w__725);
  xor g__2700(w__1016 ,w__688 ,w__12877);
  xnor g__2701(w__1015 ,w__632 ,w__625);
  xor g__2702(w__1014 ,w__761 ,w__662);
  xnor g__2703(w__1013 ,w__713 ,w__658);
  xnor g__2704(w__1012 ,w__686 ,w__12886);
  xnor g__2705(w__1011 ,w__646 ,w__655);
  xnor g__2706(w__1010 ,w__732 ,w__728);
  xor g__2707(w__1009 ,w__758 ,w__718);
  xor g__2708(w__1008 ,w__680 ,w__714);
  xnor g__2709(w__1007 ,w__743 ,w__627);
  xnor g__2710(w__1006 ,w__737 ,w__12881);
  xor g__2711(w__1005 ,w__759 ,w__647);
  xnor g__2712(w__1004 ,w__642 ,w__648);
  xnor g__2713(w__1084 ,w__692 ,w__618);
  xnor g__2714(w__1082 ,w__477 ,w__617);
  or g__2715(w__1081 ,w__702 ,w__902);
  not g__2716(w__1003 ,w__1002);
  not g__2717(w__999 ,w__998);
  not g__2718(w__982 ,w__981);
  not g__2719(w__979 ,w__980);
  not g__2720(w__977 ,w__978);
  not g__2721(w__974 ,w__975);
  not g__2722(w__971 ,w__972);
  or g__2723(w__966 ,w__645 ,w__654);
  and g__2724(w__965 ,w__631 ,w__651);
  and g__2725(w__964 ,w__12884 ,w__731);
  or g__2726(w__963 ,w__12884 ,w__731);
  or g__2727(w__962 ,w__474 ,w__750);
  and g__2728(w__961 ,w__744 ,w__739);
  nor g__2729(w__960 ,w__634 ,w__635);
  or g__2730(w__959 ,w__744 ,w__739);
  and g__2731(w__958 ,w__710 ,w__745);
  or g__2732(w__957 ,w__19 ,w__753);
  nor g__2733(w__956 ,w__710 ,w__745);
  nor g__2734(w__955 ,w__12883 ,w__754);
  and g__2735(w__954 ,w__743 ,w__627);
  or g__2736(w__953 ,w__729 ,w__726);
  nor g__2737(w__952 ,w__730 ,w__727);
  or g__2738(w__951 ,w__738 ,w__717);
  and g__2739(w__950 ,w__713 ,w__658);
  and g__2740(w__949 ,w__12882 ,w__747);
  nor g__2741(w__948 ,w__12882 ,w__747);
  or g__2742(w__947 ,w__17 ,w__639);
  or g__2743(w__946 ,w__643 ,w__633);
  and g__2744(w__945 ,w__12886 ,w__742);
  or g__2745(w__944 ,w__740 ,w__659);
  and g__2746(w__943 ,w__734 ,w__733);
  nor g__2747(w__942 ,w__741 ,w__660);
  or g__2748(w__941 ,w__734 ,w__733);
  or g__2749(w__940 ,w__78 ,w__736);
  nor g__2750(w__939 ,w__356 ,w__708);
  and g__2751(w__938 ,w__732 ,w__728);
  nor g__2752(w__937 ,w__12881 ,w__737);
  and g__2753(w__936 ,w__12880 ,w__711);
  and g__2754(w__935 ,w__644 ,w__656);
  nor g__2755(w__934 ,w__12880 ,w__711);
  and g__2756(w__933 ,w__557 ,w__692);
  or g__2757(w__932 ,w__242 ,w__707);
  or g__2758(w__931 ,w__664 ,w__720);
  nor g__2759(w__930 ,w__665 ,w__721);
  or g__2760(w__929 ,w__732 ,w__728);
  or g__2761(w__928 ,w__18 ,w__715);
  nor g__2762(w__927 ,w__12886 ,w__742);
  nor g__2763(w__926 ,w__12879 ,w__716);
  or g__2764(w__925 ,w__644 ,w__656);
  and g__2765(w__924 ,w__634 ,w__635);
  nor g__2766(w__923 ,w__12878 ,w__663);
  and g__2767(w__922 ,w__669 ,w__626);
  or g__2768(w__921 ,w__669 ,w__626);
  nor g__2769(w__920 ,w__241 ,w__705);
  nor g__2770(w__919 ,w__12759 ,w__640);
  or g__2771(w__918 ,w__743 ,w__627);
  and g__2772(w__917 ,w__12877 ,w__641);
  or g__2773(w__916 ,w__631 ,w__651);
  nor g__2774(w__915 ,w__12877 ,w__641);
  and g__2775(w__914 ,w__756 ,w__703);
  and g__2776(w__913 ,w__642 ,w__648);
  nor g__2777(w__912 ,w__646 ,w__655);
  nor g__2778(w__911 ,w__475 ,w__749);
  and g__2779(w__910 ,w__643 ,w__633);
  and g__2780(w__909 ,w__12878 ,w__663);
  and g__2781(w__908 ,w__12887 ,w__748);
  and g__2782(w__907 ,w__632 ,w__625);
  nor g__2783(w__906 ,w__12887 ,w__748);
  or g__2784(w__905 ,w__632 ,w__625);
  or g__2785(w__904 ,w__642 ,w__648);
  and g__2786(w__903 ,w__738 ,w__717);
  nor g__2787(w__902 ,w__357 ,w__701);
  nor g__2788(w__901 ,w__240 ,w__699);
  and g__2789(w__900 ,w__650 ,w__649);
  or g__2790(w__899 ,w__650 ,w__649);
  or g__2791(w__898 ,w__713 ,w__658);
  xnor g__2792(w__897 ,w__383 ,w__12934);
  xnor g__2793(w__896 ,w__487 ,w__12956);
  or g__2794(w__895 ,w__506 ,w__621);
  or g__2795(w__1002 ,w__539 ,w__620);
  xor g__2796(w__1001 ,w__445 ,w__12829);
  and g__2797(w__1000 ,w__574 ,w__697);
  xnor g__2798(w__998 ,w__394 ,w__12788);
  xor g__2799(w__997 ,w__457 ,w__12820);
  xor g__2800(w__996 ,w__377 ,w__12695);
  xor g__2801(w__995 ,w__406 ,w__12690);
  xnor g__2802(w__994 ,w__453 ,w__12789);
  xnor g__2803(w__993 ,w__399 ,w__12708);
  and g__2804(w__992 ,w__180 ,w__696);
  xnor g__2805(w__991 ,w__466 ,w__12821);
  xnor g__2806(w__990 ,w__467 ,w__12852);
  xnor g__2807(w__989 ,w__463 ,w__12834);
  xnor g__2808(w__988 ,w__465 ,w__12991);
  xnor g__2809(w__987 ,w__420 ,w__12743);
  xnor g__2810(w__986 ,w__455 ,w__12709);
  xnor g__2811(w__985 ,w__395 ,w__12816);
  xnor g__2812(w__984 ,w__460 ,w__12694);
  xnor g__2813(w__983 ,w__459 ,w__12851);
  or g__2814(w__981 ,w__510 ,w__695);
  xnor g__2815(w__980 ,w__407 ,w__12845);
  xnor g__2816(w__978 ,w__451 ,w__12703);
  or g__2817(w__976 ,w__528 ,w__624);
  xnor g__2818(w__975 ,w__448 ,w__12986);
  or g__2819(w__973 ,w__585 ,w__694);
  xnor g__2820(w__972 ,w__444 ,w__12716);
  or g__2821(w__970 ,w__556 ,w__622);
  xnor g__2822(w__969 ,w__381 ,w__12787);
  or g__2823(w__968 ,w__609 ,w__693);
  or g__2824(w__967 ,w__576 ,w__623);
  not g__2825(w__883 ,w__882);
  not g__2826(w__872 ,w__871);
  not g__2827(w__870 ,w__869);
  not g__2828(w__866 ,w__865);
  not g__2829(w__855 ,w__856);
  not g__2830(w__853 ,w__854);
  not g__2831(w__851 ,w__852);
  not g__2832(w__844 ,w__845);
  not g__2833(w__840 ,w__841);
  not g__2834(w__836 ,w__837);
  not g__2835(w__832 ,w__833);
  not g__2836(w__830 ,w__831);
  not g__2837(w__822 ,w__823);
  not g__2838(w__817 ,w__818);
  not g__2839(w__810 ,w__811);
  not g__2840(w__807 ,w__808);
  not g__2841(w__803 ,w__804);
  not g__2842(w__801 ,w__802);
  not g__2843(w__798 ,w__799);
  not g__2844(w__792 ,w__793);
  not g__2845(w__790 ,w__791);
  not g__2846(w__788 ,w__789);
  xnor g__2847(w__785 ,w__484 ,w__12927);
  xnor g__2848(w__784 ,w__485 ,w__12923);
  xnor g__2849(w__783 ,w__483 ,w__12957);
  xnor g__2850(w__782 ,w__480 ,w__12928);
  xnor g__2851(w__781 ,w__468 ,w__12677);
  xnor g__2852(w__780 ,w__416 ,w__12682);
  xnor g__2853(w__779 ,w__417 ,w__12714);
  xnor g__2854(w__778 ,w__404 ,w__12745);
  xnor g__2855(w__777 ,w__473 ,w__12678);
  xnor g__2856(w__776 ,w__470 ,w__12680);
  xnor g__2857(w__775 ,w__486 ,w__12922);
  xnor g__2858(w__774 ,w__482 ,w__12933);
  xnor g__2859(w__773 ,w__469 ,w__12931);
  xnor g__2860(w__772 ,w__481 ,w__12958);
  xnor g__2861(w__771 ,w__479 ,w__12952);
  xnor g__2862(w__770 ,w__472 ,w__12951);
  xnor g__2863(w__894 ,w__441 ,w__12712);
  xor g__2864(w__893 ,w__427 ,w__12692);
  xor g__2865(w__892 ,w__421 ,w__12985);
  xor g__2866(w__891 ,w__366 ,w__12819);
  xor g__2867(w__890 ,w__426 ,w__12707);
  xnor g__2868(w__889 ,w__380 ,w__12839);
  xnor g__2869(w__888 ,w__384 ,w__12929);
  xnor g__2870(w__887 ,w__450 ,w__12854);
  xor g__2871(w__886 ,w__432 ,w__12994);
  xor g__2872(w__885 ,w__401 ,w__12817);
  xor g__2873(w__884 ,w__379 ,w__12750);
  xnor g__2874(w__882 ,w__392 ,w__12768);
  xor g__2875(w__881 ,w__382 ,w__12814);
  xnor g__2876(w__880 ,w__430 ,w__12786);
  xor g__2877(w__879 ,w__410 ,w__12715);
  xnor g__2878(w__878 ,w__443 ,w__12767);
  xnor g__2879(w__877 ,w__374 ,w__12855);
  xnor g__2880(w__876 ,w__409 ,w__12710);
  xnor g__2881(w__875 ,w__436 ,w__12948);
  xnor g__2882(w__874 ,w__464 ,w__12842);
  xor g__2883(w__873 ,w__423 ,w__12793);
  xnor g__2884(w__871 ,w__390 ,w__12930);
  xnor g__2885(w__869 ,w__454 ,w__12996);
  xnor g__2886(w__868 ,w__373 ,w__12938);
  xnor g__2887(w__867 ,w__415 ,w__12783);
  xnor g__2888(w__864 ,w__385 ,w__12763);
  xor g__2889(w__863 ,w__449 ,w__12689);
  xnor g__2890(w__862 ,w__452 ,w__12791);
  xnor g__2891(w__861 ,w__447 ,w__12798);
  xnor g__2892(w__860 ,w__361 ,w__12794);
  xnor g__2893(w__859 ,w__400 ,w__12979);
  xnor g__2894(w__858 ,w__458 ,w__12800);
  xnor g__2895(w__857 ,w__387 ,w__12826);
  xnor g__2896(w__856 ,w__456 ,w__12781);
  xnor g__2897(w__854 ,w__365 ,w__12782);
  xnor g__2898(w__852 ,w__371 ,w__12831);
  xnor g__2899(w__850 ,w__368 ,w__12853);
  xnor g__2900(w__849 ,w__375 ,w__12874);
  xnor g__2901(w__848 ,w__402 ,w__12907);
  xnor g__2902(w__847 ,w__364 ,w__12998);
  xnor g__2903(w__846 ,w__433 ,w__12837);
  xnor g__2904(w__845 ,w__461 ,w__12762);
  xnor g__2905(w__843 ,w__403 ,w__12698);
  xnor g__2906(w__842 ,w__389 ,w__12846);
  xnor g__2907(w__841 ,w__488 ,w__12654);
  xnor g__2908(w__839 ,w__396 ,w__12701);
  xnor g__2909(w__838 ,w__372 ,w__12687);
  xnor g__2910(w__837 ,w__413 ,w__12827);
  xnor g__2911(w__835 ,w__358 ,w__12769);
  xnor g__2912(w__834 ,w__398 ,w__12740);
  xnor g__2913(w__833 ,w__369 ,w__12984);
  xnor g__2914(w__831 ,w__446 ,w__12969);
  xnor g__2915(w__829 ,w__442 ,w__12824);
  xnor g__2916(w__828 ,w__397 ,w__12932);
  xnor g__2917(w__827 ,w__376 ,w__12697);
  xnor g__2918(w__826 ,w__367 ,w__12799);
  xnor g__2919(w__825 ,w__435 ,w__12684);
  xnor g__2920(w__824 ,w__405 ,w__12652);
  xnor g__2921(w__823 ,w__362 ,w__12792);
  xnor g__2922(w__821 ,w__462 ,w__12847);
  xnor g__2923(w__820 ,w__363 ,w__12747);
  xnor g__2924(w__819 ,w__360 ,w__12784);
  xnor g__2925(w__818 ,w__386 ,w__12833);
  xnor g__2926(w__816 ,w__429 ,w__12815);
  xnor g__2927(w__815 ,w__437 ,w__12711);
  xnor g__2928(w__814 ,w__412 ,w__12823);
  xnor g__2929(w__813 ,w__393 ,w__12872);
  xnor g__2930(w__812 ,w__414 ,w__12785);
  xnor g__2931(w__811 ,w__370 ,w__12741);
  xnor g__2932(w__809 ,w__408 ,w__12691);
  xnor g__2933(w__808 ,w__425 ,w__12848);
  xnor g__2934(w__806 ,w__411 ,w__12688);
  xnor g__2935(w__805 ,w__388 ,w__12713);
  xnor g__2936(w__804 ,w__378 ,w__12832);
  xnor g__2937(w__802 ,w__424 ,w__12828);
  xnor g__2938(w__800 ,w__391 ,w__12696);
  xnor g__2939(w__799 ,w__439 ,w__12702);
  xnor g__2940(w__797 ,w__422 ,w__12849);
  xnor g__2941(w__796 ,w__440 ,w__12830);
  xnor g__2942(w__795 ,w__419 ,w__12990);
  xnor g__2943(w__794 ,w__428 ,w__12818);
  xnor g__2944(w__793 ,w__418 ,w__12825);
  xnor g__2945(w__791 ,w__438 ,w__12850);
  xnor g__2946(w__789 ,w__355 ,w__359);
  xnor g__2947(w__787 ,w__478 ,w__434);
  xnor g__2948(w__786 ,w__431 ,w__12693);
  not g__2949(w__765 ,w__764);
  not g__2950(w__753 ,w__754);
  not g__2951(w__751 ,w__752);
  not g__2952(w__749 ,w__750);
  not g__2953(w__740 ,w__741);
  not g__2954(w__736 ,w__737);
  not g__2955(w__729 ,w__730);
  not g__2956(w__726 ,w__727);
  not g__2957(w__725 ,w__724);
  not g__2958(w__722 ,w__723);
  not g__2959(w__720 ,w__721);
  not g__2960(w__715 ,w__716);
  nor g__2961(w__709 ,w__75 ,w__469);
  and g__2962(w__708 ,w__75 ,w__469);
  nor g__2963(w__707 ,w__12921 ,w__476);
  nor g__2964(w__706 ,w__43 ,w__473);
  and g__2965(w__705 ,w__43 ,w__473);
  nor g__2966(w__704 ,w__21 ,w__472);
  or g__2967(w__703 ,w__12951 ,w__471);
  nor g__2968(w__702 ,w__83 ,w__470);
  and g__2969(w__701 ,w__83 ,w__470);
  nor g__2970(w__700 ,w__73 ,w__468);
  and g__2971(w__699 ,w__73 ,w__468);
  or g__2972(w__698 ,w__89 ,w__477);
  or g__2973(w__697 ,w__560 ,w__479);
  or g__2974(w__696 ,w__276 ,w__478);
  nor g__2975(w__695 ,w__520 ,w__484);
  nor g__2976(w__694 ,w__540 ,w__486);
  nor g__2977(w__693 ,w__607 ,w__485);
  and g__2978(w__769 ,w__255 ,w__601);
  and g__2979(w__768 ,w__190 ,w__598);
  and g__2980(w__767 ,w__343 ,w__613);
  or g__2981(w__766 ,w__348 ,w__499);
  or g__2982(w__764 ,w__340 ,w__579);
  and g__2983(w__763 ,w__136 ,w__586);
  or g__2984(w__762 ,w__338 ,w__611);
  and g__2985(w__761 ,w__146 ,w__534);
  and g__2986(w__760 ,w__337 ,w__583);
  and g__2987(w__759 ,w__347 ,w__522);
  and g__2988(w__758 ,w__191 ,w__566);
  and g__2989(w__757 ,w__216 ,w__545);
  or g__2990(w__756 ,w__315 ,w__494);
  or g__2991(w__755 ,w__318 ,w__591);
  or g__2992(w__754 ,w__138 ,w__600);
  or g__2993(w__752 ,w__174 ,w__584);
  or g__2994(w__750 ,w__291 ,w__614);
  or g__2995(w__748 ,w__127 ,w__516);
  or g__2996(w__747 ,w__285 ,w__588);
  or g__2997(w__746 ,w__345 ,w__605);
  or g__2998(w__745 ,w__162 ,w__526);
  or g__2999(w__744 ,w__170 ,w__610);
  or g__3000(w__743 ,w__196 ,w__587);
  or g__3001(w__742 ,w__323 ,w__525);
  or g__3002(w__741 ,w__269 ,w__536);
  or g__3003(w__739 ,w__332 ,w__608);
  or g__3004(w__738 ,w__258 ,w__593);
  or g__3005(w__737 ,w__260 ,w__580);
  or g__3006(w__735 ,w__327 ,w__563);
  or g__3007(w__734 ,w__286 ,w__582);
  or g__3008(w__733 ,w__297 ,w__581);
  or g__3009(w__732 ,w__252 ,w__537);
  or g__3010(w__731 ,w__311 ,w__612);
  or g__3011(w__730 ,w__344 ,w__594);
  or g__3012(w__728 ,w__163 ,w__570);
  or g__3013(w__727 ,w__307 ,w__564);
  or g__3014(w__724 ,w__176 ,w__572);
  or g__3015(w__723 ,w__204 ,w__515);
  or g__3016(w__721 ,w__222 ,w__568);
  or g__3017(w__719 ,w__248 ,w__553);
  or g__3018(w__718 ,w__182 ,w__565);
  or g__3019(w__717 ,w__278 ,w__596);
  or g__3020(w__716 ,w__141 ,w__546);
  or g__3021(w__713 ,w__230 ,w__491);
  or g__3022(w__712 ,w__342 ,w__595);
  or g__3023(w__711 ,w__201 ,w__577);
  or g__3024(w__710 ,w__300 ,w__604);
  not g__3025(w__687 ,w__686);
  not g__3026(w__685 ,w__684);
  not g__3027(w__675 ,w__674);
  not g__3028(w__671 ,w__670);
  not g__3029(w__667 ,w__668);
  not g__3030(w__664 ,w__665);
  not g__3031(w__661 ,w__662);
  not g__3032(w__659 ,w__660);
  not g__3033(w__654 ,w__655);
  not g__3034(w__653 ,w__652);
  not g__3035(w__645 ,w__646);
  not g__3036(w__639 ,w__640);
  not g__3037(w__637 ,w__638);
  nor g__3038(w__624 ,w__514 ,w__487);
  nor g__3039(w__623 ,w__501 ,w__480);
  nor g__3040(w__622 ,w__606 ,w__481);
  nor g__3041(w__621 ,w__530 ,w__482);
  nor g__3042(w__620 ,w__590 ,w__483);
  or g__3043(w__619 ,w__275 ,w__507);
  xnor g__3044(w__618 ,w__352 ,w__12655);
  xnor g__3045(w__617 ,w__242 ,w__12921);
  or g__3046(w__616 ,w__339 ,w__513);
  or g__3047(w__615 ,w__132 ,w__504);
  or g__3048(w__692 ,w__200 ,w__544);
  and g__3049(w__691 ,w__264 ,w__492);
  and g__3050(w__690 ,w__321 ,w__589);
  and g__3051(w__689 ,w__229 ,w__552);
  and g__3052(w__688 ,w__173 ,w__602);
  or g__3053(w__686 ,w__217 ,w__512);
  or g__3054(w__684 ,w__158 ,w__567);
  and g__3055(w__683 ,w__147 ,w__489);
  or g__3056(w__682 ,w__202 ,w__517);
  and g__3057(w__681 ,w__326 ,w__569);
  and g__3058(w__680 ,w__254 ,w__518);
  or g__3059(w__679 ,w__143 ,w__538);
  and g__3060(w__678 ,w__292 ,w__495);
  and g__3061(w__677 ,w__166 ,w__561);
  and g__3062(w__676 ,w__233 ,w__603);
  or g__3063(w__674 ,w__129 ,w__533);
  or g__3064(w__673 ,w__140 ,w__490);
  and g__3065(w__672 ,w__329 ,w__549);
  or g__3066(w__670 ,w__301 ,w__496);
  or g__3067(w__669 ,w__295 ,w__555);
  or g__3068(w__668 ,w__279 ,w__541);
  or g__3069(w__666 ,w__296 ,w__599);
  or g__3070(w__665 ,w__310 ,w__571);
  or g__3071(w__663 ,w__157 ,w__558);
  or g__3072(w__662 ,w__302 ,w__592);
  or g__3073(w__660 ,w__193 ,w__575);
  or g__3074(w__658 ,w__265 ,w__531);
  or g__3075(w__657 ,w__189 ,w__559);
  or g__3076(w__656 ,w__268 ,w__498);
  or g__3077(w__655 ,w__181 ,w__508);
  or g__3078(w__652 ,w__160 ,w__551);
  or g__3079(w__651 ,w__284 ,w__550);
  or g__3080(w__650 ,w__220 ,w__523);
  or g__3081(w__649 ,w__197 ,w__597);
  or g__3082(w__648 ,w__188 ,w__542);
  or g__3083(w__647 ,w__212 ,w__573);
  or g__3084(w__646 ,w__346 ,w__543);
  or g__3085(w__644 ,w__317 ,w__505);
  or g__3086(w__643 ,w__294 ,w__497);
  or g__3087(w__642 ,w__149 ,w__524);
  or g__3088(w__641 ,w__224 ,w__547);
  or g__3089(w__640 ,w__156 ,w__521);
  or g__3090(w__638 ,w__214 ,w__535);
  or g__3091(w__636 ,w__309 ,w__548);
  or g__3092(w__635 ,w__251 ,w__500);
  or g__3093(w__634 ,w__205 ,w__578);
  or g__3094(w__633 ,w__130 ,w__502);
  or g__3095(w__632 ,w__178 ,w__529);
  or g__3096(w__631 ,w__303 ,w__511);
  or g__3097(w__630 ,w__324 ,w__532);
  or g__3098(w__629 ,w__128 ,w__493);
  or g__3099(w__628 ,w__304 ,w__509);
  or g__3100(w__627 ,w__246 ,w__562);
  or g__3101(w__626 ,w__261 ,w__554);
  or g__3102(w__625 ,w__263 ,w__503);
  and g__3103(w__614 ,w__12842 ,w__199);
  or g__3104(w__613 ,w__116 ,w__316);
  and g__3105(w__612 ,w__12662 ,w__135);
  and g__3106(w__611 ,w__13009 ,w__322);
  and g__3107(w__610 ,w__12977 ,w__247);
  nor g__3108(w__609 ,w__72 ,w__234);
  and g__3109(w__608 ,w__12946 ,w__331);
  and g__3110(w__607 ,w__72 ,w__234);
  and g__3111(w__606 ,w__12 ,w__237);
  and g__3112(w__605 ,w__12960 ,w__228);
  and g__3113(w__604 ,w__12796 ,w__223);
  or g__3114(w__603 ,w__111 ,w__257);
  or g__3115(w__602 ,w__107 ,w__244);
  or g__3116(w__601 ,w__61 ,w__183);
  and g__3117(w__600 ,w__13008 ,w__221);
  and g__3118(w__599 ,w__12867 ,w__336);
  or g__3119(w__598 ,w__58 ,w__175);
  and g__3120(w__597 ,w__13011 ,w__210);
  and g__3121(w__596 ,w__12963 ,w__288);
  and g__3122(w__595 ,w__12924 ,w__306);
  and g__3123(w__594 ,w__12976 ,w__308);
  and g__3124(w__593 ,w__12774 ,w__250);
  and g__3125(w__592 ,w__12980 ,w__232);
  and g__3126(w__591 ,w__12944 ,w__148);
  and g__3127(w__590 ,w__84 ,w__353);
  or g__3128(w__589 ,w__120 ,w__305);
  and g__3129(w__588 ,w__13007 ,w__177);
  and g__3130(w__587 ,w__12699 ,w__172);
  or g__3131(w__586 ,w__105 ,w__209);
  nor g__3132(w__585 ,w__97 ,w__350);
  and g__3133(w__584 ,w__12866 ,w__341);
  or g__3134(w__583 ,w__110 ,w__281);
  and g__3135(w__582 ,w__12974 ,w__277);
  and g__3136(w__581 ,w__12943 ,w__165);
  and g__3137(w__580 ,w__12659 ,w__159);
  and g__3138(w__579 ,w__13006 ,w__267);
  and g__3139(w__578 ,w__12770 ,w__272);
  and g__3140(w__577 ,w__13005 ,w__131);
  nor g__3141(w__576 ,w__33 ,w__349);
  and g__3142(w__575 ,w__12764 ,w__325);
  or g__3143(w__574 ,w__34 ,w__239);
  and g__3144(w__573 ,w__12973 ,w__169);
  and g__3145(w__572 ,w__12926 ,w__195);
  and g__3146(w__571 ,w__12920 ,w__270);
  and g__3147(w__570 ,w__12961 ,w__249);
  or g__3148(w__569 ,w__67 ,w__231);
  and g__3149(w__568 ,w__13015 ,w__298);
  and g__3150(w__567 ,w__12700 ,w__253);
  or g__3151(w__566 ,w__109 ,w__313);
  and g__3152(w__565 ,w__12783 ,w__274);
  and g__3153(w__564 ,w__12945 ,w__282);
  and g__3154(w__563 ,w__12706 ,w__208);
  and g__3155(w__562 ,w__12919 ,w__161);
  or g__3156(w__561 ,w__119 ,w__289);
  nor g__3157(w__560 ,w__12952 ,w__238);
  and g__3158(w__559 ,w__12995 ,w__271);
  and g__3159(w__558 ,w__12814 ,w__283);
  or g__3160(w__557 ,w__12655 ,w__351);
  nor g__3161(w__556 ,w__12 ,w__237);
  and g__3162(w__555 ,w__12688 ,w__150);
  and g__3163(w__554 ,w__12782 ,w__259);
  and g__3164(w__553 ,w__12993 ,w__133);
  or g__3165(w__552 ,w__51 ,w__335);
  and g__3166(w__551 ,w__12781 ,w__213);
  and g__3167(w__550 ,w__12925 ,w__218);
  or g__3168(w__549 ,w__102 ,w__215);
  and g__3169(w__548 ,w__13014 ,w__192);
  and g__3170(w__547 ,w__12687 ,w__184);
  and g__3171(w__546 ,w__12815 ,w__280);
  or g__3172(w__545 ,w__47 ,w__243);
  and g__3173(w__544 ,w__12938 ,w__154);
  and g__3174(w__543 ,w__12654 ,w__152);
  and g__3175(w__542 ,w__12950 ,w__145);
  and g__3176(w__541 ,w__13020 ,w__226);
  and g__3177(w__540 ,w__97 ,w__350);
  nor g__3178(w__539 ,w__84 ,w__353);
  and g__3179(w__538 ,w__12874 ,w__155);
  and g__3180(w__537 ,w__12992 ,w__320);
  and g__3181(w__536 ,w__12795 ,w__273);
  and g__3182(w__535 ,w__12716 ,w__312);
  or g__3183(w__534 ,w__115 ,w__151);
  and g__3184(w__533 ,w__12978 ,w__194);
  and g__3185(w__532 ,w__12715 ,w__333);
  and g__3186(w__531 ,w__12964 ,w__262);
  and g__3187(w__530 ,w__74 ,w__235);
  and g__3188(w__529 ,w__12747 ,w__134);
  nor g__3189(w__528 ,w__20 ,w__236);
  nor g__3190(w__527 ,w__77 ,w__352);
  and g__3191(w__526 ,w__12765 ,w__293);
  and g__3192(w__525 ,w__12727 ,w__185);
  and g__3193(w__524 ,w__12666 ,w__187);
  and g__3194(w__523 ,w__12885 ,w__328);
  or g__3195(w__522 ,w__59 ,w__211);
  and g__3196(w__521 ,w__13010 ,w__290);
  and g__3197(w__520 ,w__26 ,w__354);
  and g__3198(w__519 ,w__12998 ,w__225);
  or g__3199(w__518 ,w__60 ,w__266);
  and g__3200(w__517 ,w__12981 ,w__245);
  and g__3201(w__516 ,w__13012 ,w__139);
  and g__3202(w__515 ,w__13019 ,w__167);
  and g__3203(w__514 ,w__20 ,w__236);
  and g__3204(w__513 ,w__12807 ,w__198);
  and g__3205(w__512 ,w__12664 ,w__144);
  and g__3206(w__511 ,w__12705 ,w__153);
  nor g__3207(w__510 ,w__26 ,w__354);
  and g__3208(w__509 ,w__12802 ,w__319);
  and g__3209(w__508 ,w__12969 ,w__203);
  and g__3210(w__507 ,w__12965 ,w__142);
  nor g__3211(w__506 ,w__74 ,w__235);
  and g__3212(w__505 ,w__12663 ,w__164);
  and g__3213(w__504 ,w__12744 ,w__206);
  and g__3214(w__503 ,in5[1] ,w__299);
  and g__3215(w__502 ,w__12955 ,w__186);
  and g__3216(w__501 ,w__33 ,w__349);
  and g__3217(w__500 ,w__12959 ,w__330);
  and g__3218(w__499 ,w__12771 ,w__287);
  and g__3219(w__498 ,w__12947 ,w__227);
  and g__3220(w__497 ,w__12766 ,w__168);
  and g__3221(w__496 ,w__12665 ,w__171);
  or g__3222(w__495 ,w__49 ,w__207);
  and g__3223(w__494 ,w__13013 ,w__179);
  and g__3224(w__493 ,w__12797 ,w__137);
  or g__3225(w__492 ,w__123 ,w__256);
  and g__3226(w__491 ,w__12869 ,w__334);
  and g__3227(w__490 ,w__12652 ,w__219);
  or g__3228(w__489 ,w__355 ,w__314);
  xnor g__3229(w__488 ,w__12906 ,w__12812);
  not g__3230(w__476 ,w__477);
  not g__3231(w__474 ,w__475);
  not g__3232(w__471 ,w__472);
  xnor g__3233(w__467 ,w__12915 ,w__12663);
  xnor g__3234(w__466 ,w__13010 ,in5[12]);
  xnor g__3235(w__465 ,w__12897 ,w__12802);
  xnor g__3236(w__464 ,w__12937 ,w__12748);
  xnor g__3237(w__463 ,w__12771 ,w__12739);
  xnor g__3238(w__462 ,w__12910 ,w__12658);
  xnor g__3239(w__461 ,w__13014 ,w__12982);
  xnor g__3240(w__460 ,w__12946 ,w__12757);
  xnor g__3241(w__459 ,w__12914 ,w__12662);
  xnor g__3242(w__458 ,w__12926 ,w__12863);
  xnor g__3243(w__457 ,w__13009 ,in5[11]);
  xnor g__3244(w__456 ,w__12970 ,w__12718);
  xnor g__3245(w__455 ,w__12961 ,w__12898);
  xnor g__3246(w__454 ,w__12902 ,w__12807);
  xnor g__3247(w__453 ,w__12978 ,w__12726);
  xnor g__3248(w__452 ,w__12980 ,w__12728);
  xnor g__3249(w__451 ,w__12955 ,w__12860);
  xnor g__3250(w__450 ,w__12917 ,w__12665);
  xnor g__3251(w__449 ,w__12941 ,w__12752);
  xnor g__3252(w__448 ,w__12892 ,w__12797);
  xnor g__3253(w__447 ,w__12924 ,w__12861);
  xnor g__3254(w__446 ,w__12717 ,w__12686);
  xnor g__3255(w__445 ,w__12766 ,w__12734);
  xnor g__3256(w__444 ,w__12968 ,w__12905);
  xnor g__3257(w__443 ,w__13019 ,w__12987);
  xnor g__3258(w__442 ,w__13013 ,in5[15]);
  xnor g__3259(w__441 ,w__12964 ,w__12901);
  xnor g__3260(w__440 ,w__12893 ,w__12704);
  xnor g__3261(w__439 ,w__12954 ,w__12859);
  xnor g__3262(w__438 ,w__12913 ,w__12661);
  xnor g__3263(w__437 ,w__12963 ,w__12868);
  xnor g__3264(w__436 ,w__12885 ,w__12790);
  xnor g__3265(w__435 ,w__12999 ,in5[1]);
  xnor g__3266(w__434 ,w__12779 ,w__12653);
  xnor g__3267(w__433 ,w__12774 ,w__12742);
  xnor g__3268(w__432 ,w__12900 ,w__12805);
  xnor g__3269(w__431 ,w__12945 ,w__12756);
  xnor g__3270(w__430 ,w__12975 ,w__12723);
  xnor g__3271(w__429 ,w__13004 ,in5[6]);
  xnor g__3272(w__428 ,w__13007 ,in5[9]);
  xnor g__3273(w__427 ,w__12944 ,w__12755);
  xnor g__3274(w__426 ,w__12959 ,w__12864);
  xnor g__3275(w__425 ,w__12911 ,w__12659);
  xnor g__3276(w__424 ,w__12765 ,w__12733);
  xnor g__3277(w__423 ,w__12919 ,w__12856);
  xnor g__3278(w__422 ,w__12912 ,w__12660);
  xnor g__3279(w__421 ,w__12891 ,w__12796);
  xnor g__3280(w__420 ,w__12995 ,w__12806);
  xnor g__3281(w__419 ,w__12896 ,w__12801);
  xnor g__3282(w__418 ,w__12888 ,w__12699);
  xnor g__3283(w__417 ,w__12966 ,w__12903);
  xnor g__3284(w__416 ,w__13029 ,w__12777);
  xnor g__3285(w__415 ,w__12972 ,w__12720);
  xnor g__3286(w__414 ,w__12974 ,w__12722);
  xnor g__3287(w__413 ,w__12764 ,w__12732);
  xnor g__3288(w__412 ,w__13012 ,in5[14]);
  xnor g__3289(w__411 ,w__12940 ,w__12751);
  xnor g__3290(w__410 ,w__12936 ,w__12841);
  xnor g__3291(w__409 ,w__12962 ,w__12899);
  xnor g__3292(w__408 ,w__12943 ,w__12754);
  xnor g__3293(w__407 ,w__12908 ,w__12656);
  xnor g__3294(w__406 ,w__12942 ,w__12753);
  xnor g__3295(w__405 ,w__12967 ,w__12904);
  xnor g__3296(w__404 ,w__12997 ,w__12808);
  xnor g__3297(w__403 ,w__12950 ,w__12761);
  xnor g__3298(w__402 ,w__12939 ,w__12844);
  xnor g__3299(w__401 ,w__13006 ,in5[8]);
  xnor g__3300(w__400 ,w__12916 ,w__12664);
  xnor g__3301(w__399 ,w__12960 ,w__12865);
  xnor g__3302(w__398 ,w__12992 ,w__12803);
  xnor g__3303(w__397 ,w__12869 ,w__12838);
  xnor g__3304(w__396 ,w__12953 ,w__12858);
  xnor g__3305(w__395 ,w__13005 ,in5[7]);
  xnor g__3306(w__394 ,w__12977 ,w__12725);
  xnor g__3307(w__393 ,w__12935 ,w__12683);
  xnor g__3308(w__392 ,w__13020 ,w__12988);
  xnor g__3309(w__391 ,w__13011 ,w__12822);
  xnor g__3310(w__390 ,w__12867 ,w__12836);
  xnor g__3311(w__389 ,w__12909 ,w__12657);
  xnor g__3312(w__388 ,w__12965 ,w__12870);
  xnor g__3313(w__387 ,w__12889 ,w__12700);
  xnor g__3314(w__386 ,w__12770 ,w__12738);
  xnor g__3315(w__385 ,w__13015 ,w__12983);
  xnor g__3316(w__384 ,w__12866 ,w__12835);
  xnor g__3317(w__383 ,w__12871 ,w__12840);
  xnor g__3318(w__382 ,w__13003 ,in5[5]);
  xnor g__3319(w__381 ,w__12976 ,w__12724);
  xnor g__3320(w__380 ,w__12776 ,w__12744);
  xnor g__3321(w__379 ,w__12876 ,w__12813);
  xnor g__3322(w__378 ,w__12895 ,w__12706);
  xnor g__3323(w__377 ,w__12947 ,w__12758);
  xnor g__3324(w__376 ,w__12949 ,w__12760);
  xnor g__3325(w__375 ,w__12811 ,w__12685);
  xnor g__3326(w__374 ,w__12918 ,w__12666);
  xnor g__3327(w__373 ,w__12843 ,w__12749);
  xnor g__3328(w__372 ,w__13002 ,in5[4]);
  xnor g__3329(w__371 ,w__12894 ,w__12705);
  xnor g__3330(w__370 ,w__12993 ,w__12804);
  xnor g__3331(w__369 ,w__12890 ,w__12795);
  xnor g__3332(w__368 ,w__12727 ,in5[13]);
  xnor g__3333(w__367 ,w__12925 ,w__12862);
  xnor g__3334(w__366 ,w__13008 ,in5[10]);
  xnor g__3335(w__365 ,w__12971 ,w__12719);
  xnor g__3336(w__363 ,w__12873 ,w__12810);
  xnor g__3337(w__362 ,w__12981 ,w__12729);
  xnor g__3338(w__361 ,w__12920 ,w__12857);
  xnor g__3339(w__360 ,w__12973 ,w__12721);
  xnor g__3340(w__359 ,w__12875 ,w__12780);
  xnor g__3341(w__358 ,w__13021 ,w__12989);
  xnor g__3342(w__487 ,w__12735 ,w__12672);
  xnor g__3343(w__486 ,w__13017 ,w__12670);
  xnor g__3344(w__485 ,w__13018 ,w__12671);
  xnor g__3345(w__484 ,w__13022 ,w__12675);
  xnor g__3346(w__483 ,w__12736 ,w__12673);
  xnor g__3347(w__482 ,w__13028 ,w__12681);
  xnor g__3348(w__481 ,w__12737 ,w__12674);
  xnor g__3349(w__480 ,w__13023 ,w__12676);
  xnor g__3350(w__479 ,w__12731 ,w__12668);
  xnor g__3351(w__478 ,w__13000 ,in5[2]);
  xnor g__3352(w__477 ,w__13016 ,w__12669);
  xnor g__3353(w__475 ,w__13001 ,in5[3]);
  xnor g__3354(w__473 ,w__13025 ,w__12773);
  xnor g__3355(w__472 ,w__12730 ,w__12667);
  xnor g__3356(w__470 ,w__13027 ,w__12775);
  xnor g__3357(w__469 ,w__13026 ,w__12679);
  xnor g__3358(w__468 ,w__13024 ,w__12772);
  not g__3359(w__351 ,w__352);
  and g__3360(w__348 ,w__12834 ,w__12739);
  or g__3361(w__347 ,w__28 ,w__88);
  and g__3362(w__346 ,w__12906 ,w__12812);
  and g__3363(w__345 ,w__12865 ,w__12708);
  and g__3364(w__344 ,w__12787 ,w__12724);
  or g__3365(w__343 ,w__32 ,w__87);
  and g__3366(w__342 ,w__12861 ,w__12798);
  or g__3367(w__341 ,w__12929 ,w__12835);
  and g__3368(w__340 ,in5[8] ,w__12817);
  and g__3369(w__339 ,w__12996 ,w__12902);
  and g__3370(w__338 ,in5[11] ,w__12820);
  or g__3371(w__337 ,w__96 ,w__31);
  or g__3372(w__336 ,w__12930 ,w__12836);
  nor g__3373(w__335 ,w__12908 ,w__12656);
  or g__3374(w__334 ,w__12932 ,w__12838);
  or g__3375(w__333 ,w__12936 ,w__12841);
  and g__3376(w__332 ,w__12757 ,w__12694);
  or g__3377(w__331 ,w__12757 ,w__12694);
  or g__3378(w__330 ,w__12864 ,w__12707);
  or g__3379(w__329 ,w__41 ,w__76);
  or g__3380(w__328 ,w__12948 ,w__12790);
  and g__3381(w__327 ,w__12895 ,w__12832);
  or g__3382(w__326 ,w__11 ,w__14);
  or g__3383(w__325 ,w__12827 ,w__12732);
  and g__3384(w__324 ,w__12936 ,w__12841);
  and g__3385(w__323 ,in5[13] ,w__12853);
  or g__3386(w__322 ,in5[11] ,w__12820);
  or g__3387(w__321 ,w__79 ,w__37);
  or g__3388(w__320 ,w__12803 ,w__12740);
  or g__3389(w__319 ,w__12991 ,w__12897);
  and g__3390(w__318 ,w__12755 ,w__12692);
  and g__3391(w__317 ,w__12915 ,w__12852);
  nor g__3392(w__316 ,w__12994 ,w__12900);
  and g__3393(w__315 ,in5[15] ,w__12824);
  nor g__3394(w__314 ,w__12875 ,w__12780);
  nor g__3395(w__313 ,w__12941 ,w__12752);
  or g__3396(w__312 ,w__12968 ,w__12905);
  and g__3397(w__311 ,w__12914 ,w__12851);
  and g__3398(w__310 ,w__12857 ,w__12794);
  and g__3399(w__309 ,w__12982 ,w__12762);
  or g__3400(w__308 ,w__12787 ,w__12724);
  and g__3401(w__307 ,w__12756 ,w__12693);
  or g__3402(w__306 ,w__12861 ,w__12798);
  nor g__3403(w__305 ,w__12786 ,w__12723);
  and g__3404(w__304 ,w__12991 ,w__12897);
  and g__3405(w__303 ,w__12894 ,w__12831);
  and g__3406(w__302 ,w__12791 ,w__12728);
  and g__3407(w__301 ,w__12917 ,w__12854);
  and g__3408(w__300 ,w__12985 ,w__12891);
  or g__3409(w__299 ,w__12999 ,w__12684);
  or g__3410(w__298 ,w__12983 ,w__12763);
  and g__3411(w__297 ,w__12754 ,w__12691);
  and g__3412(w__296 ,w__12930 ,w__12836);
  and g__3413(w__295 ,w__12940 ,w__12751);
  and g__3414(w__294 ,w__12829 ,w__12734);
  or g__3415(w__293 ,w__12828 ,w__12733);
  or g__3416(w__292 ,w__80 ,w__13);
  and g__3417(w__291 ,w__12937 ,w__12748);
  or g__3418(w__290 ,in5[12] ,w__12821);
  nor g__3419(w__289 ,w__12909 ,w__12657);
  or g__3420(w__288 ,w__12868 ,w__12711);
  or g__3421(w__287 ,w__12834 ,w__12739);
  and g__3422(w__286 ,w__12785 ,w__12722);
  and g__3423(w__285 ,in5[9] ,w__12818);
  and g__3424(w__284 ,w__12862 ,w__12799);
  or g__3425(w__283 ,in5[5] ,w__13003);
  or g__3426(w__282 ,w__12756 ,w__12693);
  nor g__3427(w__281 ,w__12858 ,w__12701);
  or g__3428(w__280 ,in5[6] ,w__13004);
  and g__3429(w__279 ,w__12988 ,w__12768);
  and g__3430(w__278 ,w__12868 ,w__12711);
  or g__3431(w__277 ,w__12785 ,w__12722);
  nor g__3432(w__276 ,w__12779 ,w__12653);
  and g__3433(w__275 ,w__12870 ,w__12713);
  or g__3434(w__274 ,w__12972 ,w__12720);
  or g__3435(w__273 ,w__12984 ,w__12890);
  or g__3436(w__272 ,w__12833 ,w__12738);
  or g__3437(w__271 ,w__12806 ,w__12743);
  or g__3438(w__270 ,w__12857 ,w__12794);
  and g__3439(w__269 ,w__12984 ,w__12890);
  and g__3440(w__268 ,w__12758 ,w__12695);
  or g__3441(w__267 ,in5[8] ,w__12817);
  nor g__3442(w__266 ,w__12935 ,w__12683);
  and g__3443(w__265 ,w__12901 ,w__12712);
  or g__3444(w__264 ,w__86 ,w__29);
  and g__3445(w__263 ,w__12999 ,w__12684);
  or g__3446(w__262 ,w__12901 ,w__12712);
  and g__3447(w__261 ,w__12971 ,w__12719);
  and g__3448(w__260 ,w__12911 ,w__12848);
  or g__3449(w__259 ,w__12971 ,w__12719);
  and g__3450(w__258 ,w__12837 ,w__12742);
  nor g__3451(w__257 ,w__12899 ,w__12710);
  nor g__3452(w__256 ,w__12990 ,w__12896);
  or g__3453(w__255 ,w__92 ,w__27);
  or g__3454(w__254 ,w__39 ,w__81);
  or g__3455(w__253 ,w__12889 ,w__12826);
  and g__3456(w__252 ,w__12803 ,w__12740);
  and g__3457(w__251 ,w__12864 ,w__12707);
  or g__3458(w__250 ,w__12837 ,w__12742);
  or g__3459(w__249 ,w__12898 ,w__12709);
  and g__3460(w__248 ,w__12804 ,w__12741);
  or g__3461(w__247 ,w__12788 ,w__12725);
  and g__3462(w__246 ,w__12856 ,w__12793);
  or g__3463(w__245 ,w__12792 ,w__12729);
  nor g__3464(w__244 ,w__12876 ,w__12813);
  nor g__3465(w__243 ,w__12989 ,w__12769);
  or g__3466(w__357 ,w__104 ,w__55);
  or g__3467(w__356 ,w__118 ,w__108);
  or g__3468(w__355 ,w__114 ,w__98);
  or g__3469(w__354 ,w__68 ,w__50);
  or g__3470(w__353 ,w__64 ,w__100);
  or g__3471(w__352 ,w__66 ,w__122);
  or g__3472(w__350 ,w__117 ,w__65);
  or g__3473(w__349 ,w__48 ,w__63);
  not g__3474(w__238 ,w__239);
  or g__3475(w__233 ,w__36 ,w__38);
  or g__3476(w__232 ,w__12791 ,w__12728);
  nor g__3477(w__231 ,w__12910 ,w__12847);
  and g__3478(w__230 ,w__12932 ,w__12838);
  or g__3479(w__229 ,w__95 ,w__23);
  or g__3480(w__228 ,w__12865 ,w__12708);
  or g__3481(w__227 ,w__12758 ,w__12695);
  or g__3482(w__226 ,w__12988 ,w__12768);
  and g__3483(w__224 ,in5[4] ,w__13002);
  or g__3484(w__223 ,w__12985 ,w__12891);
  and g__3485(w__222 ,w__12983 ,w__12763);
  or g__3486(w__221 ,in5[10] ,w__12819);
  and g__3487(w__220 ,w__12948 ,w__12790);
  or g__3488(w__219 ,w__12967 ,w__12904);
  or g__3489(w__218 ,w__12862 ,w__12799);
  and g__3490(w__217 ,w__12979 ,w__12916);
  or g__3491(w__216 ,w__16 ,w__91);
  nor g__3492(w__215 ,w__12907 ,w__12844);
  and g__3493(w__214 ,w__12968 ,w__12905);
  or g__3494(w__213 ,w__12970 ,w__12718);
  and g__3495(w__212 ,w__12784 ,w__12721);
  nor g__3496(w__211 ,w__12753 ,w__12690);
  or g__3497(w__210 ,w__12822 ,w__12696);
  nor g__3498(w__209 ,w__12912 ,w__12849);
  or g__3499(w__208 ,w__12895 ,w__12832);
  nor g__3500(w__207 ,w__12893 ,w__12830);
  or g__3501(w__206 ,w__12839 ,w__12776);
  and g__3502(w__205 ,w__12833 ,w__12738);
  and g__3503(w__204 ,w__12987 ,w__12767);
  or g__3504(w__203 ,w__12717 ,w__12686);
  and g__3505(w__202 ,w__12792 ,w__12729);
  and g__3506(w__201 ,in5[7] ,w__12816);
  and g__3507(w__200 ,w__12843 ,w__12749);
  or g__3508(w__199 ,w__12937 ,w__12748);
  or g__3509(w__198 ,w__12996 ,w__12902);
  and g__3510(w__197 ,w__12822 ,w__12696);
  and g__3511(w__196 ,w__12888 ,w__12825);
  or g__3512(w__195 ,w__12863 ,w__12800);
  or g__3513(w__194 ,w__12789 ,w__12726);
  and g__3514(w__193 ,w__12827 ,w__12732);
  or g__3515(w__192 ,w__12982 ,w__12762);
  or g__3516(w__191 ,w__71 ,w__25);
  or g__3517(w__190 ,w__85 ,w__93);
  and g__3518(w__189 ,w__12806 ,w__12743);
  and g__3519(w__188 ,w__12761 ,w__12698);
  or g__3520(w__187 ,w__12918 ,w__12855);
  or g__3521(w__186 ,w__12860 ,w__12703);
  or g__3522(w__185 ,in5[13] ,w__12853);
  or g__3523(w__184 ,in5[4] ,w__13002);
  nor g__3524(w__183 ,w__12859 ,w__12702);
  and g__3525(w__182 ,w__12972 ,w__12720);
  and g__3526(w__181 ,w__12717 ,w__12686);
  or g__3527(w__180 ,w__15 ,w__70);
  or g__3528(w__179 ,in5[15] ,w__12824);
  and g__3529(w__178 ,w__12873 ,w__12810);
  or g__3530(w__177 ,in5[9] ,w__12818);
  and g__3531(w__176 ,w__12863 ,w__12800);
  nor g__3532(w__175 ,w__12913 ,w__12850);
  and g__3533(w__174 ,w__12929 ,w__12835);
  or g__3534(w__173 ,w__22 ,w__40);
  or g__3535(w__172 ,w__12888 ,w__12825);
  or g__3536(w__171 ,w__12917 ,w__12854);
  and g__3537(w__170 ,w__12788 ,w__12725);
  or g__3538(w__169 ,w__12784 ,w__12721);
  or g__3539(w__168 ,w__12829 ,w__12734);
  or g__3540(w__167 ,w__12987 ,w__12767);
  or g__3541(w__166 ,w__90 ,w__24);
  or g__3542(w__165 ,w__12754 ,w__12691);
  or g__3543(w__164 ,w__12915 ,w__12852);
  and g__3544(w__163 ,w__12898 ,w__12709);
  and g__3545(w__162 ,w__12828 ,w__12733);
  or g__3546(w__161 ,w__12856 ,w__12793);
  and g__3547(w__160 ,w__12970 ,w__12718);
  or g__3548(w__159 ,w__12911 ,w__12848);
  and g__3549(w__158 ,w__12889 ,w__12826);
  and g__3550(w__157 ,in5[5] ,w__13003);
  and g__3551(w__156 ,in5[12] ,w__12821);
  or g__3552(w__155 ,w__12811 ,w__12685);
  or g__3553(w__154 ,w__12843 ,w__12749);
  or g__3554(w__153 ,w__12894 ,w__12831);
  or g__3555(w__152 ,w__12906 ,w__12812);
  nor g__3556(w__151 ,w__12760 ,w__12697);
  or g__3557(w__150 ,w__12940 ,w__12751);
  and g__3558(w__149 ,w__12918 ,w__12855);
  or g__3559(w__148 ,w__12755 ,w__12692);
  or g__3560(w__147 ,w__42 ,w__44);
  or g__3561(w__146 ,w__94 ,w__30);
  or g__3562(w__145 ,w__12761 ,w__12698);
  or g__3563(w__144 ,w__12979 ,w__12916);
  and g__3564(w__143 ,w__12811 ,w__12685);
  or g__3565(w__142 ,w__12870 ,w__12713);
  and g__3566(w__141 ,in5[6] ,w__13004);
  and g__3567(w__140 ,w__12967 ,w__12904);
  or g__3568(w__139 ,in5[14] ,w__12823);
  and g__3569(w__138 ,in5[10] ,w__12819);
  or g__3570(w__137 ,w__12986 ,w__12892);
  or g__3571(w__136 ,w__82 ,w__35);
  or g__3572(w__135 ,w__12914 ,w__12851);
  or g__3573(w__134 ,w__12873 ,w__12810);
  or g__3574(w__133 ,w__12804 ,w__12741);
  and g__3575(w__132 ,w__12839 ,w__12776);
  or g__3576(w__131 ,in5[7] ,w__12816);
  and g__3577(w__130 ,w__12860 ,w__12703);
  and g__3578(w__129 ,w__12789 ,w__12726);
  and g__3579(w__128 ,w__12986 ,w__12892);
  and g__3580(w__127 ,in5[14] ,w__12823);
  or g__3581(w__126 ,w__45 ,w__53);
  or g__3582(w__242 ,w__112 ,w__121);
  or g__3583(w__241 ,w__101 ,w__46);
  or g__3584(w__240 ,w__57 ,w__113);
  or g__3585(w__239 ,w__125 ,w__103);
  or g__3586(w__237 ,w__54 ,w__62);
  or g__3587(w__236 ,w__106 ,w__69);
  or g__3588(w__235 ,w__99 ,w__52);
  or g__3589(w__234 ,w__124 ,w__56);
  not g__3590(w__125 ,w__12730);
  not g__3591(w__124 ,w__13017);
  not g__3592(w__123 ,w__12801);
  not g__3593(w__122 ,w__13001);
  not g__3594(w__121 ,w__12668);
  not g__3595(w__120 ,w__12975);
  not g__3596(w__119 ,w__12846);
  not g__3597(w__118 ,w__13025);
  not g__3598(w__117 ,w__13016);
  not g__3599(w__116 ,w__12805);
  not g__3600(w__115 ,w__12949);
  not g__3601(w__114 ,in5[2]);
  not g__3602(w__113 ,w__12676);
  not g__3603(w__112 ,w__12731);
  not g__3604(w__111 ,w__12962);
  not g__3605(w__110 ,w__12953);
  not g__3606(w__109 ,w__12689);
  not g__3607(w__108 ,w__12773);
  not g__3608(w__107 ,w__12750);
  not g__3609(w__106 ,w__13018);
  not g__3610(w__105 ,w__12660);
  not g__3611(w__104 ,w__13026);
  not g__3612(w__103 ,w__12667);
  not g__3613(w__102 ,w__12939);
  not g__3614(w__101 ,w__13024);
  not g__3615(w__100 ,w__12672);
  not g__3616(w__99 ,w__13027);
  not g__3617(w__98 ,w__13000);
  not g__3618(w__97 ,w__12922);
  not g__3619(w__96 ,w__12858);
  not g__3620(w__95 ,w__12908);
  not g__3621(w__94 ,w__12760);
  not g__3622(w__93 ,w__12850);
  not g__3623(w__92 ,w__12859);
  not g__3624(w__91 ,w__12769);
  not g__3625(w__90 ,w__12909);
  not g__3626(w__89 ,w__12921);
  not g__3627(w__88 ,w__12690);
  not g__3628(w__87 ,w__12900);
  not g__3629(w__86 ,w__12990);
  not g__3630(w__85 ,w__12913);
  not g__3631(w__84 ,w__12957);
  not g__3632(w__83 ,w__12680);
  not g__3633(w__82 ,w__12912);
  not g__3634(w__81 ,w__12683);
  not g__3635(w__80 ,w__12893);
  not g__3636(w__79 ,w__12786);
  not g__3637(w__78 ,w__12881);
  not g__3638(w__77 ,w__12655);
  not g__3639(w__76 ,w__12844);
  not g__3640(w__75 ,w__12931);
  not g__3641(w__74 ,w__12933);
  not g__3642(w__73 ,w__12677);
  not g__3643(w__72 ,w__12923);
  not g__3644(w__71 ,w__12941);
  not g__3645(w__70 ,w__12653);
  not g__3646(w__69 ,w__12671);
  not g__3647(w__68 ,w__12737);
  not g__3648(w__67 ,w__12658);
  not g__3649(w__66 ,in5[3]);
  not g__3650(w__65 ,w__12669);
  not g__3651(w__64 ,w__12735);
  not g__3652(w__63 ,w__12675);
  not g__3653(w__62 ,w__12673);
  not g__3654(w__61 ,w__12954);
  not g__3655(w__60 ,w__12872);
  not g__3656(w__59 ,w__12942);
  not g__3657(w__58 ,w__12661);
  not g__3658(w__57 ,w__13023);
  not g__3659(w__56 ,w__12670);
  not g__3660(w__55 ,w__12679);
  not g__3661(w__54 ,w__12736);
  not g__3662(w__53 ,w__12681);
  not g__3663(w__52 ,w__12775);
  not g__3664(w__51 ,w__12845);
  not g__3665(w__50 ,w__12674);
  not g__3666(w__49 ,w__12704);
  not g__3667(w__48 ,w__13022);
  not g__3668(w__47 ,w__13021);
  not g__3669(w__46 ,w__12772);
  not g__3670(w__45 ,w__13028);
  not g__3671(w__44 ,w__12780);
  not g__3672(w__43 ,w__12678);
  not g__3673(w__42 ,w__12875);
  not g__3674(w__41 ,w__12907);
  not g__3675(w__40 ,w__12813);
  not g__3676(w__39 ,w__12935);
  not g__3677(w__38 ,w__12710);
  not g__3678(w__37 ,w__12723);
  not g__3679(w__36 ,w__12899);
  not g__3680(w__35 ,w__12849);
  not g__3681(w__34 ,w__12952);
  not g__3682(w__33 ,w__12928);
  not g__3683(w__32 ,w__12994);
  not g__3684(w__31 ,w__12701);
  not g__3685(w__30 ,w__12697);
  not g__3686(w__29 ,w__12896);
  not g__3687(w__28 ,w__12753);
  not g__3688(w__27 ,w__12702);
  not g__3689(w__26 ,w__12927);
  not g__3690(w__25 ,w__12752);
  not g__3691(w__24 ,w__12657);
  not g__3692(w__23 ,w__12656);
  not g__3693(w__22 ,w__12876);
  not g__3694(w__21 ,w__12951);
  not g__3695(w__20 ,w__12956);
  not g__3696(w__19 ,w__12883);
  not g__3697(w__18 ,w__12879);
  not g__3698(w__17 ,w__12759);
  not g__3699(w__16 ,w__12989);
  not g__3700(w__15 ,w__12779);
  not g__3701(w__14 ,w__12847);
  not g__3702(w__13 ,w__12830);
  not g__3703(w__12 ,w__12958);
  not g__3704(w__11 ,w__12910);
  not g__3705(w__5 ,w__8);
  not g__3706(w__8 ,w__809);
  not g__3707(w__4 ,w__6);
  not g__3708(w__6 ,w__786);
  not g__3709(w__3 ,w__7);
  not g__3710(w__7 ,w__806);
  not g__3711(w__2 ,w__10);
  not g__3712(w__10 ,w__1706);
  not g__3713(w__9 ,w__1335);
  xor g__3714(out1[28] ,w__2391 ,w__2338);
  xor g__3715(out1[26] ,w__2387 ,w__2336);
  xor g__3716(out1[24] ,w__2383 ,w__2333);
  xor g__3717(out1[22] ,w__2379 ,w__2326);
  xor g__3718(out1[20] ,w__2375 ,w__2330);
  xor g__3719(out1[15] ,w__2364 ,w__2274);
  xor g__3720(out1[14] ,w__2362 ,w__2327);
  xor g__3721(out1[13] ,w__2360 ,w__2332);
  xor g__3722(out1[12] ,w__2358 ,w__2325);
  xor g__3723(out1[11] ,w__2356 ,w__2324);
  xor g__3724(out1[10] ,w__2354 ,w__2323);
  xor g__3725(out1[9] ,w__2352 ,w__2322);
  xor g__3726(out1[8] ,w__2350 ,w__2321);
  xor g__3727(out1[6] ,w__2346 ,w__2276);
  xor g__3728(out1[5] ,w__2344 ,w__2275);
  xor g__3729(w__1 ,w__1423 ,w__9);
  xnor g__3730(w__13606 ,w__4071 ,w__4106);
  xnor g__3731(w__13607 ,w__4074 ,w__2406);
  xnor g__3732(w__13609 ,w__4084 ,w__4098);
  xnor g__3733(w__13608 ,w__4080 ,w__4097);
  xnor g__3734(w__13605 ,w__4064 ,w__4099);
  or g__3735(w__13546 ,w__4069 ,w__4105);
  or g__3736(w__13545 ,w__4092 ,w__4104);
  or g__3737(w__13542 ,w__4087 ,w__4101);
  or g__3738(w__13541 ,w__4096 ,w__4103);
  or g__3739(w__13543 ,w__4085 ,w__4102);
  or g__3740(w__13544 ,w__4094 ,w__4100);
  xnor g__3741(w__13604 ,w__4050 ,w__4078);
  xnor g__3742(w__13610 ,w__4081 ,w__4077);
  xnor g__3743(w__13603 ,w__4052 ,w__4076);
  xnor g__3744(w__4106 ,w__3966 ,w__4082);
  and g__3745(w__4105 ,w__4058 ,w__4081);
  and g__3746(w__4104 ,w__4091 ,w__4084);
  or g__3747(w__13539 ,w__4066 ,w__4086);
  and g__3748(w__4103 ,w__4064 ,w__4088);
  nor g__3749(w__4102 ,w__4095 ,w__4083);
  or g__3750(w__13547 ,w__4048 ,w__4089);
  or g__3751(w__13540 ,w__4068 ,w__4090);
  and g__3752(w__4101 ,w__4079 ,w__4082);
  xnor g__3753(w__13611 ,w__4063 ,w__4055);
  xnor g__3754(w__13602 ,w__4051 ,w__4054);
  xnor g__3755(w__13612 ,w__3969 ,w__4056);
  nor g__3756(w__4100 ,w__4093 ,w__4080);
  xnor g__3757(w__4099 ,w__4060 ,w__3986);
  xnor g__3758(w__4098 ,w__4073 ,w__3987);
  xnor g__3759(w__4097 ,w__4061 ,w__4075);
  nor g__3760(w__4096 ,w__2594 ,w__4060);
  and g__3761(w__4095 ,w__3988 ,w__4074);
  nor g__3762(w__4094 ,w__4062 ,w__4075);
  and g__3763(w__4093 ,w__4062 ,w__4075);
  nor g__3764(w__4092 ,w__2592 ,w__4073);
  or g__3765(w__4091 ,w__2744 ,w__4072);
  nor g__3766(w__4090 ,w__4050 ,w__4067);
  and g__3767(w__4089 ,w__4047 ,w__4063);
  or g__3768(w__4088 ,w__2743 ,w__4059);
  nor g__3769(w__4087 ,w__3966 ,w__4071);
  nor g__3770(w__4086 ,w__4052 ,w__4065);
  nor g__3771(w__4085 ,w__3988 ,w__4074);
  or g__3772(w__4079 ,w__3965 ,w__4070);
  or g__3773(w__13601 ,w__4041 ,w__4057);
  xnor g__3774(w__13613 ,w__3995 ,w__2405);
  xnor g__3775(w__13615 ,w__3905 ,w__4025);
  xnor g__3776(w__13537 ,w__3973 ,w__4026);
  xnor g__3777(w__4078 ,w__3937 ,w__4032);
  xnor g__3778(w__4077 ,w__4035 ,w__3990);
  xnor g__3779(w__4076 ,w__3927 ,w__4036);
  xnor g__3780(w__4084 ,w__3972 ,w__4028);
  xnor g__3781(w__4083 ,w__4021 ,w__4024);
  xnor g__3782(w__4082 ,w__3998 ,w__4027);
  xnor g__3783(w__4081 ,w__3970 ,w__4022);
  xnor g__3784(w__4080 ,w__3994 ,w__4023);
  not g__3785(w__4072 ,w__4073);
  not g__3786(w__4070 ,w__4071);
  nor g__3787(w__4069 ,w__3990 ,w__4035);
  nor g__3788(w__4068 ,w__3937 ,w__4033);
  and g__3789(w__4067 ,w__3937 ,w__4033);
  or g__3790(w__13548 ,w__4012 ,w__4046);
  nor g__3791(w__4066 ,w__3927 ,w__4037);
  or g__3792(w__13549 ,w__4010 ,w__4045);
  or g__3793(w__13551 ,w__4006 ,w__4044);
  or g__3794(w__13600 ,w__4004 ,w__4042);
  and g__3795(w__4065 ,w__3927 ,w__4037);
  and g__3796(w__4075 ,w__4018 ,w__4038);
  and g__3797(w__4074 ,w__4001 ,w__4039);
  and g__3798(w__4073 ,w__4016 ,w__4049);
  and g__3799(w__4071 ,w__4007 ,w__4043);
  not g__3800(w__4062 ,w__4061);
  not g__3801(w__4059 ,w__4060);
  or g__3802(w__4058 ,w__3989 ,w__4034);
  nor g__3803(w__4057 ,w__4051 ,w__4040);
  or g__3804(w__13599 ,w__4000 ,w__4029);
  xnor g__3805(w__13614 ,w__3997 ,w__3978);
  or g__3806(w__13550 ,w__3958 ,w__4031);
  xnor g__3807(w__4056 ,w__3941 ,w__3993);
  xnor g__3808(w__4055 ,w__3985 ,w__3983);
  xnor g__3809(w__4054 ,w__3922 ,w__3991);
  xnor g__3810(w__4053 ,w__3996 ,w__3881);
  or g__3811(w__4064 ,w__4013 ,w__4030);
  xnor g__3812(w__4063 ,w__3924 ,w__3976);
  xnor g__3813(w__4061 ,w__3804 ,w__3975);
  xnor g__3814(w__4060 ,w__3971 ,w__3977);
  or g__3815(w__4049 ,w__3970 ,w__4014);
  nor g__3816(w__4048 ,w__3983 ,w__3985);
  or g__3817(w__4047 ,w__3982 ,w__3984);
  and g__3818(w__4046 ,w__4011 ,w__3993);
  nor g__3819(w__4045 ,w__4020 ,w__3995);
  and g__3820(w__4044 ,w__3905 ,w__4005);
  or g__3821(w__13552 ,w__3907 ,w__4003);
  or g__3822(w__4043 ,w__4021 ,w__4002);
  nor g__3823(w__4042 ,w__3979 ,w__3996);
  nor g__3824(w__4041 ,w__3922 ,w__3992);
  and g__3825(w__4040 ,w__3922 ,w__3992);
  or g__3826(w__4039 ,w__3994 ,w__4019);
  or g__3827(w__4038 ,w__3972 ,w__4017);
  and g__3828(w__4052 ,w__3899 ,w__4008);
  and g__3829(w__4051 ,w__3834 ,w__3981);
  and g__3830(w__4050 ,w__3962 ,w__4015);
  not g__3831(w__4037 ,w__4036);
  not g__3832(w__4034 ,w__4035);
  not g__3833(w__4033 ,w__4032);
  nor g__3834(w__4031 ,w__3959 ,w__3997);
  nor g__3835(w__4030 ,w__4009 ,w__3998);
  nor g__3836(w__4029 ,w__3973 ,w__3999);
  xnor g__3837(w__13616 ,w__3953 ,w__3933);
  xnor g__3838(w__13536 ,w__3902 ,w__3931);
  xnor g__3839(w__4028 ,w__3807 ,w__3939);
  xnor g__3840(w__4027 ,w__3926 ,w__3950);
  xnor g__3841(w__4026 ,w__3707 ,w__3948);
  xnor g__3842(w__4025 ,w__3945 ,w__3746);
  xnor g__3843(w__4024 ,w__3947 ,w__3921);
  xnor g__3844(w__4023 ,w__3936 ,w__3677);
  xnor g__3845(w__4022 ,w__3876 ,w__3943);
  xnor g__3846(w__4036 ,w__3952 ,w__3891);
  and g__3847(w__4035 ,w__3934 ,w__3980);
  xnor g__3848(w__4032 ,w__3974 ,w__3932);
  and g__3849(w__4020 ,w__3946 ,w__3967);
  and g__3850(w__4019 ,w__3677 ,w__3936);
  or g__3851(w__4018 ,w__3806 ,w__3939);
  nor g__3852(w__4017 ,w__3807 ,w__3938);
  or g__3853(w__4016 ,w__3876 ,w__3942);
  or g__3854(w__4015 ,w__3960 ,w__3971);
  nor g__3855(w__4014 ,w__3875 ,w__3943);
  nor g__3856(w__4013 ,w__3926 ,w__3951);
  nor g__3857(w__4012 ,w__3969 ,w__3941);
  or g__3858(w__4011 ,w__3968 ,w__3940);
  nor g__3859(w__4010 ,w__3946 ,w__3967);
  and g__3860(w__4009 ,w__3926 ,w__3951);
  or g__3861(w__4008 ,w__3909 ,w__3974);
  or g__3862(w__4007 ,w__3921 ,w__3947);
  nor g__3863(w__4006 ,w__2595 ,w__3945);
  or g__3864(w__4005 ,w__2742 ,w__3944);
  nor g__3865(w__4004 ,w__3881 ,w__3964);
  and g__3866(w__4003 ,w__3908 ,w__3953);
  and g__3867(w__4002 ,w__3921 ,w__3947);
  or g__3868(w__13597 ,w__3913 ,w__3955);
  or g__3869(w__13598 ,w__3916 ,w__3954);
  or g__3870(w__4001 ,w__3677 ,w__3936);
  nor g__3871(w__4000 ,w__3707 ,w__3949);
  and g__3872(w__3999 ,w__3707 ,w__3949);
  and g__3873(w__4021 ,w__3824 ,w__3963);
  not g__3874(w__3992 ,w__3991);
  not g__3875(w__3990 ,w__3989);
  not g__3876(w__3984 ,w__3985);
  not g__3877(w__3982 ,w__3983);
  xnor g__3878(w__13534 ,w__3675 ,w__3897);
  xnor g__3879(w__13617 ,w__3903 ,w__3890);
  or g__3880(w__3981 ,w__3868 ,w__3952);
  or g__3881(w__3980 ,w__3904 ,w__3935);
  and g__3882(w__3979 ,w__3881 ,w__3964);
  or g__3883(w__13553 ,w__3827 ,w__3961);
  xnor g__3884(w__13618 ,w__3799 ,w__3888);
  xnor g__3885(w__13535 ,w__3880 ,w__3894);
  xnor g__3886(w__3978 ,w__3838 ,w__3928);
  xnor g__3887(w__3977 ,w__3925 ,w__3837);
  xnor g__3888(w__3976 ,w__3712 ,w__3904);
  xnor g__3889(w__3975 ,w__3930 ,w__3740);
  xnor g__3890(w__3998 ,w__3705 ,w__3886);
  xnor g__3891(w__3997 ,w__3809 ,w__3887);
  xnor g__3892(w__3996 ,w__2403 ,w__3889);
  xnor g__3893(w__3995 ,w__3842 ,w__3896);
  and g__3894(w__3994 ,w__3833 ,w__3956);
  xnor g__3895(w__3993 ,w__3929 ,w__3895);
  xnor g__3896(w__3991 ,w__3843 ,w__3893);
  xnor g__3897(w__3989 ,w__3743 ,w__3892);
  xnor g__3898(w__3988 ,w__3669 ,w__3885);
  xnor g__3899(w__3987 ,w__3901 ,w__3882);
  xnor g__3900(w__3986 ,w__3744 ,w__3883);
  xnor g__3901(w__3985 ,w__3738 ,w__3884);
  and g__3902(w__3983 ,w__3862 ,w__3957);
  not g__3903(w__3968 ,w__3969);
  not g__3904(w__3965 ,w__3966);
  or g__3905(w__3963 ,w__3823 ,w__3930);
  or g__3906(w__3962 ,w__3837 ,w__3925);
  nor g__3907(w__3961 ,w__3826 ,w__3903);
  and g__3908(w__3960 ,w__3837 ,w__3925);
  and g__3909(w__3959 ,w__3839 ,w__3928);
  nor g__3910(w__3958 ,w__3839 ,w__3928);
  or g__3911(w__3957 ,w__3929 ,w__3859);
  or g__3912(w__3956 ,w__3831 ,w__3901);
  and g__3913(w__3955 ,w__3808 ,w__3915);
  and g__3914(w__3954 ,w__3902 ,w__3911);
  and g__3915(w__3974 ,w__3874 ,w__3918);
  and g__3916(w__3973 ,w__3847 ,w__3898);
  and g__3917(w__3972 ,w__3873 ,w__3919);
  and g__3918(w__3971 ,w__3829 ,w__3912);
  and g__3919(w__3970 ,w__3867 ,w__3917);
  and g__3920(w__3969 ,w__3858 ,w__3910);
  and g__3921(w__3967 ,w__3854 ,w__3920);
  and g__3922(w__3966 ,w__3852 ,w__3906);
  and g__3923(w__3964 ,w__3872 ,w__3914);
  not g__3924(w__3951 ,w__3950);
  not g__3925(w__3949 ,w__3948);
  not g__3926(w__3944 ,w__3945);
  not g__3927(w__3942 ,w__3943);
  not g__3928(w__3940 ,w__3941);
  not g__3929(w__3938 ,w__3939);
  xnor g__3930(w__13619 ,w__3755 ,w__2404);
  or g__3931(w__13554 ,w__3845 ,w__3900);
  nor g__3932(w__3935 ,w__3712 ,w__3923);
  or g__3933(w__3934 ,w__3711 ,w__3924);
  xnor g__3934(w__3933 ,w__3878 ,w__3729);
  xnor g__3935(w__3932 ,w__2401 ,w__3836);
  xnor g__3936(w__3931 ,w__3841 ,w__3730);
  xnor g__3937(w__3953 ,w__3762 ,w__3816);
  xnor g__3938(w__3952 ,w__3757 ,w__3813);
  xnor g__3939(w__3950 ,w__3714 ,w__2400);
  xnor g__3940(w__3948 ,w__3758 ,w__2402);
  xnor g__3941(w__3947 ,w__3751 ,w__3812);
  xnor g__3942(w__3946 ,w__3716 ,w__3810);
  xnor g__3943(w__3945 ,w__3756 ,w__3811);
  xnor g__3944(w__3943 ,w__3690 ,w__3818);
  xnor g__3945(w__3941 ,w__3763 ,w__3819);
  xnor g__3946(w__3939 ,w__3667 ,w__3815);
  xnor g__3947(w__3937 ,w__3748 ,w__3817);
  xnor g__3948(w__3936 ,w__3749 ,w__3814);
  not g__3949(w__3923 ,w__3924);
  or g__3950(w__3920 ,w__3809 ,w__3853);
  or g__3951(w__3919 ,w__3754 ,w__3871);
  or g__3952(w__3918 ,w__3753 ,w__3870);
  or g__3953(w__3917 ,w__3752 ,w__3865);
  nor g__3954(w__3916 ,w__2596 ,w__3841);
  or g__3955(w__3915 ,w__3701 ,w__3879);
  or g__3956(w__3914 ,w__3864 ,w__3844);
  nor g__3957(w__3913 ,w__3702 ,w__3880);
  or g__3958(w__13596 ,w__3764 ,w__3832);
  or g__3959(w__3912 ,w__3759 ,w__3828);
  or g__3960(w__3911 ,w__2741 ,w__3840);
  or g__3961(w__3910 ,w__3842 ,w__3856);
  or g__3962(w__13555 ,w__3772 ,w__3857);
  nor g__3963(w__3909 ,w__2401 ,w__3835);
  or g__3964(w__3908 ,w__2740 ,w__3877);
  nor g__3965(w__3907 ,w__2593 ,w__3878);
  or g__3966(w__3906 ,w__3750 ,w__3850);
  and g__3967(w__3930 ,w__3773 ,w__3860);
  and g__3968(w__3929 ,w__3791 ,w__3861);
  and g__3969(w__3928 ,w__3783 ,w__3851);
  and g__3970(w__3927 ,w__3787 ,w__3846);
  and g__3971(w__3926 ,w__3788 ,w__3855);
  and g__3972(w__3925 ,w__3796 ,w__3866);
  and g__3973(w__3924 ,w__3795 ,w__3863);
  and g__3974(w__3922 ,w__3780 ,w__3820);
  and g__3975(w__3921 ,w__3779 ,w__3848);
  or g__3976(w__13556 ,w__3620 ,w__3821);
  nor g__3977(w__3900 ,w__3761 ,w__3849);
  or g__3978(w__3899 ,w__3805 ,w__3836);
  xnor g__3979(w__13620 ,w__3760 ,w__3663);
  or g__3980(w__3898 ,w__2403 ,w__3869);
  xnor g__3981(w__3897 ,w__3747 ,w__3375);
  xnor g__3982(w__3896 ,w__3732 ,w__3733);
  xnor g__3983(w__3895 ,w__3735 ,w__3802);
  xnor g__3984(w__3894 ,w__3702 ,w__3808);
  xnor g__3985(w__3893 ,w__3736 ,w__3710);
  xnor g__3986(w__3892 ,w__3722 ,w__3754);
  xnor g__3987(w__3891 ,w__3682 ,w__3726);
  xnor g__3988(w__3890 ,w__3673 ,w__3728);
  xnor g__3989(w__3889 ,w__3724 ,w__3668);
  xnor g__3990(w__3888 ,w__3761 ,w__3685);
  xnor g__3991(w__3887 ,w__3731 ,w__3727);
  xnor g__3992(w__3886 ,w__3745 ,w__3759);
  xnor g__3993(w__3885 ,w__3741 ,w__3750);
  xnor g__3994(w__3884 ,w__3752 ,w__3698);
  xnor g__3995(w__3883 ,w__3753 ,w__3704);
  xnor g__3996(w__3882 ,w__3737 ,w__3723);
  or g__3997(w__3905 ,w__3778 ,w__3822);
  xnor g__3998(w__3904 ,w__3713 ,w__3720);
  xnor g__3999(w__3903 ,w__3688 ,w__3719);
  or g__4000(w__3902 ,w__3794 ,w__3825);
  and g__4001(w__3901 ,w__3766 ,w__3830);
  not g__4002(w__3879 ,w__3880);
  not g__4003(w__3877 ,w__3878);
  not g__4004(w__3875 ,w__3876);
  or g__4005(w__13595 ,w__3491 ,w__3769);
  or g__4006(w__3874 ,w__3704 ,w__3744);
  or g__4007(w__3873 ,w__3721 ,w__3743);
  or g__4008(w__3872 ,w__3710 ,w__3736);
  nor g__4009(w__3871 ,w__3722 ,w__3742);
  and g__4010(w__3870 ,w__3704 ,w__3744);
  and g__4011(w__3869 ,w__3668 ,w__3724);
  nor g__4012(w__3868 ,w__3682 ,w__3725);
  or g__4013(w__3867 ,w__3698 ,w__3738);
  or g__4014(w__3866 ,w__3714 ,w__3793);
  and g__4015(w__3865 ,w__3698 ,w__3738);
  and g__4016(w__3864 ,w__3710 ,w__3736);
  or g__4017(w__3863 ,w__3763 ,w__3792);
  or g__4018(w__3862 ,w__3735 ,w__3801);
  or g__4019(w__3861 ,w__3716 ,w__3790);
  or g__4020(w__3860 ,w__3686 ,w__3770);
  nor g__4021(w__3859 ,w__3734 ,w__3802);
  or g__4022(w__3858 ,w__3733 ,w__3732);
  nor g__4023(w__3857 ,w__3771 ,w__3755);
  and g__4024(w__3856 ,w__3733 ,w__3732);
  or g__4025(w__3855 ,w__3786 ,w__3751);
  or g__4026(w__3854 ,w__3727 ,w__3731);
  and g__4027(w__3853 ,w__3727 ,w__3731);
  or g__4028(w__3852 ,w__3669 ,w__3741);
  or g__4029(w__3851 ,w__3782 ,w__3756);
  and g__4030(w__3850 ,w__3669 ,w__3741);
  and g__4031(w__3849 ,w__3685 ,w__3800);
  or g__4032(w__3848 ,w__3775 ,w__3749);
  or g__4033(w__3847 ,w__3668 ,w__3724);
  or g__4034(w__3846 ,w__3774 ,w__3748);
  nor g__4035(w__3845 ,w__3685 ,w__3800);
  and g__4036(w__3881 ,w__3466 ,w__3789);
  and g__4037(w__3880 ,w__3507 ,w__3781);
  and g__4038(w__3878 ,w__3664 ,w__3776);
  and g__4039(w__3876 ,w__3691 ,w__3797);
  not g__4040(w__3844 ,w__3843);
  not g__4041(w__3840 ,w__3841);
  not g__4042(w__3839 ,w__3838);
  not g__4043(w__3835 ,w__3836);
  xnor g__4044(w__13533 ,w__3718 ,w__3612);
  or g__4045(w__3834 ,w__3681 ,w__3726);
  or g__4046(w__3833 ,w__3723 ,w__3737);
  nor g__4047(w__3832 ,w__3784 ,w__3747);
  and g__4048(w__3831 ,w__3723 ,w__3737);
  or g__4049(w__3830 ,w__3690 ,w__3777);
  or g__4050(w__3829 ,w__3705 ,w__3745);
  and g__4051(w__3828 ,w__3705 ,w__3745);
  nor g__4052(w__3827 ,w__3674 ,w__3728);
  and g__4053(w__3826 ,w__3674 ,w__3728);
  nor g__4054(w__3825 ,w__3785 ,w__3758);
  or g__4055(w__3824 ,w__3740 ,w__3803);
  nor g__4056(w__3823 ,w__3739 ,w__3804);
  nor g__4057(w__3822 ,w__3798 ,w__3762);
  nor g__4058(w__3821 ,w__3618 ,w__3760);
  or g__4059(w__3820 ,w__3768 ,w__3757);
  xnor g__4060(w__3819 ,w__3706 ,w__3708);
  xnor g__4061(w__3818 ,w__3498 ,w__3672);
  xnor g__4062(w__3817 ,w__3680 ,w__3697);
  xnor g__4063(w__3816 ,w__3495 ,w__3670);
  xnor g__4064(w__3815 ,w__3686 ,w__3684);
  xnor g__4065(w__3814 ,w__3678 ,w__3679);
  xnor g__4066(w__3813 ,w__3676 ,w__3295);
  xnor g__4067(w__3812 ,w__3699 ,w__3700);
  xnor g__4068(w__3811 ,w__3694 ,w__3695);
  xnor g__4069(w__3810 ,w__3703 ,w__3604);
  xnor g__4070(w__3843 ,w__3717 ,w__3610);
  and g__4071(w__3842 ,w__3640 ,w__3765);
  xnor g__4072(w__3841 ,w__3687 ,w__3597);
  xnor g__4073(w__3838 ,w__3715 ,w__3662);
  xnor g__4074(w__3837 ,w__3689 ,w__3598);
  and g__4075(w__3836 ,w__3445 ,w__3767);
  not g__4076(w__3806 ,w__3807);
  not g__4077(w__3805 ,w__2401);
  not g__4078(w__3803 ,w__3804);
  not g__4079(w__3801 ,w__3802);
  not g__4080(w__3800 ,w__3799);
  and g__4081(w__3798 ,w__3496 ,w__3670);
  or g__4082(w__3797 ,w__3692 ,w__3713);
  or g__4083(w__3796 ,w__3292 ,w__3696);
  or g__4084(w__3795 ,w__3708 ,w__3706);
  nor g__4085(w__3794 ,w__3371 ,w__3709);
  and g__4086(w__3793 ,w__3292 ,w__3696);
  and g__4087(w__3792 ,w__3708 ,w__3706);
  or g__4088(w__3791 ,w__3604 ,w__3703);
  and g__4089(w__3790 ,w__3604 ,w__3703);
  or g__4090(w__3789 ,w__3470 ,w__3717);
  or g__4091(w__3788 ,w__3700 ,w__3699);
  or g__4092(w__3787 ,w__3697 ,w__3680);
  and g__4093(w__3786 ,w__3700 ,w__3699);
  and g__4094(w__3785 ,w__3371 ,w__3709);
  nor g__4095(w__3784 ,w__3374 ,w__3675);
  or g__4096(w__3783 ,w__3695 ,w__3694);
  and g__4097(w__3782 ,w__3695 ,w__3694);
  or g__4098(w__3781 ,w__3462 ,w__3687);
  or g__4099(w__3780 ,w__3295 ,w__3676);
  or g__4100(w__3779 ,w__3679 ,w__3678);
  nor g__4101(w__3778 ,w__3496 ,w__3670);
  nor g__4102(w__3777 ,w__3498 ,w__3671);
  or g__4103(w__3776 ,w__3688 ,w__3665);
  and g__4104(w__3775 ,w__3679 ,w__3678);
  and g__4105(w__3774 ,w__3697 ,w__3680);
  or g__4106(w__3773 ,w__3667 ,w__3684);
  nor g__4107(w__3772 ,w__3605 ,w__3683);
  and g__4108(w__3771 ,w__3605 ,w__3683);
  or g__4109(w__13557 ,w__3458 ,w__3666);
  and g__4110(w__3770 ,w__3667 ,w__3684);
  nor g__4111(w__3769 ,w__3484 ,w__3718);
  and g__4112(w__3768 ,w__2550 ,w__3676);
  or g__4113(w__3767 ,w__3444 ,w__3689);
  or g__4114(w__3766 ,w__3497 ,w__3672);
  or g__4115(w__3765 ,w__3639 ,w__3715);
  and g__4116(w__3764 ,w__2598 ,w__3675);
  and g__4117(w__3809 ,w__3500 ,w__3693);
  xnor g__4118(w__3808 ,w__3590 ,w__3375);
  xnor g__4119(w__3807 ,w__3576 ,w__2617);
  xnor g__4120(w__3804 ,w__3609 ,w__3376);
  xnor g__4121(w__3802 ,w__3554 ,w__3568);
  xnor g__4122(w__3799 ,w__3499 ,w__3555);
  not g__4123(w__3742 ,w__3743);
  not g__4124(w__3739 ,w__3740);
  not g__4125(w__3734 ,w__3735);
  not g__4126(w__3725 ,w__3726);
  not g__4127(w__3721 ,w__3722);
  xnor g__4128(w__13622 ,w__3342 ,w__3595);
  xnor g__4129(w__13532 ,w__3565 ,w__2784);
  xnor g__4130(w__13621 ,w__3607 ,w__3585);
  xnor g__4131(w__3720 ,w__3603 ,w__3410);
  xnor g__4132(w__3719 ,w__3606 ,w__3327);
  xnor g__4133(w__3763 ,w__3408 ,w__3594);
  xnor g__4134(w__3762 ,w__3377 ,w__3596);
  xnor g__4135(w__3761 ,w__3421 ,w__3591);
  xnor g__4136(w__3760 ,w__3303 ,w__3592);
  xnor g__4137(w__3759 ,w__3567 ,w__2813);
  xnor g__4138(w__3758 ,w__3357 ,w__3587);
  xnor g__4139(w__3757 ,w__3580 ,w__2817);
  xnor g__4140(w__3756 ,w__3348 ,w__3560);
  xnor g__4141(w__3755 ,w__3424 ,w__3578);
  xnor g__4142(w__3754 ,w__3432 ,w__3573);
  xnor g__4143(w__3753 ,w__3355 ,w__3572);
  xnor g__4144(w__3752 ,w__3423 ,w__3570);
  xnor g__4145(w__3751 ,w__3422 ,w__3562);
  xnor g__4146(w__3750 ,w__3431 ,w__3601);
  xnor g__4147(w__3749 ,w__3425 ,w__3557);
  xnor g__4148(w__3748 ,w__3317 ,w__3556);
  xnor g__4149(w__3747 ,w__3566 ,w__2794);
  xnor g__4150(w__3746 ,w__3608 ,w__3559);
  xnor g__4151(w__3745 ,w__3354 ,w__3589);
  xnor g__4152(w__3744 ,w__3427 ,w__3574);
  xnor g__4153(w__3743 ,w__3329 ,w__3602);
  xnor g__4154(w__3741 ,w__3561 ,w__3373);
  xnor g__4155(w__3740 ,w__3395 ,w__3586);
  xnor g__4156(w__3738 ,w__3323 ,w__3571);
  xnor g__4157(w__3737 ,w__3442 ,w__3584);
  xnor g__4158(w__3736 ,w__3320 ,w__3575);
  xnor g__4159(w__3735 ,w__3390 ,w__3569);
  xnor g__4160(w__3733 ,w__3411 ,w__3564);
  xnor g__4161(w__3732 ,w__3429 ,w__3563);
  xnor g__4162(w__3731 ,w__3399 ,w__3583);
  xnor g__4163(w__3730 ,w__3558 ,w__2815);
  xnor g__4164(w__3729 ,w__3407 ,w__3582);
  xnor g__4165(w__3728 ,w__3345 ,w__3577);
  xnor g__4166(w__3727 ,w__3330 ,w__3593);
  xnor g__4167(w__3726 ,w__3391 ,w__3579);
  xnor g__4168(w__3724 ,w__3397 ,w__3581);
  xnor g__4169(w__3723 ,w__3310 ,w__3600);
  xnor g__4170(w__3722 ,w__3366 ,w__3611);
  not g__4171(w__3711 ,w__3712);
  not g__4172(w__3701 ,w__3702);
  or g__4173(w__3693 ,w__3508 ,w__3608);
  and g__4174(w__3692 ,w__3410 ,w__3603);
  or g__4175(w__3691 ,w__3410 ,w__3603);
  and g__4176(w__3718 ,w__3546 ,w__3630);
  and g__4177(w__3717 ,w__3551 ,w__3645);
  and g__4178(w__3716 ,w__3514 ,w__3642);
  and g__4179(w__3715 ,w__3505 ,w__3636);
  and g__4180(w__3714 ,w__3534 ,w__3649);
  and g__4181(w__3713 ,w__3542 ,w__3655);
  or g__4182(w__3712 ,w__3537 ,w__3650);
  and g__4183(w__3710 ,w__3544 ,w__3653);
  and g__4184(w__3709 ,w__3526 ,w__3638);
  and g__4185(w__3708 ,w__3531 ,w__3648);
  and g__4186(w__3707 ,w__3447 ,w__3660);
  and g__4187(w__3706 ,w__3527 ,w__3646);
  and g__4188(w__3705 ,w__3525 ,w__3644);
  and g__4189(w__3704 ,w__3549 ,w__3659);
  and g__4190(w__3703 ,w__3517 ,w__3643);
  and g__4191(w__3702 ,w__3545 ,w__3656);
  and g__4192(w__3700 ,w__3511 ,w__3641);
  and g__4193(w__3699 ,w__3506 ,w__3637);
  and g__4194(w__3698 ,w__3540 ,w__3654);
  and g__4195(w__3697 ,w__3504 ,w__3633);
  and g__4196(w__3696 ,w__3539 ,w__3652);
  and g__4197(w__3695 ,w__3490 ,w__3661);
  and g__4198(w__3694 ,w__3548 ,w__3632);
  not g__4199(w__3681 ,w__3682);
  not g__4200(w__3674 ,w__3673);
  not g__4201(w__3671 ,w__3672);
  and g__4202(w__3666 ,w__3465 ,w__3607);
  or g__4203(w__13558 ,w__3468 ,w__3616);
  and g__4204(w__3665 ,w__3327 ,w__3606);
  or g__4205(w__3664 ,w__3327 ,w__3606);
  xnor g__4206(w__3663 ,w__3301 ,w__3493);
  xnor g__4207(w__3662 ,w__3394 ,w__3553);
  and g__4208(w__3690 ,w__3521 ,w__3634);
  and g__4209(w__3689 ,w__3457 ,w__3614);
  and g__4210(w__3688 ,w__3486 ,w__3626);
  and g__4211(w__3687 ,w__3451 ,w__3615);
  and g__4212(w__3686 ,w__3464 ,w__3617);
  and g__4213(w__3685 ,w__3473 ,w__3624);
  and g__4214(w__3684 ,w__3513 ,w__3621);
  and g__4215(w__3683 ,w__3472 ,w__3623);
  or g__4216(w__3682 ,w__3450 ,w__3622);
  and g__4217(w__3680 ,w__3454 ,w__3627);
  and g__4218(w__3679 ,w__3485 ,w__3631);
  and g__4219(w__3678 ,w__3481 ,w__3628);
  and g__4220(w__3677 ,w__3463 ,w__3651);
  and g__4221(w__3676 ,w__3455 ,w__3657);
  or g__4222(w__3675 ,w__3449 ,w__3647);
  or g__4223(w__3673 ,w__3476 ,w__3635);
  and g__4224(w__3672 ,w__3460 ,w__3658);
  and g__4225(w__3670 ,w__3483 ,w__3629);
  and g__4226(w__3669 ,w__3492 ,w__3613);
  and g__4227(w__3668 ,w__3474 ,w__3619);
  and g__4228(w__3667 ,w__3443 ,w__3625);
  or g__4229(w__3661 ,w__3440 ,w__3489);
  or g__4230(w__3660 ,w__3441 ,w__3446);
  or g__4231(w__3659 ,w__3439 ,w__3547);
  or g__4232(w__3658 ,w__3438 ,w__3522);
  or g__4233(w__3657 ,w__3365 ,w__3456);
  or g__4234(w__3656 ,w__3543 ,w__3437);
  or g__4235(w__3655 ,w__3353 ,w__3541);
  or g__4236(w__3654 ,w__3436 ,w__3538);
  or g__4237(w__3653 ,w__3435 ,w__3535);
  or g__4238(w__3652 ,w__3433 ,w__3536);
  or g__4239(w__3651 ,w__2739 ,w__3533);
  and g__4240(w__3650 ,w__3554 ,w__3532);
  or g__4241(w__3649 ,w__3431 ,w__3529);
  or g__4242(w__3648 ,w__3430 ,w__3528);
  nor g__4243(w__3647 ,w__3452 ,w__2598);
  or g__4244(w__3646 ,w__3429 ,w__3523);
  or g__4245(w__3645 ,w__3367 ,w__3516);
  or g__4246(w__3644 ,w__2619 ,w__3520);
  or g__4247(w__3643 ,w__3428 ,w__3515);
  or g__4248(w__3642 ,w__3351 ,w__3512);
  or g__4249(w__3641 ,w__3356 ,w__3509);
  or g__4250(w__3640 ,w__3394 ,w__3552);
  nor g__4251(w__3639 ,w__3393 ,w__3553);
  or g__4252(w__3638 ,w__3426 ,w__3502);
  or g__4253(w__3637 ,w__3425 ,w__3501);
  or g__4254(w__3636 ,w__3348 ,w__3503);
  and g__4255(w__3635 ,w__3499 ,w__3530);
  or g__4256(w__3634 ,w__3423 ,w__3550);
  or g__4257(w__3633 ,w__3427 ,w__3518);
  or g__4258(w__3632 ,w__3344 ,w__3487);
  or g__4259(w__3631 ,w__3341 ,w__3482);
  or g__4260(w__3630 ,w__3479 ,w__3364);
  or g__4261(w__3629 ,w__3345 ,w__3480);
  or g__4262(w__3628 ,w__3442 ,w__3478);
  or g__4263(w__3627 ,w__3355 ,w__3475);
  or g__4264(w__3626 ,w__3360 ,w__3477);
  or g__4265(w__3625 ,w__3459 ,w__3366);
  or g__4266(w__3624 ,w__3424 ,w__3461);
  or g__4267(w__3623 ,w__3352 ,w__3471);
  and g__4268(w__3622 ,w__3453 ,w__2550);
  or g__4269(w__3621 ,w__3432 ,w__3469);
  nor g__4270(w__3620 ,w__3301 ,w__3494);
  or g__4271(w__3619 ,w__3434 ,w__3519);
  and g__4272(w__3618 ,w__3301 ,w__3494);
  or g__4273(w__3617 ,w__3363 ,w__3467);
  nor g__4274(w__3616 ,w__3342 ,w__3510);
  or g__4275(w__3615 ,w__3448 ,w__3357);
  or g__4276(w__3614 ,w__3354 ,w__3524);
  or g__4277(w__3613 ,w__2617 ,w__3488);
  xnor g__4278(w__13623 ,w__3368 ,w__3289);
  xnor g__4279(w__3612 ,w__3300 ,w__2600);
  xnor g__4280(w__3611 ,w__3334 ,w__2792);
  xnor g__4281(w__3610 ,w__3314 ,w__3293);
  xnor g__4282(w__3609 ,w__3379 ,w__2619);
  xnor g__4283(w__3602 ,w__3296 ,w__3363);
  xnor g__4284(w__3601 ,w__3413 ,w__2812);
  xnor g__4285(w__3600 ,w__3341 ,w__2786);
  xnor g__4286(w__3599 ,w__3441 ,w__2818);
  xnor g__4287(w__3598 ,w__2548 ,w__2788);
  xnor g__4288(w__3597 ,w__3383 ,w__3370);
  xnor g__4289(w__3596 ,w__3440 ,w__3047);
  xnor g__4290(w__3595 ,w__3052 ,w__3336);
  xnor g__4291(w__3594 ,w__3353 ,w__3050);
  xnor g__4292(w__3593 ,w__3428 ,w__3048);
  xnor g__4293(w__3592 ,w__3352 ,w__3051);
  xnor g__4294(w__3591 ,w__3360 ,w__3049);
  xnor g__4295(w__3590 ,w__3316 ,w__2814);
  xnor g__4296(w__3589 ,w__3378 ,w__3315);
  xnor g__4297(w__3588 ,w__3313 ,w__2790);
  xnor g__4298(w__3587 ,w__3311 ,w__2816);
  xnor g__4299(w__3586 ,w__3356 ,w__2787);
  xnor g__4300(w__3585 ,w__3338 ,w__3298);
  xnor g__4301(w__3584 ,w__3331 ,w__3306);
  xnor g__4302(w__3583 ,w__3398 ,w__3351);
  xnor g__4303(w__3582 ,w__3402 ,w__3344);
  xnor g__4304(w__3581 ,w__3426 ,w__3403);
  xnor g__4305(w__3580 ,w__3401 ,w__3367);
  xnor g__4306(w__3579 ,w__3435 ,w__3412);
  xnor g__4307(w__3578 ,w__3307 ,w__3309);
  xnor g__4308(w__3577 ,w__3299 ,w__3332);
  xnor g__4309(w__3576 ,w__3322 ,w__3318);
  xnor g__4310(w__3575 ,w__3434 ,w__2791);
  xnor g__4311(w__3574 ,w__3382 ,w__3386);
  xnor g__4312(w__3573 ,w__3302 ,w__3384);
  xnor g__4313(w__3572 ,w__3335 ,w__3319);
  xnor g__4314(w__3571 ,w__3321 ,w__3438);
  xnor g__4315(w__3570 ,w__3326 ,w__3396);
  xnor g__4316(w__3569 ,w__3405 ,w__3436);
  xnor g__4317(w__3568 ,w__3416 ,w__3418);
  xnor g__4318(w__3567 ,w__3439 ,w__3420);
  xnor g__4319(w__3566 ,w__3364 ,w__3414);
  xnor g__4320(w__3565 ,w__2796 ,w__3369);
  xnor g__4321(w__3564 ,w__3430 ,w__3409);
  xnor g__4322(w__3563 ,w__3328 ,w__3400);
  xnor g__4323(w__3562 ,w__3433 ,w__3385);
  xnor g__4324(w__3561 ,w__3404 ,w__3406);
  xnor g__4325(w__3560 ,w__3387 ,w__3389);
  xnor g__4326(w__3559 ,w__3380 ,w__3381);
  xnor g__4327(w__3558 ,w__3437 ,w__3419);
  xnor g__4328(w__3557 ,w__3388 ,w__3392);
  xnor g__4329(w__3556 ,w__3308 ,w__3365);
  xnor g__4330(w__3555 ,w__3325 ,w__3305);
  xnor g__4331(w__3608 ,w__3361 ,w__3283);
  xnor g__4332(w__3607 ,w__3277 ,w__3343);
  xnor g__4333(w__3606 ,w__3285 ,w__3339);
  xnor g__4334(w__3605 ,w__3287 ,w__3349);
  xnor g__4335(w__3604 ,w__3281 ,w__3346);
  xnor g__4336(w__3603 ,w__3279 ,w__3358);
  not g__4337(w__3552 ,w__3553);
  or g__4338(w__3551 ,w__2620 ,w__3401);
  and g__4339(w__3550 ,w__3396 ,w__3326);
  or g__4340(w__3549 ,w__2621 ,w__3420);
  or g__4341(w__3548 ,w__3402 ,w__3407);
  and g__4342(w__3547 ,w__2813 ,w__3420);
  or g__4343(w__3546 ,w__2630 ,w__3414);
  or g__4344(w__3545 ,w__2628 ,w__3419);
  or g__4345(w__3544 ,w__3412 ,w__3391);
  and g__4346(w__3543 ,w__2815 ,w__3419);
  or g__4347(w__3542 ,w__3050 ,w__3408);
  and g__4348(w__3541 ,w__3050 ,w__3408);
  or g__4349(w__3540 ,w__3405 ,w__3390);
  or g__4350(w__3539 ,w__3385 ,w__3422);
  and g__4351(w__3538 ,w__3405 ,w__3390);
  nor g__4352(w__3537 ,w__3418 ,w__3416);
  and g__4353(w__3536 ,w__3385 ,w__3422);
  and g__4354(w__3535 ,w__3412 ,w__3391);
  or g__4355(w__3534 ,w__2626 ,w__3413);
  and g__4356(w__3533 ,w__3318 ,w__3322);
  or g__4357(w__3532 ,w__3417 ,w__3415);
  or g__4358(w__3531 ,w__3411 ,w__3409);
  or g__4359(w__3530 ,w__3304 ,w__3324);
  and g__4360(w__3529 ,w__2812 ,w__3413);
  and g__4361(w__3528 ,w__3411 ,w__3409);
  or g__4362(w__3527 ,w__3400 ,w__3328);
  or g__4363(w__3526 ,w__3403 ,w__3397);
  or g__4364(w__3525 ,w__3406 ,w__3404);
  and g__4365(w__3524 ,w__3315 ,w__3378);
  and g__4366(w__3523 ,w__3400 ,w__3328);
  and g__4367(w__3522 ,w__3323 ,w__3321);
  or g__4368(w__3521 ,w__3396 ,w__3326);
  and g__4369(w__3520 ,w__3406 ,w__3404);
  and g__4370(w__3519 ,w__2625 ,w__3320);
  and g__4371(w__3518 ,w__3386 ,w__3382);
  or g__4372(w__3517 ,w__3048 ,w__3330);
  and g__4373(w__3516 ,w__2817 ,w__3401);
  and g__4374(w__3515 ,w__3048 ,w__3330);
  or g__4375(w__3514 ,w__3399 ,w__3398);
  or g__4376(w__3513 ,w__3384 ,w__3302);
  and g__4377(w__3512 ,w__3399 ,w__3398);
  or g__4378(w__3511 ,w__2624 ,w__3395);
  and g__4379(w__3510 ,w__3053 ,w__3336);
  and g__4380(w__3509 ,w__2787 ,w__3395);
  and g__4381(w__3508 ,w__3381 ,w__3380);
  or g__4382(w__3507 ,w__2552 ,w__3383);
  or g__4383(w__3506 ,w__3392 ,w__3388);
  or g__4384(w__3505 ,w__3389 ,w__3387);
  or g__4385(w__3504 ,w__3386 ,w__3382);
  and g__4386(w__3503 ,w__3389 ,w__3387);
  and g__4387(w__3502 ,w__3403 ,w__3397);
  and g__4388(w__3501 ,w__3392 ,w__3388);
  or g__4389(w__3500 ,w__3381 ,w__3380);
  and g__4390(w__3554 ,w__3282 ,w__3347);
  and g__4391(w__3553 ,w__3284 ,w__3362);
  not g__4392(w__3497 ,w__3498);
  not g__4393(w__3496 ,w__3495);
  not g__4394(w__3494 ,w__3493);
  or g__4395(w__3492 ,w__3372 ,w__3379);
  and g__4396(w__3491 ,w__2785 ,w__3300);
  or g__4397(w__3490 ,w__3047 ,w__3377);
  and g__4398(w__3489 ,w__3047 ,w__3377);
  and g__4399(w__3488 ,w__3372 ,w__3379);
  and g__4400(w__3487 ,w__3402 ,w__3407);
  or g__4401(w__3486 ,w__3049 ,w__3421);
  or g__4402(w__3485 ,w__2622 ,w__3310);
  nor g__4403(w__3484 ,w__2785 ,w__3300);
  or g__4404(w__3483 ,w__3332 ,w__3299);
  and g__4405(w__3482 ,w__2786 ,w__3310);
  or g__4406(w__3481 ,w__3306 ,w__3331);
  and g__4407(w__3480 ,w__3332 ,w__3299);
  and g__4408(w__3479 ,w__2794 ,w__3414);
  and g__4409(w__3478 ,w__3306 ,w__3331);
  and g__4410(w__3477 ,w__3049 ,w__3421);
  nor g__4411(w__3476 ,w__3305 ,w__3325);
  and g__4412(w__3475 ,w__3319 ,w__3335);
  or g__4413(w__3474 ,w__2791 ,w__3320);
  or g__4414(w__3473 ,w__3309 ,w__3307);
  or g__4415(w__3472 ,w__3051 ,w__3303);
  and g__4416(w__3471 ,w__3051 ,w__3303);
  and g__4417(w__3470 ,w__3314 ,w__3294);
  and g__4418(w__3469 ,w__3384 ,w__3302);
  nor g__4419(w__3468 ,w__3053 ,w__3336);
  and g__4420(w__3467 ,w__3329 ,w__3296);
  or g__4421(w__3466 ,w__3314 ,w__3294);
  or g__4422(w__3465 ,w__3297 ,w__3337);
  or g__4423(w__3464 ,w__3329 ,w__3296);
  or g__4424(w__3463 ,w__3318 ,w__3322);
  and g__4425(w__3462 ,w__2552 ,w__3383);
  and g__4426(w__3461 ,w__3309 ,w__3307);
  or g__4427(w__3460 ,w__3323 ,w__3321);
  nor g__4428(w__3459 ,w__2793 ,w__3334);
  nor g__4429(w__3458 ,w__3298 ,w__3338);
  or g__4430(w__3457 ,w__3315 ,w__3378);
  and g__4431(w__3456 ,w__3317 ,w__3308);
  or g__4432(w__3455 ,w__3317 ,w__3308);
  or g__4433(w__3454 ,w__3319 ,w__3335);
  or g__4434(w__3453 ,w__2789 ,w__3312);
  and g__4435(w__3452 ,w__2631 ,w__3316);
  or g__4436(w__3451 ,w__2627 ,w__3311);
  nor g__4437(w__3450 ,w__2790 ,w__3313);
  nor g__4438(w__3449 ,w__2631 ,w__3316);
  and g__4439(w__3448 ,w__2816 ,w__3311);
  or g__4440(w__3447 ,w__2629 ,w__2554);
  and g__4441(w__3446 ,w__2818 ,w__2554);
  or g__4442(w__3445 ,w__2623 ,w__2548);
  and g__4443(w__3444 ,w__2788 ,w__3291);
  or g__4444(w__3443 ,w__2792 ,w__3333);
  and g__4445(w__13559 ,w__3290 ,w__3368);
  and g__4446(w__3499 ,w__3288 ,w__3350);
  and g__4447(w__3498 ,w__3280 ,w__3359);
  and g__4448(w__3495 ,w__3286 ,w__3340);
  and g__4449(w__3493 ,w__3278 ,w__3343);
  not g__4450(w__3417 ,w__3418);
  not g__4451(w__3415 ,w__3416);
  not g__4452(w__3393 ,w__3394);
  not g__4453(w__3374 ,w__3375);
  not g__4454(w__3372 ,w__3373);
  not g__4455(w__3371 ,w__3370);
  or g__4456(w__3369 ,w__3060 ,w__3163);
  and g__4457(w__3442 ,w__3088 ,w__3192);
  and g__4458(w__3441 ,w__3111 ,w__3166);
  and g__4459(w__3440 ,w__3122 ,w__3205);
  and g__4460(w__3439 ,w__2999 ,w__3156);
  and g__4461(w__3438 ,w__3011 ,w__3169);
  and g__4462(w__3437 ,w__3110 ,w__3238);
  and g__4463(w__3436 ,w__3107 ,w__3239);
  and g__4464(w__3435 ,w__3106 ,w__3234);
  and g__4465(w__3434 ,w__2993 ,w__3144);
  and g__4466(w__3433 ,w__3104 ,w__3165);
  and g__4467(w__3432 ,w__3096 ,w__3220);
  and g__4468(w__3431 ,w__3098 ,w__3227);
  and g__4469(w__3430 ,w__3117 ,w__3225);
  and g__4470(w__3429 ,w__3093 ,w__3223);
  and g__4471(w__3428 ,w__3067 ,w__3218);
  and g__4472(w__3427 ,w__3102 ,w__3202);
  and g__4473(w__3426 ,w__3078 ,w__3275);
  and g__4474(w__3425 ,w__3082 ,w__3211);
  and g__4475(w__3424 ,w__3087 ,w__3184);
  and g__4476(w__3423 ,w__3037 ,w__3251);
  and g__4477(w__3422 ,w__3109 ,w__3237);
  and g__4478(w__3421 ,w__3030 ,w__3190);
  and g__4479(w__3420 ,w__3074 ,w__3249);
  or g__4480(w__3419 ,w__3056 ,w__3162);
  and g__4481(w__3418 ,w__3021 ,w__3232);
  and g__4482(w__3416 ,w__3023 ,w__3231);
  or g__4483(w__3414 ,w__3065 ,w__3159);
  and g__4484(w__3413 ,w__3100 ,w__3228);
  or g__4485(w__3412 ,w__3063 ,w__3161);
  and g__4486(w__3411 ,w__3115 ,w__3229);
  and g__4487(w__3410 ,w__3116 ,w__3246);
  and g__4488(w__3409 ,w__3099 ,w__3226);
  and g__4489(w__3408 ,w__3113 ,w__3245);
  and g__4490(w__3407 ,w__3079 ,w__3203);
  and g__4491(w__3406 ,w__3094 ,w__3170);
  and g__4492(w__3405 ,w__3008 ,w__3242);
  and g__4493(w__3404 ,w__2994 ,w__3152);
  or g__4494(w__3403 ,w__3058 ,w__3160);
  and g__4495(w__3402 ,w__3075 ,w__3204);
  and g__4496(w__3401 ,w__3003 ,w__3151);
  and g__4497(w__3400 ,w__3009 ,w__3224);
  and g__4498(w__3399 ,w__3086 ,w__3216);
  and g__4499(w__3398 ,w__3085 ,w__3215);
  and g__4500(w__3397 ,w__3001 ,w__3153);
  and g__4501(w__3396 ,w__3013 ,w__3188);
  and g__4502(w__3395 ,w__3024 ,w__3254);
  and g__4503(w__3394 ,w__3080 ,w__3262);
  and g__4504(w__3392 ,w__3027 ,w__3268);
  and g__4505(w__3391 ,w__3108 ,w__3240);
  and g__4506(w__3390 ,w__3083 ,w__3276);
  and g__4507(w__3389 ,w__3070 ,w__3250);
  and g__4508(w__3388 ,w__3077 ,w__3272);
  and g__4509(w__3387 ,w__3040 ,w__3141);
  or g__4510(w__3386 ,w__3054 ,w__3158);
  or g__4511(w__3385 ,w__3061 ,w__3157);
  and g__4512(w__3384 ,w__3039 ,w__3172);
  and g__4513(w__3383 ,w__2995 ,w__3155);
  and g__4514(w__3382 ,w__3068 ,w__3208);
  and g__4515(w__3381 ,w__3031 ,w__3201);
  and g__4516(w__3380 ,w__3069 ,w__3209);
  and g__4517(w__3379 ,w__3000 ,w__3148);
  and g__4518(w__3378 ,w__3026 ,w__3213);
  and g__4519(w__3377 ,w__3119 ,w__3207);
  and g__4520(w__3376 ,w__3114 ,w__3206);
  and g__4521(w__3375 ,w__3005 ,w__3154);
  and g__4522(w__3373 ,w__3091 ,w__3222);
  and g__4523(w__3370 ,w__3072 ,w__3210);
  not g__4524(w__3362 ,w__3361);
  not g__4525(w__3359 ,w__3358);
  not g__4526(w__3350 ,w__3349);
  not g__4527(w__3347 ,w__3346);
  not g__4528(w__3340 ,w__3339);
  not g__4529(w__3337 ,w__3338);
  not g__4530(w__3333 ,w__3334);
  not g__4531(w__3324 ,w__3325);
  not g__4532(w__3312 ,w__3313);
  not g__4533(w__3304 ,w__3305);
  not g__4534(w__3297 ,w__3298);
  not g__4535(w__3294 ,w__3293);
  not g__4536(w__3292 ,w__3291);
  or g__4537(w__13624 ,w__3134 ,w__3265);
  or g__4538(w__13625 ,w__3128 ,w__3241);
  or g__4539(w__13560 ,w__3120 ,w__3175);
  or g__4540(w__3368 ,w__3135 ,w__3257);
  and g__4541(w__3367 ,w__3089 ,w__3221);
  and g__4542(w__3366 ,w__3081 ,w__3185);
  and g__4543(w__3365 ,w__3138 ,w__3247);
  and g__4544(w__3364 ,w__2997 ,w__3150);
  and g__4545(w__3363 ,w__3018 ,w__3176);
  and g__4546(w__3361 ,w__3032 ,w__3267);
  and g__4547(w__3360 ,w__3125 ,w__3263);
  and g__4548(w__3358 ,w__3124 ,w__3256);
  and g__4549(w__3357 ,w__3007 ,w__3147);
  and g__4550(w__3356 ,w__3062 ,w__3260);
  and g__4551(w__3355 ,w__2996 ,w__3145);
  and g__4552(w__3354 ,w__3090 ,w__3253);
  and g__4553(w__3353 ,w__3136 ,w__3273);
  and g__4554(w__3352 ,w__3137 ,w__3261);
  and g__4555(w__3351 ,w__3132 ,w__3270);
  and g__4556(w__3349 ,w__3131 ,w__3269);
  and g__4557(w__3348 ,w__3133 ,w__3264);
  and g__4558(w__3346 ,w__3129 ,w__3271);
  and g__4559(w__3345 ,w__3127 ,w__3266);
  and g__4560(w__3344 ,w__3126 ,w__3274);
  or g__4561(w__3343 ,w__3101 ,w__3259);
  and g__4562(w__3342 ,w__3130 ,w__3258);
  and g__4563(w__3341 ,w__2998 ,w__3146);
  and g__4564(w__3339 ,w__3071 ,w__3198);
  and g__4565(w__3338 ,w__3076 ,w__3177);
  and g__4566(w__3336 ,w__3020 ,w__3179);
  and g__4567(w__3335 ,w__3084 ,w__3243);
  or g__4568(w__3334 ,w__2795 ,w__3255);
  and g__4569(w__3332 ,w__3092 ,w__3197);
  and g__4570(w__3331 ,w__3112 ,w__3233);
  and g__4571(w__3330 ,w__3038 ,w__3219);
  and g__4572(w__3329 ,w__3010 ,w__3230);
  and g__4573(w__3328 ,w__3033 ,w__3193);
  and g__4574(w__3327 ,w__3034 ,w__3191);
  and g__4575(w__3326 ,w__3118 ,w__3195);
  and g__4576(w__3325 ,w__3022 ,w__3194);
  and g__4577(w__3323 ,w__3019 ,w__3167);
  and g__4578(w__3322 ,w__3014 ,w__3248);
  and g__4579(w__3321 ,w__3004 ,w__3212);
  and g__4580(w__3320 ,w__3028 ,w__3171);
  and g__4581(w__3319 ,w__3017 ,w__3199);
  and g__4582(w__3318 ,w__3012 ,w__3168);
  and g__4583(w__3317 ,w__3097 ,w__3244);
  and g__4584(w__3316 ,w__3066 ,w__3252);
  and g__4585(w__3315 ,w__3055 ,w__3236);
  and g__4586(w__3314 ,w__3059 ,w__3217);
  and g__4587(w__3313 ,w__3064 ,w__3235);
  and g__4588(w__3311 ,w__3057 ,w__3174);
  and g__4589(w__3310 ,w__3036 ,w__3200);
  and g__4590(w__3309 ,w__3121 ,w__3187);
  and g__4591(w__3308 ,w__3006 ,w__3142);
  and g__4592(w__3307 ,w__3035 ,w__3186);
  or g__4593(w__3306 ,w__2795 ,w__3164);
  and g__4594(w__3305 ,w__3029 ,w__3189);
  and g__4595(w__3303 ,w__3095 ,w__3182);
  and g__4596(w__3302 ,w__3073 ,w__3181);
  and g__4597(w__3301 ,w__3103 ,w__3180);
  or g__4598(w__3300 ,w__3060 ,w__3149);
  and g__4599(w__3299 ,w__3105 ,w__3196);
  and g__4600(w__3298 ,w__3123 ,w__3178);
  and g__4601(w__3296 ,w__3002 ,w__3143);
  and g__4602(w__3295 ,w__3015 ,w__3183);
  and g__4603(w__3293 ,w__3016 ,w__3214);
  and g__4604(w__3291 ,w__3025 ,w__3173);
  not g__4605(w__3290 ,w__3289);
  not g__4606(w__3288 ,w__3287);
  not g__4607(w__3286 ,w__3285);
  not g__4608(w__3284 ,w__3283);
  not g__4609(w__3282 ,w__3281);
  not g__4610(w__3280 ,w__3279);
  not g__4611(w__3278 ,w__3277);
  or g__4612(w__3276 ,w__2880 ,w__2466);
  or g__4613(w__3275 ,w__2894 ,w__2451);
  or g__4614(w__3274 ,w__2856 ,w__2425);
  or g__4615(w__3273 ,w__2844 ,w__2517);
  or g__4616(w__3272 ,w__2952 ,w__2448);
  or g__4617(w__3271 ,w__2849 ,w__2425);
  or g__4618(w__3270 ,w__2851 ,w__2492);
  or g__4619(w__3269 ,w__2845 ,w__2513);
  or g__4620(w__3268 ,w__2842 ,w__2508);
  or g__4621(w__3267 ,w__2877 ,w__2444);
  or g__4622(w__3266 ,w__2853 ,w__2514);
  nor g__4623(w__3265 ,w__2516 ,w__2846);
  or g__4624(w__3264 ,w__2847 ,w__2492);
  or g__4625(w__3263 ,w__2852 ,w__2493);
  or g__4626(w__3262 ,w__2848 ,w__2505);
  or g__4627(w__3261 ,w__2854 ,w__2516);
  or g__4628(w__3260 ,w__2903 ,w__2510);
  nor g__4629(w__3259 ,w__2514 ,w__2858);
  or g__4630(w__3258 ,w__2855 ,w__2544);
  nor g__4631(w__3257 ,w__2517 ,w__2857);
  or g__4632(w__3256 ,w__2850 ,w__2543);
  nor g__4633(w__3255 ,w__2513 ,w__2843);
  or g__4634(w__3254 ,w__2973 ,w__2457);
  or g__4635(w__3253 ,w__2929 ,w__2436);
  or g__4636(w__3252 ,w__2930 ,w__2484);
  or g__4637(w__3251 ,w__2975 ,w__2463);
  or g__4638(w__3250 ,w__2939 ,w__2460);
  or g__4639(w__3249 ,w__2904 ,w__2478);
  or g__4640(w__3248 ,w__2862 ,w__2507);
  or g__4641(w__3247 ,w__2867 ,w__2439);
  or g__4642(w__3246 ,w__2934 ,w__2483);
  or g__4643(w__3245 ,w__2956 ,w__2525);
  or g__4644(w__3244 ,w__2891 ,w__2519);
  or g__4645(w__3243 ,w__2945 ,w__2442);
  or g__4646(w__3242 ,w__2970 ,w__2481);
  nor g__4647(w__3241 ,w__2493 ,w__2820);
  or g__4648(w__3240 ,w__2951 ,w__2537);
  or g__4649(w__3239 ,w__2935 ,w__2477);
  or g__4650(w__3238 ,w__2899 ,w__2438);
  or g__4651(w__3237 ,w__2869 ,w__2522);
  or g__4652(w__3236 ,w__2961 ,w__2504);
  or g__4653(w__3235 ,w__2953 ,w__2433);
  or g__4654(w__3234 ,w__2946 ,w__2441);
  or g__4655(w__3233 ,w__2955 ,w__2460);
  or g__4656(w__3232 ,w__2976 ,w__2436);
  or g__4657(w__3231 ,w__2947 ,w__2462);
  or g__4658(w__3230 ,w__2879 ,w__2459);
  or g__4659(w__3229 ,w__2822 ,w__2435);
  or g__4660(w__3228 ,w__2943 ,w__2451);
  or g__4661(w__3227 ,w__2944 ,w__2480);
  or g__4662(w__3226 ,w__2948 ,w__2450);
  or g__4663(w__3225 ,w__2938 ,w__2534);
  or g__4664(w__3224 ,w__2974 ,w__2528);
  or g__4665(w__3223 ,w__2936 ,w__2459);
  or g__4666(w__3222 ,w__2933 ,w__2442);
  or g__4667(w__3221 ,w__2887 ,w__2450);
  or g__4668(w__3220 ,w__2885 ,w__2435);
  or g__4669(w__3219 ,w__2895 ,w__2432);
  or g__4670(w__3218 ,w__2897 ,w__2510);
  or g__4671(w__3217 ,w__2861 ,w__2477);
  or g__4672(w__3216 ,w__2940 ,w__2463);
  or g__4673(w__3215 ,w__2959 ,w__2522);
  or g__4674(w__3214 ,w__2937 ,w__2507);
  or g__4675(w__3213 ,w__2900 ,w__2448);
  or g__4676(w__3289 ,w__2780 ,w__2991);
  or g__4677(w__3287 ,w__2805 ,w__2988);
  or g__4678(w__3285 ,w__2773 ,w__2989);
  or g__4679(w__3283 ,w__2778 ,w__2987);
  or g__4680(w__3281 ,w__2776 ,w__2986);
  or g__4681(w__3279 ,w__2781 ,w__2992);
  or g__4682(w__3277 ,w__2770 ,w__2990);
  or g__4683(w__3212 ,w__2915 ,w__2468);
  or g__4684(w__3211 ,w__2876 ,w__2439);
  or g__4685(w__3210 ,w__2882 ,w__2483);
  or g__4686(w__3209 ,w__2892 ,w__2456);
  or g__4687(w__3208 ,w__2884 ,w__2447);
  or g__4688(w__3207 ,w__2962 ,w__2447);
  or g__4689(w__3206 ,w__2957 ,w__2433);
  or g__4690(w__3205 ,w__2905 ,w__2419);
  or g__4691(w__3204 ,w__2893 ,w__2441);
  or g__4692(w__3203 ,w__2965 ,w__2466);
  or g__4693(w__3202 ,w__2870 ,w__2519);
  or g__4694(w__3201 ,w__2823 ,w__2462);
  or g__4695(w__3200 ,w__2890 ,w__2526);
  or g__4696(w__3199 ,w__2941 ,w__2537);
  or g__4697(w__3198 ,w__2963 ,w__2445);
  or g__4698(w__3197 ,w__2910 ,w__2421);
  or g__4699(w__3196 ,w__2860 ,w__2480);
  or g__4700(w__3195 ,w__2968 ,w__2465);
  or g__4701(w__3194 ,w__2875 ,w__2419);
  or g__4702(w__3193 ,w__2859 ,w__2495);
  or g__4703(w__3192 ,w__2901 ,w__2465);
  or g__4704(w__3191 ,w__2883 ,w__2457);
  or g__4705(w__3190 ,w__2872 ,w__2528);
  or g__4706(w__3189 ,w__2889 ,w__2504);
  or g__4707(w__3188 ,w__2871 ,w__2421);
  or g__4708(w__3187 ,w__2819 ,w__2432);
  or g__4709(w__3186 ,w__2972 ,w__2496);
  or g__4710(w__3185 ,w__2873 ,w__2495);
  or g__4711(w__3184 ,w__2865 ,w__2534);
  or g__4712(w__3183 ,w__2932 ,w__2523);
  or g__4713(w__3182 ,w__2886 ,w__2445);
  or g__4714(w__3181 ,w__2942 ,w__2456);
  or g__4715(w__3180 ,w__2950 ,w__2413);
  or g__4716(w__3179 ,w__2881 ,w__2511);
  or g__4717(w__3178 ,w__2907 ,w__2413);
  or g__4718(w__3177 ,w__2971 ,w__2444);
  or g__4719(w__3176 ,w__2866 ,w__2417);
  nor g__4720(w__3175 ,w__2511 ,w__2912);
  or g__4721(w__3174 ,w__2896 ,w__2423);
  or g__4722(w__3173 ,w__2969 ,w__2423);
  or g__4723(w__3172 ,w__2898 ,w__2520);
  or g__4724(w__3171 ,w__2888 ,w__2438);
  or g__4725(w__3170 ,w__2864 ,w__2411);
  or g__4726(w__3169 ,w__2863 ,w__2525);
  or g__4727(w__3168 ,w__2978 ,w__2411);
  or g__4728(w__3167 ,w__2874 ,w__2417);
  or g__4729(w__3166 ,w__2878 ,w__2538);
  or g__4730(w__3165 ,w__2868 ,w__2535);
  nor g__4731(w__3164 ,w__2544 ,w__2746);
  nor g__4732(w__3163 ,w__2502 ,w__2472);
  nor g__4733(w__3162 ,w__2508 ,w__2757);
  nor g__4734(w__3161 ,w__2481 ,w__2760);
  nor g__4735(w__3160 ,w__2478 ,w__2758);
  nor g__4736(w__3159 ,w__2484 ,w__2745);
  nor g__4737(w__3158 ,w__2505 ,w__2759);
  nor g__4738(w__3157 ,w__2496 ,w__2761);
  or g__4739(w__3156 ,w__2967 ,w__2469);
  or g__4740(w__3155 ,w__2964 ,w__2474);
  or g__4741(w__3154 ,w__2958 ,w__2471);
  or g__4742(w__3153 ,w__2966 ,w__2468);
  or g__4743(w__3152 ,w__2954 ,w__2469);
  or g__4744(w__3151 ,w__2980 ,w__2409);
  or g__4745(w__3150 ,w__2931 ,w__2541);
  nor g__4746(w__3149 ,w__2475 ,w__2949);
  or g__4747(w__3148 ,w__2960 ,w__2474);
  or g__4748(w__3147 ,w__2977 ,w__2471);
  or g__4749(w__3146 ,w__2982 ,w__2475);
  or g__4750(w__3145 ,w__2983 ,w__2540);
  or g__4751(w__3144 ,w__2981 ,w__2540);
  or g__4752(w__3143 ,w__2984 ,w__2472);
  or g__4753(w__3142 ,w__2979 ,w__2409);
  or g__4754(w__3141 ,w__2902 ,w__2529);
  or g__4755(w__3138 ,w__2951 ,w__2669);
  or g__4756(w__3137 ,w__2499 ,w__2845);
  or g__4757(w__3136 ,w__2487 ,w__2850);
  nor g__4758(w__3135 ,w__2499 ,w__2855);
  nor g__4759(w__3134 ,w__2487 ,w__2857);
  or g__4760(w__3133 ,w__2486 ,w__2851);
  or g__4761(w__3132 ,w__2498 ,w__2849);
  or g__4762(w__3131 ,w__2489 ,w__2852);
  or g__4763(w__3130 ,w__2498 ,w__2858);
  or g__4764(w__3129 ,w__2486 ,w__2844);
  nor g__4765(w__3128 ,w__2490 ,w__2846);
  or g__4766(w__3127 ,w__2489 ,w__2856);
  or g__4767(w__3126 ,w__2490 ,w__2847);
  or g__4768(w__3125 ,w__2427 ,w__2853);
  or g__4769(w__3124 ,w__2427 ,w__2843);
  or g__4770(w__3123 ,w__2950 ,w__2708);
  or g__4771(w__3122 ,w__2877 ,w__2693);
  or g__4772(w__3121 ,w__2872 ,w__2657);
  nor g__4773(w__3120 ,w__2881 ,w__2700);
  or g__4774(w__3119 ,w__2902 ,w__2666);
  or g__4775(w__3118 ,w__2942 ,w__2711);
  or g__4776(w__3117 ,w__2880 ,w__2711);
  or g__4777(w__3116 ,w__2885 ,w__2678);
  or g__4778(w__3115 ,w__2976 ,w__2678);
  or g__4779(w__3114 ,w__2952 ,w__2666);
  or g__4780(w__3113 ,w__2863 ,w__2699);
  or g__4781(w__3112 ,w__2933 ,w__2681);
  or g__4782(w__3111 ,w__2882 ,w__2670);
  or g__4783(w__3110 ,w__2930 ,w__2673);
  or g__4784(w__3109 ,w__2904 ,w__2687);
  or g__4785(w__3108 ,w__2888 ,w__2669);
  or g__4786(w__3107 ,w__2871 ,w__2687);
  or g__4787(w__3106 ,w__2861 ,w__2682);
  or g__4788(w__3105 ,w__2962 ,w__2658);
  or g__4789(w__3104 ,w__2961 ,w__2709);
  or g__4790(w__3103 ,w__2865 ,w__2708);
  or g__4791(w__3102 ,w__2891 ,w__2633);
  nor g__4792(w__3101 ,w__2572 ,w__2854);
  or g__4793(w__3100 ,w__2969 ,w__2642);
  or g__4794(w__3099 ,w__2947 ,w__2642);
  or g__4795(w__3098 ,w__2900 ,w__2661);
  or g__4796(w__3097 ,w__2887 ,w__2634);
  or g__4797(w__3096 ,w__2978 ,w__2672);
  or g__4798(w__3095 ,w__2972 ,w__2694);
  or g__4799(w__3094 ,w__2929 ,w__2675);
  or g__4800(w__3093 ,w__2935 ,w__2685);
  or g__4801(w__3092 ,w__2893 ,w__2681);
  or g__4802(w__3091 ,w__2869 ,w__2684);
  or g__4803(w__3090 ,w__2941 ,w__2675);
  or g__4804(w__3089 ,w__2937 ,w__2637);
  or g__4805(w__3088 ,w__2973 ,w__2705);
  or g__4806(w__3087 ,w__2889 ,w__2836);
  or g__4807(w__3086 ,w__2948 ,w__2633);
  or g__4808(w__3085 ,w__2936 ,w__2690);
  or g__4809(w__3084 ,w__2932 ,w__2690);
  or g__4810(w__3083 ,w__2968 ,w__2705);
  or g__4811(w__3082 ,w__2864 ,w__2672);
  or g__4812(w__3081 ,w__2890 ,w__2697);
  or g__4813(w__3080 ,w__2938 ,w__2706);
  or g__4814(w__3079 ,w__2892 ,w__2709);
  or g__4815(w__3078 ,w__2896 ,w__2636);
  or g__4816(w__3077 ,w__2944 ,w__2657);
  or g__4817(w__3076 ,w__2886 ,w__2693);
  or g__4818(w__3075 ,w__2939 ,w__2684);
  or g__4819(w__3074 ,w__2945 ,w__2688);
  or g__4820(w__3073 ,w__2901 ,w__2712);
  or g__4821(w__3072 ,w__2899 ,w__2679);
  or g__4822(w__3071 ,w__2905 ,w__2696);
  or g__4823(w__3070 ,w__2959 ,w__2685);
  or g__4824(w__3069 ,w__2848 ,w__2602);
  or g__4825(w__3068 ,w__2953 ,w__2660);
  or g__4826(w__3067 ,w__2859 ,w__2703);
  or g__4827(w__3140 ,w__2825 ,w__2561);
  or g__4828(w__3139 ,in2[0] ,w__2914);
  not g__4829(w__3066 ,w__3065);
  not g__4830(w__3064 ,w__3063);
  not g__4831(w__3062 ,w__3061);
  not g__4832(w__3059 ,w__3058);
  not g__4833(w__3057 ,w__3056);
  not g__4834(w__3055 ,w__3054);
  not g__4835(w__3053 ,w__3052);
  or g__4836(w__3040 ,w__2895 ,w__2663);
  or g__4837(w__3039 ,w__2862 ,w__2639);
  or g__4838(w__3038 ,w__2974 ,w__2663);
  or g__4839(w__3037 ,w__2898 ,w__2639);
  or g__4840(w__3036 ,w__2903 ,w__2702);
  or g__4841(w__3035 ,w__2875 ,w__2696);
  or g__4842(w__3034 ,w__2965 ,w__2602);
  or g__4843(w__3033 ,w__2956 ,w__2699);
  or g__4844(w__3032 ,w__2897 ,w__2697);
  or g__4845(w__3031 ,w__2940 ,w__2636);
  or g__4846(w__3030 ,w__2860 ,w__2660);
  or g__4847(w__3029 ,w__2883 ,w__2712);
  or g__4848(w__3028 ,w__2878 ,w__2673);
  or g__4849(w__3027 ,w__2943 ,w__2643);
  or g__4850(w__3026 ,w__2884 ,w__2667);
  or g__4851(w__3025 ,w__2870 ,w__2637);
  or g__4852(w__3024 ,w__2868 ,w__2706);
  or g__4853(w__3023 ,w__2975 ,w__2640);
  or g__4854(w__3022 ,w__2963 ,w__2702);
  or g__4855(w__3021 ,w__2934 ,w__2676);
  or g__4856(w__3020 ,w__2971 ,w__2694);
  or g__4857(w__3019 ,w__2866 ,w__2661);
  or g__4858(w__3018 ,w__2957 ,w__2664);
  or g__4859(w__3017 ,w__2867 ,w__2670);
  or g__4860(w__3016 ,w__2894 ,w__2634);
  or g__4861(w__3015 ,w__2946 ,w__2691);
  or g__4862(w__3014 ,w__2842 ,w__2643);
  or g__4863(w__3013 ,w__2879 ,w__2682);
  or g__4864(w__3012 ,w__2876 ,w__2679);
  or g__4865(w__3011 ,w__2873 ,w__2700);
  or g__4866(w__3010 ,w__2955 ,w__2688);
  or g__4867(w__3009 ,w__2970 ,w__2658);
  or g__4868(w__3008 ,w__2874 ,w__2667);
  or g__4869(w__3007 ,w__2645 ,w__2964);
  or g__4870(w__3006 ,w__2654 ,w__2980);
  or g__4871(w__3005 ,w__2654 ,w__2931);
  or g__4872(w__3004 ,w__2646 ,w__2984);
  or g__4873(w__3003 ,w__2649 ,w__2981);
  or g__4874(w__3002 ,w__2645 ,w__2982);
  or g__4875(w__3001 ,w__2648 ,w__2977);
  or g__4876(w__3000 ,w__2651 ,w__2954);
  or g__4877(w__2999 ,w__2651 ,w__2983);
  or g__4878(w__2998 ,w__2648 ,w__2960);
  or g__4879(w__2997 ,w__2655 ,w__2949);
  or g__4880(w__2996 ,w__2649 ,w__2979);
  or g__4881(w__2995 ,w__2652 ,w__2958);
  or g__4882(w__2994 ,w__2646 ,w__2967);
  or g__4883(w__2993 ,w__2655 ,w__2966);
  or g__4884(w__2992 ,w__2532 ,w__2918);
  or g__4885(w__2991 ,w__2761 ,w__2921);
  or g__4886(w__2990 ,w__2759 ,w__2922);
  or g__4887(w__2989 ,w__2758 ,w__2920);
  or g__4888(w__2988 ,w__2760 ,w__2916);
  or g__4889(w__2987 ,w__2757 ,w__2917);
  or g__4890(w__2986 ,w__2745 ,w__2919);
  nor g__4891(w__2985 ,w__2703 ,w__2398);
  and g__4892(w__3065 ,in2[13] ,w__2564);
  and g__4893(w__3063 ,in2[7] ,w__2562);
  and g__4894(w__3061 ,in2[3] ,w__2555);
  and g__4895(w__3060 ,in2[15] ,w__2563);
  and g__4896(w__3058 ,in2[9] ,w__2566);
  and g__4897(w__3056 ,in2[11] ,w__2560);
  and g__4898(w__3054 ,in2[5] ,w__2556);
  and g__4899(w__3052 ,in1[0] ,w__2570);
  or g__4900(w__3051 ,w__2546 ,w__2664);
  or g__4901(w__3050 ,w__2546 ,w__2652);
  or g__4902(w__3049 ,w__2762 ,w__2691);
  or g__4903(w__3048 ,w__2545 ,w__2676);
  or g__4904(w__3047 ,w__2545 ,w__2640);
  or g__4905(w__3046 ,w__2913 ,w__2558);
  or g__4906(w__3045 ,w__2908 ,w__2567);
  or g__4907(w__3044 ,w__2906 ,w__2557);
  or g__4908(w__3043 ,w__2821 ,w__2569);
  or g__4909(w__3042 ,w__2909 ,w__2565);
  or g__4910(w__3041 ,w__2824 ,w__2559);
  not g__4911(w__2928 ,w__2562);
  not g__4912(w__2927 ,w__2567);
  not g__4913(w__2925 ,w__2561);
  not g__4914(w__2924 ,w__2563);
  nor g__4915(w__2922 ,w__2610 ,w__2808);
  nor g__4916(w__2921 ,w__2746 ,w__2771);
  nor g__4917(w__2920 ,w__2608 ,w__2777);
  nor g__4918(w__2919 ,w__2606 ,w__2810);
  nor g__4919(w__2918 ,w__2604 ,w__2772);
  nor g__4920(w__2917 ,w__2612 ,w__2797);
  nor g__4921(w__2916 ,w__2614 ,w__2802);
  or g__4922(w__2915 ,w__2793 ,w__2782);
  xnor g__4923(w__2913 ,in2[13] ,in2[12]);
  xnor g__4924(w__2912 ,in1[0] ,in2[3]);
  nor g__4925(w__2911 ,w__13563 ,w__2616);
  xnor g__4926(w__2910 ,in1[0] ,in2[9]);
  xnor g__4927(w__2909 ,in2[9] ,in2[8]);
  xnor g__4928(w__2908 ,in2[7] ,in2[6]);
  xnor g__4929(w__2907 ,in1[0] ,in2[5]);
  xnor g__4930(w__2906 ,in2[3] ,in2[2]);
  or g__4931(w__2984 ,w__2714 ,w__2801);
  or g__4932(w__2983 ,w__2789 ,w__2798);
  or g__4933(w__2982 ,w__2715 ,w__2811);
  or g__4934(w__2981 ,w__2725 ,w__2806);
  or g__4935(w__2980 ,w__2717 ,w__2803);
  or g__4936(w__2979 ,w__2724 ,w__2799);
  xnor g__4937(w__2978 ,in1[4] ,in2[13]);
  or g__4938(w__2977 ,w__2722 ,w__2774);
  xnor g__4939(w__2976 ,in1[1] ,in2[13]);
  xnor g__4940(w__2975 ,in1[4] ,in2[11]);
  xnor g__4941(w__2974 ,in1[6] ,in2[7]);
  xnor g__4942(w__2973 ,in1[13] ,in2[5]);
  xnor g__4943(w__2972 ,in1[4] ,in2[3]);
  xnor g__4944(w__2971 ,in1[2] ,in2[3]);
  xnor g__4945(w__2970 ,in1[7] ,in2[7]);
  xnor g__4946(w__2969 ,in1[9] ,in2[11]);
  xnor g__4947(w__2968 ,in1[10] ,in2[5]);
  or g__4948(w__2967 ,w__2716 ,w__2807);
  or g__4949(w__2966 ,w__2723 ,w__2775);
  xnor g__4950(w__2965 ,in1[5] ,in2[5]);
  or g__4951(w__2964 ,w__2721 ,w__2779);
  xnor g__4952(w__2963 ,in1[6] ,in2[3]);
  xnor g__4953(w__2962 ,in1[3] ,in2[7]);
  xnor g__4954(w__2961 ,in1[15] ,in2[5]);
  or g__4955(w__2960 ,w__2719 ,w__2800);
  xnor g__4956(w__2959 ,in1[3] ,in2[9]);
  or g__4957(w__2958 ,w__2718 ,w__2804);
  xnor g__4958(w__2957 ,in1[10] ,in2[7]);
  xnor g__4959(w__2956 ,in1[11] ,in2[3]);
  xnor g__4960(w__2955 ,in1[8] ,in2[9]);
  or g__4961(w__2954 ,w__2720 ,w__2809);
  xnor g__4962(w__2953 ,in1[15] ,in2[7]);
  xnor g__4963(w__2952 ,in1[11] ,in2[7]);
  xnor g__4964(w__2951 ,in1[10] ,in2[13]);
  xnor g__4965(w__2950 ,in1[1] ,in2[5]);
  xnor g__4966(w__2949 ,in1[15] ,in2[15]);
  xnor g__4967(w__2948 ,in1[2] ,in2[11]);
  xnor g__4968(w__2947 ,in1[3] ,in2[11]);
  xnor g__4969(w__2946 ,in1[14] ,in2[9]);
  xnor g__4970(w__2945 ,in1[12] ,in2[9]);
  xnor g__4971(w__2944 ,in1[12] ,in2[7]);
  xnor g__4972(w__2943 ,in1[8] ,in2[11]);
  xnor g__4973(w__2942 ,in1[11] ,in2[5]);
  xnor g__4974(w__2941 ,in1[8] ,in2[13]);
  xnor g__4975(w__2940 ,in1[1] ,in2[11]);
  xnor g__4976(w__2939 ,in1[2] ,in2[9]);
  xnor g__4977(w__2938 ,in1[8] ,in2[5]);
  xnor g__4978(w__2937 ,in1[13] ,in2[11]);
  xnor g__4979(w__2936 ,in1[4] ,in2[9]);
  xnor g__4980(w__2935 ,in1[5] ,in2[9]);
  xnor g__4981(w__2934 ,in1[2] ,in2[13]);
  xnor g__4982(w__2933 ,in1[9] ,in2[9]);
  xnor g__4983(w__2932 ,in1[13] ,in2[9]);
  or g__4984(w__2931 ,w__2600 ,w__2783);
  xnor g__4985(w__2930 ,in1[15] ,in2[13]);
  xnor g__4986(w__2929 ,in1[7] ,in2[13]);
  xnor g__4987(w__2926 ,w__2614 ,in2[6]);
  xnor g__4988(w__2923 ,w__2604 ,in2[14]);
  not g__4989(w__2841 ,w__2560);
  not g__4990(w__2840 ,w__2559);
  not g__4991(w__2838 ,w__2570);
  not g__4992(w__2836 ,w__2556);
  not g__4993(w__2835 ,w__2569);
  not g__4994(w__2834 ,w__2555);
  not g__4995(w__2833 ,w__2557);
  not g__4996(w__2831 ,w__2566);
  not g__4997(w__2830 ,w__2565);
  not g__4998(w__2828 ,w__2564);
  not g__4999(w__2827 ,w__2558);
  xnor g__5000(w__2825 ,in2[15] ,in2[14]);
  xnor g__5001(w__2824 ,in2[11] ,in2[10]);
  xnor g__5002(w__2823 ,in1[0] ,in2[11]);
  xnor g__5003(w__2822 ,in1[0] ,in2[13]);
  xnor g__5004(w__2821 ,in2[5] ,in2[4]);
  xnor g__5005(w__2820 ,in1[0] ,in2[1]);
  xnor g__5006(w__2819 ,in1[0] ,in2[7]);
  xnor g__5007(w__2905 ,in1[7] ,in2[3]);
  xnor g__5008(w__2904 ,in1[11] ,in2[9]);
  xnor g__5009(w__2903 ,in1[15] ,in2[3]);
  xnor g__5010(w__2902 ,in1[4] ,in2[7]);
  xnor g__5011(w__2901 ,in1[12] ,in2[5]);
  xnor g__5012(w__2900 ,in1[13] ,in2[7]);
  xnor g__5013(w__2899 ,in1[14] ,in2[13]);
  xnor g__5014(w__2898 ,in1[5] ,in2[11]);
  xnor g__5015(w__2897 ,in1[9] ,in2[3]);
  xnor g__5016(w__2896 ,in1[15] ,in2[11]);
  xnor g__5017(w__2895 ,in1[5] ,in2[7]);
  xnor g__5018(w__2894 ,in1[14] ,in2[11]);
  xnor g__5019(w__2893 ,in1[1] ,in2[9]);
  xnor g__5020(w__2892 ,in1[6] ,in2[5]);
  xnor g__5021(w__2891 ,in1[11] ,in2[11]);
  xnor g__5022(w__2890 ,in1[14] ,in2[3]);
  xnor g__5023(w__2889 ,in1[3] ,in2[5]);
  xnor g__5024(w__2888 ,in1[11] ,in2[13]);
  xnor g__5025(w__2887 ,in1[12] ,in2[11]);
  xnor g__5026(w__2886 ,in1[3] ,in2[3]);
  xnor g__5027(w__2885 ,in1[3] ,in2[13]);
  xnor g__5028(w__2884 ,in1[14] ,in2[7]);
  xnor g__5029(w__2883 ,in1[4] ,in2[5]);
  xnor g__5030(w__2882 ,in1[13] ,in2[13]);
  xnor g__5031(w__2881 ,in1[1] ,in2[3]);
  xnor g__5032(w__2880 ,in1[9] ,in2[5]);
  xnor g__5033(w__2879 ,in1[7] ,in2[9]);
  xnor g__5034(w__2878 ,in1[12] ,in2[13]);
  xnor g__5035(w__2877 ,in1[8] ,in2[3]);
  xnor g__5036(w__2876 ,in1[5] ,in2[13]);
  xnor g__5037(w__2875 ,in1[5] ,in2[3]);
  xnor g__5038(w__2874 ,in1[8] ,in2[7]);
  xnor g__5039(w__2873 ,in1[13] ,in2[3]);
  xnor g__5040(w__2872 ,in1[1] ,in2[7]);
  xnor g__5041(w__2871 ,in1[6] ,in2[9]);
  xnor g__5042(w__2870 ,in1[10] ,in2[11]);
  xnor g__5043(w__2869 ,in1[10] ,in2[9]);
  xnor g__5044(w__2868 ,in1[14] ,in2[5]);
  xnor g__5045(w__2867 ,in1[9] ,in2[13]);
  xnor g__5046(w__2866 ,in1[9] ,in2[7]);
  xnor g__5047(w__2865 ,in1[2] ,in2[5]);
  xnor g__5048(w__2864 ,in1[6] ,in2[13]);
  xnor g__5049(w__2863 ,in1[12] ,in2[3]);
  xnor g__5050(w__2862 ,in1[6] ,in2[11]);
  xnor g__5051(w__2861 ,in1[15] ,in2[9]);
  xnor g__5052(w__2860 ,in1[2] ,in2[7]);
  xnor g__5053(w__2859 ,in1[10] ,in2[3]);
  xnor g__5054(w__2858 ,in1[4] ,in2[1]);
  xnor g__5055(w__2857 ,in1[2] ,in2[1]);
  xnor g__5056(w__2856 ,in1[9] ,in2[1]);
  xnor g__5057(w__2855 ,in1[3] ,in2[1]);
  xnor g__5058(w__2854 ,in1[5] ,in2[1]);
  xnor g__5059(w__2853 ,in1[8] ,in2[1]);
  xnor g__5060(w__2852 ,in1[7] ,in2[1]);
  xnor g__5061(w__2851 ,in1[11] ,in2[1]);
  xnor g__5062(w__2850 ,in1[14] ,in2[1]);
  xnor g__5063(w__2849 ,in1[12] ,in2[1]);
  xnor g__5064(w__2848 ,in1[7] ,in2[5]);
  xnor g__5065(w__2847 ,in1[10] ,in2[1]);
  xnor g__5066(w__2846 ,in1[1] ,in2[1]);
  xnor g__5067(w__2845 ,in1[6] ,in2[1]);
  xnor g__5068(w__2844 ,in1[13] ,in2[1]);
  xnor g__5069(w__2843 ,in1[15] ,in2[1]);
  xnor g__5070(w__2842 ,in1[7] ,in2[11]);
  xnor g__5071(w__2839 ,w__2612 ,in2[10]);
  xnor g__5072(w__2837 ,w__2610 ,in2[4]);
  xnor g__5073(w__2832 ,w__2616 ,in2[2]);
  xnor g__5074(w__2829 ,w__2608 ,in2[8]);
  xnor g__5075(w__2826 ,w__2606 ,in2[12]);
  nor g__5076(w__2811 ,in1[2] ,in2[15]);
  nor g__5077(w__2810 ,in1[0] ,in2[12]);
  nor g__5078(w__2809 ,in1[4] ,in2[15]);
  nor g__5079(w__2808 ,in1[0] ,in2[4]);
  nor g__5080(w__2807 ,in1[5] ,in2[15]);
  nor g__5081(w__2806 ,in1[9] ,in2[15]);
  and g__5082(w__2805 ,in1[0] ,in2[6]);
  nor g__5083(w__2804 ,in1[13] ,in2[15]);
  nor g__5084(w__2803 ,in1[8] ,in2[15]);
  nor g__5085(w__2802 ,in1[0] ,in2[6]);
  nor g__5086(w__2801 ,in1[1] ,in2[15]);
  nor g__5087(w__2800 ,in1[3] ,in2[15]);
  nor g__5088(w__2799 ,in1[7] ,in2[15]);
  nor g__5089(w__2798 ,in1[6] ,in2[15]);
  nor g__5090(w__2797 ,in1[0] ,in2[10]);
  or g__5091(w__2796 ,w__2766 ,w__2429);
  or g__5092(w__2818 ,w__2768 ,w__2453);
  or g__5093(w__2817 ,w__2769 ,w__2531);
  or g__5094(w__2816 ,w__2751 ,w__2501);
  or g__5095(w__2815 ,w__2755 ,w__2430);
  or g__5096(w__2814 ,w__2764 ,w__2454);
  or g__5097(w__2813 ,w__2763 ,w__2415);
  or g__5098(w__2812 ,w__2754 ,w__2501);
  not g__5099(w__2792 ,w__2793);
  not g__5100(w__2789 ,w__2790);
  not g__5101(w__2784 ,w__2785);
  nor g__5102(w__2783 ,in1[14] ,in2[15]);
  nor g__5103(w__2782 ,in1[0] ,in2[15]);
  and g__5104(w__2781 ,in1[0] ,in2[14]);
  and g__5105(w__2780 ,in1[0] ,in2[2]);
  nor g__5106(w__2779 ,in1[12] ,in2[15]);
  and g__5107(w__2778 ,in1[0] ,in2[10]);
  nor g__5108(w__2777 ,in1[0] ,in2[8]);
  and g__5109(w__2776 ,in1[0] ,in2[12]);
  nor g__5110(w__2775 ,in1[10] ,in2[15]);
  nor g__5111(w__2774 ,in1[11] ,in2[15]);
  and g__5112(w__2773 ,in1[0] ,in2[8]);
  nor g__5113(w__2772 ,in1[0] ,in2[14]);
  nor g__5114(w__2771 ,in1[0] ,in2[2]);
  and g__5115(w__2770 ,in1[0] ,in2[4]);
  and g__5116(w__13563 ,in1[0] ,in2[0]);
  and g__5117(w__2795 ,in2[1] ,in2[0]);
  or g__5118(w__2794 ,w__2752 ,w__2429);
  and g__5119(w__2793 ,in1[0] ,in2[15]);
  or g__5120(w__2791 ,w__2750 ,w__2453);
  or g__5121(w__2790 ,w__2765 ,w__2531);
  or g__5122(w__2788 ,w__2756 ,w__2454);
  or g__5123(w__2787 ,w__2749 ,w__2430);
  or g__5124(w__2786 ,w__2767 ,w__2415);
  or g__5125(w__2785 ,w__2753 ,w__2502);
  not g__5126(w__2769 ,in1[7]);
  not g__5127(w__2768 ,in1[9]);
  not g__5128(w__2767 ,in1[1]);
  not g__5129(w__2766 ,in1[15]);
  not g__5130(w__2765 ,in1[6]);
  not g__5131(w__2764 ,in1[12]);
  not g__5132(w__2763 ,in1[4]);
  not g__5133(w__2762 ,in1[0]);
  not g__5134(w__2761 ,in2[3]);
  not g__5135(w__2760 ,in2[7]);
  not g__5136(w__2759 ,in2[5]);
  not g__5137(w__2758 ,in2[9]);
  not g__5138(w__2757 ,in2[11]);
  not g__5139(w__2756 ,in1[5]);
  not g__5140(w__2755 ,in1[11]);
  not g__5141(w__2754 ,in1[3]);
  not g__5142(w__2753 ,in1[14]);
  not g__5143(w__2752 ,in1[13]);
  not g__5144(w__2751 ,in1[10]);
  not g__5145(w__2750 ,in1[8]);
  not g__5146(w__2749 ,in1[2]);
  not g__5147(w__2748 ,in2[0]);
  not g__5148(w__2747 ,in2[15]);
  not g__5149(w__2746 ,in2[1]);
  not g__5150(w__2745 ,in2[13]);
  not g__5151(w__2399 ,w__2713);
  not g__5152(w__2713 ,w__2762);
  not g__5153(w__2712 ,w__2710);
  not g__5154(w__2711 ,w__2710);
  not g__5155(w__2710 ,w__2732);
  not g__5156(w__2709 ,w__2707);
  not g__5157(w__2708 ,w__2707);
  not g__5158(w__2707 ,w__2838);
  not g__5159(w__2706 ,w__2704);
  not g__5160(w__2705 ,w__2704);
  not g__5161(w__2704 ,w__2835);
  not g__5162(w__2703 ,w__2701);
  not g__5163(w__2702 ,w__2701);
  not g__5164(w__2701 ,w__2833);
  not g__5165(w__2700 ,w__2698);
  not g__5166(w__2699 ,w__2698);
  not g__5167(w__2698 ,w__2834);
  not g__5168(w__2697 ,w__2695);
  not g__5169(w__2696 ,w__2695);
  not g__5170(w__2695 ,w__2731);
  not g__5171(w__2694 ,w__2692);
  not g__5172(w__2693 ,w__2692);
  not g__5173(w__2692 ,w__2730);
  not g__5174(w__2691 ,w__2689);
  not g__5175(w__2690 ,w__2689);
  not g__5176(w__2689 ,w__2830);
  not g__5177(w__2688 ,w__2686);
  not g__5178(w__2687 ,w__2686);
  not g__5179(w__2686 ,w__2831);
  not g__5180(w__2685 ,w__2683);
  not g__5181(w__2684 ,w__2683);
  not g__5182(w__2683 ,w__2729);
  not g__5183(w__2682 ,w__2680);
  not g__5184(w__2681 ,w__2680);
  not g__5185(w__2680 ,w__2728);
  not g__5186(w__2679 ,w__2677);
  not g__5187(w__2678 ,w__2677);
  not g__5188(w__2677 ,w__2828);
  not g__5189(w__2676 ,w__2674);
  not g__5190(w__2675 ,w__2674);
  not g__5191(w__2674 ,w__2827);
  not g__5192(w__2673 ,w__2671);
  not g__5193(w__2672 ,w__2671);
  not g__5194(w__2671 ,w__2727);
  not g__5195(w__2670 ,w__2668);
  not g__5196(w__2669 ,w__2668);
  not g__5197(w__2668 ,w__2726);
  not g__5198(w__2667 ,w__2665);
  not g__5199(w__2666 ,w__2665);
  not g__5200(w__2665 ,w__2928);
  not g__5201(w__2664 ,w__2662);
  not g__5202(w__2663 ,w__2662);
  not g__5203(w__2662 ,w__2927);
  not g__5204(w__2661 ,w__2659);
  not g__5205(w__2660 ,w__2659);
  not g__5206(w__2659 ,w__2738);
  not g__5207(w__2658 ,w__2656);
  not g__5208(w__2657 ,w__2656);
  not g__5209(w__2656 ,w__2737);
  not g__5210(w__2655 ,w__2653);
  not g__5211(w__2654 ,w__2653);
  not g__5212(w__2653 ,w__2925);
  not g__5213(w__2652 ,w__2650);
  not g__5214(w__2651 ,w__2650);
  not g__5215(w__2650 ,w__2924);
  not g__5216(w__2649 ,w__2647);
  not g__5217(w__2648 ,w__2647);
  not g__5218(w__2647 ,w__2736);
  not g__5219(w__2646 ,w__2644);
  not g__5220(w__2645 ,w__2644);
  not g__5221(w__2644 ,w__2735);
  not g__5222(w__2643 ,w__2641);
  not g__5223(w__2642 ,w__2641);
  not g__5224(w__2641 ,w__2841);
  not g__5225(w__2640 ,w__2638);
  not g__5226(w__2639 ,w__2638);
  not g__5227(w__2638 ,w__2840);
  not g__5228(w__2637 ,w__2635);
  not g__5229(w__2636 ,w__2635);
  not g__5230(w__2635 ,w__2734);
  not g__5231(w__2634 ,w__2632);
  not g__5232(w__2633 ,w__2632);
  not g__5233(w__2632 ,w__2733);
  not g__5234(w__2631 ,w__2721);
  not g__5235(w__2721 ,w__2814);
  not g__5236(w__2630 ,w__2718);
  not g__5237(w__2718 ,w__2794);
  not g__5238(w__2629 ,w__2725);
  not g__5239(w__2725 ,w__2818);
  not g__5240(w__2628 ,w__2722);
  not g__5241(w__2722 ,w__2815);
  not g__5242(w__2627 ,w__2723);
  not g__5243(w__2723 ,w__2816);
  not g__5244(w__2626 ,w__2719);
  not g__5245(w__2719 ,w__2812);
  not g__5246(w__2625 ,w__2717);
  not g__5247(w__2717 ,w__2791);
  not g__5248(w__2624 ,w__2715);
  not g__5249(w__2715 ,w__2787);
  not g__5250(w__2623 ,w__2716);
  not g__5251(w__2716 ,w__2788);
  not g__5252(w__2622 ,w__2714);
  not g__5253(w__2714 ,w__2786);
  not g__5254(w__2621 ,w__2720);
  not g__5255(w__2720 ,w__2813);
  not g__5256(w__2620 ,w__2724);
  not g__5257(w__2724 ,w__2817);
  not g__5258(w__2619 ,w__2618);
  not g__5259(w__2618 ,w__3373);
  not g__5260(w__2617 ,w__2739);
  not g__5261(w__2739 ,w__3376);
  not g__5262(w__2616 ,w__2615);
  not g__5263(w__2615 ,w__2746);
  not g__5264(w__2614 ,w__2613);
  not g__5265(w__2613 ,w__2759);
  not g__5266(w__2612 ,w__2611);
  not g__5267(w__2611 ,w__2758);
  not g__5268(w__2610 ,w__2609);
  not g__5269(w__2609 ,w__2761);
  not g__5270(w__2608 ,w__2607);
  not g__5271(w__2607 ,w__2760);
  not g__5272(w__2606 ,w__2605);
  not g__5273(w__2605 ,w__2757);
  not g__5274(w__2604 ,w__2603);
  not g__5275(w__2603 ,w__2745);
  not g__5276(w__2602 ,w__2601);
  not g__5277(w__2601 ,w__2836);
  buf g__5278(w__13561 ,w__2985);
  buf g__5279(w__13562 ,w__2911);
  not g__5280(w__2600 ,w__2599);
  not g__5281(w__2599 ,w__2784);
  not g__5282(w__2598 ,w__2597);
  not g__5283(w__2597 ,w__3374);
  not g__5284(w__2596 ,w__2741);
  not g__5285(w__2741 ,w__3730);
  not g__5286(w__2595 ,w__2742);
  not g__5287(w__2742 ,w__3746);
  not g__5288(w__2594 ,w__2743);
  not g__5289(w__2743 ,w__3986);
  not g__5290(w__2593 ,w__2740);
  not g__5291(w__2740 ,w__3729);
  not g__5292(w__2592 ,w__2744);
  not g__5293(w__2744 ,w__3987);
  not g__5294(w__2591 ,w__2590);
  not g__5295(w__2590 ,w__3139);
  not g__5296(w__2589 ,w__2588);
  not g__5297(w__2588 ,w__3046);
  not g__5298(w__2587 ,w__2586);
  not g__5299(w__2586 ,w__3045);
  not g__5300(w__2585 ,w__2584);
  not g__5301(w__2584 ,w__3042);
  not g__5302(w__2583 ,w__2582);
  not g__5303(w__2582 ,w__3041);
  not g__5304(w__2581 ,w__2580);
  not g__5305(w__2580 ,w__3044);
  not g__5306(w__2579 ,w__2578);
  not g__5307(w__2578 ,w__3043);
  not g__5308(w__2577 ,w__2576);
  not g__5309(w__2576 ,w__2747);
  not g__5310(w__2575 ,w__2574);
  not g__5311(w__2574 ,w__3140);
  not g__5312(w__2573 ,w__2571);
  not g__5313(w__2572 ,w__2571);
  not g__5314(w__2571 ,w__2748);
  not g__5315(w__2570 ,w__2568);
  not g__5316(w__2569 ,w__2568);
  not g__5317(w__2568 ,w__2837);
  not g__5318(w__2567 ,w__2737);
  not g__5319(w__2737 ,w__2926);
  not g__5320(w__2566 ,w__2729);
  not g__5321(w__2729 ,w__2829);
  not g__5322(w__2565 ,w__2728);
  not g__5323(w__2728 ,w__2829);
  not g__5324(w__2564 ,w__2727);
  not g__5325(w__2727 ,w__2826);
  not g__5326(w__2563 ,w__2735);
  not g__5327(w__2735 ,w__2923);
  not g__5328(w__2562 ,w__2738);
  not g__5329(w__2738 ,w__2926);
  not g__5330(w__2561 ,w__2736);
  not g__5331(w__2736 ,w__2923);
  not g__5332(w__2560 ,w__2734);
  not g__5333(w__2734 ,w__2839);
  not g__5334(w__2559 ,w__2733);
  not g__5335(w__2733 ,w__2839);
  not g__5336(w__2558 ,w__2726);
  not g__5337(w__2726 ,w__2826);
  not g__5338(w__2557 ,w__2730);
  not g__5339(w__2730 ,w__2832);
  not g__5340(w__2556 ,w__2732);
  not g__5341(w__2732 ,w__2837);
  not g__5342(w__2555 ,w__2731);
  not g__5343(w__2731 ,w__2832);
  not g__5344(w__2554 ,w__2553);
  not g__5345(w__2553 ,w__3293);
  not g__5346(w__2552 ,w__2551);
  not g__5347(w__2551 ,w__3370);
  not g__5348(w__2550 ,w__2549);
  not g__5349(w__2549 ,w__3295);
  not g__5350(w__2548 ,w__2547);
  not g__5351(w__2547 ,w__3291);
  not g__5352(w__2398 ,w__2407);
  not g__5353(w__2546 ,w__2407);
  not g__5354(w__2407 ,w__2399);
  not g__5355(w__2545 ,w__2713);
  not g__5356(w__2544 ,w__2542);
  not g__5357(w__2543 ,w__2542);
  not g__5358(w__2542 ,w__3139);
  not g__5359(w__2541 ,w__2539);
  not g__5360(w__2540 ,w__2539);
  not g__5361(w__2539 ,w__3140);
  not g__5362(w__2538 ,w__2536);
  not g__5363(w__2537 ,w__2536);
  not g__5364(w__2536 ,w__3046);
  not g__5365(w__2535 ,w__2533);
  not g__5366(w__2534 ,w__2533);
  not g__5367(w__2533 ,w__3043);
  not g__5368(w__2532 ,w__2530);
  not g__5369(w__2531 ,w__2530);
  not g__5370(w__2530 ,w__2747);
  not g__5371(w__2529 ,w__2527);
  not g__5372(w__2528 ,w__2527);
  not g__5373(w__2527 ,w__3045);
  not g__5374(w__2526 ,w__2524);
  not g__5375(w__2525 ,w__2524);
  not g__5376(w__2524 ,w__3044);
  not g__5377(w__2523 ,w__2521);
  not g__5378(w__2522 ,w__2521);
  not g__5379(w__2521 ,w__3042);
  not g__5380(w__2520 ,w__2518);
  not g__5381(w__2519 ,w__2518);
  not g__5382(w__2518 ,w__3041);
  not g__5383(w__2517 ,w__2515);
  not g__5384(w__2516 ,w__2515);
  not g__5385(w__2515 ,w__3139);
  not g__5386(w__2514 ,w__2512);
  not g__5387(w__2513 ,w__2512);
  not g__5388(w__2512 ,w__2591);
  not g__5389(w__2511 ,w__2509);
  not g__5390(w__2510 ,w__2509);
  not g__5391(w__2509 ,w__2581);
  not g__5392(w__2508 ,w__2506);
  not g__5393(w__2507 ,w__2506);
  not g__5394(w__2506 ,w__2583);
  not g__5395(w__2505 ,w__2503);
  not g__5396(w__2504 ,w__2503);
  not g__5397(w__2503 ,w__2579);
  not g__5398(w__2502 ,w__2500);
  not g__5399(w__2501 ,w__2500);
  not g__5400(w__2500 ,w__2577);
  not g__5401(w__2499 ,w__2497);
  not g__5402(w__2498 ,w__2497);
  not g__5403(w__2497 ,w__2573);
  not g__5404(w__2496 ,w__2494);
  not g__5405(w__2495 ,w__2494);
  not g__5406(w__2494 ,w__3044);
  not g__5407(w__2493 ,w__2491);
  not g__5408(w__2492 ,w__2491);
  not g__5409(w__2491 ,w__2591);
  not g__5410(w__2490 ,w__2488);
  not g__5411(w__2489 ,w__2488);
  not g__5412(w__2488 ,w__2748);
  not g__5413(w__2487 ,w__2485);
  not g__5414(w__2486 ,w__2485);
  not g__5415(w__2485 ,w__2748);
  not g__5416(w__2484 ,w__2482);
  not g__5417(w__2483 ,w__2482);
  not g__5418(w__2482 ,w__2589);
  not g__5419(w__2481 ,w__2479);
  not g__5420(w__2480 ,w__2479);
  not g__5421(w__2479 ,w__2587);
  not g__5422(w__2478 ,w__2476);
  not g__5423(w__2477 ,w__2476);
  not g__5424(w__2476 ,w__2585);
  not g__5425(w__2475 ,w__2473);
  not g__5426(w__2474 ,w__2473);
  not g__5427(w__2473 ,w__3140);
  not g__5428(w__2472 ,w__2470);
  not g__5429(w__2471 ,w__2470);
  not g__5430(w__2470 ,w__2575);
  not g__5431(w__2469 ,w__2467);
  not g__5432(w__2468 ,w__2467);
  not g__5433(w__2467 ,w__2575);
  not g__5434(w__2466 ,w__2464);
  not g__5435(w__2465 ,w__2464);
  not g__5436(w__2464 ,w__3043);
  not g__5437(w__2463 ,w__2461);
  not g__5438(w__2462 ,w__2461);
  not g__5439(w__2461 ,w__2583);
  not g__5440(w__2460 ,w__2458);
  not g__5441(w__2459 ,w__2458);
  not g__5442(w__2458 ,w__3042);
  not g__5443(w__2457 ,w__2455);
  not g__5444(w__2456 ,w__2455);
  not g__5445(w__2455 ,w__2579);
  not g__5446(w__2454 ,w__2452);
  not g__5447(w__2453 ,w__2452);
  not g__5448(w__2452 ,w__2577);
  not g__5449(w__2451 ,w__2449);
  not g__5450(w__2450 ,w__2449);
  not g__5451(w__2449 ,w__3041);
  not g__5452(w__2448 ,w__2446);
  not g__5453(w__2447 ,w__2446);
  not g__5454(w__2446 ,w__3045);
  not g__5455(w__2445 ,w__2443);
  not g__5456(w__2444 ,w__2443);
  not g__5457(w__2443 ,w__2581);
  not g__5458(w__2442 ,w__2440);
  not g__5459(w__2441 ,w__2440);
  not g__5460(w__2440 ,w__2585);
  not g__5461(w__2439 ,w__2437);
  not g__5462(w__2438 ,w__2437);
  not g__5463(w__2437 ,w__2589);
  not g__5464(w__2436 ,w__2434);
  not g__5465(w__2435 ,w__2434);
  not g__5466(w__2434 ,w__3046);
  not g__5467(w__2433 ,w__2431);
  not g__5468(w__2432 ,w__2431);
  not g__5469(w__2431 ,w__2587);
  not g__5470(w__2430 ,w__2428);
  not g__5471(w__2429 ,w__2428);
  not g__5472(w__2428 ,w__2747);
  not g__5473(w__2427 ,w__2426);
  not g__5474(w__2426 ,w__2572);
  not g__5475(w__2425 ,w__2424);
  not g__5476(w__2424 ,w__2543);
  not g__5477(w__2423 ,w__2422);
  not g__5478(w__2422 ,w__2520);
  not g__5479(w__2421 ,w__2420);
  not g__5480(w__2420 ,w__2523);
  not g__5481(w__2419 ,w__2418);
  not g__5482(w__2418 ,w__2526);
  not g__5483(w__2417 ,w__2416);
  not g__5484(w__2416 ,w__2529);
  not g__5485(w__2415 ,w__2414);
  not g__5486(w__2414 ,w__2532);
  not g__5487(w__2413 ,w__2412);
  not g__5488(w__2412 ,w__2535);
  not g__5489(w__2411 ,w__2410);
  not g__5490(w__2410 ,w__2538);
  not g__5491(w__2409 ,w__2408);
  not g__5492(w__2408 ,w__2541);
  xor g__5493(w__2406 ,w__3988 ,w__4083);
  xor g__5494(w__13538 ,w__3964 ,w__4053);
  xor g__5495(w__2405 ,w__3946 ,w__3967);
  xor g__5496(w__2404 ,w__3605 ,w__3683);
  xor g__5497(w__2403 ,w__3599 ,w__2553);
  xor g__5498(w__2402 ,w__3709 ,w__2551);
  xor g__5499(w__2401 ,w__3588 ,w__2549);
  xor g__5500(w__2400 ,w__3696 ,w__2547);
  xnor g__5501(w__13734 ,w__5780 ,w__5815);
  xnor g__5502(w__13735 ,w__5783 ,w__4115);
  xnor g__5503(w__13737 ,w__5793 ,w__5807);
  xnor g__5504(w__13736 ,w__5789 ,w__5806);
  xnor g__5505(w__13733 ,w__5773 ,w__5808);
  or g__5506(w__13673 ,w__5778 ,w__5814);
  or g__5507(w__13672 ,w__5801 ,w__5813);
  or g__5508(w__13669 ,w__5796 ,w__5810);
  or g__5509(w__13668 ,w__5805 ,w__5812);
  or g__5510(w__13670 ,w__5794 ,w__5811);
  or g__5511(w__13671 ,w__5803 ,w__5809);
  xnor g__5512(w__13732 ,w__5759 ,w__5787);
  xnor g__5513(w__13738 ,w__5790 ,w__5786);
  xnor g__5514(w__13731 ,w__5761 ,w__5785);
  xnor g__5515(w__5815 ,w__5675 ,w__5791);
  and g__5516(w__5814 ,w__5767 ,w__5790);
  and g__5517(w__5813 ,w__5800 ,w__5793);
  or g__5518(w__13666 ,w__5775 ,w__5795);
  and g__5519(w__5812 ,w__5773 ,w__5797);
  nor g__5520(w__5811 ,w__5804 ,w__5792);
  or g__5521(w__13674 ,w__5757 ,w__5798);
  or g__5522(w__13667 ,w__5777 ,w__5799);
  and g__5523(w__5810 ,w__5788 ,w__5791);
  xnor g__5524(w__13739 ,w__5772 ,w__5764);
  xnor g__5525(w__13730 ,w__5760 ,w__5763);
  xnor g__5526(w__13740 ,w__5678 ,w__5765);
  nor g__5527(w__5809 ,w__5802 ,w__5789);
  xnor g__5528(w__5808 ,w__5769 ,w__5695);
  xnor g__5529(w__5807 ,w__5782 ,w__5696);
  xnor g__5530(w__5806 ,w__5770 ,w__5784);
  nor g__5531(w__5805 ,w__4303 ,w__5769);
  and g__5532(w__5804 ,w__5697 ,w__5783);
  nor g__5533(w__5803 ,w__5771 ,w__5784);
  and g__5534(w__5802 ,w__5771 ,w__5784);
  nor g__5535(w__5801 ,w__4301 ,w__5782);
  or g__5536(w__5800 ,w__4453 ,w__5781);
  nor g__5537(w__5799 ,w__5759 ,w__5776);
  and g__5538(w__5798 ,w__5756 ,w__5772);
  or g__5539(w__5797 ,w__4452 ,w__5768);
  nor g__5540(w__5796 ,w__5675 ,w__5780);
  nor g__5541(w__5795 ,w__5761 ,w__5774);
  nor g__5542(w__5794 ,w__5697 ,w__5783);
  or g__5543(w__5788 ,w__5674 ,w__5779);
  or g__5544(w__13729 ,w__5750 ,w__5766);
  xnor g__5545(w__13741 ,w__5704 ,w__4114);
  xnor g__5546(w__13743 ,w__5614 ,w__5734);
  xnor g__5547(w__13664 ,w__5682 ,w__5735);
  xnor g__5548(w__5787 ,w__5646 ,w__5741);
  xnor g__5549(w__5786 ,w__5744 ,w__5699);
  xnor g__5550(w__5785 ,w__5636 ,w__5745);
  xnor g__5551(w__5793 ,w__5681 ,w__5737);
  xnor g__5552(w__5792 ,w__5730 ,w__5733);
  xnor g__5553(w__5791 ,w__5707 ,w__5736);
  xnor g__5554(w__5790 ,w__5679 ,w__5731);
  xnor g__5555(w__5789 ,w__5703 ,w__5732);
  not g__5556(w__5781 ,w__5782);
  not g__5557(w__5779 ,w__5780);
  nor g__5558(w__5778 ,w__5699 ,w__5744);
  nor g__5559(w__5777 ,w__5646 ,w__5742);
  and g__5560(w__5776 ,w__5646 ,w__5742);
  or g__5561(w__13675 ,w__5721 ,w__5755);
  nor g__5562(w__5775 ,w__5636 ,w__5746);
  or g__5563(w__13676 ,w__5719 ,w__5754);
  or g__5564(w__13678 ,w__5715 ,w__5753);
  or g__5565(w__13728 ,w__5713 ,w__5751);
  and g__5566(w__5774 ,w__5636 ,w__5746);
  and g__5567(w__5784 ,w__5727 ,w__5747);
  and g__5568(w__5783 ,w__5710 ,w__5748);
  and g__5569(w__5782 ,w__5725 ,w__5758);
  and g__5570(w__5780 ,w__5716 ,w__5752);
  not g__5571(w__5771 ,w__5770);
  not g__5572(w__5768 ,w__5769);
  or g__5573(w__5767 ,w__5698 ,w__5743);
  nor g__5574(w__5766 ,w__5760 ,w__5749);
  or g__5575(w__13727 ,w__5709 ,w__5738);
  xnor g__5576(w__13742 ,w__5706 ,w__5687);
  or g__5577(w__13677 ,w__5667 ,w__5740);
  xnor g__5578(w__5765 ,w__5650 ,w__5702);
  xnor g__5579(w__5764 ,w__5694 ,w__5692);
  xnor g__5580(w__5763 ,w__5631 ,w__5700);
  xnor g__5581(w__5762 ,w__5705 ,w__5590);
  or g__5582(w__5773 ,w__5722 ,w__5739);
  xnor g__5583(w__5772 ,w__5633 ,w__5685);
  xnor g__5584(w__5770 ,w__5513 ,w__5684);
  xnor g__5585(w__5769 ,w__5680 ,w__5686);
  or g__5586(w__5758 ,w__5679 ,w__5723);
  nor g__5587(w__5757 ,w__5692 ,w__5694);
  or g__5588(w__5756 ,w__5691 ,w__5693);
  and g__5589(w__5755 ,w__5720 ,w__5702);
  nor g__5590(w__5754 ,w__5729 ,w__5704);
  and g__5591(w__5753 ,w__5614 ,w__5714);
  or g__5592(w__13679 ,w__5616 ,w__5712);
  or g__5593(w__5752 ,w__5730 ,w__5711);
  nor g__5594(w__5751 ,w__5688 ,w__5705);
  nor g__5595(w__5750 ,w__5631 ,w__5701);
  and g__5596(w__5749 ,w__5631 ,w__5701);
  or g__5597(w__5748 ,w__5703 ,w__5728);
  or g__5598(w__5747 ,w__5681 ,w__5726);
  and g__5599(w__5761 ,w__5608 ,w__5717);
  and g__5600(w__5760 ,w__5543 ,w__5690);
  and g__5601(w__5759 ,w__5671 ,w__5724);
  not g__5602(w__5746 ,w__5745);
  not g__5603(w__5743 ,w__5744);
  not g__5604(w__5742 ,w__5741);
  nor g__5605(w__5740 ,w__5668 ,w__5706);
  nor g__5606(w__5739 ,w__5718 ,w__5707);
  nor g__5607(w__5738 ,w__5682 ,w__5708);
  xnor g__5608(w__13744 ,w__5662 ,w__5642);
  xnor g__5609(w__13663 ,w__5611 ,w__5640);
  xnor g__5610(w__5737 ,w__5516 ,w__5648);
  xnor g__5611(w__5736 ,w__5635 ,w__5659);
  xnor g__5612(w__5735 ,w__5416 ,w__5657);
  xnor g__5613(w__5734 ,w__5654 ,w__5455);
  xnor g__5614(w__5733 ,w__5656 ,w__5630);
  xnor g__5615(w__5732 ,w__5645 ,w__5386);
  xnor g__5616(w__5731 ,w__5585 ,w__5652);
  xnor g__5617(w__5745 ,w__5661 ,w__5600);
  and g__5618(w__5744 ,w__5643 ,w__5689);
  xnor g__5619(w__5741 ,w__5683 ,w__5641);
  and g__5620(w__5729 ,w__5655 ,w__5676);
  and g__5621(w__5728 ,w__5386 ,w__5645);
  or g__5622(w__5727 ,w__5515 ,w__5648);
  nor g__5623(w__5726 ,w__5516 ,w__5647);
  or g__5624(w__5725 ,w__5585 ,w__5651);
  or g__5625(w__5724 ,w__5669 ,w__5680);
  nor g__5626(w__5723 ,w__5584 ,w__5652);
  nor g__5627(w__5722 ,w__5635 ,w__5660);
  nor g__5628(w__5721 ,w__5678 ,w__5650);
  or g__5629(w__5720 ,w__5677 ,w__5649);
  nor g__5630(w__5719 ,w__5655 ,w__5676);
  and g__5631(w__5718 ,w__5635 ,w__5660);
  or g__5632(w__5717 ,w__5618 ,w__5683);
  or g__5633(w__5716 ,w__5630 ,w__5656);
  nor g__5634(w__5715 ,w__4304 ,w__5654);
  or g__5635(w__5714 ,w__4451 ,w__5653);
  nor g__5636(w__5713 ,w__5590 ,w__5673);
  and g__5637(w__5712 ,w__5617 ,w__5662);
  and g__5638(w__5711 ,w__5630 ,w__5656);
  or g__5639(w__13725 ,w__5622 ,w__5664);
  or g__5640(w__13726 ,w__5625 ,w__5663);
  or g__5641(w__5710 ,w__5386 ,w__5645);
  nor g__5642(w__5709 ,w__5416 ,w__5658);
  and g__5643(w__5708 ,w__5416 ,w__5658);
  and g__5644(w__5730 ,w__5533 ,w__5672);
  not g__5645(w__5701 ,w__5700);
  not g__5646(w__5699 ,w__5698);
  not g__5647(w__5693 ,w__5694);
  not g__5648(w__5691 ,w__5692);
  xnor g__5649(w__13661 ,w__5384 ,w__5606);
  xnor g__5650(w__13745 ,w__5612 ,w__5599);
  or g__5651(w__5690 ,w__5577 ,w__5661);
  or g__5652(w__5689 ,w__5613 ,w__5644);
  and g__5653(w__5688 ,w__5590 ,w__5673);
  or g__5654(w__13680 ,w__5536 ,w__5670);
  xnor g__5655(w__13746 ,w__5508 ,w__5597);
  xnor g__5656(w__13662 ,w__5589 ,w__5603);
  xnor g__5657(w__5687 ,w__5547 ,w__5637);
  xnor g__5658(w__5686 ,w__5634 ,w__5546);
  xnor g__5659(w__5685 ,w__5421 ,w__5613);
  xnor g__5660(w__5684 ,w__5639 ,w__5449);
  xnor g__5661(w__5707 ,w__5414 ,w__5595);
  xnor g__5662(w__5706 ,w__5518 ,w__5596);
  xnor g__5663(w__5705 ,w__4112 ,w__5598);
  xnor g__5664(w__5704 ,w__5551 ,w__5605);
  and g__5665(w__5703 ,w__5542 ,w__5665);
  xnor g__5666(w__5702 ,w__5638 ,w__5604);
  xnor g__5667(w__5700 ,w__5552 ,w__5602);
  xnor g__5668(w__5698 ,w__5452 ,w__5601);
  xnor g__5669(w__5697 ,w__5378 ,w__5594);
  xnor g__5670(w__5696 ,w__5610 ,w__5591);
  xnor g__5671(w__5695 ,w__5453 ,w__5592);
  xnor g__5672(w__5694 ,w__5447 ,w__5593);
  and g__5673(w__5692 ,w__5571 ,w__5666);
  not g__5674(w__5677 ,w__5678);
  not g__5675(w__5674 ,w__5675);
  or g__5676(w__5672 ,w__5532 ,w__5639);
  or g__5677(w__5671 ,w__5546 ,w__5634);
  nor g__5678(w__5670 ,w__5535 ,w__5612);
  and g__5679(w__5669 ,w__5546 ,w__5634);
  and g__5680(w__5668 ,w__5548 ,w__5637);
  nor g__5681(w__5667 ,w__5548 ,w__5637);
  or g__5682(w__5666 ,w__5638 ,w__5568);
  or g__5683(w__5665 ,w__5540 ,w__5610);
  and g__5684(w__5664 ,w__5517 ,w__5624);
  and g__5685(w__5663 ,w__5611 ,w__5620);
  and g__5686(w__5683 ,w__5583 ,w__5627);
  and g__5687(w__5682 ,w__5556 ,w__5607);
  and g__5688(w__5681 ,w__5582 ,w__5628);
  and g__5689(w__5680 ,w__5538 ,w__5621);
  and g__5690(w__5679 ,w__5576 ,w__5626);
  and g__5691(w__5678 ,w__5567 ,w__5619);
  and g__5692(w__5676 ,w__5563 ,w__5629);
  and g__5693(w__5675 ,w__5561 ,w__5615);
  and g__5694(w__5673 ,w__5581 ,w__5623);
  not g__5695(w__5660 ,w__5659);
  not g__5696(w__5658 ,w__5657);
  not g__5697(w__5653 ,w__5654);
  not g__5698(w__5651 ,w__5652);
  not g__5699(w__5649 ,w__5650);
  not g__5700(w__5647 ,w__5648);
  xnor g__5701(w__13747 ,w__5464 ,w__4113);
  or g__5702(w__13681 ,w__5554 ,w__5609);
  nor g__5703(w__5644 ,w__5421 ,w__5632);
  or g__5704(w__5643 ,w__5420 ,w__5633);
  xnor g__5705(w__5642 ,w__5587 ,w__5438);
  xnor g__5706(w__5641 ,w__4110 ,w__5545);
  xnor g__5707(w__5640 ,w__5550 ,w__5439);
  xnor g__5708(w__5662 ,w__5471 ,w__5525);
  xnor g__5709(w__5661 ,w__5466 ,w__5522);
  xnor g__5710(w__5659 ,w__5423 ,w__4109);
  xnor g__5711(w__5657 ,w__5467 ,w__4111);
  xnor g__5712(w__5656 ,w__5460 ,w__5521);
  xnor g__5713(w__5655 ,w__5425 ,w__5519);
  xnor g__5714(w__5654 ,w__5465 ,w__5520);
  xnor g__5715(w__5652 ,w__5399 ,w__5527);
  xnor g__5716(w__5650 ,w__5472 ,w__5528);
  xnor g__5717(w__5648 ,w__5376 ,w__5524);
  xnor g__5718(w__5646 ,w__5457 ,w__5526);
  xnor g__5719(w__5645 ,w__5458 ,w__5523);
  not g__5720(w__5632 ,w__5633);
  or g__5721(w__5629 ,w__5518 ,w__5562);
  or g__5722(w__5628 ,w__5463 ,w__5580);
  or g__5723(w__5627 ,w__5462 ,w__5579);
  or g__5724(w__5626 ,w__5461 ,w__5574);
  nor g__5725(w__5625 ,w__4305 ,w__5550);
  or g__5726(w__5624 ,w__5410 ,w__5588);
  or g__5727(w__5623 ,w__5573 ,w__5553);
  nor g__5728(w__5622 ,w__5411 ,w__5589);
  or g__5729(w__13724 ,w__5473 ,w__5541);
  or g__5730(w__5621 ,w__5468 ,w__5537);
  or g__5731(w__5620 ,w__4450 ,w__5549);
  or g__5732(w__5619 ,w__5551 ,w__5565);
  or g__5733(w__13682 ,w__5481 ,w__5566);
  nor g__5734(w__5618 ,w__4110 ,w__5544);
  or g__5735(w__5617 ,w__4449 ,w__5586);
  nor g__5736(w__5616 ,w__4302 ,w__5587);
  or g__5737(w__5615 ,w__5459 ,w__5559);
  and g__5738(w__5639 ,w__5482 ,w__5569);
  and g__5739(w__5638 ,w__5500 ,w__5570);
  and g__5740(w__5637 ,w__5492 ,w__5560);
  and g__5741(w__5636 ,w__5496 ,w__5555);
  and g__5742(w__5635 ,w__5497 ,w__5564);
  and g__5743(w__5634 ,w__5505 ,w__5575);
  and g__5744(w__5633 ,w__5504 ,w__5572);
  and g__5745(w__5631 ,w__5489 ,w__5529);
  and g__5746(w__5630 ,w__5488 ,w__5557);
  or g__5747(w__13683 ,w__5329 ,w__5530);
  nor g__5748(w__5609 ,w__5470 ,w__5558);
  or g__5749(w__5608 ,w__5514 ,w__5545);
  xnor g__5750(w__13748 ,w__5469 ,w__5372);
  or g__5751(w__5607 ,w__4112 ,w__5578);
  xnor g__5752(w__5606 ,w__5456 ,w__5084);
  xnor g__5753(w__5605 ,w__5441 ,w__5442);
  xnor g__5754(w__5604 ,w__5444 ,w__5511);
  xnor g__5755(w__5603 ,w__5411 ,w__5517);
  xnor g__5756(w__5602 ,w__5445 ,w__5419);
  xnor g__5757(w__5601 ,w__5431 ,w__5463);
  xnor g__5758(w__5600 ,w__5391 ,w__5435);
  xnor g__5759(w__5599 ,w__5382 ,w__5437);
  xnor g__5760(w__5598 ,w__5433 ,w__5377);
  xnor g__5761(w__5597 ,w__5470 ,w__5394);
  xnor g__5762(w__5596 ,w__5440 ,w__5436);
  xnor g__5763(w__5595 ,w__5454 ,w__5468);
  xnor g__5764(w__5594 ,w__5450 ,w__5459);
  xnor g__5765(w__5593 ,w__5461 ,w__5407);
  xnor g__5766(w__5592 ,w__5462 ,w__5413);
  xnor g__5767(w__5591 ,w__5446 ,w__5432);
  or g__5768(w__5614 ,w__5487 ,w__5531);
  xnor g__5769(w__5613 ,w__5422 ,w__5429);
  xnor g__5770(w__5612 ,w__5397 ,w__5428);
  or g__5771(w__5611 ,w__5503 ,w__5534);
  and g__5772(w__5610 ,w__5475 ,w__5539);
  not g__5773(w__5588 ,w__5589);
  not g__5774(w__5586 ,w__5587);
  not g__5775(w__5584 ,w__5585);
  or g__5776(w__13723 ,w__5200 ,w__5478);
  or g__5777(w__5583 ,w__5413 ,w__5453);
  or g__5778(w__5582 ,w__5430 ,w__5452);
  or g__5779(w__5581 ,w__5419 ,w__5445);
  nor g__5780(w__5580 ,w__5431 ,w__5451);
  and g__5781(w__5579 ,w__5413 ,w__5453);
  and g__5782(w__5578 ,w__5377 ,w__5433);
  nor g__5783(w__5577 ,w__5391 ,w__5434);
  or g__5784(w__5576 ,w__5407 ,w__5447);
  or g__5785(w__5575 ,w__5423 ,w__5502);
  and g__5786(w__5574 ,w__5407 ,w__5447);
  and g__5787(w__5573 ,w__5419 ,w__5445);
  or g__5788(w__5572 ,w__5472 ,w__5501);
  or g__5789(w__5571 ,w__5444 ,w__5510);
  or g__5790(w__5570 ,w__5425 ,w__5499);
  or g__5791(w__5569 ,w__5395 ,w__5479);
  nor g__5792(w__5568 ,w__5443 ,w__5511);
  or g__5793(w__5567 ,w__5442 ,w__5441);
  nor g__5794(w__5566 ,w__5480 ,w__5464);
  and g__5795(w__5565 ,w__5442 ,w__5441);
  or g__5796(w__5564 ,w__5495 ,w__5460);
  or g__5797(w__5563 ,w__5436 ,w__5440);
  and g__5798(w__5562 ,w__5436 ,w__5440);
  or g__5799(w__5561 ,w__5378 ,w__5450);
  or g__5800(w__5560 ,w__5491 ,w__5465);
  and g__5801(w__5559 ,w__5378 ,w__5450);
  and g__5802(w__5558 ,w__5394 ,w__5509);
  or g__5803(w__5557 ,w__5484 ,w__5458);
  or g__5804(w__5556 ,w__5377 ,w__5433);
  or g__5805(w__5555 ,w__5483 ,w__5457);
  nor g__5806(w__5554 ,w__5394 ,w__5509);
  and g__5807(w__5590 ,w__5175 ,w__5498);
  and g__5808(w__5589 ,w__5216 ,w__5490);
  and g__5809(w__5587 ,w__5373 ,w__5485);
  and g__5810(w__5585 ,w__5400 ,w__5506);
  not g__5811(w__5553 ,w__5552);
  not g__5812(w__5549 ,w__5550);
  not g__5813(w__5548 ,w__5547);
  not g__5814(w__5544 ,w__5545);
  xnor g__5815(w__13660 ,w__5427 ,w__5321);
  or g__5816(w__5543 ,w__5390 ,w__5435);
  or g__5817(w__5542 ,w__5432 ,w__5446);
  nor g__5818(w__5541 ,w__5493 ,w__5456);
  and g__5819(w__5540 ,w__5432 ,w__5446);
  or g__5820(w__5539 ,w__5399 ,w__5486);
  or g__5821(w__5538 ,w__5414 ,w__5454);
  and g__5822(w__5537 ,w__5414 ,w__5454);
  nor g__5823(w__5536 ,w__5383 ,w__5437);
  and g__5824(w__5535 ,w__5383 ,w__5437);
  nor g__5825(w__5534 ,w__5494 ,w__5467);
  or g__5826(w__5533 ,w__5449 ,w__5512);
  nor g__5827(w__5532 ,w__5448 ,w__5513);
  nor g__5828(w__5531 ,w__5507 ,w__5471);
  nor g__5829(w__5530 ,w__5327 ,w__5469);
  or g__5830(w__5529 ,w__5477 ,w__5466);
  xnor g__5831(w__5528 ,w__5415 ,w__5417);
  xnor g__5832(w__5527 ,w__5207 ,w__5381);
  xnor g__5833(w__5526 ,w__5389 ,w__5406);
  xnor g__5834(w__5525 ,w__5204 ,w__5379);
  xnor g__5835(w__5524 ,w__5395 ,w__5393);
  xnor g__5836(w__5523 ,w__5387 ,w__5388);
  xnor g__5837(w__5522 ,w__5385 ,w__5004);
  xnor g__5838(w__5521 ,w__5408 ,w__5409);
  xnor g__5839(w__5520 ,w__5403 ,w__5404);
  xnor g__5840(w__5519 ,w__5412 ,w__5313);
  xnor g__5841(w__5552 ,w__5426 ,w__5319);
  and g__5842(w__5551 ,w__5349 ,w__5474);
  xnor g__5843(w__5550 ,w__5396 ,w__5306);
  xnor g__5844(w__5547 ,w__5424 ,w__5371);
  xnor g__5845(w__5546 ,w__5398 ,w__5307);
  and g__5846(w__5545 ,w__5154 ,w__5476);
  not g__5847(w__5515 ,w__5516);
  not g__5848(w__5514 ,w__4110);
  not g__5849(w__5512 ,w__5513);
  not g__5850(w__5510 ,w__5511);
  not g__5851(w__5509 ,w__5508);
  and g__5852(w__5507 ,w__5205 ,w__5379);
  or g__5853(w__5506 ,w__5401 ,w__5422);
  or g__5854(w__5505 ,w__5001 ,w__5405);
  or g__5855(w__5504 ,w__5417 ,w__5415);
  nor g__5856(w__5503 ,w__5080 ,w__5418);
  and g__5857(w__5502 ,w__5001 ,w__5405);
  and g__5858(w__5501 ,w__5417 ,w__5415);
  or g__5859(w__5500 ,w__5313 ,w__5412);
  and g__5860(w__5499 ,w__5313 ,w__5412);
  or g__5861(w__5498 ,w__5179 ,w__5426);
  or g__5862(w__5497 ,w__5409 ,w__5408);
  or g__5863(w__5496 ,w__5406 ,w__5389);
  and g__5864(w__5495 ,w__5409 ,w__5408);
  and g__5865(w__5494 ,w__5080 ,w__5418);
  nor g__5866(w__5493 ,w__5083 ,w__5384);
  or g__5867(w__5492 ,w__5404 ,w__5403);
  and g__5868(w__5491 ,w__5404 ,w__5403);
  or g__5869(w__5490 ,w__5171 ,w__5396);
  or g__5870(w__5489 ,w__5004 ,w__5385);
  or g__5871(w__5488 ,w__5388 ,w__5387);
  nor g__5872(w__5487 ,w__5205 ,w__5379);
  nor g__5873(w__5486 ,w__5207 ,w__5380);
  or g__5874(w__5485 ,w__5397 ,w__5374);
  and g__5875(w__5484 ,w__5388 ,w__5387);
  and g__5876(w__5483 ,w__5406 ,w__5389);
  or g__5877(w__5482 ,w__5376 ,w__5393);
  nor g__5878(w__5481 ,w__5314 ,w__5392);
  and g__5879(w__5480 ,w__5314 ,w__5392);
  or g__5880(w__13684 ,w__5167 ,w__5375);
  and g__5881(w__5479 ,w__5376 ,w__5393);
  nor g__5882(w__5478 ,w__5193 ,w__5427);
  and g__5883(w__5477 ,w__4259 ,w__5385);
  or g__5884(w__5476 ,w__5153 ,w__5398);
  or g__5885(w__5475 ,w__5206 ,w__5381);
  or g__5886(w__5474 ,w__5348 ,w__5424);
  and g__5887(w__5473 ,w__4307 ,w__5384);
  and g__5888(w__5518 ,w__5209 ,w__5402);
  xnor g__5889(w__5517 ,w__5299 ,w__5084);
  xnor g__5890(w__5516 ,w__5285 ,w__4326);
  xnor g__5891(w__5513 ,w__5318 ,w__5085);
  xnor g__5892(w__5511 ,w__5263 ,w__5277);
  xnor g__5893(w__5508 ,w__5208 ,w__5264);
  not g__5894(w__5451 ,w__5452);
  not g__5895(w__5448 ,w__5449);
  not g__5896(w__5443 ,w__5444);
  not g__5897(w__5434 ,w__5435);
  not g__5898(w__5430 ,w__5431);
  xnor g__5899(w__13750 ,w__5051 ,w__5304);
  xnor g__5900(w__13659 ,w__5274 ,w__4493);
  xnor g__5901(w__13749 ,w__5316 ,w__5294);
  xnor g__5902(w__5429 ,w__5312 ,w__5119);
  xnor g__5903(w__5428 ,w__5315 ,w__5036);
  xnor g__5904(w__5472 ,w__5117 ,w__5303);
  xnor g__5905(w__5471 ,w__5086 ,w__5305);
  xnor g__5906(w__5470 ,w__5130 ,w__5300);
  xnor g__5907(w__5469 ,w__5012 ,w__5301);
  xnor g__5908(w__5468 ,w__5276 ,w__4522);
  xnor g__5909(w__5467 ,w__5066 ,w__5296);
  xnor g__5910(w__5466 ,w__5289 ,w__4526);
  xnor g__5911(w__5465 ,w__5057 ,w__5269);
  xnor g__5912(w__5464 ,w__5133 ,w__5287);
  xnor g__5913(w__5463 ,w__5141 ,w__5282);
  xnor g__5914(w__5462 ,w__5064 ,w__5281);
  xnor g__5915(w__5461 ,w__5132 ,w__5279);
  xnor g__5916(w__5460 ,w__5131 ,w__5271);
  xnor g__5917(w__5459 ,w__5140 ,w__5310);
  xnor g__5918(w__5458 ,w__5134 ,w__5266);
  xnor g__5919(w__5457 ,w__5026 ,w__5265);
  xnor g__5920(w__5456 ,w__5275 ,w__4503);
  xnor g__5921(w__5455 ,w__5317 ,w__5268);
  xnor g__5922(w__5454 ,w__5063 ,w__5298);
  xnor g__5923(w__5453 ,w__5136 ,w__5283);
  xnor g__5924(w__5452 ,w__5038 ,w__5311);
  xnor g__5925(w__5450 ,w__5270 ,w__5082);
  xnor g__5926(w__5449 ,w__5104 ,w__5295);
  xnor g__5927(w__5447 ,w__5032 ,w__5280);
  xnor g__5928(w__5446 ,w__5151 ,w__5293);
  xnor g__5929(w__5445 ,w__5029 ,w__5284);
  xnor g__5930(w__5444 ,w__5099 ,w__5278);
  xnor g__5931(w__5442 ,w__5120 ,w__5273);
  xnor g__5932(w__5441 ,w__5138 ,w__5272);
  xnor g__5933(w__5440 ,w__5108 ,w__5292);
  xnor g__5934(w__5439 ,w__5267 ,w__4524);
  xnor g__5935(w__5438 ,w__5116 ,w__5291);
  xnor g__5936(w__5437 ,w__5054 ,w__5286);
  xnor g__5937(w__5436 ,w__5039 ,w__5302);
  xnor g__5938(w__5435 ,w__5100 ,w__5288);
  xnor g__5939(w__5433 ,w__5106 ,w__5290);
  xnor g__5940(w__5432 ,w__5019 ,w__5309);
  xnor g__5941(w__5431 ,w__5075 ,w__5320);
  not g__5942(w__5420 ,w__5421);
  not g__5943(w__5410 ,w__5411);
  or g__5944(w__5402 ,w__5217 ,w__5317);
  and g__5945(w__5401 ,w__5119 ,w__5312);
  or g__5946(w__5400 ,w__5119 ,w__5312);
  and g__5947(w__5427 ,w__5255 ,w__5339);
  and g__5948(w__5426 ,w__5260 ,w__5354);
  and g__5949(w__5425 ,w__5223 ,w__5351);
  and g__5950(w__5424 ,w__5214 ,w__5345);
  and g__5951(w__5423 ,w__5243 ,w__5358);
  and g__5952(w__5422 ,w__5251 ,w__5364);
  or g__5953(w__5421 ,w__5246 ,w__5359);
  and g__5954(w__5419 ,w__5253 ,w__5362);
  and g__5955(w__5418 ,w__5235 ,w__5347);
  and g__5956(w__5417 ,w__5240 ,w__5357);
  and g__5957(w__5416 ,w__5156 ,w__5369);
  and g__5958(w__5415 ,w__5236 ,w__5355);
  and g__5959(w__5414 ,w__5234 ,w__5353);
  and g__5960(w__5413 ,w__5258 ,w__5368);
  and g__5961(w__5412 ,w__5226 ,w__5352);
  and g__5962(w__5411 ,w__5254 ,w__5365);
  and g__5963(w__5409 ,w__5220 ,w__5350);
  and g__5964(w__5408 ,w__5215 ,w__5346);
  and g__5965(w__5407 ,w__5249 ,w__5363);
  and g__5966(w__5406 ,w__5213 ,w__5342);
  and g__5967(w__5405 ,w__5248 ,w__5361);
  and g__5968(w__5404 ,w__5199 ,w__5370);
  and g__5969(w__5403 ,w__5257 ,w__5341);
  not g__5970(w__5390 ,w__5391);
  not g__5971(w__5383 ,w__5382);
  not g__5972(w__5380 ,w__5381);
  and g__5973(w__5375 ,w__5174 ,w__5316);
  or g__5974(w__13685 ,w__5177 ,w__5325);
  and g__5975(w__5374 ,w__5036 ,w__5315);
  or g__5976(w__5373 ,w__5036 ,w__5315);
  xnor g__5977(w__5372 ,w__5010 ,w__5202);
  xnor g__5978(w__5371 ,w__5103 ,w__5262);
  and g__5979(w__5399 ,w__5230 ,w__5343);
  and g__5980(w__5398 ,w__5166 ,w__5323);
  and g__5981(w__5397 ,w__5195 ,w__5335);
  and g__5982(w__5396 ,w__5160 ,w__5324);
  and g__5983(w__5395 ,w__5173 ,w__5326);
  and g__5984(w__5394 ,w__5182 ,w__5333);
  and g__5985(w__5393 ,w__5222 ,w__5330);
  and g__5986(w__5392 ,w__5181 ,w__5332);
  or g__5987(w__5391 ,w__5159 ,w__5331);
  and g__5988(w__5389 ,w__5163 ,w__5336);
  and g__5989(w__5388 ,w__5194 ,w__5340);
  and g__5990(w__5387 ,w__5190 ,w__5337);
  and g__5991(w__5386 ,w__5172 ,w__5360);
  and g__5992(w__5385 ,w__5164 ,w__5366);
  or g__5993(w__5384 ,w__5158 ,w__5356);
  or g__5994(w__5382 ,w__5185 ,w__5344);
  and g__5995(w__5381 ,w__5169 ,w__5367);
  and g__5996(w__5379 ,w__5192 ,w__5338);
  and g__5997(w__5378 ,w__5201 ,w__5322);
  and g__5998(w__5377 ,w__5183 ,w__5328);
  and g__5999(w__5376 ,w__5152 ,w__5334);
  or g__6000(w__5370 ,w__5149 ,w__5198);
  or g__6001(w__5369 ,w__5150 ,w__5155);
  or g__6002(w__5368 ,w__5148 ,w__5256);
  or g__6003(w__5367 ,w__5147 ,w__5231);
  or g__6004(w__5366 ,w__5074 ,w__5165);
  or g__6005(w__5365 ,w__5252 ,w__5146);
  or g__6006(w__5364 ,w__5062 ,w__5250);
  or g__6007(w__5363 ,w__5145 ,w__5247);
  or g__6008(w__5362 ,w__5144 ,w__5244);
  or g__6009(w__5361 ,w__5142 ,w__5245);
  or g__6010(w__5360 ,w__4448 ,w__5242);
  and g__6011(w__5359 ,w__5263 ,w__5241);
  or g__6012(w__5358 ,w__5140 ,w__5238);
  or g__6013(w__5357 ,w__5139 ,w__5237);
  nor g__6014(w__5356 ,w__5161 ,w__4307);
  or g__6015(w__5355 ,w__5138 ,w__5232);
  or g__6016(w__5354 ,w__5076 ,w__5225);
  or g__6017(w__5353 ,w__4328 ,w__5229);
  or g__6018(w__5352 ,w__5137 ,w__5224);
  or g__6019(w__5351 ,w__5060 ,w__5221);
  or g__6020(w__5350 ,w__5065 ,w__5218);
  or g__6021(w__5349 ,w__5103 ,w__5261);
  nor g__6022(w__5348 ,w__5102 ,w__5262);
  or g__6023(w__5347 ,w__5135 ,w__5211);
  or g__6024(w__5346 ,w__5134 ,w__5210);
  or g__6025(w__5345 ,w__5057 ,w__5212);
  and g__6026(w__5344 ,w__5208 ,w__5239);
  or g__6027(w__5343 ,w__5132 ,w__5259);
  or g__6028(w__5342 ,w__5136 ,w__5227);
  or g__6029(w__5341 ,w__5053 ,w__5196);
  or g__6030(w__5340 ,w__5050 ,w__5191);
  or g__6031(w__5339 ,w__5188 ,w__5073);
  or g__6032(w__5338 ,w__5054 ,w__5189);
  or g__6033(w__5337 ,w__5151 ,w__5187);
  or g__6034(w__5336 ,w__5064 ,w__5184);
  or g__6035(w__5335 ,w__5069 ,w__5186);
  or g__6036(w__5334 ,w__5168 ,w__5075);
  or g__6037(w__5333 ,w__5133 ,w__5170);
  or g__6038(w__5332 ,w__5061 ,w__5180);
  and g__6039(w__5331 ,w__5162 ,w__4259);
  or g__6040(w__5330 ,w__5141 ,w__5178);
  nor g__6041(w__5329 ,w__5010 ,w__5203);
  or g__6042(w__5328 ,w__5143 ,w__5228);
  and g__6043(w__5327 ,w__5010 ,w__5203);
  or g__6044(w__5326 ,w__5072 ,w__5176);
  nor g__6045(w__5325 ,w__5051 ,w__5219);
  or g__6046(w__5324 ,w__5157 ,w__5066);
  or g__6047(w__5323 ,w__5063 ,w__5233);
  or g__6048(w__5322 ,w__4326 ,w__5197);
  xnor g__6049(w__13751 ,w__5077 ,w__4998);
  xnor g__6050(w__5321 ,w__5009 ,w__4309);
  xnor g__6051(w__5320 ,w__5043 ,w__4501);
  xnor g__6052(w__5319 ,w__5023 ,w__5002);
  xnor g__6053(w__5318 ,w__5088 ,w__4328);
  xnor g__6054(w__5311 ,w__5005 ,w__5072);
  xnor g__6055(w__5310 ,w__5122 ,w__4521);
  xnor g__6056(w__5309 ,w__5050 ,w__4495);
  xnor g__6057(w__5308 ,w__5150 ,w__4527);
  xnor g__6058(w__5307 ,w__4257 ,w__4497);
  xnor g__6059(w__5306 ,w__5092 ,w__5079);
  xnor g__6060(w__5305 ,w__5149 ,w__4756);
  xnor g__6061(w__5304 ,w__4761 ,w__5045);
  xnor g__6062(w__5303 ,w__5062 ,w__4759);
  xnor g__6063(w__5302 ,w__5137 ,w__4757);
  xnor g__6064(w__5301 ,w__5061 ,w__4760);
  xnor g__6065(w__5300 ,w__5069 ,w__4758);
  xnor g__6066(w__5299 ,w__5025 ,w__4523);
  xnor g__6067(w__5298 ,w__5087 ,w__5024);
  xnor g__6068(w__5297 ,w__5022 ,w__4499);
  xnor g__6069(w__5296 ,w__5020 ,w__4525);
  xnor g__6070(w__5295 ,w__5065 ,w__4496);
  xnor g__6071(w__5294 ,w__5047 ,w__5007);
  xnor g__6072(w__5293 ,w__5040 ,w__5015);
  xnor g__6073(w__5292 ,w__5107 ,w__5060);
  xnor g__6074(w__5291 ,w__5111 ,w__5053);
  xnor g__6075(w__5290 ,w__5135 ,w__5112);
  xnor g__6076(w__5289 ,w__5110 ,w__5076);
  xnor g__6077(w__5288 ,w__5144 ,w__5121);
  xnor g__6078(w__5287 ,w__5016 ,w__5018);
  xnor g__6079(w__5286 ,w__5008 ,w__5041);
  xnor g__6080(w__5285 ,w__5031 ,w__5027);
  xnor g__6081(w__5284 ,w__5143 ,w__4500);
  xnor g__6082(w__5283 ,w__5091 ,w__5095);
  xnor g__6083(w__5282 ,w__5011 ,w__5093);
  xnor g__6084(w__5281 ,w__5044 ,w__5028);
  xnor g__6085(w__5280 ,w__5030 ,w__5147);
  xnor g__6086(w__5279 ,w__5035 ,w__5105);
  xnor g__6087(w__5278 ,w__5114 ,w__5145);
  xnor g__6088(w__5277 ,w__5125 ,w__5127);
  xnor g__6089(w__5276 ,w__5148 ,w__5129);
  xnor g__6090(w__5275 ,w__5073 ,w__5123);
  xnor g__6091(w__5274 ,w__4505 ,w__5078);
  xnor g__6092(w__5273 ,w__5139 ,w__5118);
  xnor g__6093(w__5272 ,w__5037 ,w__5109);
  xnor g__6094(w__5271 ,w__5142 ,w__5094);
  xnor g__6095(w__5270 ,w__5113 ,w__5115);
  xnor g__6096(w__5269 ,w__5096 ,w__5098);
  xnor g__6097(w__5268 ,w__5089 ,w__5090);
  xnor g__6098(w__5267 ,w__5146 ,w__5128);
  xnor g__6099(w__5266 ,w__5097 ,w__5101);
  xnor g__6100(w__5265 ,w__5017 ,w__5074);
  xnor g__6101(w__5264 ,w__5034 ,w__5014);
  xnor g__6102(w__5317 ,w__5070 ,w__4992);
  xnor g__6103(w__5316 ,w__4986 ,w__5052);
  xnor g__6104(w__5315 ,w__4994 ,w__5048);
  xnor g__6105(w__5314 ,w__4996 ,w__5058);
  xnor g__6106(w__5313 ,w__4990 ,w__5055);
  xnor g__6107(w__5312 ,w__4988 ,w__5067);
  not g__6108(w__5261 ,w__5262);
  or g__6109(w__5260 ,w__4329 ,w__5110);
  and g__6110(w__5259 ,w__5105 ,w__5035);
  or g__6111(w__5258 ,w__4330 ,w__5129);
  or g__6112(w__5257 ,w__5111 ,w__5116);
  and g__6113(w__5256 ,w__4522 ,w__5129);
  or g__6114(w__5255 ,w__4339 ,w__5123);
  or g__6115(w__5254 ,w__4337 ,w__5128);
  or g__6116(w__5253 ,w__5121 ,w__5100);
  and g__6117(w__5252 ,w__4524 ,w__5128);
  or g__6118(w__5251 ,w__4759 ,w__5117);
  and g__6119(w__5250 ,w__4759 ,w__5117);
  or g__6120(w__5249 ,w__5114 ,w__5099);
  or g__6121(w__5248 ,w__5094 ,w__5131);
  and g__6122(w__5247 ,w__5114 ,w__5099);
  nor g__6123(w__5246 ,w__5127 ,w__5125);
  and g__6124(w__5245 ,w__5094 ,w__5131);
  and g__6125(w__5244 ,w__5121 ,w__5100);
  or g__6126(w__5243 ,w__4335 ,w__5122);
  and g__6127(w__5242 ,w__5027 ,w__5031);
  or g__6128(w__5241 ,w__5126 ,w__5124);
  or g__6129(w__5240 ,w__5120 ,w__5118);
  or g__6130(w__5239 ,w__5013 ,w__5033);
  and g__6131(w__5238 ,w__4521 ,w__5122);
  and g__6132(w__5237 ,w__5120 ,w__5118);
  or g__6133(w__5236 ,w__5109 ,w__5037);
  or g__6134(w__5235 ,w__5112 ,w__5106);
  or g__6135(w__5234 ,w__5115 ,w__5113);
  and g__6136(w__5233 ,w__5024 ,w__5087);
  and g__6137(w__5232 ,w__5109 ,w__5037);
  and g__6138(w__5231 ,w__5032 ,w__5030);
  or g__6139(w__5230 ,w__5105 ,w__5035);
  and g__6140(w__5229 ,w__5115 ,w__5113);
  and g__6141(w__5228 ,w__4334 ,w__5029);
  and g__6142(w__5227 ,w__5095 ,w__5091);
  or g__6143(w__5226 ,w__4757 ,w__5039);
  and g__6144(w__5225 ,w__4526 ,w__5110);
  and g__6145(w__5224 ,w__4757 ,w__5039);
  or g__6146(w__5223 ,w__5108 ,w__5107);
  or g__6147(w__5222 ,w__5093 ,w__5011);
  and g__6148(w__5221 ,w__5108 ,w__5107);
  or g__6149(w__5220 ,w__4333 ,w__5104);
  and g__6150(w__5219 ,w__4762 ,w__5045);
  and g__6151(w__5218 ,w__4496 ,w__5104);
  and g__6152(w__5217 ,w__5090 ,w__5089);
  or g__6153(w__5216 ,w__4261 ,w__5092);
  or g__6154(w__5215 ,w__5101 ,w__5097);
  or g__6155(w__5214 ,w__5098 ,w__5096);
  or g__6156(w__5213 ,w__5095 ,w__5091);
  and g__6157(w__5212 ,w__5098 ,w__5096);
  and g__6158(w__5211 ,w__5112 ,w__5106);
  and g__6159(w__5210 ,w__5101 ,w__5097);
  or g__6160(w__5209 ,w__5090 ,w__5089);
  and g__6161(w__5263 ,w__4991 ,w__5056);
  and g__6162(w__5262 ,w__4993 ,w__5071);
  not g__6163(w__5206 ,w__5207);
  not g__6164(w__5205 ,w__5204);
  not g__6165(w__5203 ,w__5202);
  or g__6166(w__5201 ,w__5081 ,w__5088);
  and g__6167(w__5200 ,w__4494 ,w__5009);
  or g__6168(w__5199 ,w__4756 ,w__5086);
  and g__6169(w__5198 ,w__4756 ,w__5086);
  and g__6170(w__5197 ,w__5081 ,w__5088);
  and g__6171(w__5196 ,w__5111 ,w__5116);
  or g__6172(w__5195 ,w__4758 ,w__5130);
  or g__6173(w__5194 ,w__4331 ,w__5019);
  nor g__6174(w__5193 ,w__4494 ,w__5009);
  or g__6175(w__5192 ,w__5041 ,w__5008);
  and g__6176(w__5191 ,w__4495 ,w__5019);
  or g__6177(w__5190 ,w__5015 ,w__5040);
  and g__6178(w__5189 ,w__5041 ,w__5008);
  and g__6179(w__5188 ,w__4503 ,w__5123);
  and g__6180(w__5187 ,w__5015 ,w__5040);
  and g__6181(w__5186 ,w__4758 ,w__5130);
  nor g__6182(w__5185 ,w__5014 ,w__5034);
  and g__6183(w__5184 ,w__5028 ,w__5044);
  or g__6184(w__5183 ,w__4500 ,w__5029);
  or g__6185(w__5182 ,w__5018 ,w__5016);
  or g__6186(w__5181 ,w__4760 ,w__5012);
  and g__6187(w__5180 ,w__4760 ,w__5012);
  and g__6188(w__5179 ,w__5023 ,w__5003);
  and g__6189(w__5178 ,w__5093 ,w__5011);
  nor g__6190(w__5177 ,w__4762 ,w__5045);
  and g__6191(w__5176 ,w__5038 ,w__5005);
  or g__6192(w__5175 ,w__5023 ,w__5003);
  or g__6193(w__5174 ,w__5006 ,w__5046);
  or g__6194(w__5173 ,w__5038 ,w__5005);
  or g__6195(w__5172 ,w__5027 ,w__5031);
  and g__6196(w__5171 ,w__4261 ,w__5092);
  and g__6197(w__5170 ,w__5018 ,w__5016);
  or g__6198(w__5169 ,w__5032 ,w__5030);
  nor g__6199(w__5168 ,w__4502 ,w__5043);
  nor g__6200(w__5167 ,w__5007 ,w__5047);
  or g__6201(w__5166 ,w__5024 ,w__5087);
  and g__6202(w__5165 ,w__5026 ,w__5017);
  or g__6203(w__5164 ,w__5026 ,w__5017);
  or g__6204(w__5163 ,w__5028 ,w__5044);
  or g__6205(w__5162 ,w__4498 ,w__5021);
  and g__6206(w__5161 ,w__4340 ,w__5025);
  or g__6207(w__5160 ,w__4336 ,w__5020);
  nor g__6208(w__5159 ,w__4499 ,w__5022);
  nor g__6209(w__5158 ,w__4340 ,w__5025);
  and g__6210(w__5157 ,w__4525 ,w__5020);
  or g__6211(w__5156 ,w__4338 ,w__4263);
  and g__6212(w__5155 ,w__4527 ,w__4263);
  or g__6213(w__5154 ,w__4332 ,w__4257);
  and g__6214(w__5153 ,w__4497 ,w__5000);
  or g__6215(w__5152 ,w__4501 ,w__5042);
  and g__6216(w__13686 ,w__4999 ,w__5077);
  and g__6217(w__5208 ,w__4997 ,w__5059);
  and g__6218(w__5207 ,w__4989 ,w__5068);
  and g__6219(w__5204 ,w__4995 ,w__5049);
  and g__6220(w__5202 ,w__4987 ,w__5052);
  not g__6221(w__5126 ,w__5127);
  not g__6222(w__5124 ,w__5125);
  not g__6223(w__5102 ,w__5103);
  not g__6224(w__5083 ,w__5084);
  not g__6225(w__5081 ,w__5082);
  not g__6226(w__5080 ,w__5079);
  or g__6227(w__5078 ,w__4769 ,w__4872);
  and g__6228(w__5151 ,w__4797 ,w__4901);
  and g__6229(w__5150 ,w__4820 ,w__4875);
  and g__6230(w__5149 ,w__4831 ,w__4914);
  and g__6231(w__5148 ,w__4708 ,w__4865);
  and g__6232(w__5147 ,w__4720 ,w__4878);
  and g__6233(w__5146 ,w__4819 ,w__4947);
  and g__6234(w__5145 ,w__4816 ,w__4948);
  and g__6235(w__5144 ,w__4815 ,w__4943);
  and g__6236(w__5143 ,w__4702 ,w__4853);
  and g__6237(w__5142 ,w__4813 ,w__4874);
  and g__6238(w__5141 ,w__4805 ,w__4929);
  and g__6239(w__5140 ,w__4807 ,w__4936);
  and g__6240(w__5139 ,w__4826 ,w__4934);
  and g__6241(w__5138 ,w__4802 ,w__4932);
  and g__6242(w__5137 ,w__4776 ,w__4927);
  and g__6243(w__5136 ,w__4811 ,w__4911);
  and g__6244(w__5135 ,w__4787 ,w__4984);
  and g__6245(w__5134 ,w__4791 ,w__4920);
  and g__6246(w__5133 ,w__4796 ,w__4893);
  and g__6247(w__5132 ,w__4746 ,w__4960);
  and g__6248(w__5131 ,w__4818 ,w__4946);
  and g__6249(w__5130 ,w__4739 ,w__4899);
  and g__6250(w__5129 ,w__4783 ,w__4958);
  or g__6251(w__5128 ,w__4765 ,w__4871);
  and g__6252(w__5127 ,w__4730 ,w__4941);
  and g__6253(w__5125 ,w__4732 ,w__4940);
  or g__6254(w__5123 ,w__4774 ,w__4868);
  and g__6255(w__5122 ,w__4809 ,w__4937);
  or g__6256(w__5121 ,w__4772 ,w__4870);
  and g__6257(w__5120 ,w__4824 ,w__4938);
  and g__6258(w__5119 ,w__4825 ,w__4955);
  and g__6259(w__5118 ,w__4808 ,w__4935);
  and g__6260(w__5117 ,w__4822 ,w__4954);
  and g__6261(w__5116 ,w__4788 ,w__4912);
  and g__6262(w__5115 ,w__4803 ,w__4879);
  and g__6263(w__5114 ,w__4717 ,w__4951);
  and g__6264(w__5113 ,w__4703 ,w__4861);
  or g__6265(w__5112 ,w__4767 ,w__4869);
  and g__6266(w__5111 ,w__4784 ,w__4913);
  and g__6267(w__5110 ,w__4712 ,w__4860);
  and g__6268(w__5109 ,w__4718 ,w__4933);
  and g__6269(w__5108 ,w__4795 ,w__4925);
  and g__6270(w__5107 ,w__4794 ,w__4924);
  and g__6271(w__5106 ,w__4710 ,w__4862);
  and g__6272(w__5105 ,w__4722 ,w__4897);
  and g__6273(w__5104 ,w__4733 ,w__4963);
  and g__6274(w__5103 ,w__4789 ,w__4971);
  and g__6275(w__5101 ,w__4736 ,w__4977);
  and g__6276(w__5100 ,w__4817 ,w__4949);
  and g__6277(w__5099 ,w__4792 ,w__4985);
  and g__6278(w__5098 ,w__4779 ,w__4959);
  and g__6279(w__5097 ,w__4786 ,w__4981);
  and g__6280(w__5096 ,w__4749 ,w__4850);
  or g__6281(w__5095 ,w__4763 ,w__4867);
  or g__6282(w__5094 ,w__4770 ,w__4866);
  and g__6283(w__5093 ,w__4748 ,w__4881);
  and g__6284(w__5092 ,w__4704 ,w__4864);
  and g__6285(w__5091 ,w__4777 ,w__4917);
  and g__6286(w__5090 ,w__4740 ,w__4910);
  and g__6287(w__5089 ,w__4778 ,w__4918);
  and g__6288(w__5088 ,w__4709 ,w__4857);
  and g__6289(w__5087 ,w__4735 ,w__4922);
  and g__6290(w__5086 ,w__4828 ,w__4916);
  and g__6291(w__5085 ,w__4823 ,w__4915);
  and g__6292(w__5084 ,w__4714 ,w__4863);
  and g__6293(w__5082 ,w__4800 ,w__4931);
  and g__6294(w__5079 ,w__4781 ,w__4919);
  not g__6295(w__5071 ,w__5070);
  not g__6296(w__5068 ,w__5067);
  not g__6297(w__5059 ,w__5058);
  not g__6298(w__5056 ,w__5055);
  not g__6299(w__5049 ,w__5048);
  not g__6300(w__5046 ,w__5047);
  not g__6301(w__5042 ,w__5043);
  not g__6302(w__5033 ,w__5034);
  not g__6303(w__5021 ,w__5022);
  not g__6304(w__5013 ,w__5014);
  not g__6305(w__5006 ,w__5007);
  not g__6306(w__5003 ,w__5002);
  not g__6307(w__5001 ,w__5000);
  or g__6308(w__13752 ,w__4843 ,w__4974);
  or g__6309(w__13753 ,w__4837 ,w__4950);
  or g__6310(w__13687 ,w__4829 ,w__4884);
  or g__6311(w__5077 ,w__4844 ,w__4966);
  and g__6312(w__5076 ,w__4798 ,w__4930);
  and g__6313(w__5075 ,w__4790 ,w__4894);
  and g__6314(w__5074 ,w__4847 ,w__4956);
  and g__6315(w__5073 ,w__4706 ,w__4859);
  and g__6316(w__5072 ,w__4727 ,w__4885);
  and g__6317(w__5070 ,w__4741 ,w__4976);
  and g__6318(w__5069 ,w__4834 ,w__4972);
  and g__6319(w__5067 ,w__4833 ,w__4965);
  and g__6320(w__5066 ,w__4716 ,w__4856);
  and g__6321(w__5065 ,w__4771 ,w__4969);
  and g__6322(w__5064 ,w__4705 ,w__4854);
  and g__6323(w__5063 ,w__4799 ,w__4962);
  and g__6324(w__5062 ,w__4845 ,w__4982);
  and g__6325(w__5061 ,w__4846 ,w__4970);
  and g__6326(w__5060 ,w__4841 ,w__4979);
  and g__6327(w__5058 ,w__4840 ,w__4978);
  and g__6328(w__5057 ,w__4842 ,w__4973);
  and g__6329(w__5055 ,w__4838 ,w__4980);
  and g__6330(w__5054 ,w__4836 ,w__4975);
  and g__6331(w__5053 ,w__4835 ,w__4983);
  or g__6332(w__5052 ,w__4810 ,w__4968);
  and g__6333(w__5051 ,w__4839 ,w__4967);
  and g__6334(w__5050 ,w__4707 ,w__4855);
  and g__6335(w__5048 ,w__4780 ,w__4907);
  and g__6336(w__5047 ,w__4785 ,w__4886);
  and g__6337(w__5045 ,w__4729 ,w__4888);
  and g__6338(w__5044 ,w__4793 ,w__4952);
  or g__6339(w__5043 ,w__4504 ,w__4964);
  and g__6340(w__5041 ,w__4801 ,w__4906);
  and g__6341(w__5040 ,w__4821 ,w__4942);
  and g__6342(w__5039 ,w__4747 ,w__4928);
  and g__6343(w__5038 ,w__4719 ,w__4939);
  and g__6344(w__5037 ,w__4742 ,w__4902);
  and g__6345(w__5036 ,w__4743 ,w__4900);
  and g__6346(w__5035 ,w__4827 ,w__4904);
  and g__6347(w__5034 ,w__4731 ,w__4903);
  and g__6348(w__5032 ,w__4728 ,w__4876);
  and g__6349(w__5031 ,w__4723 ,w__4957);
  and g__6350(w__5030 ,w__4713 ,w__4921);
  and g__6351(w__5029 ,w__4737 ,w__4880);
  and g__6352(w__5028 ,w__4726 ,w__4908);
  and g__6353(w__5027 ,w__4721 ,w__4877);
  and g__6354(w__5026 ,w__4806 ,w__4953);
  and g__6355(w__5025 ,w__4775 ,w__4961);
  and g__6356(w__5024 ,w__4764 ,w__4945);
  and g__6357(w__5023 ,w__4768 ,w__4926);
  and g__6358(w__5022 ,w__4773 ,w__4944);
  and g__6359(w__5020 ,w__4766 ,w__4883);
  and g__6360(w__5019 ,w__4745 ,w__4909);
  and g__6361(w__5018 ,w__4830 ,w__4896);
  and g__6362(w__5017 ,w__4715 ,w__4851);
  and g__6363(w__5016 ,w__4744 ,w__4895);
  and g__6364(w__5014 ,w__4738 ,w__4898);
  and g__6365(w__5012 ,w__4804 ,w__4891);
  and g__6366(w__5011 ,w__4782 ,w__4890);
  and g__6367(w__5010 ,w__4812 ,w__4889);
  or g__6368(w__5009 ,w__4769 ,w__4858);
  and g__6369(w__5008 ,w__4814 ,w__4905);
  and g__6370(w__5007 ,w__4832 ,w__4887);
  and g__6371(w__5005 ,w__4711 ,w__4852);
  and g__6372(w__5004 ,w__4724 ,w__4892);
  and g__6373(w__5002 ,w__4725 ,w__4923);
  and g__6374(w__5000 ,w__4734 ,w__4882);
  not g__6375(w__4999 ,w__4998);
  not g__6376(w__4997 ,w__4996);
  not g__6377(w__4995 ,w__4994);
  not g__6378(w__4993 ,w__4992);
  not g__6379(w__4991 ,w__4990);
  not g__6380(w__4989 ,w__4988);
  not g__6381(w__4987 ,w__4986);
  or g__6382(w__4985 ,w__4589 ,w__4175);
  or g__6383(w__4984 ,w__4603 ,w__4160);
  or g__6384(w__4983 ,w__4565 ,w__4134);
  or g__6385(w__4982 ,w__4553 ,w__4226);
  or g__6386(w__4981 ,w__4661 ,w__4157);
  or g__6387(w__4980 ,w__4558 ,w__4134);
  or g__6388(w__4979 ,w__4560 ,w__4201);
  or g__6389(w__4978 ,w__4554 ,w__4222);
  or g__6390(w__4977 ,w__4551 ,w__4217);
  or g__6391(w__4976 ,w__4586 ,w__4153);
  or g__6392(w__4975 ,w__4562 ,w__4223);
  nor g__6393(w__4974 ,w__4225 ,w__4555);
  or g__6394(w__4973 ,w__4556 ,w__4201);
  or g__6395(w__4972 ,w__4561 ,w__4202);
  or g__6396(w__4971 ,w__4557 ,w__4214);
  or g__6397(w__4970 ,w__4563 ,w__4225);
  or g__6398(w__4969 ,w__4612 ,w__4219);
  nor g__6399(w__4968 ,w__4223 ,w__4567);
  or g__6400(w__4967 ,w__4564 ,w__4253);
  nor g__6401(w__4966 ,w__4226 ,w__4566);
  or g__6402(w__4965 ,w__4559 ,w__4252);
  nor g__6403(w__4964 ,w__4222 ,w__4552);
  or g__6404(w__4963 ,w__4682 ,w__4166);
  or g__6405(w__4962 ,w__4638 ,w__4145);
  or g__6406(w__4961 ,w__4639 ,w__4193);
  or g__6407(w__4960 ,w__4684 ,w__4172);
  or g__6408(w__4959 ,w__4648 ,w__4169);
  or g__6409(w__4958 ,w__4613 ,w__4187);
  or g__6410(w__4957 ,w__4571 ,w__4216);
  or g__6411(w__4956 ,w__4576 ,w__4148);
  or g__6412(w__4955 ,w__4643 ,w__4192);
  or g__6413(w__4954 ,w__4665 ,w__4234);
  or g__6414(w__4953 ,w__4600 ,w__4228);
  or g__6415(w__4952 ,w__4654 ,w__4151);
  or g__6416(w__4951 ,w__4679 ,w__4190);
  nor g__6417(w__4950 ,w__4202 ,w__4529);
  or g__6418(w__4949 ,w__4660 ,w__4246);
  or g__6419(w__4948 ,w__4644 ,w__4186);
  or g__6420(w__4947 ,w__4608 ,w__4147);
  or g__6421(w__4946 ,w__4578 ,w__4231);
  or g__6422(w__4945 ,w__4670 ,w__4213);
  or g__6423(w__4944 ,w__4662 ,w__4142);
  or g__6424(w__4943 ,w__4655 ,w__4150);
  or g__6425(w__4942 ,w__4664 ,w__4169);
  or g__6426(w__4941 ,w__4685 ,w__4145);
  or g__6427(w__4940 ,w__4656 ,w__4171);
  or g__6428(w__4939 ,w__4588 ,w__4168);
  or g__6429(w__4938 ,w__4531 ,w__4144);
  or g__6430(w__4937 ,w__4652 ,w__4160);
  or g__6431(w__4936 ,w__4653 ,w__4189);
  or g__6432(w__4935 ,w__4657 ,w__4159);
  or g__6433(w__4934 ,w__4647 ,w__4243);
  or g__6434(w__4933 ,w__4683 ,w__4237);
  or g__6435(w__4932 ,w__4645 ,w__4168);
  or g__6436(w__4931 ,w__4642 ,w__4151);
  or g__6437(w__4930 ,w__4596 ,w__4159);
  or g__6438(w__4929 ,w__4594 ,w__4144);
  or g__6439(w__4928 ,w__4604 ,w__4141);
  or g__6440(w__4927 ,w__4606 ,w__4219);
  or g__6441(w__4926 ,w__4570 ,w__4186);
  or g__6442(w__4925 ,w__4649 ,w__4172);
  or g__6443(w__4924 ,w__4668 ,w__4231);
  or g__6444(w__4923 ,w__4646 ,w__4216);
  or g__6445(w__4922 ,w__4609 ,w__4157);
  or g__6446(w__4998 ,w__4489 ,w__4700);
  or g__6447(w__4996 ,w__4514 ,w__4697);
  or g__6448(w__4994 ,w__4482 ,w__4698);
  or g__6449(w__4992 ,w__4487 ,w__4696);
  or g__6450(w__4990 ,w__4485 ,w__4695);
  or g__6451(w__4988 ,w__4490 ,w__4701);
  or g__6452(w__4986 ,w__4479 ,w__4699);
  or g__6453(w__4921 ,w__4624 ,w__4177);
  or g__6454(w__4920 ,w__4585 ,w__4148);
  or g__6455(w__4919 ,w__4591 ,w__4192);
  or g__6456(w__4918 ,w__4601 ,w__4165);
  or g__6457(w__4917 ,w__4593 ,w__4156);
  or g__6458(w__4916 ,w__4671 ,w__4156);
  or g__6459(w__4915 ,w__4666 ,w__4142);
  or g__6460(w__4914 ,w__4614 ,w__4128);
  or g__6461(w__4913 ,w__4602 ,w__4150);
  or g__6462(w__4912 ,w__4674 ,w__4175);
  or g__6463(w__4911 ,w__4579 ,w__4228);
  or g__6464(w__4910 ,w__4532 ,w__4171);
  or g__6465(w__4909 ,w__4599 ,w__4235);
  or g__6466(w__4908 ,w__4650 ,w__4246);
  or g__6467(w__4907 ,w__4672 ,w__4154);
  or g__6468(w__4906 ,w__4619 ,w__4130);
  or g__6469(w__4905 ,w__4569 ,w__4189);
  or g__6470(w__4904 ,w__4677 ,w__4174);
  or g__6471(w__4903 ,w__4584 ,w__4128);
  or g__6472(w__4902 ,w__4568 ,w__4204);
  or g__6473(w__4901 ,w__4610 ,w__4174);
  or g__6474(w__4900 ,w__4592 ,w__4166);
  or g__6475(w__4899 ,w__4581 ,w__4237);
  or g__6476(w__4898 ,w__4598 ,w__4213);
  or g__6477(w__4897 ,w__4580 ,w__4130);
  or g__6478(w__4896 ,w__4528 ,w__4141);
  or g__6479(w__4895 ,w__4681 ,w__4205);
  or g__6480(w__4894 ,w__4582 ,w__4204);
  or g__6481(w__4893 ,w__4574 ,w__4243);
  or g__6482(w__4892 ,w__4641 ,w__4232);
  or g__6483(w__4891 ,w__4595 ,w__4154);
  or g__6484(w__4890 ,w__4651 ,w__4165);
  or g__6485(w__4889 ,w__4659 ,w__4122);
  or g__6486(w__4888 ,w__4590 ,w__4220);
  or g__6487(w__4887 ,w__4616 ,w__4122);
  or g__6488(w__4886 ,w__4680 ,w__4153);
  or g__6489(w__4885 ,w__4575 ,w__4126);
  nor g__6490(w__4884 ,w__4220 ,w__4621);
  or g__6491(w__4883 ,w__4605 ,w__4132);
  or g__6492(w__4882 ,w__4678 ,w__4132);
  or g__6493(w__4881 ,w__4607 ,w__4229);
  or g__6494(w__4880 ,w__4597 ,w__4147);
  or g__6495(w__4879 ,w__4573 ,w__4120);
  or g__6496(w__4878 ,w__4572 ,w__4234);
  or g__6497(w__4877 ,w__4687 ,w__4120);
  or g__6498(w__4876 ,w__4583 ,w__4126);
  or g__6499(w__4875 ,w__4587 ,w__4247);
  or g__6500(w__4874 ,w__4577 ,w__4244);
  nor g__6501(w__4872 ,w__4211 ,w__4181);
  nor g__6502(w__4871 ,w__4217 ,w__4466);
  nor g__6503(w__4870 ,w__4190 ,w__4469);
  nor g__6504(w__4869 ,w__4187 ,w__4467);
  nor g__6505(w__4868 ,w__4193 ,w__4454);
  nor g__6506(w__4867 ,w__4214 ,w__4468);
  nor g__6507(w__4866 ,w__4205 ,w__4470);
  or g__6508(w__4865 ,w__4676 ,w__4178);
  or g__6509(w__4864 ,w__4673 ,w__4183);
  or g__6510(w__4863 ,w__4667 ,w__4180);
  or g__6511(w__4862 ,w__4675 ,w__4177);
  or g__6512(w__4861 ,w__4663 ,w__4178);
  or g__6513(w__4860 ,w__4689 ,w__4118);
  or g__6514(w__4859 ,w__4640 ,w__4250);
  nor g__6515(w__4858 ,w__4184 ,w__4658);
  or g__6516(w__4857 ,w__4669 ,w__4183);
  or g__6517(w__4856 ,w__4686 ,w__4180);
  or g__6518(w__4855 ,w__4691 ,w__4184);
  or g__6519(w__4854 ,w__4692 ,w__4249);
  or g__6520(w__4853 ,w__4690 ,w__4249);
  or g__6521(w__4852 ,w__4693 ,w__4181);
  or g__6522(w__4851 ,w__4688 ,w__4118);
  or g__6523(w__4850 ,w__4611 ,w__4238);
  or g__6524(w__4847 ,w__4660 ,w__4378);
  or g__6525(w__4846 ,w__4208 ,w__4554);
  or g__6526(w__4845 ,w__4196 ,w__4559);
  nor g__6527(w__4844 ,w__4208 ,w__4564);
  nor g__6528(w__4843 ,w__4196 ,w__4566);
  or g__6529(w__4842 ,w__4195 ,w__4560);
  or g__6530(w__4841 ,w__4207 ,w__4558);
  or g__6531(w__4840 ,w__4198 ,w__4561);
  or g__6532(w__4839 ,w__4207 ,w__4567);
  or g__6533(w__4838 ,w__4195 ,w__4553);
  nor g__6534(w__4837 ,w__4199 ,w__4555);
  or g__6535(w__4836 ,w__4198 ,w__4565);
  or g__6536(w__4835 ,w__4199 ,w__4556);
  or g__6537(w__4834 ,w__4136 ,w__4562);
  or g__6538(w__4833 ,w__4136 ,w__4552);
  or g__6539(w__4832 ,w__4659 ,w__4417);
  or g__6540(w__4831 ,w__4586 ,w__4402);
  or g__6541(w__4830 ,w__4581 ,w__4366);
  nor g__6542(w__4829 ,w__4590 ,w__4409);
  or g__6543(w__4828 ,w__4611 ,w__4375);
  or g__6544(w__4827 ,w__4651 ,w__4420);
  or g__6545(w__4826 ,w__4589 ,w__4420);
  or g__6546(w__4825 ,w__4594 ,w__4387);
  or g__6547(w__4824 ,w__4685 ,w__4387);
  or g__6548(w__4823 ,w__4661 ,w__4375);
  or g__6549(w__4822 ,w__4572 ,w__4408);
  or g__6550(w__4821 ,w__4642 ,w__4390);
  or g__6551(w__4820 ,w__4591 ,w__4379);
  or g__6552(w__4819 ,w__4639 ,w__4382);
  or g__6553(w__4818 ,w__4613 ,w__4396);
  or g__6554(w__4817 ,w__4597 ,w__4378);
  or g__6555(w__4816 ,w__4580 ,w__4396);
  or g__6556(w__4815 ,w__4570 ,w__4391);
  or g__6557(w__4814 ,w__4671 ,w__4367);
  or g__6558(w__4813 ,w__4670 ,w__4418);
  or g__6559(w__4812 ,w__4574 ,w__4417);
  or g__6560(w__4811 ,w__4600 ,w__4342);
  nor g__6561(w__4810 ,w__4281 ,w__4563);
  or g__6562(w__4809 ,w__4678 ,w__4351);
  or g__6563(w__4808 ,w__4656 ,w__4351);
  or g__6564(w__4807 ,w__4609 ,w__4370);
  or g__6565(w__4806 ,w__4596 ,w__4343);
  or g__6566(w__4805 ,w__4687 ,w__4381);
  or g__6567(w__4804 ,w__4681 ,w__4403);
  or g__6568(w__4803 ,w__4638 ,w__4384);
  or g__6569(w__4802 ,w__4644 ,w__4394);
  or g__6570(w__4801 ,w__4602 ,w__4390);
  or g__6571(w__4800 ,w__4578 ,w__4393);
  or g__6572(w__4799 ,w__4650 ,w__4384);
  or g__6573(w__4798 ,w__4646 ,w__4346);
  or g__6574(w__4797 ,w__4682 ,w__4414);
  or g__6575(w__4796 ,w__4598 ,w__4545);
  or g__6576(w__4795 ,w__4657 ,w__4342);
  or g__6577(w__4794 ,w__4645 ,w__4399);
  or g__6578(w__4793 ,w__4641 ,w__4399);
  or g__6579(w__4792 ,w__4677 ,w__4414);
  or g__6580(w__4791 ,w__4573 ,w__4381);
  or g__6581(w__4790 ,w__4599 ,w__4406);
  or g__6582(w__4789 ,w__4647 ,w__4415);
  or g__6583(w__4788 ,w__4601 ,w__4418);
  or g__6584(w__4787 ,w__4605 ,w__4345);
  or g__6585(w__4786 ,w__4653 ,w__4366);
  or g__6586(w__4785 ,w__4595 ,w__4402);
  or g__6587(w__4784 ,w__4648 ,w__4393);
  or g__6588(w__4783 ,w__4654 ,w__4397);
  or g__6589(w__4782 ,w__4610 ,w__4421);
  or g__6590(w__4781 ,w__4608 ,w__4388);
  or g__6591(w__4780 ,w__4614 ,w__4405);
  or g__6592(w__4779 ,w__4668 ,w__4394);
  or g__6593(w__4778 ,w__4557 ,w__4311);
  or g__6594(w__4777 ,w__4662 ,w__4369);
  or g__6595(w__4776 ,w__4568 ,w__4412);
  or g__6596(w__4849 ,w__4534 ,w__4270);
  or g__6597(w__4848 ,in9[0] ,w__4623);
  not g__6598(w__4775 ,w__4774);
  not g__6599(w__4773 ,w__4772);
  not g__6600(w__4771 ,w__4770);
  not g__6601(w__4768 ,w__4767);
  not g__6602(w__4766 ,w__4765);
  not g__6603(w__4764 ,w__4763);
  not g__6604(w__4762 ,w__4761);
  or g__6605(w__4749 ,w__4604 ,w__4372);
  or g__6606(w__4748 ,w__4571 ,w__4348);
  or g__6607(w__4747 ,w__4683 ,w__4372);
  or g__6608(w__4746 ,w__4607 ,w__4348);
  or g__6609(w__4745 ,w__4612 ,w__4411);
  or g__6610(w__4744 ,w__4584 ,w__4405);
  or g__6611(w__4743 ,w__4674 ,w__4311);
  or g__6612(w__4742 ,w__4665 ,w__4408);
  or g__6613(w__4741 ,w__4606 ,w__4406);
  or g__6614(w__4740 ,w__4649 ,w__4345);
  or g__6615(w__4739 ,w__4569 ,w__4369);
  or g__6616(w__4738 ,w__4592 ,w__4421);
  or g__6617(w__4737 ,w__4587 ,w__4382);
  or g__6618(w__4736 ,w__4652 ,w__4352);
  or g__6619(w__4735 ,w__4593 ,w__4376);
  or g__6620(w__4734 ,w__4579 ,w__4346);
  or g__6621(w__4733 ,w__4577 ,w__4415);
  or g__6622(w__4732 ,w__4684 ,w__4349);
  or g__6623(w__4731 ,w__4672 ,w__4411);
  or g__6624(w__4730 ,w__4643 ,w__4385);
  or g__6625(w__4729 ,w__4680 ,w__4403);
  or g__6626(w__4728 ,w__4575 ,w__4370);
  or g__6627(w__4727 ,w__4666 ,w__4373);
  or g__6628(w__4726 ,w__4576 ,w__4379);
  or g__6629(w__4725 ,w__4603 ,w__4343);
  or g__6630(w__4724 ,w__4655 ,w__4400);
  or g__6631(w__4723 ,w__4551 ,w__4352);
  or g__6632(w__4722 ,w__4588 ,w__4391);
  or g__6633(w__4721 ,w__4585 ,w__4388);
  or g__6634(w__4720 ,w__4582 ,w__4409);
  or g__6635(w__4719 ,w__4664 ,w__4397);
  or g__6636(w__4718 ,w__4679 ,w__4367);
  or g__6637(w__4717 ,w__4583 ,w__4376);
  or g__6638(w__4716 ,w__4354 ,w__4673);
  or g__6639(w__4715 ,w__4363 ,w__4689);
  or g__6640(w__4714 ,w__4363 ,w__4640);
  or g__6641(w__4713 ,w__4355 ,w__4693);
  or g__6642(w__4712 ,w__4358 ,w__4690);
  or g__6643(w__4711 ,w__4354 ,w__4691);
  or g__6644(w__4710 ,w__4357 ,w__4686);
  or g__6645(w__4709 ,w__4360 ,w__4663);
  or g__6646(w__4708 ,w__4360 ,w__4692);
  or g__6647(w__4707 ,w__4357 ,w__4669);
  or g__6648(w__4706 ,w__4364 ,w__4658);
  or g__6649(w__4705 ,w__4358 ,w__4688);
  or g__6650(w__4704 ,w__4361 ,w__4667);
  or g__6651(w__4703 ,w__4355 ,w__4676);
  or g__6652(w__4702 ,w__4364 ,w__4675);
  or g__6653(w__4701 ,w__4241 ,w__4627);
  or g__6654(w__4700 ,w__4470 ,w__4630);
  or g__6655(w__4699 ,w__4468 ,w__4631);
  or g__6656(w__4698 ,w__4467 ,w__4629);
  or g__6657(w__4697 ,w__4469 ,w__4625);
  or g__6658(w__4696 ,w__4466 ,w__4626);
  or g__6659(w__4695 ,w__4454 ,w__4628);
  nor g__6660(w__4694 ,w__4412 ,w__4107);
  and g__6661(w__4774 ,in9[13] ,w__4273);
  and g__6662(w__4772 ,in9[7] ,w__4271);
  and g__6663(w__4770 ,in9[3] ,w__4264);
  and g__6664(w__4769 ,in9[15] ,w__4272);
  and g__6665(w__4767 ,in9[9] ,w__4275);
  and g__6666(w__4765 ,in9[11] ,w__4269);
  and g__6667(w__4763 ,in9[5] ,w__4265);
  and g__6668(w__4761 ,in8[0] ,w__4279);
  or g__6669(w__4760 ,w__4255 ,w__4373);
  or g__6670(w__4759 ,w__4255 ,w__4361);
  or g__6671(w__4758 ,w__4471 ,w__4400);
  or g__6672(w__4757 ,w__4254 ,w__4385);
  or g__6673(w__4756 ,w__4254 ,w__4349);
  or g__6674(w__4755 ,w__4622 ,w__4267);
  or g__6675(w__4754 ,w__4617 ,w__4276);
  or g__6676(w__4753 ,w__4615 ,w__4266);
  or g__6677(w__4752 ,w__4530 ,w__4278);
  or g__6678(w__4751 ,w__4618 ,w__4274);
  or g__6679(w__4750 ,w__4533 ,w__4268);
  not g__6680(w__4637 ,w__4271);
  not g__6681(w__4636 ,w__4276);
  not g__6682(w__4634 ,w__4270);
  not g__6683(w__4633 ,w__4272);
  nor g__6684(w__4631 ,w__4319 ,w__4517);
  nor g__6685(w__4630 ,w__4455 ,w__4480);
  nor g__6686(w__4629 ,w__4317 ,w__4486);
  nor g__6687(w__4628 ,w__4315 ,w__4519);
  nor g__6688(w__4627 ,w__4313 ,w__4481);
  nor g__6689(w__4626 ,w__4321 ,w__4506);
  nor g__6690(w__4625 ,w__4323 ,w__4511);
  or g__6691(w__4624 ,w__4502 ,w__4491);
  xnor g__6692(w__4622 ,in9[13] ,in9[12]);
  xnor g__6693(w__4621 ,in8[0] ,in9[3]);
  nor g__6694(w__4620 ,w__13690 ,w__4325);
  xnor g__6695(w__4619 ,in8[0] ,in9[9]);
  xnor g__6696(w__4618 ,in9[9] ,in9[8]);
  xnor g__6697(w__4617 ,in9[7] ,in9[6]);
  xnor g__6698(w__4616 ,in8[0] ,in9[5]);
  xnor g__6699(w__4615 ,in9[3] ,in9[2]);
  or g__6700(w__4693 ,w__4423 ,w__4510);
  or g__6701(w__4692 ,w__4498 ,w__4507);
  or g__6702(w__4691 ,w__4424 ,w__4520);
  or g__6703(w__4690 ,w__4434 ,w__4515);
  or g__6704(w__4689 ,w__4426 ,w__4512);
  or g__6705(w__4688 ,w__4433 ,w__4508);
  xnor g__6706(w__4687 ,in8[4] ,in9[13]);
  or g__6707(w__4686 ,w__4431 ,w__4483);
  xnor g__6708(w__4685 ,in8[1] ,in9[13]);
  xnor g__6709(w__4684 ,in8[4] ,in9[11]);
  xnor g__6710(w__4683 ,in8[6] ,in9[7]);
  xnor g__6711(w__4682 ,in8[13] ,in9[5]);
  xnor g__6712(w__4681 ,in8[4] ,in9[3]);
  xnor g__6713(w__4680 ,in8[2] ,in9[3]);
  xnor g__6714(w__4679 ,in8[7] ,in9[7]);
  xnor g__6715(w__4678 ,in8[9] ,in9[11]);
  xnor g__6716(w__4677 ,in8[10] ,in9[5]);
  or g__6717(w__4676 ,w__4425 ,w__4516);
  or g__6718(w__4675 ,w__4432 ,w__4484);
  xnor g__6719(w__4674 ,in8[5] ,in9[5]);
  or g__6720(w__4673 ,w__4430 ,w__4488);
  xnor g__6721(w__4672 ,in8[6] ,in9[3]);
  xnor g__6722(w__4671 ,in8[3] ,in9[7]);
  xnor g__6723(w__4670 ,in8[15] ,in9[5]);
  or g__6724(w__4669 ,w__4428 ,w__4509);
  xnor g__6725(w__4668 ,in8[3] ,in9[9]);
  or g__6726(w__4667 ,w__4427 ,w__4513);
  xnor g__6727(w__4666 ,in8[10] ,in9[7]);
  xnor g__6728(w__4665 ,in8[11] ,in9[3]);
  xnor g__6729(w__4664 ,in8[8] ,in9[9]);
  or g__6730(w__4663 ,w__4429 ,w__4518);
  xnor g__6731(w__4662 ,in8[15] ,in9[7]);
  xnor g__6732(w__4661 ,in8[11] ,in9[7]);
  xnor g__6733(w__4660 ,in8[10] ,in9[13]);
  xnor g__6734(w__4659 ,in8[1] ,in9[5]);
  xnor g__6735(w__4658 ,in8[15] ,in9[15]);
  xnor g__6736(w__4657 ,in8[2] ,in9[11]);
  xnor g__6737(w__4656 ,in8[3] ,in9[11]);
  xnor g__6738(w__4655 ,in8[14] ,in9[9]);
  xnor g__6739(w__4654 ,in8[12] ,in9[9]);
  xnor g__6740(w__4653 ,in8[12] ,in9[7]);
  xnor g__6741(w__4652 ,in8[8] ,in9[11]);
  xnor g__6742(w__4651 ,in8[11] ,in9[5]);
  xnor g__6743(w__4650 ,in8[8] ,in9[13]);
  xnor g__6744(w__4649 ,in8[1] ,in9[11]);
  xnor g__6745(w__4648 ,in8[2] ,in9[9]);
  xnor g__6746(w__4647 ,in8[8] ,in9[5]);
  xnor g__6747(w__4646 ,in8[13] ,in9[11]);
  xnor g__6748(w__4645 ,in8[4] ,in9[9]);
  xnor g__6749(w__4644 ,in8[5] ,in9[9]);
  xnor g__6750(w__4643 ,in8[2] ,in9[13]);
  xnor g__6751(w__4642 ,in8[9] ,in9[9]);
  xnor g__6752(w__4641 ,in8[13] ,in9[9]);
  or g__6753(w__4640 ,w__4309 ,w__4492);
  xnor g__6754(w__4639 ,in8[15] ,in9[13]);
  xnor g__6755(w__4638 ,in8[7] ,in9[13]);
  xnor g__6756(w__4635 ,w__4323 ,in9[6]);
  xnor g__6757(w__4632 ,w__4313 ,in9[14]);
  not g__6758(w__4550 ,w__4269);
  not g__6759(w__4549 ,w__4268);
  not g__6760(w__4547 ,w__4279);
  not g__6761(w__4545 ,w__4265);
  not g__6762(w__4544 ,w__4278);
  not g__6763(w__4543 ,w__4264);
  not g__6764(w__4542 ,w__4266);
  not g__6765(w__4540 ,w__4275);
  not g__6766(w__4539 ,w__4274);
  not g__6767(w__4537 ,w__4273);
  not g__6768(w__4536 ,w__4267);
  xnor g__6769(w__4534 ,in9[15] ,in9[14]);
  xnor g__6770(w__4533 ,in9[11] ,in9[10]);
  xnor g__6771(w__4532 ,in8[0] ,in9[11]);
  xnor g__6772(w__4531 ,in8[0] ,in9[13]);
  xnor g__6773(w__4530 ,in9[5] ,in9[4]);
  xnor g__6774(w__4529 ,in8[0] ,in9[1]);
  xnor g__6775(w__4528 ,in8[0] ,in9[7]);
  xnor g__6776(w__4614 ,in8[7] ,in9[3]);
  xnor g__6777(w__4613 ,in8[11] ,in9[9]);
  xnor g__6778(w__4612 ,in8[15] ,in9[3]);
  xnor g__6779(w__4611 ,in8[4] ,in9[7]);
  xnor g__6780(w__4610 ,in8[12] ,in9[5]);
  xnor g__6781(w__4609 ,in8[13] ,in9[7]);
  xnor g__6782(w__4608 ,in8[14] ,in9[13]);
  xnor g__6783(w__4607 ,in8[5] ,in9[11]);
  xnor g__6784(w__4606 ,in8[9] ,in9[3]);
  xnor g__6785(w__4605 ,in8[15] ,in9[11]);
  xnor g__6786(w__4604 ,in8[5] ,in9[7]);
  xnor g__6787(w__4603 ,in8[14] ,in9[11]);
  xnor g__6788(w__4602 ,in8[1] ,in9[9]);
  xnor g__6789(w__4601 ,in8[6] ,in9[5]);
  xnor g__6790(w__4600 ,in8[11] ,in9[11]);
  xnor g__6791(w__4599 ,in8[14] ,in9[3]);
  xnor g__6792(w__4598 ,in8[3] ,in9[5]);
  xnor g__6793(w__4597 ,in8[11] ,in9[13]);
  xnor g__6794(w__4596 ,in8[12] ,in9[11]);
  xnor g__6795(w__4595 ,in8[3] ,in9[3]);
  xnor g__6796(w__4594 ,in8[3] ,in9[13]);
  xnor g__6797(w__4593 ,in8[14] ,in9[7]);
  xnor g__6798(w__4592 ,in8[4] ,in9[5]);
  xnor g__6799(w__4591 ,in8[13] ,in9[13]);
  xnor g__6800(w__4590 ,in8[1] ,in9[3]);
  xnor g__6801(w__4589 ,in8[9] ,in9[5]);
  xnor g__6802(w__4588 ,in8[7] ,in9[9]);
  xnor g__6803(w__4587 ,in8[12] ,in9[13]);
  xnor g__6804(w__4586 ,in8[8] ,in9[3]);
  xnor g__6805(w__4585 ,in8[5] ,in9[13]);
  xnor g__6806(w__4584 ,in8[5] ,in9[3]);
  xnor g__6807(w__4583 ,in8[8] ,in9[7]);
  xnor g__6808(w__4582 ,in8[13] ,in9[3]);
  xnor g__6809(w__4581 ,in8[1] ,in9[7]);
  xnor g__6810(w__4580 ,in8[6] ,in9[9]);
  xnor g__6811(w__4579 ,in8[10] ,in9[11]);
  xnor g__6812(w__4578 ,in8[10] ,in9[9]);
  xnor g__6813(w__4577 ,in8[14] ,in9[5]);
  xnor g__6814(w__4576 ,in8[9] ,in9[13]);
  xnor g__6815(w__4575 ,in8[9] ,in9[7]);
  xnor g__6816(w__4574 ,in8[2] ,in9[5]);
  xnor g__6817(w__4573 ,in8[6] ,in9[13]);
  xnor g__6818(w__4572 ,in8[12] ,in9[3]);
  xnor g__6819(w__4571 ,in8[6] ,in9[11]);
  xnor g__6820(w__4570 ,in8[15] ,in9[9]);
  xnor g__6821(w__4569 ,in8[2] ,in9[7]);
  xnor g__6822(w__4568 ,in8[10] ,in9[3]);
  xnor g__6823(w__4567 ,in8[4] ,in9[1]);
  xnor g__6824(w__4566 ,in8[2] ,in9[1]);
  xnor g__6825(w__4565 ,in8[9] ,in9[1]);
  xnor g__6826(w__4564 ,in8[3] ,in9[1]);
  xnor g__6827(w__4563 ,in8[5] ,in9[1]);
  xnor g__6828(w__4562 ,in8[8] ,in9[1]);
  xnor g__6829(w__4561 ,in8[7] ,in9[1]);
  xnor g__6830(w__4560 ,in8[11] ,in9[1]);
  xnor g__6831(w__4559 ,in8[14] ,in9[1]);
  xnor g__6832(w__4558 ,in8[12] ,in9[1]);
  xnor g__6833(w__4557 ,in8[7] ,in9[5]);
  xnor g__6834(w__4556 ,in8[10] ,in9[1]);
  xnor g__6835(w__4555 ,in8[1] ,in9[1]);
  xnor g__6836(w__4554 ,in8[6] ,in9[1]);
  xnor g__6837(w__4553 ,in8[13] ,in9[1]);
  xnor g__6838(w__4552 ,in8[15] ,in9[1]);
  xnor g__6839(w__4551 ,in8[7] ,in9[11]);
  xnor g__6840(w__4548 ,w__4321 ,in9[10]);
  xnor g__6841(w__4546 ,w__4319 ,in9[4]);
  xnor g__6842(w__4541 ,w__4325 ,in9[2]);
  xnor g__6843(w__4538 ,w__4317 ,in9[8]);
  xnor g__6844(w__4535 ,w__4315 ,in9[12]);
  nor g__6845(w__4520 ,in8[2] ,in9[15]);
  nor g__6846(w__4519 ,in8[0] ,in9[12]);
  nor g__6847(w__4518 ,in8[4] ,in9[15]);
  nor g__6848(w__4517 ,in8[0] ,in9[4]);
  nor g__6849(w__4516 ,in8[5] ,in9[15]);
  nor g__6850(w__4515 ,in8[9] ,in9[15]);
  and g__6851(w__4514 ,in8[0] ,in9[6]);
  nor g__6852(w__4513 ,in8[13] ,in9[15]);
  nor g__6853(w__4512 ,in8[8] ,in9[15]);
  nor g__6854(w__4511 ,in8[0] ,in9[6]);
  nor g__6855(w__4510 ,in8[1] ,in9[15]);
  nor g__6856(w__4509 ,in8[3] ,in9[15]);
  nor g__6857(w__4508 ,in8[7] ,in9[15]);
  nor g__6858(w__4507 ,in8[6] ,in9[15]);
  nor g__6859(w__4506 ,in8[0] ,in9[10]);
  or g__6860(w__4505 ,w__4475 ,w__4138);
  or g__6861(w__4527 ,w__4477 ,w__4162);
  or g__6862(w__4526 ,w__4478 ,w__4240);
  or g__6863(w__4525 ,w__4460 ,w__4210);
  or g__6864(w__4524 ,w__4464 ,w__4139);
  or g__6865(w__4523 ,w__4473 ,w__4163);
  or g__6866(w__4522 ,w__4472 ,w__4124);
  or g__6867(w__4521 ,w__4463 ,w__4210);
  not g__6868(w__4501 ,w__4502);
  not g__6869(w__4498 ,w__4499);
  not g__6870(w__4493 ,w__4494);
  nor g__6871(w__4492 ,in8[14] ,in9[15]);
  nor g__6872(w__4491 ,in8[0] ,in9[15]);
  and g__6873(w__4490 ,in8[0] ,in9[14]);
  and g__6874(w__4489 ,in8[0] ,in9[2]);
  nor g__6875(w__4488 ,in8[12] ,in9[15]);
  and g__6876(w__4487 ,in8[0] ,in9[10]);
  nor g__6877(w__4486 ,in8[0] ,in9[8]);
  and g__6878(w__4485 ,in8[0] ,in9[12]);
  nor g__6879(w__4484 ,in8[10] ,in9[15]);
  nor g__6880(w__4483 ,in8[11] ,in9[15]);
  and g__6881(w__4482 ,in8[0] ,in9[8]);
  nor g__6882(w__4481 ,in8[0] ,in9[14]);
  nor g__6883(w__4480 ,in8[0] ,in9[2]);
  and g__6884(w__4479 ,in8[0] ,in9[4]);
  and g__6885(w__13690 ,in8[0] ,in9[0]);
  and g__6886(w__4504 ,in9[1] ,in9[0]);
  or g__6887(w__4503 ,w__4461 ,w__4138);
  and g__6888(w__4502 ,in8[0] ,in9[15]);
  or g__6889(w__4500 ,w__4459 ,w__4162);
  or g__6890(w__4499 ,w__4474 ,w__4240);
  or g__6891(w__4497 ,w__4465 ,w__4163);
  or g__6892(w__4496 ,w__4458 ,w__4139);
  or g__6893(w__4495 ,w__4476 ,w__4124);
  or g__6894(w__4494 ,w__4462 ,w__4211);
  not g__6895(w__4478 ,in8[7]);
  not g__6896(w__4477 ,in8[9]);
  not g__6897(w__4476 ,in8[1]);
  not g__6898(w__4475 ,in8[15]);
  not g__6899(w__4474 ,in8[6]);
  not g__6900(w__4473 ,in8[12]);
  not g__6901(w__4472 ,in8[4]);
  not g__6902(w__4471 ,in8[0]);
  not g__6903(w__4470 ,in9[3]);
  not g__6904(w__4469 ,in9[7]);
  not g__6905(w__4468 ,in9[5]);
  not g__6906(w__4467 ,in9[9]);
  not g__6907(w__4466 ,in9[11]);
  not g__6908(w__4465 ,in8[5]);
  not g__6909(w__4464 ,in8[11]);
  not g__6910(w__4463 ,in8[3]);
  not g__6911(w__4462 ,in8[14]);
  not g__6912(w__4461 ,in8[13]);
  not g__6913(w__4460 ,in8[10]);
  not g__6914(w__4459 ,in8[8]);
  not g__6915(w__4458 ,in8[2]);
  not g__6916(w__4457 ,in9[0]);
  not g__6917(w__4456 ,in9[15]);
  not g__6918(w__4455 ,in9[1]);
  not g__6919(w__4454 ,in9[13]);
  not g__6920(w__4108 ,w__4422);
  not g__6921(w__4422 ,w__4471);
  not g__6922(w__4421 ,w__4419);
  not g__6923(w__4420 ,w__4419);
  not g__6924(w__4419 ,w__4441);
  not g__6925(w__4418 ,w__4416);
  not g__6926(w__4417 ,w__4416);
  not g__6927(w__4416 ,w__4547);
  not g__6928(w__4415 ,w__4413);
  not g__6929(w__4414 ,w__4413);
  not g__6930(w__4413 ,w__4544);
  not g__6931(w__4412 ,w__4410);
  not g__6932(w__4411 ,w__4410);
  not g__6933(w__4410 ,w__4542);
  not g__6934(w__4409 ,w__4407);
  not g__6935(w__4408 ,w__4407);
  not g__6936(w__4407 ,w__4543);
  not g__6937(w__4406 ,w__4404);
  not g__6938(w__4405 ,w__4404);
  not g__6939(w__4404 ,w__4440);
  not g__6940(w__4403 ,w__4401);
  not g__6941(w__4402 ,w__4401);
  not g__6942(w__4401 ,w__4439);
  not g__6943(w__4400 ,w__4398);
  not g__6944(w__4399 ,w__4398);
  not g__6945(w__4398 ,w__4539);
  not g__6946(w__4397 ,w__4395);
  not g__6947(w__4396 ,w__4395);
  not g__6948(w__4395 ,w__4540);
  not g__6949(w__4394 ,w__4392);
  not g__6950(w__4393 ,w__4392);
  not g__6951(w__4392 ,w__4438);
  not g__6952(w__4391 ,w__4389);
  not g__6953(w__4390 ,w__4389);
  not g__6954(w__4389 ,w__4437);
  not g__6955(w__4388 ,w__4386);
  not g__6956(w__4387 ,w__4386);
  not g__6957(w__4386 ,w__4537);
  not g__6958(w__4385 ,w__4383);
  not g__6959(w__4384 ,w__4383);
  not g__6960(w__4383 ,w__4536);
  not g__6961(w__4382 ,w__4380);
  not g__6962(w__4381 ,w__4380);
  not g__6963(w__4380 ,w__4436);
  not g__6964(w__4379 ,w__4377);
  not g__6965(w__4378 ,w__4377);
  not g__6966(w__4377 ,w__4435);
  not g__6967(w__4376 ,w__4374);
  not g__6968(w__4375 ,w__4374);
  not g__6969(w__4374 ,w__4637);
  not g__6970(w__4373 ,w__4371);
  not g__6971(w__4372 ,w__4371);
  not g__6972(w__4371 ,w__4636);
  not g__6973(w__4370 ,w__4368);
  not g__6974(w__4369 ,w__4368);
  not g__6975(w__4368 ,w__4447);
  not g__6976(w__4367 ,w__4365);
  not g__6977(w__4366 ,w__4365);
  not g__6978(w__4365 ,w__4446);
  not g__6979(w__4364 ,w__4362);
  not g__6980(w__4363 ,w__4362);
  not g__6981(w__4362 ,w__4634);
  not g__6982(w__4361 ,w__4359);
  not g__6983(w__4360 ,w__4359);
  not g__6984(w__4359 ,w__4633);
  not g__6985(w__4358 ,w__4356);
  not g__6986(w__4357 ,w__4356);
  not g__6987(w__4356 ,w__4445);
  not g__6988(w__4355 ,w__4353);
  not g__6989(w__4354 ,w__4353);
  not g__6990(w__4353 ,w__4444);
  not g__6991(w__4352 ,w__4350);
  not g__6992(w__4351 ,w__4350);
  not g__6993(w__4350 ,w__4550);
  not g__6994(w__4349 ,w__4347);
  not g__6995(w__4348 ,w__4347);
  not g__6996(w__4347 ,w__4549);
  not g__6997(w__4346 ,w__4344);
  not g__6998(w__4345 ,w__4344);
  not g__6999(w__4344 ,w__4443);
  not g__7000(w__4343 ,w__4341);
  not g__7001(w__4342 ,w__4341);
  not g__7002(w__4341 ,w__4442);
  not g__7003(w__4340 ,w__4430);
  not g__7004(w__4430 ,w__4523);
  not g__7005(w__4339 ,w__4427);
  not g__7006(w__4427 ,w__4503);
  not g__7007(w__4338 ,w__4434);
  not g__7008(w__4434 ,w__4527);
  not g__7009(w__4337 ,w__4431);
  not g__7010(w__4431 ,w__4524);
  not g__7011(w__4336 ,w__4432);
  not g__7012(w__4432 ,w__4525);
  not g__7013(w__4335 ,w__4428);
  not g__7014(w__4428 ,w__4521);
  not g__7015(w__4334 ,w__4426);
  not g__7016(w__4426 ,w__4500);
  not g__7017(w__4333 ,w__4424);
  not g__7018(w__4424 ,w__4496);
  not g__7019(w__4332 ,w__4425);
  not g__7020(w__4425 ,w__4497);
  not g__7021(w__4331 ,w__4423);
  not g__7022(w__4423 ,w__4495);
  not g__7023(w__4330 ,w__4429);
  not g__7024(w__4429 ,w__4522);
  not g__7025(w__4329 ,w__4433);
  not g__7026(w__4433 ,w__4526);
  not g__7027(w__4328 ,w__4327);
  not g__7028(w__4327 ,w__5082);
  not g__7029(w__4326 ,w__4448);
  not g__7030(w__4448 ,w__5085);
  not g__7031(w__4325 ,w__4324);
  not g__7032(w__4324 ,w__4455);
  not g__7033(w__4323 ,w__4322);
  not g__7034(w__4322 ,w__4468);
  not g__7035(w__4321 ,w__4320);
  not g__7036(w__4320 ,w__4467);
  not g__7037(w__4319 ,w__4318);
  not g__7038(w__4318 ,w__4470);
  not g__7039(w__4317 ,w__4316);
  not g__7040(w__4316 ,w__4469);
  not g__7041(w__4315 ,w__4314);
  not g__7042(w__4314 ,w__4466);
  not g__7043(w__4313 ,w__4312);
  not g__7044(w__4312 ,w__4454);
  not g__7045(w__4311 ,w__4310);
  not g__7046(w__4310 ,w__4545);
  buf g__7047(w__13688 ,w__4694);
  buf g__7048(w__13689 ,w__4620);
  not g__7049(w__4309 ,w__4308);
  not g__7050(w__4308 ,w__4493);
  not g__7051(w__4307 ,w__4306);
  not g__7052(w__4306 ,w__5083);
  not g__7053(w__4305 ,w__4450);
  not g__7054(w__4450 ,w__5439);
  not g__7055(w__4304 ,w__4451);
  not g__7056(w__4451 ,w__5455);
  not g__7057(w__4303 ,w__4452);
  not g__7058(w__4452 ,w__5695);
  not g__7059(w__4302 ,w__4449);
  not g__7060(w__4449 ,w__5438);
  not g__7061(w__4301 ,w__4453);
  not g__7062(w__4453 ,w__5696);
  not g__7063(w__4300 ,w__4299);
  not g__7064(w__4299 ,w__4848);
  not g__7065(w__4298 ,w__4297);
  not g__7066(w__4297 ,w__4755);
  not g__7067(w__4296 ,w__4295);
  not g__7068(w__4295 ,w__4754);
  not g__7069(w__4294 ,w__4293);
  not g__7070(w__4293 ,w__4751);
  not g__7071(w__4292 ,w__4291);
  not g__7072(w__4291 ,w__4750);
  not g__7073(w__4290 ,w__4289);
  not g__7074(w__4289 ,w__4753);
  not g__7075(w__4288 ,w__4287);
  not g__7076(w__4287 ,w__4752);
  not g__7077(w__4286 ,w__4285);
  not g__7078(w__4285 ,w__4456);
  not g__7079(w__4284 ,w__4283);
  not g__7080(w__4283 ,w__4849);
  not g__7081(w__4282 ,w__4280);
  not g__7082(w__4281 ,w__4280);
  not g__7083(w__4280 ,w__4457);
  not g__7084(w__4279 ,w__4277);
  not g__7085(w__4278 ,w__4277);
  not g__7086(w__4277 ,w__4546);
  not g__7087(w__4276 ,w__4446);
  not g__7088(w__4446 ,w__4635);
  not g__7089(w__4275 ,w__4438);
  not g__7090(w__4438 ,w__4538);
  not g__7091(w__4274 ,w__4437);
  not g__7092(w__4437 ,w__4538);
  not g__7093(w__4273 ,w__4436);
  not g__7094(w__4436 ,w__4535);
  not g__7095(w__4272 ,w__4444);
  not g__7096(w__4444 ,w__4632);
  not g__7097(w__4271 ,w__4447);
  not g__7098(w__4447 ,w__4635);
  not g__7099(w__4270 ,w__4445);
  not g__7100(w__4445 ,w__4632);
  not g__7101(w__4269 ,w__4443);
  not g__7102(w__4443 ,w__4548);
  not g__7103(w__4268 ,w__4442);
  not g__7104(w__4442 ,w__4548);
  not g__7105(w__4267 ,w__4435);
  not g__7106(w__4435 ,w__4535);
  not g__7107(w__4266 ,w__4439);
  not g__7108(w__4439 ,w__4541);
  not g__7109(w__4265 ,w__4441);
  not g__7110(w__4441 ,w__4546);
  not g__7111(w__4264 ,w__4440);
  not g__7112(w__4440 ,w__4541);
  not g__7113(w__4263 ,w__4262);
  not g__7114(w__4262 ,w__5002);
  not g__7115(w__4261 ,w__4260);
  not g__7116(w__4260 ,w__5079);
  not g__7117(w__4259 ,w__4258);
  not g__7118(w__4258 ,w__5004);
  not g__7119(w__4257 ,w__4256);
  not g__7120(w__4256 ,w__5000);
  not g__7121(w__4107 ,w__4116);
  not g__7122(w__4255 ,w__4116);
  not g__7123(w__4116 ,w__4108);
  not g__7124(w__4254 ,w__4422);
  not g__7125(w__4253 ,w__4251);
  not g__7126(w__4252 ,w__4251);
  not g__7127(w__4251 ,w__4848);
  not g__7128(w__4250 ,w__4248);
  not g__7129(w__4249 ,w__4248);
  not g__7130(w__4248 ,w__4849);
  not g__7131(w__4247 ,w__4245);
  not g__7132(w__4246 ,w__4245);
  not g__7133(w__4245 ,w__4755);
  not g__7134(w__4244 ,w__4242);
  not g__7135(w__4243 ,w__4242);
  not g__7136(w__4242 ,w__4752);
  not g__7137(w__4241 ,w__4239);
  not g__7138(w__4240 ,w__4239);
  not g__7139(w__4239 ,w__4456);
  not g__7140(w__4238 ,w__4236);
  not g__7141(w__4237 ,w__4236);
  not g__7142(w__4236 ,w__4754);
  not g__7143(w__4235 ,w__4233);
  not g__7144(w__4234 ,w__4233);
  not g__7145(w__4233 ,w__4753);
  not g__7146(w__4232 ,w__4230);
  not g__7147(w__4231 ,w__4230);
  not g__7148(w__4230 ,w__4751);
  not g__7149(w__4229 ,w__4227);
  not g__7150(w__4228 ,w__4227);
  not g__7151(w__4227 ,w__4750);
  not g__7152(w__4226 ,w__4224);
  not g__7153(w__4225 ,w__4224);
  not g__7154(w__4224 ,w__4848);
  not g__7155(w__4223 ,w__4221);
  not g__7156(w__4222 ,w__4221);
  not g__7157(w__4221 ,w__4300);
  not g__7158(w__4220 ,w__4218);
  not g__7159(w__4219 ,w__4218);
  not g__7160(w__4218 ,w__4290);
  not g__7161(w__4217 ,w__4215);
  not g__7162(w__4216 ,w__4215);
  not g__7163(w__4215 ,w__4292);
  not g__7164(w__4214 ,w__4212);
  not g__7165(w__4213 ,w__4212);
  not g__7166(w__4212 ,w__4288);
  not g__7167(w__4211 ,w__4209);
  not g__7168(w__4210 ,w__4209);
  not g__7169(w__4209 ,w__4286);
  not g__7170(w__4208 ,w__4206);
  not g__7171(w__4207 ,w__4206);
  not g__7172(w__4206 ,w__4282);
  not g__7173(w__4205 ,w__4203);
  not g__7174(w__4204 ,w__4203);
  not g__7175(w__4203 ,w__4753);
  not g__7176(w__4202 ,w__4200);
  not g__7177(w__4201 ,w__4200);
  not g__7178(w__4200 ,w__4300);
  not g__7179(w__4199 ,w__4197);
  not g__7180(w__4198 ,w__4197);
  not g__7181(w__4197 ,w__4457);
  not g__7182(w__4196 ,w__4194);
  not g__7183(w__4195 ,w__4194);
  not g__7184(w__4194 ,w__4457);
  not g__7185(w__4193 ,w__4191);
  not g__7186(w__4192 ,w__4191);
  not g__7187(w__4191 ,w__4298);
  not g__7188(w__4190 ,w__4188);
  not g__7189(w__4189 ,w__4188);
  not g__7190(w__4188 ,w__4296);
  not g__7191(w__4187 ,w__4185);
  not g__7192(w__4186 ,w__4185);
  not g__7193(w__4185 ,w__4294);
  not g__7194(w__4184 ,w__4182);
  not g__7195(w__4183 ,w__4182);
  not g__7196(w__4182 ,w__4849);
  not g__7197(w__4181 ,w__4179);
  not g__7198(w__4180 ,w__4179);
  not g__7199(w__4179 ,w__4284);
  not g__7200(w__4178 ,w__4176);
  not g__7201(w__4177 ,w__4176);
  not g__7202(w__4176 ,w__4284);
  not g__7203(w__4175 ,w__4173);
  not g__7204(w__4174 ,w__4173);
  not g__7205(w__4173 ,w__4752);
  not g__7206(w__4172 ,w__4170);
  not g__7207(w__4171 ,w__4170);
  not g__7208(w__4170 ,w__4292);
  not g__7209(w__4169 ,w__4167);
  not g__7210(w__4168 ,w__4167);
  not g__7211(w__4167 ,w__4751);
  not g__7212(w__4166 ,w__4164);
  not g__7213(w__4165 ,w__4164);
  not g__7214(w__4164 ,w__4288);
  not g__7215(w__4163 ,w__4161);
  not g__7216(w__4162 ,w__4161);
  not g__7217(w__4161 ,w__4286);
  not g__7218(w__4160 ,w__4158);
  not g__7219(w__4159 ,w__4158);
  not g__7220(w__4158 ,w__4750);
  not g__7221(w__4157 ,w__4155);
  not g__7222(w__4156 ,w__4155);
  not g__7223(w__4155 ,w__4754);
  not g__7224(w__4154 ,w__4152);
  not g__7225(w__4153 ,w__4152);
  not g__7226(w__4152 ,w__4290);
  not g__7227(w__4151 ,w__4149);
  not g__7228(w__4150 ,w__4149);
  not g__7229(w__4149 ,w__4294);
  not g__7230(w__4148 ,w__4146);
  not g__7231(w__4147 ,w__4146);
  not g__7232(w__4146 ,w__4298);
  not g__7233(w__4145 ,w__4143);
  not g__7234(w__4144 ,w__4143);
  not g__7235(w__4143 ,w__4755);
  not g__7236(w__4142 ,w__4140);
  not g__7237(w__4141 ,w__4140);
  not g__7238(w__4140 ,w__4296);
  not g__7239(w__4139 ,w__4137);
  not g__7240(w__4138 ,w__4137);
  not g__7241(w__4137 ,w__4456);
  not g__7242(w__4136 ,w__4135);
  not g__7243(w__4135 ,w__4281);
  not g__7244(w__4134 ,w__4133);
  not g__7245(w__4133 ,w__4252);
  not g__7246(w__4132 ,w__4131);
  not g__7247(w__4131 ,w__4229);
  not g__7248(w__4130 ,w__4129);
  not g__7249(w__4129 ,w__4232);
  not g__7250(w__4128 ,w__4127);
  not g__7251(w__4127 ,w__4235);
  not g__7252(w__4126 ,w__4125);
  not g__7253(w__4125 ,w__4238);
  not g__7254(w__4124 ,w__4123);
  not g__7255(w__4123 ,w__4241);
  not g__7256(w__4122 ,w__4121);
  not g__7257(w__4121 ,w__4244);
  not g__7258(w__4120 ,w__4119);
  not g__7259(w__4119 ,w__4247);
  not g__7260(w__4118 ,w__4117);
  not g__7261(w__4117 ,w__4250);
  xor g__7262(w__4115 ,w__5697 ,w__5792);
  xor g__7263(w__13665 ,w__5673 ,w__5762);
  xor g__7264(w__4114 ,w__5655 ,w__5676);
  xor g__7265(w__4113 ,w__5314 ,w__5392);
  xor g__7266(w__4112 ,w__5308 ,w__4262);
  xor g__7267(w__4111 ,w__5418 ,w__4260);
  xor g__7268(w__4110 ,w__5297 ,w__4258);
  xor g__7269(w__4109 ,w__5405 ,w__4256);
  xnor g__7270(w__13479 ,w__7489 ,w__7524);
  xnor g__7271(w__13480 ,w__7492 ,w__5824);
  xnor g__7272(w__13482 ,w__7502 ,w__7516);
  xnor g__7273(w__13481 ,w__7498 ,w__7515);
  xnor g__7274(w__13478 ,w__7482 ,w__7517);
  or g__7275(w__13418 ,w__7487 ,w__7523);
  or g__7276(w__13417 ,w__7510 ,w__7522);
  or g__7277(w__13414 ,w__7505 ,w__7519);
  or g__7278(w__13413 ,w__7514 ,w__7521);
  or g__7279(w__13415 ,w__7503 ,w__7520);
  or g__7280(w__13416 ,w__7512 ,w__7518);
  xnor g__7281(w__13477 ,w__7468 ,w__7496);
  xnor g__7282(w__13483 ,w__7499 ,w__7495);
  xnor g__7283(w__13476 ,w__7470 ,w__7494);
  xnor g__7284(w__7524 ,w__7384 ,w__7500);
  and g__7285(w__7523 ,w__7476 ,w__7499);
  and g__7286(w__7522 ,w__7509 ,w__7502);
  or g__7287(w__13411 ,w__7484 ,w__7504);
  and g__7288(w__7521 ,w__7482 ,w__7506);
  nor g__7289(w__7520 ,w__7513 ,w__7501);
  or g__7290(w__13419 ,w__7466 ,w__7507);
  or g__7291(w__13412 ,w__7486 ,w__7508);
  and g__7292(w__7519 ,w__7497 ,w__7500);
  xnor g__7293(w__13484 ,w__7481 ,w__7473);
  xnor g__7294(w__13475 ,w__7469 ,w__7472);
  xnor g__7295(w__13485 ,w__7387 ,w__7474);
  nor g__7296(w__7518 ,w__7511 ,w__7498);
  xnor g__7297(w__7517 ,w__7478 ,w__7404);
  xnor g__7298(w__7516 ,w__7491 ,w__7405);
  xnor g__7299(w__7515 ,w__7479 ,w__7493);
  nor g__7300(w__7514 ,w__6012 ,w__7478);
  and g__7301(w__7513 ,w__7406 ,w__7492);
  nor g__7302(w__7512 ,w__7480 ,w__7493);
  and g__7303(w__7511 ,w__7480 ,w__7493);
  nor g__7304(w__7510 ,w__6010 ,w__7491);
  or g__7305(w__7509 ,w__6162 ,w__7490);
  nor g__7306(w__7508 ,w__7468 ,w__7485);
  and g__7307(w__7507 ,w__7465 ,w__7481);
  or g__7308(w__7506 ,w__6161 ,w__7477);
  nor g__7309(w__7505 ,w__7384 ,w__7489);
  nor g__7310(w__7504 ,w__7470 ,w__7483);
  nor g__7311(w__7503 ,w__7406 ,w__7492);
  or g__7312(w__7497 ,w__7383 ,w__7488);
  or g__7313(w__13474 ,w__7459 ,w__7475);
  xnor g__7314(w__13486 ,w__7413 ,w__5823);
  xnor g__7315(w__13488 ,w__7323 ,w__7443);
  xnor g__7316(w__13409 ,w__7391 ,w__7444);
  xnor g__7317(w__7496 ,w__7355 ,w__7450);
  xnor g__7318(w__7495 ,w__7453 ,w__7408);
  xnor g__7319(w__7494 ,w__7345 ,w__7454);
  xnor g__7320(w__7502 ,w__7390 ,w__7446);
  xnor g__7321(w__7501 ,w__7439 ,w__7442);
  xnor g__7322(w__7500 ,w__7416 ,w__7445);
  xnor g__7323(w__7499 ,w__7388 ,w__7440);
  xnor g__7324(w__7498 ,w__7412 ,w__7441);
  not g__7325(w__7490 ,w__7491);
  not g__7326(w__7488 ,w__7489);
  nor g__7327(w__7487 ,w__7408 ,w__7453);
  nor g__7328(w__7486 ,w__7355 ,w__7451);
  and g__7329(w__7485 ,w__7355 ,w__7451);
  or g__7330(w__13420 ,w__7430 ,w__7464);
  nor g__7331(w__7484 ,w__7345 ,w__7455);
  or g__7332(w__13421 ,w__7428 ,w__7463);
  or g__7333(w__13423 ,w__7424 ,w__7462);
  or g__7334(w__13473 ,w__7422 ,w__7460);
  and g__7335(w__7483 ,w__7345 ,w__7455);
  and g__7336(w__7493 ,w__7436 ,w__7456);
  and g__7337(w__7492 ,w__7419 ,w__7457);
  and g__7338(w__7491 ,w__7434 ,w__7467);
  and g__7339(w__7489 ,w__7425 ,w__7461);
  not g__7340(w__7480 ,w__7479);
  not g__7341(w__7477 ,w__7478);
  or g__7342(w__7476 ,w__7407 ,w__7452);
  nor g__7343(w__7475 ,w__7469 ,w__7458);
  or g__7344(w__13472 ,w__7418 ,w__7447);
  xnor g__7345(w__13487 ,w__7415 ,w__7396);
  or g__7346(w__13422 ,w__7376 ,w__7449);
  xnor g__7347(w__7474 ,w__7359 ,w__7411);
  xnor g__7348(w__7473 ,w__7403 ,w__7401);
  xnor g__7349(w__7472 ,w__7340 ,w__7409);
  xnor g__7350(w__7471 ,w__7414 ,w__7299);
  or g__7351(w__7482 ,w__7431 ,w__7448);
  xnor g__7352(w__7481 ,w__7342 ,w__7394);
  xnor g__7353(w__7479 ,w__7222 ,w__7393);
  xnor g__7354(w__7478 ,w__7389 ,w__7395);
  or g__7355(w__7467 ,w__7388 ,w__7432);
  nor g__7356(w__7466 ,w__7401 ,w__7403);
  or g__7357(w__7465 ,w__7400 ,w__7402);
  and g__7358(w__7464 ,w__7429 ,w__7411);
  nor g__7359(w__7463 ,w__7438 ,w__7413);
  and g__7360(w__7462 ,w__7323 ,w__7423);
  or g__7361(w__13424 ,w__7325 ,w__7421);
  or g__7362(w__7461 ,w__7439 ,w__7420);
  nor g__7363(w__7460 ,w__7397 ,w__7414);
  nor g__7364(w__7459 ,w__7340 ,w__7410);
  and g__7365(w__7458 ,w__7340 ,w__7410);
  or g__7366(w__7457 ,w__7412 ,w__7437);
  or g__7367(w__7456 ,w__7390 ,w__7435);
  and g__7368(w__7470 ,w__7317 ,w__7426);
  and g__7369(w__7469 ,w__7252 ,w__7399);
  and g__7370(w__7468 ,w__7380 ,w__7433);
  not g__7371(w__7455 ,w__7454);
  not g__7372(w__7452 ,w__7453);
  not g__7373(w__7451 ,w__7450);
  nor g__7374(w__7449 ,w__7377 ,w__7415);
  nor g__7375(w__7448 ,w__7427 ,w__7416);
  nor g__7376(w__7447 ,w__7391 ,w__7417);
  xnor g__7377(w__13489 ,w__7371 ,w__7351);
  xnor g__7378(w__13408 ,w__7320 ,w__7349);
  xnor g__7379(w__7446 ,w__7225 ,w__7357);
  xnor g__7380(w__7445 ,w__7344 ,w__7368);
  xnor g__7381(w__7444 ,w__7125 ,w__7366);
  xnor g__7382(w__7443 ,w__7363 ,w__7164);
  xnor g__7383(w__7442 ,w__7365 ,w__7339);
  xnor g__7384(w__7441 ,w__7354 ,w__7095);
  xnor g__7385(w__7440 ,w__7294 ,w__7361);
  xnor g__7386(w__7454 ,w__7370 ,w__7309);
  and g__7387(w__7453 ,w__7352 ,w__7398);
  xnor g__7388(w__7450 ,w__7392 ,w__7350);
  and g__7389(w__7438 ,w__7364 ,w__7385);
  and g__7390(w__7437 ,w__7095 ,w__7354);
  or g__7391(w__7436 ,w__7224 ,w__7357);
  nor g__7392(w__7435 ,w__7225 ,w__7356);
  or g__7393(w__7434 ,w__7294 ,w__7360);
  or g__7394(w__7433 ,w__7378 ,w__7389);
  nor g__7395(w__7432 ,w__7293 ,w__7361);
  nor g__7396(w__7431 ,w__7344 ,w__7369);
  nor g__7397(w__7430 ,w__7387 ,w__7359);
  or g__7398(w__7429 ,w__7386 ,w__7358);
  nor g__7399(w__7428 ,w__7364 ,w__7385);
  and g__7400(w__7427 ,w__7344 ,w__7369);
  or g__7401(w__7426 ,w__7327 ,w__7392);
  or g__7402(w__7425 ,w__7339 ,w__7365);
  nor g__7403(w__7424 ,w__6013 ,w__7363);
  or g__7404(w__7423 ,w__6160 ,w__7362);
  nor g__7405(w__7422 ,w__7299 ,w__7382);
  and g__7406(w__7421 ,w__7326 ,w__7371);
  and g__7407(w__7420 ,w__7339 ,w__7365);
  or g__7408(w__13470 ,w__7331 ,w__7373);
  or g__7409(w__13471 ,w__7334 ,w__7372);
  or g__7410(w__7419 ,w__7095 ,w__7354);
  nor g__7411(w__7418 ,w__7125 ,w__7367);
  and g__7412(w__7417 ,w__7125 ,w__7367);
  and g__7413(w__7439 ,w__7242 ,w__7381);
  not g__7414(w__7410 ,w__7409);
  not g__7415(w__7408 ,w__7407);
  not g__7416(w__7402 ,w__7403);
  not g__7417(w__7400 ,w__7401);
  xnor g__7418(w__13406 ,w__7093 ,w__7315);
  xnor g__7419(w__13490 ,w__7321 ,w__7308);
  or g__7420(w__7399 ,w__7286 ,w__7370);
  or g__7421(w__7398 ,w__7322 ,w__7353);
  and g__7422(w__7397 ,w__7299 ,w__7382);
  or g__7423(w__13425 ,w__7245 ,w__7379);
  xnor g__7424(w__13491 ,w__7217 ,w__7306);
  xnor g__7425(w__13407 ,w__7298 ,w__7312);
  xnor g__7426(w__7396 ,w__7256 ,w__7346);
  xnor g__7427(w__7395 ,w__7343 ,w__7255);
  xnor g__7428(w__7394 ,w__7130 ,w__7322);
  xnor g__7429(w__7393 ,w__7348 ,w__7158);
  xnor g__7430(w__7416 ,w__7123 ,w__7304);
  xnor g__7431(w__7415 ,w__7227 ,w__7305);
  xnor g__7432(w__7414 ,w__5821 ,w__7307);
  xnor g__7433(w__7413 ,w__7260 ,w__7314);
  and g__7434(w__7412 ,w__7251 ,w__7374);
  xnor g__7435(w__7411 ,w__7347 ,w__7313);
  xnor g__7436(w__7409 ,w__7261 ,w__7311);
  xnor g__7437(w__7407 ,w__7161 ,w__7310);
  xnor g__7438(w__7406 ,w__7087 ,w__7303);
  xnor g__7439(w__7405 ,w__7319 ,w__7300);
  xnor g__7440(w__7404 ,w__7162 ,w__7301);
  xnor g__7441(w__7403 ,w__7156 ,w__7302);
  and g__7442(w__7401 ,w__7280 ,w__7375);
  not g__7443(w__7386 ,w__7387);
  not g__7444(w__7383 ,w__7384);
  or g__7445(w__7381 ,w__7241 ,w__7348);
  or g__7446(w__7380 ,w__7255 ,w__7343);
  nor g__7447(w__7379 ,w__7244 ,w__7321);
  and g__7448(w__7378 ,w__7255 ,w__7343);
  and g__7449(w__7377 ,w__7257 ,w__7346);
  nor g__7450(w__7376 ,w__7257 ,w__7346);
  or g__7451(w__7375 ,w__7347 ,w__7277);
  or g__7452(w__7374 ,w__7249 ,w__7319);
  and g__7453(w__7373 ,w__7226 ,w__7333);
  and g__7454(w__7372 ,w__7320 ,w__7329);
  and g__7455(w__7392 ,w__7292 ,w__7336);
  and g__7456(w__7391 ,w__7265 ,w__7316);
  and g__7457(w__7390 ,w__7291 ,w__7337);
  and g__7458(w__7389 ,w__7247 ,w__7330);
  and g__7459(w__7388 ,w__7285 ,w__7335);
  and g__7460(w__7387 ,w__7276 ,w__7328);
  and g__7461(w__7385 ,w__7272 ,w__7338);
  and g__7462(w__7384 ,w__7270 ,w__7324);
  and g__7463(w__7382 ,w__7290 ,w__7332);
  not g__7464(w__7369 ,w__7368);
  not g__7465(w__7367 ,w__7366);
  not g__7466(w__7362 ,w__7363);
  not g__7467(w__7360 ,w__7361);
  not g__7468(w__7358 ,w__7359);
  not g__7469(w__7356 ,w__7357);
  xnor g__7470(w__13492 ,w__7173 ,w__5822);
  or g__7471(w__13426 ,w__7263 ,w__7318);
  nor g__7472(w__7353 ,w__7130 ,w__7341);
  or g__7473(w__7352 ,w__7129 ,w__7342);
  xnor g__7474(w__7351 ,w__7296 ,w__7147);
  xnor g__7475(w__7350 ,w__5819 ,w__7254);
  xnor g__7476(w__7349 ,w__7259 ,w__7148);
  xnor g__7477(w__7371 ,w__7180 ,w__7234);
  xnor g__7478(w__7370 ,w__7175 ,w__7231);
  xnor g__7479(w__7368 ,w__7132 ,w__5818);
  xnor g__7480(w__7366 ,w__7176 ,w__5820);
  xnor g__7481(w__7365 ,w__7169 ,w__7230);
  xnor g__7482(w__7364 ,w__7134 ,w__7228);
  xnor g__7483(w__7363 ,w__7174 ,w__7229);
  xnor g__7484(w__7361 ,w__7108 ,w__7236);
  xnor g__7485(w__7359 ,w__7181 ,w__7237);
  xnor g__7486(w__7357 ,w__7085 ,w__7233);
  xnor g__7487(w__7355 ,w__7166 ,w__7235);
  xnor g__7488(w__7354 ,w__7167 ,w__7232);
  not g__7489(w__7341 ,w__7342);
  or g__7490(w__7338 ,w__7227 ,w__7271);
  or g__7491(w__7337 ,w__7172 ,w__7289);
  or g__7492(w__7336 ,w__7171 ,w__7288);
  or g__7493(w__7335 ,w__7170 ,w__7283);
  nor g__7494(w__7334 ,w__6014 ,w__7259);
  or g__7495(w__7333 ,w__7119 ,w__7297);
  or g__7496(w__7332 ,w__7282 ,w__7262);
  nor g__7497(w__7331 ,w__7120 ,w__7298);
  or g__7498(w__13469 ,w__7182 ,w__7250);
  or g__7499(w__7330 ,w__7177 ,w__7246);
  or g__7500(w__7329 ,w__6159 ,w__7258);
  or g__7501(w__7328 ,w__7260 ,w__7274);
  or g__7502(w__13427 ,w__7190 ,w__7275);
  nor g__7503(w__7327 ,w__5819 ,w__7253);
  or g__7504(w__7326 ,w__6158 ,w__7295);
  nor g__7505(w__7325 ,w__6011 ,w__7296);
  or g__7506(w__7324 ,w__7168 ,w__7268);
  and g__7507(w__7348 ,w__7191 ,w__7278);
  and g__7508(w__7347 ,w__7209 ,w__7279);
  and g__7509(w__7346 ,w__7201 ,w__7269);
  and g__7510(w__7345 ,w__7205 ,w__7264);
  and g__7511(w__7344 ,w__7206 ,w__7273);
  and g__7512(w__7343 ,w__7214 ,w__7284);
  and g__7513(w__7342 ,w__7213 ,w__7281);
  and g__7514(w__7340 ,w__7198 ,w__7238);
  and g__7515(w__7339 ,w__7197 ,w__7266);
  or g__7516(w__13428 ,w__7038 ,w__7239);
  nor g__7517(w__7318 ,w__7179 ,w__7267);
  or g__7518(w__7317 ,w__7223 ,w__7254);
  xnor g__7519(w__13493 ,w__7178 ,w__7081);
  or g__7520(w__7316 ,w__5821 ,w__7287);
  xnor g__7521(w__7315 ,w__7165 ,w__6793);
  xnor g__7522(w__7314 ,w__7150 ,w__7151);
  xnor g__7523(w__7313 ,w__7153 ,w__7220);
  xnor g__7524(w__7312 ,w__7120 ,w__7226);
  xnor g__7525(w__7311 ,w__7154 ,w__7128);
  xnor g__7526(w__7310 ,w__7140 ,w__7172);
  xnor g__7527(w__7309 ,w__7100 ,w__7144);
  xnor g__7528(w__7308 ,w__7091 ,w__7146);
  xnor g__7529(w__7307 ,w__7142 ,w__7086);
  xnor g__7530(w__7306 ,w__7179 ,w__7103);
  xnor g__7531(w__7305 ,w__7149 ,w__7145);
  xnor g__7532(w__7304 ,w__7163 ,w__7177);
  xnor g__7533(w__7303 ,w__7159 ,w__7168);
  xnor g__7534(w__7302 ,w__7170 ,w__7116);
  xnor g__7535(w__7301 ,w__7171 ,w__7122);
  xnor g__7536(w__7300 ,w__7155 ,w__7141);
  or g__7537(w__7323 ,w__7196 ,w__7240);
  xnor g__7538(w__7322 ,w__7131 ,w__7138);
  xnor g__7539(w__7321 ,w__7106 ,w__7137);
  or g__7540(w__7320 ,w__7212 ,w__7243);
  and g__7541(w__7319 ,w__7184 ,w__7248);
  not g__7542(w__7297 ,w__7298);
  not g__7543(w__7295 ,w__7296);
  not g__7544(w__7293 ,w__7294);
  or g__7545(w__13468 ,w__6909 ,w__7187);
  or g__7546(w__7292 ,w__7122 ,w__7162);
  or g__7547(w__7291 ,w__7139 ,w__7161);
  or g__7548(w__7290 ,w__7128 ,w__7154);
  nor g__7549(w__7289 ,w__7140 ,w__7160);
  and g__7550(w__7288 ,w__7122 ,w__7162);
  and g__7551(w__7287 ,w__7086 ,w__7142);
  nor g__7552(w__7286 ,w__7100 ,w__7143);
  or g__7553(w__7285 ,w__7116 ,w__7156);
  or g__7554(w__7284 ,w__7132 ,w__7211);
  and g__7555(w__7283 ,w__7116 ,w__7156);
  and g__7556(w__7282 ,w__7128 ,w__7154);
  or g__7557(w__7281 ,w__7181 ,w__7210);
  or g__7558(w__7280 ,w__7153 ,w__7219);
  or g__7559(w__7279 ,w__7134 ,w__7208);
  or g__7560(w__7278 ,w__7104 ,w__7188);
  nor g__7561(w__7277 ,w__7152 ,w__7220);
  or g__7562(w__7276 ,w__7151 ,w__7150);
  nor g__7563(w__7275 ,w__7189 ,w__7173);
  and g__7564(w__7274 ,w__7151 ,w__7150);
  or g__7565(w__7273 ,w__7204 ,w__7169);
  or g__7566(w__7272 ,w__7145 ,w__7149);
  and g__7567(w__7271 ,w__7145 ,w__7149);
  or g__7568(w__7270 ,w__7087 ,w__7159);
  or g__7569(w__7269 ,w__7200 ,w__7174);
  and g__7570(w__7268 ,w__7087 ,w__7159);
  and g__7571(w__7267 ,w__7103 ,w__7218);
  or g__7572(w__7266 ,w__7193 ,w__7167);
  or g__7573(w__7265 ,w__7086 ,w__7142);
  or g__7574(w__7264 ,w__7192 ,w__7166);
  nor g__7575(w__7263 ,w__7103 ,w__7218);
  and g__7576(w__7299 ,w__6884 ,w__7207);
  and g__7577(w__7298 ,w__6925 ,w__7199);
  and g__7578(w__7296 ,w__7082 ,w__7194);
  and g__7579(w__7294 ,w__7109 ,w__7215);
  not g__7580(w__7262 ,w__7261);
  not g__7581(w__7258 ,w__7259);
  not g__7582(w__7257 ,w__7256);
  not g__7583(w__7253 ,w__7254);
  xnor g__7584(w__13405 ,w__7136 ,w__7030);
  or g__7585(w__7252 ,w__7099 ,w__7144);
  or g__7586(w__7251 ,w__7141 ,w__7155);
  nor g__7587(w__7250 ,w__7202 ,w__7165);
  and g__7588(w__7249 ,w__7141 ,w__7155);
  or g__7589(w__7248 ,w__7108 ,w__7195);
  or g__7590(w__7247 ,w__7123 ,w__7163);
  and g__7591(w__7246 ,w__7123 ,w__7163);
  nor g__7592(w__7245 ,w__7092 ,w__7146);
  and g__7593(w__7244 ,w__7092 ,w__7146);
  nor g__7594(w__7243 ,w__7203 ,w__7176);
  or g__7595(w__7242 ,w__7158 ,w__7221);
  nor g__7596(w__7241 ,w__7157 ,w__7222);
  nor g__7597(w__7240 ,w__7216 ,w__7180);
  nor g__7598(w__7239 ,w__7036 ,w__7178);
  or g__7599(w__7238 ,w__7186 ,w__7175);
  xnor g__7600(w__7237 ,w__7124 ,w__7126);
  xnor g__7601(w__7236 ,w__6916 ,w__7090);
  xnor g__7602(w__7235 ,w__7098 ,w__7115);
  xnor g__7603(w__7234 ,w__6913 ,w__7088);
  xnor g__7604(w__7233 ,w__7104 ,w__7102);
  xnor g__7605(w__7232 ,w__7096 ,w__7097);
  xnor g__7606(w__7231 ,w__7094 ,w__6713);
  xnor g__7607(w__7230 ,w__7117 ,w__7118);
  xnor g__7608(w__7229 ,w__7112 ,w__7113);
  xnor g__7609(w__7228 ,w__7121 ,w__7022);
  xnor g__7610(w__7261 ,w__7135 ,w__7028);
  and g__7611(w__7260 ,w__7058 ,w__7183);
  xnor g__7612(w__7259 ,w__7105 ,w__7015);
  xnor g__7613(w__7256 ,w__7133 ,w__7080);
  xnor g__7614(w__7255 ,w__7107 ,w__7016);
  and g__7615(w__7254 ,w__6863 ,w__7185);
  not g__7616(w__7224 ,w__7225);
  not g__7617(w__7223 ,w__5819);
  not g__7618(w__7221 ,w__7222);
  not g__7619(w__7219 ,w__7220);
  not g__7620(w__7218 ,w__7217);
  and g__7621(w__7216 ,w__6914 ,w__7088);
  or g__7622(w__7215 ,w__7110 ,w__7131);
  or g__7623(w__7214 ,w__6710 ,w__7114);
  or g__7624(w__7213 ,w__7126 ,w__7124);
  nor g__7625(w__7212 ,w__6789 ,w__7127);
  and g__7626(w__7211 ,w__6710 ,w__7114);
  and g__7627(w__7210 ,w__7126 ,w__7124);
  or g__7628(w__7209 ,w__7022 ,w__7121);
  and g__7629(w__7208 ,w__7022 ,w__7121);
  or g__7630(w__7207 ,w__6888 ,w__7135);
  or g__7631(w__7206 ,w__7118 ,w__7117);
  or g__7632(w__7205 ,w__7115 ,w__7098);
  and g__7633(w__7204 ,w__7118 ,w__7117);
  and g__7634(w__7203 ,w__6789 ,w__7127);
  nor g__7635(w__7202 ,w__6792 ,w__7093);
  or g__7636(w__7201 ,w__7113 ,w__7112);
  and g__7637(w__7200 ,w__7113 ,w__7112);
  or g__7638(w__7199 ,w__6880 ,w__7105);
  or g__7639(w__7198 ,w__6713 ,w__7094);
  or g__7640(w__7197 ,w__7097 ,w__7096);
  nor g__7641(w__7196 ,w__6914 ,w__7088);
  nor g__7642(w__7195 ,w__6916 ,w__7089);
  or g__7643(w__7194 ,w__7106 ,w__7083);
  and g__7644(w__7193 ,w__7097 ,w__7096);
  and g__7645(w__7192 ,w__7115 ,w__7098);
  or g__7646(w__7191 ,w__7085 ,w__7102);
  nor g__7647(w__7190 ,w__7023 ,w__7101);
  and g__7648(w__7189 ,w__7023 ,w__7101);
  or g__7649(w__13429 ,w__6876 ,w__7084);
  and g__7650(w__7188 ,w__7085 ,w__7102);
  nor g__7651(w__7187 ,w__6902 ,w__7136);
  and g__7652(w__7186 ,w__5968 ,w__7094);
  or g__7653(w__7185 ,w__6862 ,w__7107);
  or g__7654(w__7184 ,w__6915 ,w__7090);
  or g__7655(w__7183 ,w__7057 ,w__7133);
  and g__7656(w__7182 ,w__6016 ,w__7093);
  and g__7657(w__7227 ,w__6918 ,w__7111);
  xnor g__7658(w__7226 ,w__7008 ,w__6793);
  xnor g__7659(w__7225 ,w__6994 ,w__6035);
  xnor g__7660(w__7222 ,w__7027 ,w__6794);
  xnor g__7661(w__7220 ,w__6972 ,w__6986);
  xnor g__7662(w__7217 ,w__6917 ,w__6973);
  not g__7663(w__7160 ,w__7161);
  not g__7664(w__7157 ,w__7158);
  not g__7665(w__7152 ,w__7153);
  not g__7666(w__7143 ,w__7144);
  not g__7667(w__7139 ,w__7140);
  xnor g__7668(w__13495 ,w__6760 ,w__7013);
  xnor g__7669(w__13404 ,w__6983 ,w__6202);
  xnor g__7670(w__13494 ,w__7025 ,w__7003);
  xnor g__7671(w__7138 ,w__7021 ,w__6828);
  xnor g__7672(w__7137 ,w__7024 ,w__6745);
  xnor g__7673(w__7181 ,w__6826 ,w__7012);
  xnor g__7674(w__7180 ,w__6795 ,w__7014);
  xnor g__7675(w__7179 ,w__6839 ,w__7009);
  xnor g__7676(w__7178 ,w__6721 ,w__7010);
  xnor g__7677(w__7177 ,w__6985 ,w__6231);
  xnor g__7678(w__7176 ,w__6775 ,w__7005);
  xnor g__7679(w__7175 ,w__6998 ,w__6235);
  xnor g__7680(w__7174 ,w__6766 ,w__6978);
  xnor g__7681(w__7173 ,w__6842 ,w__6996);
  xnor g__7682(w__7172 ,w__6850 ,w__6991);
  xnor g__7683(w__7171 ,w__6773 ,w__6990);
  xnor g__7684(w__7170 ,w__6841 ,w__6988);
  xnor g__7685(w__7169 ,w__6840 ,w__6980);
  xnor g__7686(w__7168 ,w__6849 ,w__7019);
  xnor g__7687(w__7167 ,w__6843 ,w__6975);
  xnor g__7688(w__7166 ,w__6735 ,w__6974);
  xnor g__7689(w__7165 ,w__6984 ,w__6212);
  xnor g__7690(w__7164 ,w__7026 ,w__6977);
  xnor g__7691(w__7163 ,w__6772 ,w__7007);
  xnor g__7692(w__7162 ,w__6845 ,w__6992);
  xnor g__7693(w__7161 ,w__6747 ,w__7020);
  xnor g__7694(w__7159 ,w__6979 ,w__6791);
  xnor g__7695(w__7158 ,w__6813 ,w__7004);
  xnor g__7696(w__7156 ,w__6741 ,w__6989);
  xnor g__7697(w__7155 ,w__6860 ,w__7002);
  xnor g__7698(w__7154 ,w__6738 ,w__6993);
  xnor g__7699(w__7153 ,w__6808 ,w__6987);
  xnor g__7700(w__7151 ,w__6829 ,w__6982);
  xnor g__7701(w__7150 ,w__6847 ,w__6981);
  xnor g__7702(w__7149 ,w__6817 ,w__7001);
  xnor g__7703(w__7148 ,w__6976 ,w__6233);
  xnor g__7704(w__7147 ,w__6825 ,w__7000);
  xnor g__7705(w__7146 ,w__6763 ,w__6995);
  xnor g__7706(w__7145 ,w__6748 ,w__7011);
  xnor g__7707(w__7144 ,w__6809 ,w__6997);
  xnor g__7708(w__7142 ,w__6815 ,w__6999);
  xnor g__7709(w__7141 ,w__6728 ,w__7018);
  xnor g__7710(w__7140 ,w__6784 ,w__7029);
  not g__7711(w__7129 ,w__7130);
  not g__7712(w__7119 ,w__7120);
  or g__7713(w__7111 ,w__6926 ,w__7026);
  and g__7714(w__7110 ,w__6828 ,w__7021);
  or g__7715(w__7109 ,w__6828 ,w__7021);
  and g__7716(w__7136 ,w__6964 ,w__7048);
  and g__7717(w__7135 ,w__6969 ,w__7063);
  and g__7718(w__7134 ,w__6932 ,w__7060);
  and g__7719(w__7133 ,w__6923 ,w__7054);
  and g__7720(w__7132 ,w__6952 ,w__7067);
  and g__7721(w__7131 ,w__6960 ,w__7073);
  or g__7722(w__7130 ,w__6955 ,w__7068);
  and g__7723(w__7128 ,w__6962 ,w__7071);
  and g__7724(w__7127 ,w__6944 ,w__7056);
  and g__7725(w__7126 ,w__6949 ,w__7066);
  and g__7726(w__7125 ,w__6865 ,w__7078);
  and g__7727(w__7124 ,w__6945 ,w__7064);
  and g__7728(w__7123 ,w__6943 ,w__7062);
  and g__7729(w__7122 ,w__6967 ,w__7077);
  and g__7730(w__7121 ,w__6935 ,w__7061);
  and g__7731(w__7120 ,w__6963 ,w__7074);
  and g__7732(w__7118 ,w__6929 ,w__7059);
  and g__7733(w__7117 ,w__6924 ,w__7055);
  and g__7734(w__7116 ,w__6958 ,w__7072);
  and g__7735(w__7115 ,w__6922 ,w__7051);
  and g__7736(w__7114 ,w__6957 ,w__7070);
  and g__7737(w__7113 ,w__6908 ,w__7079);
  and g__7738(w__7112 ,w__6966 ,w__7050);
  not g__7739(w__7099 ,w__7100);
  not g__7740(w__7092 ,w__7091);
  not g__7741(w__7089 ,w__7090);
  and g__7742(w__7084 ,w__6883 ,w__7025);
  or g__7743(w__13430 ,w__6886 ,w__7034);
  and g__7744(w__7083 ,w__6745 ,w__7024);
  or g__7745(w__7082 ,w__6745 ,w__7024);
  xnor g__7746(w__7081 ,w__6719 ,w__6911);
  xnor g__7747(w__7080 ,w__6812 ,w__6971);
  and g__7748(w__7108 ,w__6939 ,w__7052);
  and g__7749(w__7107 ,w__6875 ,w__7032);
  and g__7750(w__7106 ,w__6904 ,w__7044);
  and g__7751(w__7105 ,w__6869 ,w__7033);
  and g__7752(w__7104 ,w__6882 ,w__7035);
  and g__7753(w__7103 ,w__6891 ,w__7042);
  and g__7754(w__7102 ,w__6931 ,w__7039);
  and g__7755(w__7101 ,w__6890 ,w__7041);
  or g__7756(w__7100 ,w__6868 ,w__7040);
  and g__7757(w__7098 ,w__6872 ,w__7045);
  and g__7758(w__7097 ,w__6903 ,w__7049);
  and g__7759(w__7096 ,w__6899 ,w__7046);
  and g__7760(w__7095 ,w__6881 ,w__7069);
  and g__7761(w__7094 ,w__6873 ,w__7075);
  or g__7762(w__7093 ,w__6867 ,w__7065);
  or g__7763(w__7091 ,w__6894 ,w__7053);
  and g__7764(w__7090 ,w__6878 ,w__7076);
  and g__7765(w__7088 ,w__6901 ,w__7047);
  and g__7766(w__7087 ,w__6910 ,w__7031);
  and g__7767(w__7086 ,w__6892 ,w__7037);
  and g__7768(w__7085 ,w__6861 ,w__7043);
  or g__7769(w__7079 ,w__6858 ,w__6907);
  or g__7770(w__7078 ,w__6859 ,w__6864);
  or g__7771(w__7077 ,w__6857 ,w__6965);
  or g__7772(w__7076 ,w__6856 ,w__6940);
  or g__7773(w__7075 ,w__6783 ,w__6874);
  or g__7774(w__7074 ,w__6961 ,w__6855);
  or g__7775(w__7073 ,w__6771 ,w__6959);
  or g__7776(w__7072 ,w__6854 ,w__6956);
  or g__7777(w__7071 ,w__6853 ,w__6953);
  or g__7778(w__7070 ,w__6851 ,w__6954);
  or g__7779(w__7069 ,w__6157 ,w__6951);
  and g__7780(w__7068 ,w__6972 ,w__6950);
  or g__7781(w__7067 ,w__6849 ,w__6947);
  or g__7782(w__7066 ,w__6848 ,w__6946);
  nor g__7783(w__7065 ,w__6870 ,w__6016);
  or g__7784(w__7064 ,w__6847 ,w__6941);
  or g__7785(w__7063 ,w__6785 ,w__6934);
  or g__7786(w__7062 ,w__6037 ,w__6938);
  or g__7787(w__7061 ,w__6846 ,w__6933);
  or g__7788(w__7060 ,w__6769 ,w__6930);
  or g__7789(w__7059 ,w__6774 ,w__6927);
  or g__7790(w__7058 ,w__6812 ,w__6970);
  nor g__7791(w__7057 ,w__6811 ,w__6971);
  or g__7792(w__7056 ,w__6844 ,w__6920);
  or g__7793(w__7055 ,w__6843 ,w__6919);
  or g__7794(w__7054 ,w__6766 ,w__6921);
  and g__7795(w__7053 ,w__6917 ,w__6948);
  or g__7796(w__7052 ,w__6841 ,w__6968);
  or g__7797(w__7051 ,w__6845 ,w__6936);
  or g__7798(w__7050 ,w__6762 ,w__6905);
  or g__7799(w__7049 ,w__6759 ,w__6900);
  or g__7800(w__7048 ,w__6897 ,w__6782);
  or g__7801(w__7047 ,w__6763 ,w__6898);
  or g__7802(w__7046 ,w__6860 ,w__6896);
  or g__7803(w__7045 ,w__6773 ,w__6893);
  or g__7804(w__7044 ,w__6778 ,w__6895);
  or g__7805(w__7043 ,w__6877 ,w__6784);
  or g__7806(w__7042 ,w__6842 ,w__6879);
  or g__7807(w__7041 ,w__6770 ,w__6889);
  and g__7808(w__7040 ,w__6871 ,w__5968);
  or g__7809(w__7039 ,w__6850 ,w__6887);
  nor g__7810(w__7038 ,w__6719 ,w__6912);
  or g__7811(w__7037 ,w__6852 ,w__6937);
  and g__7812(w__7036 ,w__6719 ,w__6912);
  or g__7813(w__7035 ,w__6781 ,w__6885);
  nor g__7814(w__7034 ,w__6760 ,w__6928);
  or g__7815(w__7033 ,w__6866 ,w__6775);
  or g__7816(w__7032 ,w__6772 ,w__6942);
  or g__7817(w__7031 ,w__6035 ,w__6906);
  xnor g__7818(w__13496 ,w__6786 ,w__6707);
  xnor g__7819(w__7030 ,w__6718 ,w__6018);
  xnor g__7820(w__7029 ,w__6752 ,w__6210);
  xnor g__7821(w__7028 ,w__6732 ,w__6711);
  xnor g__7822(w__7027 ,w__6797 ,w__6037);
  xnor g__7823(w__7020 ,w__6714 ,w__6781);
  xnor g__7824(w__7019 ,w__6831 ,w__6230);
  xnor g__7825(w__7018 ,w__6759 ,w__6204);
  xnor g__7826(w__7017 ,w__6859 ,w__6236);
  xnor g__7827(w__7016 ,w__5966 ,w__6206);
  xnor g__7828(w__7015 ,w__6801 ,w__6788);
  xnor g__7829(w__7014 ,w__6858 ,w__6465);
  xnor g__7830(w__7013 ,w__6470 ,w__6754);
  xnor g__7831(w__7012 ,w__6771 ,w__6468);
  xnor g__7832(w__7011 ,w__6846 ,w__6466);
  xnor g__7833(w__7010 ,w__6770 ,w__6469);
  xnor g__7834(w__7009 ,w__6778 ,w__6467);
  xnor g__7835(w__7008 ,w__6734 ,w__6232);
  xnor g__7836(w__7007 ,w__6796 ,w__6733);
  xnor g__7837(w__7006 ,w__6731 ,w__6208);
  xnor g__7838(w__7005 ,w__6729 ,w__6234);
  xnor g__7839(w__7004 ,w__6774 ,w__6205);
  xnor g__7840(w__7003 ,w__6756 ,w__6716);
  xnor g__7841(w__7002 ,w__6749 ,w__6724);
  xnor g__7842(w__7001 ,w__6816 ,w__6769);
  xnor g__7843(w__7000 ,w__6820 ,w__6762);
  xnor g__7844(w__6999 ,w__6844 ,w__6821);
  xnor g__7845(w__6998 ,w__6819 ,w__6785);
  xnor g__7846(w__6997 ,w__6853 ,w__6830);
  xnor g__7847(w__6996 ,w__6725 ,w__6727);
  xnor g__7848(w__6995 ,w__6717 ,w__6750);
  xnor g__7849(w__6994 ,w__6740 ,w__6736);
  xnor g__7850(w__6993 ,w__6852 ,w__6209);
  xnor g__7851(w__6992 ,w__6800 ,w__6804);
  xnor g__7852(w__6991 ,w__6720 ,w__6802);
  xnor g__7853(w__6990 ,w__6753 ,w__6737);
  xnor g__7854(w__6989 ,w__6739 ,w__6856);
  xnor g__7855(w__6988 ,w__6744 ,w__6814);
  xnor g__7856(w__6987 ,w__6823 ,w__6854);
  xnor g__7857(w__6986 ,w__6834 ,w__6836);
  xnor g__7858(w__6985 ,w__6857 ,w__6838);
  xnor g__7859(w__6984 ,w__6782 ,w__6832);
  xnor g__7860(w__6983 ,w__6214 ,w__6787);
  xnor g__7861(w__6982 ,w__6848 ,w__6827);
  xnor g__7862(w__6981 ,w__6746 ,w__6818);
  xnor g__7863(w__6980 ,w__6851 ,w__6803);
  xnor g__7864(w__6979 ,w__6822 ,w__6824);
  xnor g__7865(w__6978 ,w__6805 ,w__6807);
  xnor g__7866(w__6977 ,w__6798 ,w__6799);
  xnor g__7867(w__6976 ,w__6855 ,w__6837);
  xnor g__7868(w__6975 ,w__6806 ,w__6810);
  xnor g__7869(w__6974 ,w__6726 ,w__6783);
  xnor g__7870(w__6973 ,w__6743 ,w__6723);
  xnor g__7871(w__7026 ,w__6779 ,w__6701);
  xnor g__7872(w__7025 ,w__6695 ,w__6761);
  xnor g__7873(w__7024 ,w__6703 ,w__6757);
  xnor g__7874(w__7023 ,w__6705 ,w__6767);
  xnor g__7875(w__7022 ,w__6699 ,w__6764);
  xnor g__7876(w__7021 ,w__6697 ,w__6776);
  not g__7877(w__6970 ,w__6971);
  or g__7878(w__6969 ,w__6038 ,w__6819);
  and g__7879(w__6968 ,w__6814 ,w__6744);
  or g__7880(w__6967 ,w__6039 ,w__6838);
  or g__7881(w__6966 ,w__6820 ,w__6825);
  and g__7882(w__6965 ,w__6231 ,w__6838);
  or g__7883(w__6964 ,w__6048 ,w__6832);
  or g__7884(w__6963 ,w__6046 ,w__6837);
  or g__7885(w__6962 ,w__6830 ,w__6809);
  and g__7886(w__6961 ,w__6233 ,w__6837);
  or g__7887(w__6960 ,w__6468 ,w__6826);
  and g__7888(w__6959 ,w__6468 ,w__6826);
  or g__7889(w__6958 ,w__6823 ,w__6808);
  or g__7890(w__6957 ,w__6803 ,w__6840);
  and g__7891(w__6956 ,w__6823 ,w__6808);
  nor g__7892(w__6955 ,w__6836 ,w__6834);
  and g__7893(w__6954 ,w__6803 ,w__6840);
  and g__7894(w__6953 ,w__6830 ,w__6809);
  or g__7895(w__6952 ,w__6044 ,w__6831);
  and g__7896(w__6951 ,w__6736 ,w__6740);
  or g__7897(w__6950 ,w__6835 ,w__6833);
  or g__7898(w__6949 ,w__6829 ,w__6827);
  or g__7899(w__6948 ,w__6722 ,w__6742);
  and g__7900(w__6947 ,w__6230 ,w__6831);
  and g__7901(w__6946 ,w__6829 ,w__6827);
  or g__7902(w__6945 ,w__6818 ,w__6746);
  or g__7903(w__6944 ,w__6821 ,w__6815);
  or g__7904(w__6943 ,w__6824 ,w__6822);
  and g__7905(w__6942 ,w__6733 ,w__6796);
  and g__7906(w__6941 ,w__6818 ,w__6746);
  and g__7907(w__6940 ,w__6741 ,w__6739);
  or g__7908(w__6939 ,w__6814 ,w__6744);
  and g__7909(w__6938 ,w__6824 ,w__6822);
  and g__7910(w__6937 ,w__6043 ,w__6738);
  and g__7911(w__6936 ,w__6804 ,w__6800);
  or g__7912(w__6935 ,w__6466 ,w__6748);
  and g__7913(w__6934 ,w__6235 ,w__6819);
  and g__7914(w__6933 ,w__6466 ,w__6748);
  or g__7915(w__6932 ,w__6817 ,w__6816);
  or g__7916(w__6931 ,w__6802 ,w__6720);
  and g__7917(w__6930 ,w__6817 ,w__6816);
  or g__7918(w__6929 ,w__6042 ,w__6813);
  and g__7919(w__6928 ,w__6471 ,w__6754);
  and g__7920(w__6927 ,w__6205 ,w__6813);
  and g__7921(w__6926 ,w__6799 ,w__6798);
  or g__7922(w__6925 ,w__5970 ,w__6801);
  or g__7923(w__6924 ,w__6810 ,w__6806);
  or g__7924(w__6923 ,w__6807 ,w__6805);
  or g__7925(w__6922 ,w__6804 ,w__6800);
  and g__7926(w__6921 ,w__6807 ,w__6805);
  and g__7927(w__6920 ,w__6821 ,w__6815);
  and g__7928(w__6919 ,w__6810 ,w__6806);
  or g__7929(w__6918 ,w__6799 ,w__6798);
  and g__7930(w__6972 ,w__6700 ,w__6765);
  and g__7931(w__6971 ,w__6702 ,w__6780);
  not g__7932(w__6915 ,w__6916);
  not g__7933(w__6914 ,w__6913);
  not g__7934(w__6912 ,w__6911);
  or g__7935(w__6910 ,w__6790 ,w__6797);
  and g__7936(w__6909 ,w__6203 ,w__6718);
  or g__7937(w__6908 ,w__6465 ,w__6795);
  and g__7938(w__6907 ,w__6465 ,w__6795);
  and g__7939(w__6906 ,w__6790 ,w__6797);
  and g__7940(w__6905 ,w__6820 ,w__6825);
  or g__7941(w__6904 ,w__6467 ,w__6839);
  or g__7942(w__6903 ,w__6040 ,w__6728);
  nor g__7943(w__6902 ,w__6203 ,w__6718);
  or g__7944(w__6901 ,w__6750 ,w__6717);
  and g__7945(w__6900 ,w__6204 ,w__6728);
  or g__7946(w__6899 ,w__6724 ,w__6749);
  and g__7947(w__6898 ,w__6750 ,w__6717);
  and g__7948(w__6897 ,w__6212 ,w__6832);
  and g__7949(w__6896 ,w__6724 ,w__6749);
  and g__7950(w__6895 ,w__6467 ,w__6839);
  nor g__7951(w__6894 ,w__6723 ,w__6743);
  and g__7952(w__6893 ,w__6737 ,w__6753);
  or g__7953(w__6892 ,w__6209 ,w__6738);
  or g__7954(w__6891 ,w__6727 ,w__6725);
  or g__7955(w__6890 ,w__6469 ,w__6721);
  and g__7956(w__6889 ,w__6469 ,w__6721);
  and g__7957(w__6888 ,w__6732 ,w__6712);
  and g__7958(w__6887 ,w__6802 ,w__6720);
  nor g__7959(w__6886 ,w__6471 ,w__6754);
  and g__7960(w__6885 ,w__6747 ,w__6714);
  or g__7961(w__6884 ,w__6732 ,w__6712);
  or g__7962(w__6883 ,w__6715 ,w__6755);
  or g__7963(w__6882 ,w__6747 ,w__6714);
  or g__7964(w__6881 ,w__6736 ,w__6740);
  and g__7965(w__6880 ,w__5970 ,w__6801);
  and g__7966(w__6879 ,w__6727 ,w__6725);
  or g__7967(w__6878 ,w__6741 ,w__6739);
  nor g__7968(w__6877 ,w__6211 ,w__6752);
  nor g__7969(w__6876 ,w__6716 ,w__6756);
  or g__7970(w__6875 ,w__6733 ,w__6796);
  and g__7971(w__6874 ,w__6735 ,w__6726);
  or g__7972(w__6873 ,w__6735 ,w__6726);
  or g__7973(w__6872 ,w__6737 ,w__6753);
  or g__7974(w__6871 ,w__6207 ,w__6730);
  and g__7975(w__6870 ,w__6049 ,w__6734);
  or g__7976(w__6869 ,w__6045 ,w__6729);
  nor g__7977(w__6868 ,w__6208 ,w__6731);
  nor g__7978(w__6867 ,w__6049 ,w__6734);
  and g__7979(w__6866 ,w__6234 ,w__6729);
  or g__7980(w__6865 ,w__6047 ,w__5972);
  and g__7981(w__6864 ,w__6236 ,w__5972);
  or g__7982(w__6863 ,w__6041 ,w__5966);
  and g__7983(w__6862 ,w__6206 ,w__6709);
  or g__7984(w__6861 ,w__6210 ,w__6751);
  and g__7985(w__13431 ,w__6708 ,w__6786);
  and g__7986(w__6917 ,w__6706 ,w__6768);
  and g__7987(w__6916 ,w__6698 ,w__6777);
  and g__7988(w__6913 ,w__6704 ,w__6758);
  and g__7989(w__6911 ,w__6696 ,w__6761);
  not g__7990(w__6835 ,w__6836);
  not g__7991(w__6833 ,w__6834);
  not g__7992(w__6811 ,w__6812);
  not g__7993(w__6792 ,w__6793);
  not g__7994(w__6790 ,w__6791);
  not g__7995(w__6789 ,w__6788);
  or g__7996(w__6787 ,w__6478 ,w__6581);
  and g__7997(w__6860 ,w__6506 ,w__6610);
  and g__7998(w__6859 ,w__6529 ,w__6584);
  and g__7999(w__6858 ,w__6540 ,w__6623);
  and g__8000(w__6857 ,w__6417 ,w__6574);
  and g__8001(w__6856 ,w__6429 ,w__6587);
  and g__8002(w__6855 ,w__6528 ,w__6656);
  and g__8003(w__6854 ,w__6525 ,w__6657);
  and g__8004(w__6853 ,w__6524 ,w__6652);
  and g__8005(w__6852 ,w__6411 ,w__6562);
  and g__8006(w__6851 ,w__6522 ,w__6583);
  and g__8007(w__6850 ,w__6514 ,w__6638);
  and g__8008(w__6849 ,w__6516 ,w__6645);
  and g__8009(w__6848 ,w__6535 ,w__6643);
  and g__8010(w__6847 ,w__6511 ,w__6641);
  and g__8011(w__6846 ,w__6485 ,w__6636);
  and g__8012(w__6845 ,w__6520 ,w__6620);
  and g__8013(w__6844 ,w__6496 ,w__6693);
  and g__8014(w__6843 ,w__6500 ,w__6629);
  and g__8015(w__6842 ,w__6505 ,w__6602);
  and g__8016(w__6841 ,w__6455 ,w__6669);
  and g__8017(w__6840 ,w__6527 ,w__6655);
  and g__8018(w__6839 ,w__6448 ,w__6608);
  and g__8019(w__6838 ,w__6492 ,w__6667);
  or g__8020(w__6837 ,w__6474 ,w__6580);
  and g__8021(w__6836 ,w__6439 ,w__6650);
  and g__8022(w__6834 ,w__6441 ,w__6649);
  or g__8023(w__6832 ,w__6483 ,w__6577);
  and g__8024(w__6831 ,w__6518 ,w__6646);
  or g__8025(w__6830 ,w__6481 ,w__6579);
  and g__8026(w__6829 ,w__6533 ,w__6647);
  and g__8027(w__6828 ,w__6534 ,w__6664);
  and g__8028(w__6827 ,w__6517 ,w__6644);
  and g__8029(w__6826 ,w__6531 ,w__6663);
  and g__8030(w__6825 ,w__6497 ,w__6621);
  and g__8031(w__6824 ,w__6512 ,w__6588);
  and g__8032(w__6823 ,w__6426 ,w__6660);
  and g__8033(w__6822 ,w__6412 ,w__6570);
  or g__8034(w__6821 ,w__6476 ,w__6578);
  and g__8035(w__6820 ,w__6493 ,w__6622);
  and g__8036(w__6819 ,w__6421 ,w__6569);
  and g__8037(w__6818 ,w__6427 ,w__6642);
  and g__8038(w__6817 ,w__6504 ,w__6634);
  and g__8039(w__6816 ,w__6503 ,w__6633);
  and g__8040(w__6815 ,w__6419 ,w__6571);
  and g__8041(w__6814 ,w__6431 ,w__6606);
  and g__8042(w__6813 ,w__6442 ,w__6672);
  and g__8043(w__6812 ,w__6498 ,w__6680);
  and g__8044(w__6810 ,w__6445 ,w__6686);
  and g__8045(w__6809 ,w__6526 ,w__6658);
  and g__8046(w__6808 ,w__6501 ,w__6694);
  and g__8047(w__6807 ,w__6488 ,w__6668);
  and g__8048(w__6806 ,w__6495 ,w__6690);
  and g__8049(w__6805 ,w__6458 ,w__6559);
  or g__8050(w__6804 ,w__6472 ,w__6576);
  or g__8051(w__6803 ,w__6479 ,w__6575);
  and g__8052(w__6802 ,w__6457 ,w__6590);
  and g__8053(w__6801 ,w__6413 ,w__6573);
  and g__8054(w__6800 ,w__6486 ,w__6626);
  and g__8055(w__6799 ,w__6449 ,w__6619);
  and g__8056(w__6798 ,w__6487 ,w__6627);
  and g__8057(w__6797 ,w__6418 ,w__6566);
  and g__8058(w__6796 ,w__6444 ,w__6631);
  and g__8059(w__6795 ,w__6537 ,w__6625);
  and g__8060(w__6794 ,w__6532 ,w__6624);
  and g__8061(w__6793 ,w__6423 ,w__6572);
  and g__8062(w__6791 ,w__6509 ,w__6640);
  and g__8063(w__6788 ,w__6490 ,w__6628);
  not g__8064(w__6780 ,w__6779);
  not g__8065(w__6777 ,w__6776);
  not g__8066(w__6768 ,w__6767);
  not g__8067(w__6765 ,w__6764);
  not g__8068(w__6758 ,w__6757);
  not g__8069(w__6755 ,w__6756);
  not g__8070(w__6751 ,w__6752);
  not g__8071(w__6742 ,w__6743);
  not g__8072(w__6730 ,w__6731);
  not g__8073(w__6722 ,w__6723);
  not g__8074(w__6715 ,w__6716);
  not g__8075(w__6712 ,w__6711);
  not g__8076(w__6710 ,w__6709);
  or g__8077(w__13497 ,w__6552 ,w__6683);
  or g__8078(w__13498 ,w__6546 ,w__6659);
  or g__8079(w__13432 ,w__6538 ,w__6593);
  or g__8080(w__6786 ,w__6553 ,w__6675);
  and g__8081(w__6785 ,w__6507 ,w__6639);
  and g__8082(w__6784 ,w__6499 ,w__6603);
  and g__8083(w__6783 ,w__6556 ,w__6665);
  and g__8084(w__6782 ,w__6415 ,w__6568);
  and g__8085(w__6781 ,w__6436 ,w__6594);
  and g__8086(w__6779 ,w__6450 ,w__6685);
  and g__8087(w__6778 ,w__6543 ,w__6681);
  and g__8088(w__6776 ,w__6542 ,w__6674);
  and g__8089(w__6775 ,w__6425 ,w__6565);
  and g__8090(w__6774 ,w__6480 ,w__6678);
  and g__8091(w__6773 ,w__6414 ,w__6563);
  and g__8092(w__6772 ,w__6508 ,w__6671);
  and g__8093(w__6771 ,w__6554 ,w__6691);
  and g__8094(w__6770 ,w__6555 ,w__6679);
  and g__8095(w__6769 ,w__6550 ,w__6688);
  and g__8096(w__6767 ,w__6549 ,w__6687);
  and g__8097(w__6766 ,w__6551 ,w__6682);
  and g__8098(w__6764 ,w__6547 ,w__6689);
  and g__8099(w__6763 ,w__6545 ,w__6684);
  and g__8100(w__6762 ,w__6544 ,w__6692);
  or g__8101(w__6761 ,w__6519 ,w__6677);
  and g__8102(w__6760 ,w__6548 ,w__6676);
  and g__8103(w__6759 ,w__6416 ,w__6564);
  and g__8104(w__6757 ,w__6489 ,w__6616);
  and g__8105(w__6756 ,w__6494 ,w__6595);
  and g__8106(w__6754 ,w__6438 ,w__6597);
  and g__8107(w__6753 ,w__6502 ,w__6661);
  or g__8108(w__6752 ,w__6213 ,w__6673);
  and g__8109(w__6750 ,w__6510 ,w__6615);
  and g__8110(w__6749 ,w__6530 ,w__6651);
  and g__8111(w__6748 ,w__6456 ,w__6637);
  and g__8112(w__6747 ,w__6428 ,w__6648);
  and g__8113(w__6746 ,w__6451 ,w__6611);
  and g__8114(w__6745 ,w__6452 ,w__6609);
  and g__8115(w__6744 ,w__6536 ,w__6613);
  and g__8116(w__6743 ,w__6440 ,w__6612);
  and g__8117(w__6741 ,w__6437 ,w__6585);
  and g__8118(w__6740 ,w__6432 ,w__6666);
  and g__8119(w__6739 ,w__6422 ,w__6630);
  and g__8120(w__6738 ,w__6446 ,w__6589);
  and g__8121(w__6737 ,w__6435 ,w__6617);
  and g__8122(w__6736 ,w__6430 ,w__6586);
  and g__8123(w__6735 ,w__6515 ,w__6662);
  and g__8124(w__6734 ,w__6484 ,w__6670);
  and g__8125(w__6733 ,w__6473 ,w__6654);
  and g__8126(w__6732 ,w__6477 ,w__6635);
  and g__8127(w__6731 ,w__6482 ,w__6653);
  and g__8128(w__6729 ,w__6475 ,w__6592);
  and g__8129(w__6728 ,w__6454 ,w__6618);
  and g__8130(w__6727 ,w__6539 ,w__6605);
  and g__8131(w__6726 ,w__6424 ,w__6560);
  and g__8132(w__6725 ,w__6453 ,w__6604);
  or g__8133(w__6724 ,w__6213 ,w__6582);
  and g__8134(w__6723 ,w__6447 ,w__6607);
  and g__8135(w__6721 ,w__6513 ,w__6600);
  and g__8136(w__6720 ,w__6491 ,w__6599);
  and g__8137(w__6719 ,w__6521 ,w__6598);
  or g__8138(w__6718 ,w__6478 ,w__6567);
  and g__8139(w__6717 ,w__6523 ,w__6614);
  and g__8140(w__6716 ,w__6541 ,w__6596);
  and g__8141(w__6714 ,w__6420 ,w__6561);
  and g__8142(w__6713 ,w__6433 ,w__6601);
  and g__8143(w__6711 ,w__6434 ,w__6632);
  and g__8144(w__6709 ,w__6443 ,w__6591);
  not g__8145(w__6708 ,w__6707);
  not g__8146(w__6706 ,w__6705);
  not g__8147(w__6704 ,w__6703);
  not g__8148(w__6702 ,w__6701);
  not g__8149(w__6700 ,w__6699);
  not g__8150(w__6698 ,w__6697);
  not g__8151(w__6696 ,w__6695);
  or g__8152(w__6694 ,w__6298 ,w__5884);
  or g__8153(w__6693 ,w__6312 ,w__5869);
  or g__8154(w__6692 ,w__6274 ,w__5843);
  or g__8155(w__6691 ,w__6262 ,w__5935);
  or g__8156(w__6690 ,w__6370 ,w__5866);
  or g__8157(w__6689 ,w__6267 ,w__5843);
  or g__8158(w__6688 ,w__6269 ,w__5910);
  or g__8159(w__6687 ,w__6263 ,w__5931);
  or g__8160(w__6686 ,w__6260 ,w__5926);
  or g__8161(w__6685 ,w__6295 ,w__5862);
  or g__8162(w__6684 ,w__6271 ,w__5932);
  nor g__8163(w__6683 ,w__5934 ,w__6264);
  or g__8164(w__6682 ,w__6265 ,w__5910);
  or g__8165(w__6681 ,w__6270 ,w__5911);
  or g__8166(w__6680 ,w__6266 ,w__5923);
  or g__8167(w__6679 ,w__6272 ,w__5934);
  or g__8168(w__6678 ,w__6321 ,w__5928);
  nor g__8169(w__6677 ,w__5932 ,w__6276);
  or g__8170(w__6676 ,w__6273 ,w__5962);
  nor g__8171(w__6675 ,w__5935 ,w__6275);
  or g__8172(w__6674 ,w__6268 ,w__5961);
  nor g__8173(w__6673 ,w__5931 ,w__6261);
  or g__8174(w__6672 ,w__6391 ,w__5875);
  or g__8175(w__6671 ,w__6347 ,w__5854);
  or g__8176(w__6670 ,w__6348 ,w__5902);
  or g__8177(w__6669 ,w__6393 ,w__5881);
  or g__8178(w__6668 ,w__6357 ,w__5878);
  or g__8179(w__6667 ,w__6322 ,w__5896);
  or g__8180(w__6666 ,w__6280 ,w__5925);
  or g__8181(w__6665 ,w__6285 ,w__5857);
  or g__8182(w__6664 ,w__6352 ,w__5901);
  or g__8183(w__6663 ,w__6374 ,w__5943);
  or g__8184(w__6662 ,w__6309 ,w__5937);
  or g__8185(w__6661 ,w__6363 ,w__5860);
  or g__8186(w__6660 ,w__6388 ,w__5899);
  nor g__8187(w__6659 ,w__5911 ,w__6238);
  or g__8188(w__6658 ,w__6369 ,w__5955);
  or g__8189(w__6657 ,w__6353 ,w__5895);
  or g__8190(w__6656 ,w__6317 ,w__5856);
  or g__8191(w__6655 ,w__6287 ,w__5940);
  or g__8192(w__6654 ,w__6379 ,w__5922);
  or g__8193(w__6653 ,w__6371 ,w__5851);
  or g__8194(w__6652 ,w__6364 ,w__5859);
  or g__8195(w__6651 ,w__6373 ,w__5878);
  or g__8196(w__6650 ,w__6394 ,w__5854);
  or g__8197(w__6649 ,w__6365 ,w__5880);
  or g__8198(w__6648 ,w__6297 ,w__5877);
  or g__8199(w__6647 ,w__6240 ,w__5853);
  or g__8200(w__6646 ,w__6361 ,w__5869);
  or g__8201(w__6645 ,w__6362 ,w__5898);
  or g__8202(w__6644 ,w__6366 ,w__5868);
  or g__8203(w__6643 ,w__6356 ,w__5952);
  or g__8204(w__6642 ,w__6392 ,w__5946);
  or g__8205(w__6641 ,w__6354 ,w__5877);
  or g__8206(w__6640 ,w__6351 ,w__5860);
  or g__8207(w__6639 ,w__6305 ,w__5868);
  or g__8208(w__6638 ,w__6303 ,w__5853);
  or g__8209(w__6637 ,w__6313 ,w__5850);
  or g__8210(w__6636 ,w__6315 ,w__5928);
  or g__8211(w__6635 ,w__6279 ,w__5895);
  or g__8212(w__6634 ,w__6358 ,w__5881);
  or g__8213(w__6633 ,w__6377 ,w__5940);
  or g__8214(w__6632 ,w__6355 ,w__5925);
  or g__8215(w__6631 ,w__6318 ,w__5866);
  or g__8216(w__6707 ,w__6198 ,w__6409);
  or g__8217(w__6705 ,w__6223 ,w__6406);
  or g__8218(w__6703 ,w__6191 ,w__6407);
  or g__8219(w__6701 ,w__6196 ,w__6405);
  or g__8220(w__6699 ,w__6194 ,w__6404);
  or g__8221(w__6697 ,w__6199 ,w__6410);
  or g__8222(w__6695 ,w__6188 ,w__6408);
  or g__8223(w__6630 ,w__6333 ,w__5886);
  or g__8224(w__6629 ,w__6294 ,w__5857);
  or g__8225(w__6628 ,w__6300 ,w__5901);
  or g__8226(w__6627 ,w__6310 ,w__5874);
  or g__8227(w__6626 ,w__6302 ,w__5865);
  or g__8228(w__6625 ,w__6380 ,w__5865);
  or g__8229(w__6624 ,w__6375 ,w__5851);
  or g__8230(w__6623 ,w__6323 ,w__5837);
  or g__8231(w__6622 ,w__6311 ,w__5859);
  or g__8232(w__6621 ,w__6383 ,w__5884);
  or g__8233(w__6620 ,w__6288 ,w__5937);
  or g__8234(w__6619 ,w__6241 ,w__5880);
  or g__8235(w__6618 ,w__6308 ,w__5944);
  or g__8236(w__6617 ,w__6359 ,w__5955);
  or g__8237(w__6616 ,w__6381 ,w__5863);
  or g__8238(w__6615 ,w__6328 ,w__5839);
  or g__8239(w__6614 ,w__6278 ,w__5898);
  or g__8240(w__6613 ,w__6386 ,w__5883);
  or g__8241(w__6612 ,w__6293 ,w__5837);
  or g__8242(w__6611 ,w__6277 ,w__5913);
  or g__8243(w__6610 ,w__6319 ,w__5883);
  or g__8244(w__6609 ,w__6301 ,w__5875);
  or g__8245(w__6608 ,w__6290 ,w__5946);
  or g__8246(w__6607 ,w__6307 ,w__5922);
  or g__8247(w__6606 ,w__6289 ,w__5839);
  or g__8248(w__6605 ,w__6237 ,w__5850);
  or g__8249(w__6604 ,w__6390 ,w__5914);
  or g__8250(w__6603 ,w__6291 ,w__5913);
  or g__8251(w__6602 ,w__6283 ,w__5952);
  or g__8252(w__6601 ,w__6350 ,w__5941);
  or g__8253(w__6600 ,w__6304 ,w__5863);
  or g__8254(w__6599 ,w__6360 ,w__5874);
  or g__8255(w__6598 ,w__6368 ,w__5831);
  or g__8256(w__6597 ,w__6299 ,w__5929);
  or g__8257(w__6596 ,w__6325 ,w__5831);
  or g__8258(w__6595 ,w__6389 ,w__5862);
  or g__8259(w__6594 ,w__6284 ,w__5835);
  nor g__8260(w__6593 ,w__5929 ,w__6330);
  or g__8261(w__6592 ,w__6314 ,w__5841);
  or g__8262(w__6591 ,w__6387 ,w__5841);
  or g__8263(w__6590 ,w__6316 ,w__5938);
  or g__8264(w__6589 ,w__6306 ,w__5856);
  or g__8265(w__6588 ,w__6282 ,w__5829);
  or g__8266(w__6587 ,w__6281 ,w__5943);
  or g__8267(w__6586 ,w__6396 ,w__5829);
  or g__8268(w__6585 ,w__6292 ,w__5835);
  or g__8269(w__6584 ,w__6296 ,w__5956);
  or g__8270(w__6583 ,w__6286 ,w__5953);
  nor g__8271(w__6582 ,w__5962 ,w__6164);
  nor g__8272(w__6581 ,w__5920 ,w__5890);
  nor g__8273(w__6580 ,w__5926 ,w__6175);
  nor g__8274(w__6579 ,w__5899 ,w__6178);
  nor g__8275(w__6578 ,w__5896 ,w__6176);
  nor g__8276(w__6577 ,w__5902 ,w__6163);
  nor g__8277(w__6576 ,w__5923 ,w__6177);
  nor g__8278(w__6575 ,w__5914 ,w__6179);
  or g__8279(w__6574 ,w__6385 ,w__5887);
  or g__8280(w__6573 ,w__6382 ,w__5892);
  or g__8281(w__6572 ,w__6376 ,w__5889);
  or g__8282(w__6571 ,w__6384 ,w__5886);
  or g__8283(w__6570 ,w__6372 ,w__5887);
  or g__8284(w__6569 ,w__6398 ,w__5827);
  or g__8285(w__6568 ,w__6349 ,w__5959);
  nor g__8286(w__6567 ,w__5893 ,w__6367);
  or g__8287(w__6566 ,w__6378 ,w__5892);
  or g__8288(w__6565 ,w__6395 ,w__5889);
  or g__8289(w__6564 ,w__6400 ,w__5893);
  or g__8290(w__6563 ,w__6401 ,w__5958);
  or g__8291(w__6562 ,w__6399 ,w__5958);
  or g__8292(w__6561 ,w__6402 ,w__5890);
  or g__8293(w__6560 ,w__6397 ,w__5827);
  or g__8294(w__6559 ,w__6320 ,w__5947);
  or g__8295(w__6556 ,w__6369 ,w__6087);
  or g__8296(w__6555 ,w__5917 ,w__6263);
  or g__8297(w__6554 ,w__5905 ,w__6268);
  nor g__8298(w__6553 ,w__5917 ,w__6273);
  nor g__8299(w__6552 ,w__5905 ,w__6275);
  or g__8300(w__6551 ,w__5904 ,w__6269);
  or g__8301(w__6550 ,w__5916 ,w__6267);
  or g__8302(w__6549 ,w__5907 ,w__6270);
  or g__8303(w__6548 ,w__5916 ,w__6276);
  or g__8304(w__6547 ,w__5904 ,w__6262);
  nor g__8305(w__6546 ,w__5908 ,w__6264);
  or g__8306(w__6545 ,w__5907 ,w__6274);
  or g__8307(w__6544 ,w__5908 ,w__6265);
  or g__8308(w__6543 ,w__5845 ,w__6271);
  or g__8309(w__6542 ,w__5845 ,w__6261);
  or g__8310(w__6541 ,w__6368 ,w__6126);
  or g__8311(w__6540 ,w__6295 ,w__6111);
  or g__8312(w__6539 ,w__6290 ,w__6075);
  nor g__8313(w__6538 ,w__6299 ,w__6118);
  or g__8314(w__6537 ,w__6320 ,w__6084);
  or g__8315(w__6536 ,w__6360 ,w__6129);
  or g__8316(w__6535 ,w__6298 ,w__6129);
  or g__8317(w__6534 ,w__6303 ,w__6096);
  or g__8318(w__6533 ,w__6394 ,w__6096);
  or g__8319(w__6532 ,w__6370 ,w__6084);
  or g__8320(w__6531 ,w__6281 ,w__6117);
  or g__8321(w__6530 ,w__6351 ,w__6099);
  or g__8322(w__6529 ,w__6300 ,w__6088);
  or g__8323(w__6528 ,w__6348 ,w__6091);
  or g__8324(w__6527 ,w__6322 ,w__6105);
  or g__8325(w__6526 ,w__6306 ,w__6087);
  or g__8326(w__6525 ,w__6289 ,w__6105);
  or g__8327(w__6524 ,w__6279 ,w__6100);
  or g__8328(w__6523 ,w__6380 ,w__6076);
  or g__8329(w__6522 ,w__6379 ,w__6127);
  or g__8330(w__6521 ,w__6283 ,w__6126);
  or g__8331(w__6520 ,w__6309 ,w__6051);
  nor g__8332(w__6519 ,w__5990 ,w__6272);
  or g__8333(w__6518 ,w__6387 ,w__6060);
  or g__8334(w__6517 ,w__6365 ,w__6060);
  or g__8335(w__6516 ,w__6318 ,w__6079);
  or g__8336(w__6515 ,w__6305 ,w__6052);
  or g__8337(w__6514 ,w__6396 ,w__6090);
  or g__8338(w__6513 ,w__6390 ,w__6112);
  or g__8339(w__6512 ,w__6347 ,w__6093);
  or g__8340(w__6511 ,w__6353 ,w__6103);
  or g__8341(w__6510 ,w__6311 ,w__6099);
  or g__8342(w__6509 ,w__6287 ,w__6102);
  or g__8343(w__6508 ,w__6359 ,w__6093);
  or g__8344(w__6507 ,w__6355 ,w__6055);
  or g__8345(w__6506 ,w__6391 ,w__6123);
  or g__8346(w__6505 ,w__6307 ,w__6254);
  or g__8347(w__6504 ,w__6366 ,w__6051);
  or g__8348(w__6503 ,w__6354 ,w__6108);
  or g__8349(w__6502 ,w__6350 ,w__6108);
  or g__8350(w__6501 ,w__6386 ,w__6123);
  or g__8351(w__6500 ,w__6282 ,w__6090);
  or g__8352(w__6499 ,w__6308 ,w__6115);
  or g__8353(w__6498 ,w__6356 ,w__6124);
  or g__8354(w__6497 ,w__6310 ,w__6127);
  or g__8355(w__6496 ,w__6314 ,w__6054);
  or g__8356(w__6495 ,w__6362 ,w__6075);
  or g__8357(w__6494 ,w__6304 ,w__6111);
  or g__8358(w__6493 ,w__6357 ,w__6102);
  or g__8359(w__6492 ,w__6363 ,w__6106);
  or g__8360(w__6491 ,w__6319 ,w__6130);
  or g__8361(w__6490 ,w__6317 ,w__6097);
  or g__8362(w__6489 ,w__6323 ,w__6114);
  or g__8363(w__6488 ,w__6377 ,w__6103);
  or g__8364(w__6487 ,w__6266 ,w__6020);
  or g__8365(w__6486 ,w__6371 ,w__6078);
  or g__8366(w__6485 ,w__6277 ,w__6121);
  or g__8367(w__6558 ,w__6243 ,w__5979);
  or g__8368(w__6557 ,in13[0] ,w__6332);
  not g__8369(w__6484 ,w__6483);
  not g__8370(w__6482 ,w__6481);
  not g__8371(w__6480 ,w__6479);
  not g__8372(w__6477 ,w__6476);
  not g__8373(w__6475 ,w__6474);
  not g__8374(w__6473 ,w__6472);
  not g__8375(w__6471 ,w__6470);
  or g__8376(w__6458 ,w__6313 ,w__6081);
  or g__8377(w__6457 ,w__6280 ,w__6057);
  or g__8378(w__6456 ,w__6392 ,w__6081);
  or g__8379(w__6455 ,w__6316 ,w__6057);
  or g__8380(w__6454 ,w__6321 ,w__6120);
  or g__8381(w__6453 ,w__6293 ,w__6114);
  or g__8382(w__6452 ,w__6383 ,w__6020);
  or g__8383(w__6451 ,w__6374 ,w__6117);
  or g__8384(w__6450 ,w__6315 ,w__6115);
  or g__8385(w__6449 ,w__6358 ,w__6054);
  or g__8386(w__6448 ,w__6278 ,w__6078);
  or g__8387(w__6447 ,w__6301 ,w__6130);
  or g__8388(w__6446 ,w__6296 ,w__6091);
  or g__8389(w__6445 ,w__6361 ,w__6061);
  or g__8390(w__6444 ,w__6302 ,w__6085);
  or g__8391(w__6443 ,w__6288 ,w__6055);
  or g__8392(w__6442 ,w__6286 ,w__6124);
  or g__8393(w__6441 ,w__6393 ,w__6058);
  or g__8394(w__6440 ,w__6381 ,w__6120);
  or g__8395(w__6439 ,w__6352 ,w__6094);
  or g__8396(w__6438 ,w__6389 ,w__6112);
  or g__8397(w__6437 ,w__6284 ,w__6079);
  or g__8398(w__6436 ,w__6375 ,w__6082);
  or g__8399(w__6435 ,w__6285 ,w__6088);
  or g__8400(w__6434 ,w__6312 ,w__6052);
  or g__8401(w__6433 ,w__6364 ,w__6109);
  or g__8402(w__6432 ,w__6260 ,w__6061);
  or g__8403(w__6431 ,w__6297 ,w__6100);
  or g__8404(w__6430 ,w__6294 ,w__6097);
  or g__8405(w__6429 ,w__6291 ,w__6118);
  or g__8406(w__6428 ,w__6373 ,w__6106);
  or g__8407(w__6427 ,w__6388 ,w__6076);
  or g__8408(w__6426 ,w__6292 ,w__6085);
  or g__8409(w__6425 ,w__6063 ,w__6382);
  or g__8410(w__6424 ,w__6072 ,w__6398);
  or g__8411(w__6423 ,w__6072 ,w__6349);
  or g__8412(w__6422 ,w__6064 ,w__6402);
  or g__8413(w__6421 ,w__6067 ,w__6399);
  or g__8414(w__6420 ,w__6063 ,w__6400);
  or g__8415(w__6419 ,w__6066 ,w__6395);
  or g__8416(w__6418 ,w__6069 ,w__6372);
  or g__8417(w__6417 ,w__6069 ,w__6401);
  or g__8418(w__6416 ,w__6066 ,w__6378);
  or g__8419(w__6415 ,w__6073 ,w__6367);
  or g__8420(w__6414 ,w__6067 ,w__6397);
  or g__8421(w__6413 ,w__6070 ,w__6376);
  or g__8422(w__6412 ,w__6064 ,w__6385);
  or g__8423(w__6411 ,w__6073 ,w__6384);
  or g__8424(w__6410 ,w__5950 ,w__6336);
  or g__8425(w__6409 ,w__6179 ,w__6339);
  or g__8426(w__6408 ,w__6177 ,w__6340);
  or g__8427(w__6407 ,w__6176 ,w__6338);
  or g__8428(w__6406 ,w__6178 ,w__6334);
  or g__8429(w__6405 ,w__6175 ,w__6335);
  or g__8430(w__6404 ,w__6163 ,w__6337);
  nor g__8431(w__6403 ,w__6121 ,w__5816);
  and g__8432(w__6483 ,in13[13] ,w__5982);
  and g__8433(w__6481 ,in13[7] ,w__5980);
  and g__8434(w__6479 ,in13[3] ,w__5973);
  and g__8435(w__6478 ,in13[15] ,w__5981);
  and g__8436(w__6476 ,in13[9] ,w__5984);
  and g__8437(w__6474 ,in13[11] ,w__5978);
  and g__8438(w__6472 ,in13[5] ,w__5974);
  and g__8439(w__6470 ,in12[0] ,w__5988);
  or g__8440(w__6469 ,w__5964 ,w__6082);
  or g__8441(w__6468 ,w__5964 ,w__6070);
  or g__8442(w__6467 ,w__6180 ,w__6109);
  or g__8443(w__6466 ,w__5963 ,w__6094);
  or g__8444(w__6465 ,w__5963 ,w__6058);
  or g__8445(w__6464 ,w__6331 ,w__5976);
  or g__8446(w__6463 ,w__6326 ,w__5985);
  or g__8447(w__6462 ,w__6324 ,w__5975);
  or g__8448(w__6461 ,w__6239 ,w__5987);
  or g__8449(w__6460 ,w__6327 ,w__5983);
  or g__8450(w__6459 ,w__6242 ,w__5977);
  not g__8451(w__6346 ,w__5980);
  not g__8452(w__6345 ,w__5985);
  not g__8453(w__6343 ,w__5979);
  not g__8454(w__6342 ,w__5981);
  nor g__8455(w__6340 ,w__6028 ,w__6226);
  nor g__8456(w__6339 ,w__6164 ,w__6189);
  nor g__8457(w__6338 ,w__6026 ,w__6195);
  nor g__8458(w__6337 ,w__6024 ,w__6228);
  nor g__8459(w__6336 ,w__6022 ,w__6190);
  nor g__8460(w__6335 ,w__6030 ,w__6215);
  nor g__8461(w__6334 ,w__6032 ,w__6220);
  or g__8462(w__6333 ,w__6211 ,w__6200);
  xnor g__8463(w__6331 ,in13[13] ,in13[12]);
  xnor g__8464(w__6330 ,in12[0] ,in13[3]);
  nor g__8465(w__6329 ,w__13435 ,w__6034);
  xnor g__8466(w__6328 ,in12[0] ,in13[9]);
  xnor g__8467(w__6327 ,in13[9] ,in13[8]);
  xnor g__8468(w__6326 ,in13[7] ,in13[6]);
  xnor g__8469(w__6325 ,in12[0] ,in13[5]);
  xnor g__8470(w__6324 ,in13[3] ,in13[2]);
  or g__8471(w__6402 ,w__6132 ,w__6219);
  or g__8472(w__6401 ,w__6207 ,w__6216);
  or g__8473(w__6400 ,w__6133 ,w__6229);
  or g__8474(w__6399 ,w__6143 ,w__6224);
  or g__8475(w__6398 ,w__6135 ,w__6221);
  or g__8476(w__6397 ,w__6142 ,w__6217);
  xnor g__8477(w__6396 ,in12[4] ,in13[13]);
  or g__8478(w__6395 ,w__6140 ,w__6192);
  xnor g__8479(w__6394 ,in12[1] ,in13[13]);
  xnor g__8480(w__6393 ,in12[4] ,in13[11]);
  xnor g__8481(w__6392 ,in12[6] ,in13[7]);
  xnor g__8482(w__6391 ,in12[13] ,in13[5]);
  xnor g__8483(w__6390 ,in12[4] ,in13[3]);
  xnor g__8484(w__6389 ,in12[2] ,in13[3]);
  xnor g__8485(w__6388 ,in12[7] ,in13[7]);
  xnor g__8486(w__6387 ,in12[9] ,in13[11]);
  xnor g__8487(w__6386 ,in12[10] ,in13[5]);
  or g__8488(w__6385 ,w__6134 ,w__6225);
  or g__8489(w__6384 ,w__6141 ,w__6193);
  xnor g__8490(w__6383 ,in12[5] ,in13[5]);
  or g__8491(w__6382 ,w__6139 ,w__6197);
  xnor g__8492(w__6381 ,in12[6] ,in13[3]);
  xnor g__8493(w__6380 ,in12[3] ,in13[7]);
  xnor g__8494(w__6379 ,in12[15] ,in13[5]);
  or g__8495(w__6378 ,w__6137 ,w__6218);
  xnor g__8496(w__6377 ,in12[3] ,in13[9]);
  or g__8497(w__6376 ,w__6136 ,w__6222);
  xnor g__8498(w__6375 ,in12[10] ,in13[7]);
  xnor g__8499(w__6374 ,in12[11] ,in13[3]);
  xnor g__8500(w__6373 ,in12[8] ,in13[9]);
  or g__8501(w__6372 ,w__6138 ,w__6227);
  xnor g__8502(w__6371 ,in12[15] ,in13[7]);
  xnor g__8503(w__6370 ,in12[11] ,in13[7]);
  xnor g__8504(w__6369 ,in12[10] ,in13[13]);
  xnor g__8505(w__6368 ,in12[1] ,in13[5]);
  xnor g__8506(w__6367 ,in12[15] ,in13[15]);
  xnor g__8507(w__6366 ,in12[2] ,in13[11]);
  xnor g__8508(w__6365 ,in12[3] ,in13[11]);
  xnor g__8509(w__6364 ,in12[14] ,in13[9]);
  xnor g__8510(w__6363 ,in12[12] ,in13[9]);
  xnor g__8511(w__6362 ,in12[12] ,in13[7]);
  xnor g__8512(w__6361 ,in12[8] ,in13[11]);
  xnor g__8513(w__6360 ,in12[11] ,in13[5]);
  xnor g__8514(w__6359 ,in12[8] ,in13[13]);
  xnor g__8515(w__6358 ,in12[1] ,in13[11]);
  xnor g__8516(w__6357 ,in12[2] ,in13[9]);
  xnor g__8517(w__6356 ,in12[8] ,in13[5]);
  xnor g__8518(w__6355 ,in12[13] ,in13[11]);
  xnor g__8519(w__6354 ,in12[4] ,in13[9]);
  xnor g__8520(w__6353 ,in12[5] ,in13[9]);
  xnor g__8521(w__6352 ,in12[2] ,in13[13]);
  xnor g__8522(w__6351 ,in12[9] ,in13[9]);
  xnor g__8523(w__6350 ,in12[13] ,in13[9]);
  or g__8524(w__6349 ,w__6018 ,w__6201);
  xnor g__8525(w__6348 ,in12[15] ,in13[13]);
  xnor g__8526(w__6347 ,in12[7] ,in13[13]);
  xnor g__8527(w__6344 ,w__6032 ,in13[6]);
  xnor g__8528(w__6341 ,w__6022 ,in13[14]);
  not g__8529(w__6259 ,w__5978);
  not g__8530(w__6258 ,w__5977);
  not g__8531(w__6256 ,w__5988);
  not g__8532(w__6254 ,w__5974);
  not g__8533(w__6253 ,w__5987);
  not g__8534(w__6252 ,w__5973);
  not g__8535(w__6251 ,w__5975);
  not g__8536(w__6249 ,w__5984);
  not g__8537(w__6248 ,w__5983);
  not g__8538(w__6246 ,w__5982);
  not g__8539(w__6245 ,w__5976);
  xnor g__8540(w__6243 ,in13[15] ,in13[14]);
  xnor g__8541(w__6242 ,in13[11] ,in13[10]);
  xnor g__8542(w__6241 ,in12[0] ,in13[11]);
  xnor g__8543(w__6240 ,in12[0] ,in13[13]);
  xnor g__8544(w__6239 ,in13[5] ,in13[4]);
  xnor g__8545(w__6237 ,in12[0] ,in13[7]);
  xnor g__8546(w__6323 ,in12[7] ,in13[3]);
  xnor g__8547(w__6322 ,in12[11] ,in13[9]);
  xnor g__8548(w__6321 ,in12[15] ,in13[3]);
  xnor g__8549(w__6320 ,in12[4] ,in13[7]);
  xnor g__8550(w__6319 ,in12[12] ,in13[5]);
  xnor g__8551(w__6318 ,in12[13] ,in13[7]);
  xnor g__8552(w__6317 ,in12[14] ,in13[13]);
  xnor g__8553(w__6316 ,in12[5] ,in13[11]);
  xnor g__8554(w__6315 ,in12[9] ,in13[3]);
  xnor g__8555(w__6314 ,in12[15] ,in13[11]);
  xnor g__8556(w__6313 ,in12[5] ,in13[7]);
  xnor g__8557(w__6312 ,in12[14] ,in13[11]);
  xnor g__8558(w__6311 ,in12[1] ,in13[9]);
  xnor g__8559(w__6310 ,in12[6] ,in13[5]);
  xnor g__8560(w__6309 ,in12[11] ,in13[11]);
  xnor g__8561(w__6308 ,in12[14] ,in13[3]);
  xnor g__8562(w__6307 ,in12[3] ,in13[5]);
  xnor g__8563(w__6306 ,in12[11] ,in13[13]);
  xnor g__8564(w__6305 ,in12[12] ,in13[11]);
  xnor g__8565(w__6304 ,in12[3] ,in13[3]);
  xnor g__8566(w__6303 ,in12[3] ,in13[13]);
  xnor g__8567(w__6302 ,in12[14] ,in13[7]);
  xnor g__8568(w__6301 ,in12[4] ,in13[5]);
  xnor g__8569(w__6300 ,in12[13] ,in13[13]);
  xnor g__8570(w__6299 ,in12[1] ,in13[3]);
  xnor g__8571(w__6298 ,in12[9] ,in13[5]);
  xnor g__8572(w__6297 ,in12[7] ,in13[9]);
  xnor g__8573(w__6296 ,in12[12] ,in13[13]);
  xnor g__8574(w__6295 ,in12[8] ,in13[3]);
  xnor g__8575(w__6294 ,in12[5] ,in13[13]);
  xnor g__8576(w__6293 ,in12[5] ,in13[3]);
  xnor g__8577(w__6292 ,in12[8] ,in13[7]);
  xnor g__8578(w__6291 ,in12[13] ,in13[3]);
  xnor g__8579(w__6290 ,in12[1] ,in13[7]);
  xnor g__8580(w__6289 ,in12[6] ,in13[9]);
  xnor g__8581(w__6288 ,in12[10] ,in13[11]);
  xnor g__8582(w__6287 ,in12[10] ,in13[9]);
  xnor g__8583(w__6286 ,in12[14] ,in13[5]);
  xnor g__8584(w__6285 ,in12[9] ,in13[13]);
  xnor g__8585(w__6284 ,in12[9] ,in13[7]);
  xnor g__8586(w__6283 ,in12[2] ,in13[5]);
  xnor g__8587(w__6282 ,in12[6] ,in13[13]);
  xnor g__8588(w__6281 ,in12[12] ,in13[3]);
  xnor g__8589(w__6280 ,in12[6] ,in13[11]);
  xnor g__8590(w__6279 ,in12[15] ,in13[9]);
  xnor g__8591(w__6278 ,in12[2] ,in13[7]);
  xnor g__8592(w__6277 ,in12[10] ,in13[3]);
  xnor g__8593(w__6276 ,in12[4] ,in13[1]);
  xnor g__8594(w__6275 ,in12[2] ,in13[1]);
  xnor g__8595(w__6274 ,in12[9] ,in13[1]);
  xnor g__8596(w__6273 ,in12[3] ,in13[1]);
  xnor g__8597(w__6272 ,in12[5] ,in13[1]);
  xnor g__8598(w__6271 ,in12[8] ,in13[1]);
  xnor g__8599(w__6270 ,in12[7] ,in13[1]);
  xnor g__8600(w__6269 ,in12[11] ,in13[1]);
  xnor g__8601(w__6268 ,in12[14] ,in13[1]);
  xnor g__8602(w__6267 ,in12[12] ,in13[1]);
  xnor g__8603(w__6266 ,in12[7] ,in13[5]);
  xnor g__8604(w__6265 ,in12[10] ,in13[1]);
  xnor g__8605(w__6264 ,in12[1] ,in13[1]);
  xnor g__8606(w__6263 ,in12[6] ,in13[1]);
  xnor g__8607(w__6262 ,in12[13] ,in13[1]);
  xnor g__8608(w__6261 ,in12[15] ,in13[1]);
  xnor g__8609(w__6260 ,in12[7] ,in13[11]);
  xnor g__8610(w__6257 ,w__6030 ,in13[10]);
  xnor g__8611(w__6255 ,w__6028 ,in13[4]);
  xnor g__8612(w__6250 ,w__6034 ,in13[2]);
  xnor g__8613(w__6247 ,w__6026 ,in13[8]);
  xnor g__8614(w__6244 ,w__6024 ,in13[12]);
  nor g__8615(w__6229 ,in12[2] ,in13[15]);
  nor g__8616(w__6228 ,in12[0] ,in13[12]);
  nor g__8617(w__6227 ,in12[4] ,in13[15]);
  nor g__8618(w__6226 ,in12[0] ,in13[4]);
  nor g__8619(w__6225 ,in12[5] ,in13[15]);
  nor g__8620(w__6224 ,in12[9] ,in13[15]);
  and g__8621(w__6223 ,in12[0] ,in13[6]);
  nor g__8622(w__6222 ,in12[13] ,in13[15]);
  nor g__8623(w__6221 ,in12[8] ,in13[15]);
  nor g__8624(w__6220 ,in12[0] ,in13[6]);
  nor g__8625(w__6219 ,in12[1] ,in13[15]);
  nor g__8626(w__6218 ,in12[3] ,in13[15]);
  nor g__8627(w__6217 ,in12[7] ,in13[15]);
  nor g__8628(w__6216 ,in12[6] ,in13[15]);
  nor g__8629(w__6215 ,in12[0] ,in13[10]);
  or g__8630(w__6214 ,w__6184 ,w__5847);
  or g__8631(w__6236 ,w__6186 ,w__5871);
  or g__8632(w__6235 ,w__6187 ,w__5949);
  or g__8633(w__6234 ,w__6169 ,w__5919);
  or g__8634(w__6233 ,w__6173 ,w__5848);
  or g__8635(w__6232 ,w__6182 ,w__5872);
  or g__8636(w__6231 ,w__6181 ,w__5833);
  or g__8637(w__6230 ,w__6172 ,w__5919);
  not g__8638(w__6210 ,w__6211);
  not g__8639(w__6207 ,w__6208);
  not g__8640(w__6202 ,w__6203);
  nor g__8641(w__6201 ,in12[14] ,in13[15]);
  nor g__8642(w__6200 ,in12[0] ,in13[15]);
  and g__8643(w__6199 ,in12[0] ,in13[14]);
  and g__8644(w__6198 ,in12[0] ,in13[2]);
  nor g__8645(w__6197 ,in12[12] ,in13[15]);
  and g__8646(w__6196 ,in12[0] ,in13[10]);
  nor g__8647(w__6195 ,in12[0] ,in13[8]);
  and g__8648(w__6194 ,in12[0] ,in13[12]);
  nor g__8649(w__6193 ,in12[10] ,in13[15]);
  nor g__8650(w__6192 ,in12[11] ,in13[15]);
  and g__8651(w__6191 ,in12[0] ,in13[8]);
  nor g__8652(w__6190 ,in12[0] ,in13[14]);
  nor g__8653(w__6189 ,in12[0] ,in13[2]);
  and g__8654(w__6188 ,in12[0] ,in13[4]);
  and g__8655(w__13435 ,in12[0] ,in13[0]);
  and g__8656(w__6213 ,in13[1] ,in13[0]);
  or g__8657(w__6212 ,w__6170 ,w__5847);
  and g__8658(w__6211 ,in12[0] ,in13[15]);
  or g__8659(w__6209 ,w__6168 ,w__5871);
  or g__8660(w__6208 ,w__6183 ,w__5949);
  or g__8661(w__6206 ,w__6174 ,w__5872);
  or g__8662(w__6205 ,w__6167 ,w__5848);
  or g__8663(w__6204 ,w__6185 ,w__5833);
  or g__8664(w__6203 ,w__6171 ,w__5920);
  not g__8665(w__6187 ,in12[7]);
  not g__8666(w__6186 ,in12[9]);
  not g__8667(w__6185 ,in12[1]);
  not g__8668(w__6184 ,in12[15]);
  not g__8669(w__6183 ,in12[6]);
  not g__8670(w__6182 ,in12[12]);
  not g__8671(w__6181 ,in12[4]);
  not g__8672(w__6180 ,in12[0]);
  not g__8673(w__6179 ,in13[3]);
  not g__8674(w__6178 ,in13[7]);
  not g__8675(w__6177 ,in13[5]);
  not g__8676(w__6176 ,in13[9]);
  not g__8677(w__6175 ,in13[11]);
  not g__8678(w__6174 ,in12[5]);
  not g__8679(w__6173 ,in12[11]);
  not g__8680(w__6172 ,in12[3]);
  not g__8681(w__6171 ,in12[14]);
  not g__8682(w__6170 ,in12[13]);
  not g__8683(w__6169 ,in12[10]);
  not g__8684(w__6168 ,in12[8]);
  not g__8685(w__6167 ,in12[2]);
  not g__8686(w__6166 ,in13[0]);
  not g__8687(w__6165 ,in13[15]);
  not g__8688(w__6164 ,in13[1]);
  not g__8689(w__6163 ,in13[13]);
  not g__8690(w__5817 ,w__6131);
  not g__8691(w__6131 ,w__6180);
  not g__8692(w__6130 ,w__6128);
  not g__8693(w__6129 ,w__6128);
  not g__8694(w__6128 ,w__6150);
  not g__8695(w__6127 ,w__6125);
  not g__8696(w__6126 ,w__6125);
  not g__8697(w__6125 ,w__6256);
  not g__8698(w__6124 ,w__6122);
  not g__8699(w__6123 ,w__6122);
  not g__8700(w__6122 ,w__6253);
  not g__8701(w__6121 ,w__6119);
  not g__8702(w__6120 ,w__6119);
  not g__8703(w__6119 ,w__6251);
  not g__8704(w__6118 ,w__6116);
  not g__8705(w__6117 ,w__6116);
  not g__8706(w__6116 ,w__6252);
  not g__8707(w__6115 ,w__6113);
  not g__8708(w__6114 ,w__6113);
  not g__8709(w__6113 ,w__6149);
  not g__8710(w__6112 ,w__6110);
  not g__8711(w__6111 ,w__6110);
  not g__8712(w__6110 ,w__6148);
  not g__8713(w__6109 ,w__6107);
  not g__8714(w__6108 ,w__6107);
  not g__8715(w__6107 ,w__6248);
  not g__8716(w__6106 ,w__6104);
  not g__8717(w__6105 ,w__6104);
  not g__8718(w__6104 ,w__6249);
  not g__8719(w__6103 ,w__6101);
  not g__8720(w__6102 ,w__6101);
  not g__8721(w__6101 ,w__6147);
  not g__8722(w__6100 ,w__6098);
  not g__8723(w__6099 ,w__6098);
  not g__8724(w__6098 ,w__6146);
  not g__8725(w__6097 ,w__6095);
  not g__8726(w__6096 ,w__6095);
  not g__8727(w__6095 ,w__6246);
  not g__8728(w__6094 ,w__6092);
  not g__8729(w__6093 ,w__6092);
  not g__8730(w__6092 ,w__6245);
  not g__8731(w__6091 ,w__6089);
  not g__8732(w__6090 ,w__6089);
  not g__8733(w__6089 ,w__6145);
  not g__8734(w__6088 ,w__6086);
  not g__8735(w__6087 ,w__6086);
  not g__8736(w__6086 ,w__6144);
  not g__8737(w__6085 ,w__6083);
  not g__8738(w__6084 ,w__6083);
  not g__8739(w__6083 ,w__6346);
  not g__8740(w__6082 ,w__6080);
  not g__8741(w__6081 ,w__6080);
  not g__8742(w__6080 ,w__6345);
  not g__8743(w__6079 ,w__6077);
  not g__8744(w__6078 ,w__6077);
  not g__8745(w__6077 ,w__6156);
  not g__8746(w__6076 ,w__6074);
  not g__8747(w__6075 ,w__6074);
  not g__8748(w__6074 ,w__6155);
  not g__8749(w__6073 ,w__6071);
  not g__8750(w__6072 ,w__6071);
  not g__8751(w__6071 ,w__6343);
  not g__8752(w__6070 ,w__6068);
  not g__8753(w__6069 ,w__6068);
  not g__8754(w__6068 ,w__6342);
  not g__8755(w__6067 ,w__6065);
  not g__8756(w__6066 ,w__6065);
  not g__8757(w__6065 ,w__6154);
  not g__8758(w__6064 ,w__6062);
  not g__8759(w__6063 ,w__6062);
  not g__8760(w__6062 ,w__6153);
  not g__8761(w__6061 ,w__6059);
  not g__8762(w__6060 ,w__6059);
  not g__8763(w__6059 ,w__6259);
  not g__8764(w__6058 ,w__6056);
  not g__8765(w__6057 ,w__6056);
  not g__8766(w__6056 ,w__6258);
  not g__8767(w__6055 ,w__6053);
  not g__8768(w__6054 ,w__6053);
  not g__8769(w__6053 ,w__6152);
  not g__8770(w__6052 ,w__6050);
  not g__8771(w__6051 ,w__6050);
  not g__8772(w__6050 ,w__6151);
  not g__8773(w__6049 ,w__6139);
  not g__8774(w__6139 ,w__6232);
  not g__8775(w__6048 ,w__6136);
  not g__8776(w__6136 ,w__6212);
  not g__8777(w__6047 ,w__6143);
  not g__8778(w__6143 ,w__6236);
  not g__8779(w__6046 ,w__6140);
  not g__8780(w__6140 ,w__6233);
  not g__8781(w__6045 ,w__6141);
  not g__8782(w__6141 ,w__6234);
  not g__8783(w__6044 ,w__6137);
  not g__8784(w__6137 ,w__6230);
  not g__8785(w__6043 ,w__6135);
  not g__8786(w__6135 ,w__6209);
  not g__8787(w__6042 ,w__6133);
  not g__8788(w__6133 ,w__6205);
  not g__8789(w__6041 ,w__6134);
  not g__8790(w__6134 ,w__6206);
  not g__8791(w__6040 ,w__6132);
  not g__8792(w__6132 ,w__6204);
  not g__8793(w__6039 ,w__6138);
  not g__8794(w__6138 ,w__6231);
  not g__8795(w__6038 ,w__6142);
  not g__8796(w__6142 ,w__6235);
  not g__8797(w__6037 ,w__6036);
  not g__8798(w__6036 ,w__6791);
  not g__8799(w__6035 ,w__6157);
  not g__8800(w__6157 ,w__6794);
  not g__8801(w__6034 ,w__6033);
  not g__8802(w__6033 ,w__6164);
  not g__8803(w__6032 ,w__6031);
  not g__8804(w__6031 ,w__6177);
  not g__8805(w__6030 ,w__6029);
  not g__8806(w__6029 ,w__6176);
  not g__8807(w__6028 ,w__6027);
  not g__8808(w__6027 ,w__6179);
  not g__8809(w__6026 ,w__6025);
  not g__8810(w__6025 ,w__6178);
  not g__8811(w__6024 ,w__6023);
  not g__8812(w__6023 ,w__6175);
  not g__8813(w__6022 ,w__6021);
  not g__8814(w__6021 ,w__6163);
  not g__8815(w__6020 ,w__6019);
  not g__8816(w__6019 ,w__6254);
  buf g__8817(w__13433 ,w__6403);
  buf g__8818(w__13434 ,w__6329);
  not g__8819(w__6018 ,w__6017);
  not g__8820(w__6017 ,w__6202);
  not g__8821(w__6016 ,w__6015);
  not g__8822(w__6015 ,w__6792);
  not g__8823(w__6014 ,w__6159);
  not g__8824(w__6159 ,w__7148);
  not g__8825(w__6013 ,w__6160);
  not g__8826(w__6160 ,w__7164);
  not g__8827(w__6012 ,w__6161);
  not g__8828(w__6161 ,w__7404);
  not g__8829(w__6011 ,w__6158);
  not g__8830(w__6158 ,w__7147);
  not g__8831(w__6010 ,w__6162);
  not g__8832(w__6162 ,w__7405);
  not g__8833(w__6009 ,w__6008);
  not g__8834(w__6008 ,w__6557);
  not g__8835(w__6007 ,w__6006);
  not g__8836(w__6006 ,w__6464);
  not g__8837(w__6005 ,w__6004);
  not g__8838(w__6004 ,w__6463);
  not g__8839(w__6003 ,w__6002);
  not g__8840(w__6002 ,w__6460);
  not g__8841(w__6001 ,w__6000);
  not g__8842(w__6000 ,w__6459);
  not g__8843(w__5999 ,w__5998);
  not g__8844(w__5998 ,w__6462);
  not g__8845(w__5997 ,w__5996);
  not g__8846(w__5996 ,w__6461);
  not g__8847(w__5995 ,w__5994);
  not g__8848(w__5994 ,w__6165);
  not g__8849(w__5993 ,w__5992);
  not g__8850(w__5992 ,w__6558);
  not g__8851(w__5991 ,w__5989);
  not g__8852(w__5990 ,w__5989);
  not g__8853(w__5989 ,w__6166);
  not g__8854(w__5988 ,w__5986);
  not g__8855(w__5987 ,w__5986);
  not g__8856(w__5986 ,w__6255);
  not g__8857(w__5985 ,w__6155);
  not g__8858(w__6155 ,w__6344);
  not g__8859(w__5984 ,w__6147);
  not g__8860(w__6147 ,w__6247);
  not g__8861(w__5983 ,w__6146);
  not g__8862(w__6146 ,w__6247);
  not g__8863(w__5982 ,w__6145);
  not g__8864(w__6145 ,w__6244);
  not g__8865(w__5981 ,w__6153);
  not g__8866(w__6153 ,w__6341);
  not g__8867(w__5980 ,w__6156);
  not g__8868(w__6156 ,w__6344);
  not g__8869(w__5979 ,w__6154);
  not g__8870(w__6154 ,w__6341);
  not g__8871(w__5978 ,w__6152);
  not g__8872(w__6152 ,w__6257);
  not g__8873(w__5977 ,w__6151);
  not g__8874(w__6151 ,w__6257);
  not g__8875(w__5976 ,w__6144);
  not g__8876(w__6144 ,w__6244);
  not g__8877(w__5975 ,w__6148);
  not g__8878(w__6148 ,w__6250);
  not g__8879(w__5974 ,w__6150);
  not g__8880(w__6150 ,w__6255);
  not g__8881(w__5973 ,w__6149);
  not g__8882(w__6149 ,w__6250);
  not g__8883(w__5972 ,w__5971);
  not g__8884(w__5971 ,w__6711);
  not g__8885(w__5970 ,w__5969);
  not g__8886(w__5969 ,w__6788);
  not g__8887(w__5968 ,w__5967);
  not g__8888(w__5967 ,w__6713);
  not g__8889(w__5966 ,w__5965);
  not g__8890(w__5965 ,w__6709);
  not g__8891(w__5816 ,w__5825);
  not g__8892(w__5964 ,w__5825);
  not g__8893(w__5825 ,w__5817);
  not g__8894(w__5963 ,w__6131);
  not g__8895(w__5962 ,w__5960);
  not g__8896(w__5961 ,w__5960);
  not g__8897(w__5960 ,w__6557);
  not g__8898(w__5959 ,w__5957);
  not g__8899(w__5958 ,w__5957);
  not g__8900(w__5957 ,w__6558);
  not g__8901(w__5956 ,w__5954);
  not g__8902(w__5955 ,w__5954);
  not g__8903(w__5954 ,w__6464);
  not g__8904(w__5953 ,w__5951);
  not g__8905(w__5952 ,w__5951);
  not g__8906(w__5951 ,w__6461);
  not g__8907(w__5950 ,w__5948);
  not g__8908(w__5949 ,w__5948);
  not g__8909(w__5948 ,w__6165);
  not g__8910(w__5947 ,w__5945);
  not g__8911(w__5946 ,w__5945);
  not g__8912(w__5945 ,w__6463);
  not g__8913(w__5944 ,w__5942);
  not g__8914(w__5943 ,w__5942);
  not g__8915(w__5942 ,w__6462);
  not g__8916(w__5941 ,w__5939);
  not g__8917(w__5940 ,w__5939);
  not g__8918(w__5939 ,w__6460);
  not g__8919(w__5938 ,w__5936);
  not g__8920(w__5937 ,w__5936);
  not g__8921(w__5936 ,w__6459);
  not g__8922(w__5935 ,w__5933);
  not g__8923(w__5934 ,w__5933);
  not g__8924(w__5933 ,w__6557);
  not g__8925(w__5932 ,w__5930);
  not g__8926(w__5931 ,w__5930);
  not g__8927(w__5930 ,w__6009);
  not g__8928(w__5929 ,w__5927);
  not g__8929(w__5928 ,w__5927);
  not g__8930(w__5927 ,w__5999);
  not g__8931(w__5926 ,w__5924);
  not g__8932(w__5925 ,w__5924);
  not g__8933(w__5924 ,w__6001);
  not g__8934(w__5923 ,w__5921);
  not g__8935(w__5922 ,w__5921);
  not g__8936(w__5921 ,w__5997);
  not g__8937(w__5920 ,w__5918);
  not g__8938(w__5919 ,w__5918);
  not g__8939(w__5918 ,w__5995);
  not g__8940(w__5917 ,w__5915);
  not g__8941(w__5916 ,w__5915);
  not g__8942(w__5915 ,w__5991);
  not g__8943(w__5914 ,w__5912);
  not g__8944(w__5913 ,w__5912);
  not g__8945(w__5912 ,w__6462);
  not g__8946(w__5911 ,w__5909);
  not g__8947(w__5910 ,w__5909);
  not g__8948(w__5909 ,w__6009);
  not g__8949(w__5908 ,w__5906);
  not g__8950(w__5907 ,w__5906);
  not g__8951(w__5906 ,w__6166);
  not g__8952(w__5905 ,w__5903);
  not g__8953(w__5904 ,w__5903);
  not g__8954(w__5903 ,w__6166);
  not g__8955(w__5902 ,w__5900);
  not g__8956(w__5901 ,w__5900);
  not g__8957(w__5900 ,w__6007);
  not g__8958(w__5899 ,w__5897);
  not g__8959(w__5898 ,w__5897);
  not g__8960(w__5897 ,w__6005);
  not g__8961(w__5896 ,w__5894);
  not g__8962(w__5895 ,w__5894);
  not g__8963(w__5894 ,w__6003);
  not g__8964(w__5893 ,w__5891);
  not g__8965(w__5892 ,w__5891);
  not g__8966(w__5891 ,w__6558);
  not g__8967(w__5890 ,w__5888);
  not g__8968(w__5889 ,w__5888);
  not g__8969(w__5888 ,w__5993);
  not g__8970(w__5887 ,w__5885);
  not g__8971(w__5886 ,w__5885);
  not g__8972(w__5885 ,w__5993);
  not g__8973(w__5884 ,w__5882);
  not g__8974(w__5883 ,w__5882);
  not g__8975(w__5882 ,w__6461);
  not g__8976(w__5881 ,w__5879);
  not g__8977(w__5880 ,w__5879);
  not g__8978(w__5879 ,w__6001);
  not g__8979(w__5878 ,w__5876);
  not g__8980(w__5877 ,w__5876);
  not g__8981(w__5876 ,w__6460);
  not g__8982(w__5875 ,w__5873);
  not g__8983(w__5874 ,w__5873);
  not g__8984(w__5873 ,w__5997);
  not g__8985(w__5872 ,w__5870);
  not g__8986(w__5871 ,w__5870);
  not g__8987(w__5870 ,w__5995);
  not g__8988(w__5869 ,w__5867);
  not g__8989(w__5868 ,w__5867);
  not g__8990(w__5867 ,w__6459);
  not g__8991(w__5866 ,w__5864);
  not g__8992(w__5865 ,w__5864);
  not g__8993(w__5864 ,w__6463);
  not g__8994(w__5863 ,w__5861);
  not g__8995(w__5862 ,w__5861);
  not g__8996(w__5861 ,w__5999);
  not g__8997(w__5860 ,w__5858);
  not g__8998(w__5859 ,w__5858);
  not g__8999(w__5858 ,w__6003);
  not g__9000(w__5857 ,w__5855);
  not g__9001(w__5856 ,w__5855);
  not g__9002(w__5855 ,w__6007);
  not g__9003(w__5854 ,w__5852);
  not g__9004(w__5853 ,w__5852);
  not g__9005(w__5852 ,w__6464);
  not g__9006(w__5851 ,w__5849);
  not g__9007(w__5850 ,w__5849);
  not g__9008(w__5849 ,w__6005);
  not g__9009(w__5848 ,w__5846);
  not g__9010(w__5847 ,w__5846);
  not g__9011(w__5846 ,w__6165);
  not g__9012(w__5845 ,w__5844);
  not g__9013(w__5844 ,w__5990);
  not g__9014(w__5843 ,w__5842);
  not g__9015(w__5842 ,w__5961);
  not g__9016(w__5841 ,w__5840);
  not g__9017(w__5840 ,w__5938);
  not g__9018(w__5839 ,w__5838);
  not g__9019(w__5838 ,w__5941);
  not g__9020(w__5837 ,w__5836);
  not g__9021(w__5836 ,w__5944);
  not g__9022(w__5835 ,w__5834);
  not g__9023(w__5834 ,w__5947);
  not g__9024(w__5833 ,w__5832);
  not g__9025(w__5832 ,w__5950);
  not g__9026(w__5831 ,w__5830);
  not g__9027(w__5830 ,w__5953);
  not g__9028(w__5829 ,w__5828);
  not g__9029(w__5828 ,w__5956);
  not g__9030(w__5827 ,w__5826);
  not g__9031(w__5826 ,w__5959);
  xor g__9032(w__5824 ,w__7406 ,w__7501);
  xor g__9033(w__13410 ,w__7382 ,w__7471);
  xor g__9034(w__5823 ,w__7364 ,w__7385);
  xor g__9035(w__5822 ,w__7023 ,w__7101);
  xor g__9036(w__5821 ,w__7017 ,w__5971);
  xor g__9037(w__5820 ,w__7127 ,w__5969);
  xor g__9038(w__5819 ,w__7006 ,w__5967);
  xor g__9039(w__5818 ,w__7114 ,w__5965);
  xnor g__9040(w__13351 ,w__9198 ,w__9233);
  xnor g__9041(w__13352 ,w__9201 ,w__7533);
  xnor g__9042(w__13354 ,w__9211 ,w__9225);
  xnor g__9043(w__13353 ,w__9207 ,w__9224);
  xnor g__9044(w__13350 ,w__9191 ,w__9226);
  or g__9045(w__13291 ,w__9196 ,w__9232);
  or g__9046(w__13290 ,w__9219 ,w__9231);
  or g__9047(w__13287 ,w__9214 ,w__9228);
  or g__9048(w__13286 ,w__9223 ,w__9230);
  or g__9049(w__13288 ,w__9212 ,w__9229);
  or g__9050(w__13289 ,w__9221 ,w__9227);
  xnor g__9051(w__13349 ,w__9177 ,w__9205);
  xnor g__9052(w__13355 ,w__9208 ,w__9204);
  xnor g__9053(w__13348 ,w__9179 ,w__9203);
  xnor g__9054(w__9233 ,w__9093 ,w__9209);
  and g__9055(w__9232 ,w__9185 ,w__9208);
  and g__9056(w__9231 ,w__9218 ,w__9211);
  or g__9057(w__13284 ,w__9193 ,w__9213);
  and g__9058(w__9230 ,w__9191 ,w__9215);
  nor g__9059(w__9229 ,w__9222 ,w__9210);
  or g__9060(w__13292 ,w__9175 ,w__9216);
  or g__9061(w__13285 ,w__9195 ,w__9217);
  and g__9062(w__9228 ,w__9206 ,w__9209);
  xnor g__9063(w__13356 ,w__9190 ,w__9182);
  xnor g__9064(w__13347 ,w__9178 ,w__9181);
  xnor g__9065(w__13357 ,w__9096 ,w__9183);
  nor g__9066(w__9227 ,w__9220 ,w__9207);
  xnor g__9067(w__9226 ,w__9187 ,w__9113);
  xnor g__9068(w__9225 ,w__9200 ,w__9114);
  xnor g__9069(w__9224 ,w__9188 ,w__9202);
  nor g__9070(w__9223 ,w__7721 ,w__9187);
  and g__9071(w__9222 ,w__9115 ,w__9201);
  nor g__9072(w__9221 ,w__9189 ,w__9202);
  and g__9073(w__9220 ,w__9189 ,w__9202);
  nor g__9074(w__9219 ,w__7719 ,w__9200);
  or g__9075(w__9218 ,w__7871 ,w__9199);
  nor g__9076(w__9217 ,w__9177 ,w__9194);
  and g__9077(w__9216 ,w__9174 ,w__9190);
  or g__9078(w__9215 ,w__7870 ,w__9186);
  nor g__9079(w__9214 ,w__9093 ,w__9198);
  nor g__9080(w__9213 ,w__9179 ,w__9192);
  nor g__9081(w__9212 ,w__9115 ,w__9201);
  or g__9082(w__9206 ,w__9092 ,w__9197);
  or g__9083(w__13346 ,w__9168 ,w__9184);
  xnor g__9084(w__13358 ,w__9122 ,w__7532);
  xnor g__9085(w__13360 ,w__9032 ,w__9152);
  xnor g__9086(w__13282 ,w__9100 ,w__9153);
  xnor g__9087(w__9205 ,w__9064 ,w__9159);
  xnor g__9088(w__9204 ,w__9162 ,w__9117);
  xnor g__9089(w__9203 ,w__9054 ,w__9163);
  xnor g__9090(w__9211 ,w__9099 ,w__9155);
  xnor g__9091(w__9210 ,w__9148 ,w__9151);
  xnor g__9092(w__9209 ,w__9125 ,w__9154);
  xnor g__9093(w__9208 ,w__9097 ,w__9149);
  xnor g__9094(w__9207 ,w__9121 ,w__9150);
  not g__9095(w__9199 ,w__9200);
  not g__9096(w__9197 ,w__9198);
  nor g__9097(w__9196 ,w__9117 ,w__9162);
  nor g__9098(w__9195 ,w__9064 ,w__9160);
  and g__9099(w__9194 ,w__9064 ,w__9160);
  or g__9100(w__13293 ,w__9139 ,w__9173);
  nor g__9101(w__9193 ,w__9054 ,w__9164);
  or g__9102(w__13294 ,w__9137 ,w__9172);
  or g__9103(w__13296 ,w__9133 ,w__9171);
  or g__9104(w__13345 ,w__9131 ,w__9169);
  and g__9105(w__9192 ,w__9054 ,w__9164);
  and g__9106(w__9202 ,w__9145 ,w__9165);
  and g__9107(w__9201 ,w__9128 ,w__9166);
  and g__9108(w__9200 ,w__9143 ,w__9176);
  and g__9109(w__9198 ,w__9134 ,w__9170);
  not g__9110(w__9189 ,w__9188);
  not g__9111(w__9186 ,w__9187);
  or g__9112(w__9185 ,w__9116 ,w__9161);
  nor g__9113(w__9184 ,w__9178 ,w__9167);
  or g__9114(w__13344 ,w__9127 ,w__9156);
  xnor g__9115(w__13359 ,w__9124 ,w__9105);
  or g__9116(w__13295 ,w__9085 ,w__9158);
  xnor g__9117(w__9183 ,w__9068 ,w__9120);
  xnor g__9118(w__9182 ,w__9112 ,w__9110);
  xnor g__9119(w__9181 ,w__9049 ,w__9118);
  xnor g__9120(w__9180 ,w__9123 ,w__9008);
  or g__9121(w__9191 ,w__9140 ,w__9157);
  xnor g__9122(w__9190 ,w__9051 ,w__9103);
  xnor g__9123(w__9188 ,w__8931 ,w__9102);
  xnor g__9124(w__9187 ,w__9098 ,w__9104);
  or g__9125(w__9176 ,w__9097 ,w__9141);
  nor g__9126(w__9175 ,w__9110 ,w__9112);
  or g__9127(w__9174 ,w__9109 ,w__9111);
  and g__9128(w__9173 ,w__9138 ,w__9120);
  nor g__9129(w__9172 ,w__9147 ,w__9122);
  and g__9130(w__9171 ,w__9032 ,w__9132);
  or g__9131(w__13297 ,w__9034 ,w__9130);
  or g__9132(w__9170 ,w__9148 ,w__9129);
  nor g__9133(w__9169 ,w__9106 ,w__9123);
  nor g__9134(w__9168 ,w__9049 ,w__9119);
  and g__9135(w__9167 ,w__9049 ,w__9119);
  or g__9136(w__9166 ,w__9121 ,w__9146);
  or g__9137(w__9165 ,w__9099 ,w__9144);
  and g__9138(w__9179 ,w__9026 ,w__9135);
  and g__9139(w__9178 ,w__8961 ,w__9108);
  and g__9140(w__9177 ,w__9089 ,w__9142);
  not g__9141(w__9164 ,w__9163);
  not g__9142(w__9161 ,w__9162);
  not g__9143(w__9160 ,w__9159);
  nor g__9144(w__9158 ,w__9086 ,w__9124);
  nor g__9145(w__9157 ,w__9136 ,w__9125);
  nor g__9146(w__9156 ,w__9100 ,w__9126);
  xnor g__9147(w__13361 ,w__9080 ,w__9060);
  xnor g__9148(w__13281 ,w__9029 ,w__9058);
  xnor g__9149(w__9155 ,w__8934 ,w__9066);
  xnor g__9150(w__9154 ,w__9053 ,w__9077);
  xnor g__9151(w__9153 ,w__8834 ,w__9075);
  xnor g__9152(w__9152 ,w__9072 ,w__8873);
  xnor g__9153(w__9151 ,w__9074 ,w__9048);
  xnor g__9154(w__9150 ,w__9063 ,w__8804);
  xnor g__9155(w__9149 ,w__9003 ,w__9070);
  xnor g__9156(w__9163 ,w__9079 ,w__9018);
  and g__9157(w__9162 ,w__9061 ,w__9107);
  xnor g__9158(w__9159 ,w__9101 ,w__9059);
  and g__9159(w__9147 ,w__9073 ,w__9094);
  and g__9160(w__9146 ,w__8804 ,w__9063);
  or g__9161(w__9145 ,w__8933 ,w__9066);
  nor g__9162(w__9144 ,w__8934 ,w__9065);
  or g__9163(w__9143 ,w__9003 ,w__9069);
  or g__9164(w__9142 ,w__9087 ,w__9098);
  nor g__9165(w__9141 ,w__9002 ,w__9070);
  nor g__9166(w__9140 ,w__9053 ,w__9078);
  nor g__9167(w__9139 ,w__9096 ,w__9068);
  or g__9168(w__9138 ,w__9095 ,w__9067);
  nor g__9169(w__9137 ,w__9073 ,w__9094);
  and g__9170(w__9136 ,w__9053 ,w__9078);
  or g__9171(w__9135 ,w__9036 ,w__9101);
  or g__9172(w__9134 ,w__9048 ,w__9074);
  nor g__9173(w__9133 ,w__7722 ,w__9072);
  or g__9174(w__9132 ,w__7869 ,w__9071);
  nor g__9175(w__9131 ,w__9008 ,w__9091);
  and g__9176(w__9130 ,w__9035 ,w__9080);
  and g__9177(w__9129 ,w__9048 ,w__9074);
  or g__9178(w__13342 ,w__9040 ,w__9082);
  or g__9179(w__13343 ,w__9043 ,w__9081);
  or g__9180(w__9128 ,w__8804 ,w__9063);
  nor g__9181(w__9127 ,w__8834 ,w__9076);
  and g__9182(w__9126 ,w__8834 ,w__9076);
  and g__9183(w__9148 ,w__8951 ,w__9090);
  not g__9184(w__9119 ,w__9118);
  not g__9185(w__9117 ,w__9116);
  not g__9186(w__9111 ,w__9112);
  not g__9187(w__9109 ,w__9110);
  xnor g__9188(w__13279 ,w__8802 ,w__9024);
  xnor g__9189(w__13362 ,w__9030 ,w__9017);
  or g__9190(w__9108 ,w__8995 ,w__9079);
  or g__9191(w__9107 ,w__9031 ,w__9062);
  and g__9192(w__9106 ,w__9008 ,w__9091);
  or g__9193(w__13298 ,w__8954 ,w__9088);
  xnor g__9194(w__13363 ,w__8926 ,w__9015);
  xnor g__9195(w__13280 ,w__9007 ,w__9021);
  xnor g__9196(w__9105 ,w__8965 ,w__9055);
  xnor g__9197(w__9104 ,w__9052 ,w__8964);
  xnor g__9198(w__9103 ,w__8839 ,w__9031);
  xnor g__9199(w__9102 ,w__9057 ,w__8867);
  xnor g__9200(w__9125 ,w__8832 ,w__9013);
  xnor g__9201(w__9124 ,w__8936 ,w__9014);
  xnor g__9202(w__9123 ,w__7530 ,w__9016);
  xnor g__9203(w__9122 ,w__8969 ,w__9023);
  and g__9204(w__9121 ,w__8960 ,w__9083);
  xnor g__9205(w__9120 ,w__9056 ,w__9022);
  xnor g__9206(w__9118 ,w__8970 ,w__9020);
  xnor g__9207(w__9116 ,w__8870 ,w__9019);
  xnor g__9208(w__9115 ,w__8796 ,w__9012);
  xnor g__9209(w__9114 ,w__9028 ,w__9009);
  xnor g__9210(w__9113 ,w__8871 ,w__9010);
  xnor g__9211(w__9112 ,w__8865 ,w__9011);
  and g__9212(w__9110 ,w__8989 ,w__9084);
  not g__9213(w__9095 ,w__9096);
  not g__9214(w__9092 ,w__9093);
  or g__9215(w__9090 ,w__8950 ,w__9057);
  or g__9216(w__9089 ,w__8964 ,w__9052);
  nor g__9217(w__9088 ,w__8953 ,w__9030);
  and g__9218(w__9087 ,w__8964 ,w__9052);
  and g__9219(w__9086 ,w__8966 ,w__9055);
  nor g__9220(w__9085 ,w__8966 ,w__9055);
  or g__9221(w__9084 ,w__9056 ,w__8986);
  or g__9222(w__9083 ,w__8958 ,w__9028);
  and g__9223(w__9082 ,w__8935 ,w__9042);
  and g__9224(w__9081 ,w__9029 ,w__9038);
  and g__9225(w__9101 ,w__9001 ,w__9045);
  and g__9226(w__9100 ,w__8974 ,w__9025);
  and g__9227(w__9099 ,w__9000 ,w__9046);
  and g__9228(w__9098 ,w__8956 ,w__9039);
  and g__9229(w__9097 ,w__8994 ,w__9044);
  and g__9230(w__9096 ,w__8985 ,w__9037);
  and g__9231(w__9094 ,w__8981 ,w__9047);
  and g__9232(w__9093 ,w__8979 ,w__9033);
  and g__9233(w__9091 ,w__8999 ,w__9041);
  not g__9234(w__9078 ,w__9077);
  not g__9235(w__9076 ,w__9075);
  not g__9236(w__9071 ,w__9072);
  not g__9237(w__9069 ,w__9070);
  not g__9238(w__9067 ,w__9068);
  not g__9239(w__9065 ,w__9066);
  xnor g__9240(w__13364 ,w__8882 ,w__7531);
  or g__9241(w__13299 ,w__8972 ,w__9027);
  nor g__9242(w__9062 ,w__8839 ,w__9050);
  or g__9243(w__9061 ,w__8838 ,w__9051);
  xnor g__9244(w__9060 ,w__9005 ,w__8856);
  xnor g__9245(w__9059 ,w__7528 ,w__8963);
  xnor g__9246(w__9058 ,w__8968 ,w__8857);
  xnor g__9247(w__9080 ,w__8889 ,w__8943);
  xnor g__9248(w__9079 ,w__8884 ,w__8940);
  xnor g__9249(w__9077 ,w__8841 ,w__7527);
  xnor g__9250(w__9075 ,w__8885 ,w__7529);
  xnor g__9251(w__9074 ,w__8878 ,w__8939);
  xnor g__9252(w__9073 ,w__8843 ,w__8937);
  xnor g__9253(w__9072 ,w__8883 ,w__8938);
  xnor g__9254(w__9070 ,w__8817 ,w__8945);
  xnor g__9255(w__9068 ,w__8890 ,w__8946);
  xnor g__9256(w__9066 ,w__8794 ,w__8942);
  xnor g__9257(w__9064 ,w__8875 ,w__8944);
  xnor g__9258(w__9063 ,w__8876 ,w__8941);
  not g__9259(w__9050 ,w__9051);
  or g__9260(w__9047 ,w__8936 ,w__8980);
  or g__9261(w__9046 ,w__8881 ,w__8998);
  or g__9262(w__9045 ,w__8880 ,w__8997);
  or g__9263(w__9044 ,w__8879 ,w__8992);
  nor g__9264(w__9043 ,w__7723 ,w__8968);
  or g__9265(w__9042 ,w__8828 ,w__9006);
  or g__9266(w__9041 ,w__8991 ,w__8971);
  nor g__9267(w__9040 ,w__8829 ,w__9007);
  or g__9268(w__13341 ,w__8891 ,w__8959);
  or g__9269(w__9039 ,w__8886 ,w__8955);
  or g__9270(w__9038 ,w__7868 ,w__8967);
  or g__9271(w__9037 ,w__8969 ,w__8983);
  or g__9272(w__13300 ,w__8899 ,w__8984);
  nor g__9273(w__9036 ,w__7528 ,w__8962);
  or g__9274(w__9035 ,w__7867 ,w__9004);
  nor g__9275(w__9034 ,w__7720 ,w__9005);
  or g__9276(w__9033 ,w__8877 ,w__8977);
  and g__9277(w__9057 ,w__8900 ,w__8987);
  and g__9278(w__9056 ,w__8918 ,w__8988);
  and g__9279(w__9055 ,w__8910 ,w__8978);
  and g__9280(w__9054 ,w__8914 ,w__8973);
  and g__9281(w__9053 ,w__8915 ,w__8982);
  and g__9282(w__9052 ,w__8923 ,w__8993);
  and g__9283(w__9051 ,w__8922 ,w__8990);
  and g__9284(w__9049 ,w__8907 ,w__8947);
  and g__9285(w__9048 ,w__8906 ,w__8975);
  or g__9286(w__13301 ,w__8747 ,w__8948);
  nor g__9287(w__9027 ,w__8888 ,w__8976);
  or g__9288(w__9026 ,w__8932 ,w__8963);
  xnor g__9289(w__13365 ,w__8887 ,w__8790);
  or g__9290(w__9025 ,w__7530 ,w__8996);
  xnor g__9291(w__9024 ,w__8874 ,w__8502);
  xnor g__9292(w__9023 ,w__8859 ,w__8860);
  xnor g__9293(w__9022 ,w__8862 ,w__8929);
  xnor g__9294(w__9021 ,w__8829 ,w__8935);
  xnor g__9295(w__9020 ,w__8863 ,w__8837);
  xnor g__9296(w__9019 ,w__8849 ,w__8881);
  xnor g__9297(w__9018 ,w__8809 ,w__8853);
  xnor g__9298(w__9017 ,w__8800 ,w__8855);
  xnor g__9299(w__9016 ,w__8851 ,w__8795);
  xnor g__9300(w__9015 ,w__8888 ,w__8812);
  xnor g__9301(w__9014 ,w__8858 ,w__8854);
  xnor g__9302(w__9013 ,w__8872 ,w__8886);
  xnor g__9303(w__9012 ,w__8868 ,w__8877);
  xnor g__9304(w__9011 ,w__8879 ,w__8825);
  xnor g__9305(w__9010 ,w__8880 ,w__8831);
  xnor g__9306(w__9009 ,w__8864 ,w__8850);
  or g__9307(w__9032 ,w__8905 ,w__8949);
  xnor g__9308(w__9031 ,w__8840 ,w__8847);
  xnor g__9309(w__9030 ,w__8815 ,w__8846);
  or g__9310(w__9029 ,w__8921 ,w__8952);
  and g__9311(w__9028 ,w__8893 ,w__8957);
  not g__9312(w__9006 ,w__9007);
  not g__9313(w__9004 ,w__9005);
  not g__9314(w__9002 ,w__9003);
  or g__9315(w__13340 ,w__8618 ,w__8896);
  or g__9316(w__9001 ,w__8831 ,w__8871);
  or g__9317(w__9000 ,w__8848 ,w__8870);
  or g__9318(w__8999 ,w__8837 ,w__8863);
  nor g__9319(w__8998 ,w__8849 ,w__8869);
  and g__9320(w__8997 ,w__8831 ,w__8871);
  and g__9321(w__8996 ,w__8795 ,w__8851);
  nor g__9322(w__8995 ,w__8809 ,w__8852);
  or g__9323(w__8994 ,w__8825 ,w__8865);
  or g__9324(w__8993 ,w__8841 ,w__8920);
  and g__9325(w__8992 ,w__8825 ,w__8865);
  and g__9326(w__8991 ,w__8837 ,w__8863);
  or g__9327(w__8990 ,w__8890 ,w__8919);
  or g__9328(w__8989 ,w__8862 ,w__8928);
  or g__9329(w__8988 ,w__8843 ,w__8917);
  or g__9330(w__8987 ,w__8813 ,w__8897);
  nor g__9331(w__8986 ,w__8861 ,w__8929);
  or g__9332(w__8985 ,w__8860 ,w__8859);
  nor g__9333(w__8984 ,w__8898 ,w__8882);
  and g__9334(w__8983 ,w__8860 ,w__8859);
  or g__9335(w__8982 ,w__8913 ,w__8878);
  or g__9336(w__8981 ,w__8854 ,w__8858);
  and g__9337(w__8980 ,w__8854 ,w__8858);
  or g__9338(w__8979 ,w__8796 ,w__8868);
  or g__9339(w__8978 ,w__8909 ,w__8883);
  and g__9340(w__8977 ,w__8796 ,w__8868);
  and g__9341(w__8976 ,w__8812 ,w__8927);
  or g__9342(w__8975 ,w__8902 ,w__8876);
  or g__9343(w__8974 ,w__8795 ,w__8851);
  or g__9344(w__8973 ,w__8901 ,w__8875);
  nor g__9345(w__8972 ,w__8812 ,w__8927);
  and g__9346(w__9008 ,w__8593 ,w__8916);
  and g__9347(w__9007 ,w__8634 ,w__8908);
  and g__9348(w__9005 ,w__8791 ,w__8903);
  and g__9349(w__9003 ,w__8818 ,w__8924);
  not g__9350(w__8971 ,w__8970);
  not g__9351(w__8967 ,w__8968);
  not g__9352(w__8966 ,w__8965);
  not g__9353(w__8962 ,w__8963);
  xnor g__9354(w__13278 ,w__8845 ,w__8739);
  or g__9355(w__8961 ,w__8808 ,w__8853);
  or g__9356(w__8960 ,w__8850 ,w__8864);
  nor g__9357(w__8959 ,w__8911 ,w__8874);
  and g__9358(w__8958 ,w__8850 ,w__8864);
  or g__9359(w__8957 ,w__8817 ,w__8904);
  or g__9360(w__8956 ,w__8832 ,w__8872);
  and g__9361(w__8955 ,w__8832 ,w__8872);
  nor g__9362(w__8954 ,w__8801 ,w__8855);
  and g__9363(w__8953 ,w__8801 ,w__8855);
  nor g__9364(w__8952 ,w__8912 ,w__8885);
  or g__9365(w__8951 ,w__8867 ,w__8930);
  nor g__9366(w__8950 ,w__8866 ,w__8931);
  nor g__9367(w__8949 ,w__8925 ,w__8889);
  nor g__9368(w__8948 ,w__8745 ,w__8887);
  or g__9369(w__8947 ,w__8895 ,w__8884);
  xnor g__9370(w__8946 ,w__8833 ,w__8835);
  xnor g__9371(w__8945 ,w__8625 ,w__8799);
  xnor g__9372(w__8944 ,w__8807 ,w__8824);
  xnor g__9373(w__8943 ,w__8622 ,w__8797);
  xnor g__9374(w__8942 ,w__8813 ,w__8811);
  xnor g__9375(w__8941 ,w__8805 ,w__8806);
  xnor g__9376(w__8940 ,w__8803 ,w__8422);
  xnor g__9377(w__8939 ,w__8826 ,w__8827);
  xnor g__9378(w__8938 ,w__8821 ,w__8822);
  xnor g__9379(w__8937 ,w__8830 ,w__8731);
  xnor g__9380(w__8970 ,w__8844 ,w__8737);
  and g__9381(w__8969 ,w__8767 ,w__8892);
  xnor g__9382(w__8968 ,w__8814 ,w__8724);
  xnor g__9383(w__8965 ,w__8842 ,w__8789);
  xnor g__9384(w__8964 ,w__8816 ,w__8725);
  and g__9385(w__8963 ,w__8572 ,w__8894);
  not g__9386(w__8933 ,w__8934);
  not g__9387(w__8932 ,w__7528);
  not g__9388(w__8930 ,w__8931);
  not g__9389(w__8928 ,w__8929);
  not g__9390(w__8927 ,w__8926);
  and g__9391(w__8925 ,w__8623 ,w__8797);
  or g__9392(w__8924 ,w__8819 ,w__8840);
  or g__9393(w__8923 ,w__8419 ,w__8823);
  or g__9394(w__8922 ,w__8835 ,w__8833);
  nor g__9395(w__8921 ,w__8498 ,w__8836);
  and g__9396(w__8920 ,w__8419 ,w__8823);
  and g__9397(w__8919 ,w__8835 ,w__8833);
  or g__9398(w__8918 ,w__8731 ,w__8830);
  and g__9399(w__8917 ,w__8731 ,w__8830);
  or g__9400(w__8916 ,w__8597 ,w__8844);
  or g__9401(w__8915 ,w__8827 ,w__8826);
  or g__9402(w__8914 ,w__8824 ,w__8807);
  and g__9403(w__8913 ,w__8827 ,w__8826);
  and g__9404(w__8912 ,w__8498 ,w__8836);
  nor g__9405(w__8911 ,w__8501 ,w__8802);
  or g__9406(w__8910 ,w__8822 ,w__8821);
  and g__9407(w__8909 ,w__8822 ,w__8821);
  or g__9408(w__8908 ,w__8589 ,w__8814);
  or g__9409(w__8907 ,w__8422 ,w__8803);
  or g__9410(w__8906 ,w__8806 ,w__8805);
  nor g__9411(w__8905 ,w__8623 ,w__8797);
  nor g__9412(w__8904 ,w__8625 ,w__8798);
  or g__9413(w__8903 ,w__8815 ,w__8792);
  and g__9414(w__8902 ,w__8806 ,w__8805);
  and g__9415(w__8901 ,w__8824 ,w__8807);
  or g__9416(w__8900 ,w__8794 ,w__8811);
  nor g__9417(w__8899 ,w__8732 ,w__8810);
  and g__9418(w__8898 ,w__8732 ,w__8810);
  or g__9419(w__13302 ,w__8585 ,w__8793);
  and g__9420(w__8897 ,w__8794 ,w__8811);
  nor g__9421(w__8896 ,w__8611 ,w__8845);
  and g__9422(w__8895 ,w__7677 ,w__8803);
  or g__9423(w__8894 ,w__8571 ,w__8816);
  or g__9424(w__8893 ,w__8624 ,w__8799);
  or g__9425(w__8892 ,w__8766 ,w__8842);
  and g__9426(w__8891 ,w__7725 ,w__8802);
  and g__9427(w__8936 ,w__8627 ,w__8820);
  xnor g__9428(w__8935 ,w__8717 ,w__8502);
  xnor g__9429(w__8934 ,w__8703 ,w__7744);
  xnor g__9430(w__8931 ,w__8736 ,w__8503);
  xnor g__9431(w__8929 ,w__8681 ,w__8695);
  xnor g__9432(w__8926 ,w__8626 ,w__8682);
  not g__9433(w__8869 ,w__8870);
  not g__9434(w__8866 ,w__8867);
  not g__9435(w__8861 ,w__8862);
  not g__9436(w__8852 ,w__8853);
  not g__9437(w__8848 ,w__8849);
  xnor g__9438(w__13367 ,w__8469 ,w__8722);
  xnor g__9439(w__13277 ,w__8692 ,w__7911);
  xnor g__9440(w__13366 ,w__8734 ,w__8712);
  xnor g__9441(w__8847 ,w__8730 ,w__8537);
  xnor g__9442(w__8846 ,w__8733 ,w__8454);
  xnor g__9443(w__8890 ,w__8535 ,w__8721);
  xnor g__9444(w__8889 ,w__8504 ,w__8723);
  xnor g__9445(w__8888 ,w__8548 ,w__8718);
  xnor g__9446(w__8887 ,w__8430 ,w__8719);
  xnor g__9447(w__8886 ,w__8694 ,w__7940);
  xnor g__9448(w__8885 ,w__8484 ,w__8714);
  xnor g__9449(w__8884 ,w__8707 ,w__7944);
  xnor g__9450(w__8883 ,w__8475 ,w__8687);
  xnor g__9451(w__8882 ,w__8551 ,w__8705);
  xnor g__9452(w__8881 ,w__8559 ,w__8700);
  xnor g__9453(w__8880 ,w__8482 ,w__8699);
  xnor g__9454(w__8879 ,w__8550 ,w__8697);
  xnor g__9455(w__8878 ,w__8549 ,w__8689);
  xnor g__9456(w__8877 ,w__8558 ,w__8728);
  xnor g__9457(w__8876 ,w__8552 ,w__8684);
  xnor g__9458(w__8875 ,w__8444 ,w__8683);
  xnor g__9459(w__8874 ,w__8693 ,w__7921);
  xnor g__9460(w__8873 ,w__8735 ,w__8686);
  xnor g__9461(w__8872 ,w__8481 ,w__8716);
  xnor g__9462(w__8871 ,w__8554 ,w__8701);
  xnor g__9463(w__8870 ,w__8456 ,w__8729);
  xnor g__9464(w__8868 ,w__8688 ,w__8500);
  xnor g__9465(w__8867 ,w__8522 ,w__8713);
  xnor g__9466(w__8865 ,w__8450 ,w__8698);
  xnor g__9467(w__8864 ,w__8569 ,w__8711);
  xnor g__9468(w__8863 ,w__8447 ,w__8702);
  xnor g__9469(w__8862 ,w__8517 ,w__8696);
  xnor g__9470(w__8860 ,w__8538 ,w__8691);
  xnor g__9471(w__8859 ,w__8556 ,w__8690);
  xnor g__9472(w__8858 ,w__8526 ,w__8710);
  xnor g__9473(w__8857 ,w__8685 ,w__7942);
  xnor g__9474(w__8856 ,w__8534 ,w__8709);
  xnor g__9475(w__8855 ,w__8472 ,w__8704);
  xnor g__9476(w__8854 ,w__8457 ,w__8720);
  xnor g__9477(w__8853 ,w__8518 ,w__8706);
  xnor g__9478(w__8851 ,w__8524 ,w__8708);
  xnor g__9479(w__8850 ,w__8437 ,w__8727);
  xnor g__9480(w__8849 ,w__8493 ,w__8738);
  not g__9481(w__8838 ,w__8839);
  not g__9482(w__8828 ,w__8829);
  or g__9483(w__8820 ,w__8635 ,w__8735);
  and g__9484(w__8819 ,w__8537 ,w__8730);
  or g__9485(w__8818 ,w__8537 ,w__8730);
  and g__9486(w__8845 ,w__8673 ,w__8757);
  and g__9487(w__8844 ,w__8678 ,w__8772);
  and g__9488(w__8843 ,w__8641 ,w__8769);
  and g__9489(w__8842 ,w__8632 ,w__8763);
  and g__9490(w__8841 ,w__8661 ,w__8776);
  and g__9491(w__8840 ,w__8669 ,w__8782);
  or g__9492(w__8839 ,w__8664 ,w__8777);
  and g__9493(w__8837 ,w__8671 ,w__8780);
  and g__9494(w__8836 ,w__8653 ,w__8765);
  and g__9495(w__8835 ,w__8658 ,w__8775);
  and g__9496(w__8834 ,w__8574 ,w__8787);
  and g__9497(w__8833 ,w__8654 ,w__8773);
  and g__9498(w__8832 ,w__8652 ,w__8771);
  and g__9499(w__8831 ,w__8676 ,w__8786);
  and g__9500(w__8830 ,w__8644 ,w__8770);
  and g__9501(w__8829 ,w__8672 ,w__8783);
  and g__9502(w__8827 ,w__8638 ,w__8768);
  and g__9503(w__8826 ,w__8633 ,w__8764);
  and g__9504(w__8825 ,w__8667 ,w__8781);
  and g__9505(w__8824 ,w__8631 ,w__8760);
  and g__9506(w__8823 ,w__8666 ,w__8779);
  and g__9507(w__8822 ,w__8617 ,w__8788);
  and g__9508(w__8821 ,w__8675 ,w__8759);
  not g__9509(w__8808 ,w__8809);
  not g__9510(w__8801 ,w__8800);
  not g__9511(w__8798 ,w__8799);
  and g__9512(w__8793 ,w__8592 ,w__8734);
  or g__9513(w__13303 ,w__8595 ,w__8743);
  and g__9514(w__8792 ,w__8454 ,w__8733);
  or g__9515(w__8791 ,w__8454 ,w__8733);
  xnor g__9516(w__8790 ,w__8428 ,w__8620);
  xnor g__9517(w__8789 ,w__8521 ,w__8680);
  and g__9518(w__8817 ,w__8648 ,w__8761);
  and g__9519(w__8816 ,w__8584 ,w__8741);
  and g__9520(w__8815 ,w__8613 ,w__8753);
  and g__9521(w__8814 ,w__8578 ,w__8742);
  and g__9522(w__8813 ,w__8591 ,w__8744);
  and g__9523(w__8812 ,w__8600 ,w__8751);
  and g__9524(w__8811 ,w__8640 ,w__8748);
  and g__9525(w__8810 ,w__8599 ,w__8750);
  or g__9526(w__8809 ,w__8577 ,w__8749);
  and g__9527(w__8807 ,w__8581 ,w__8754);
  and g__9528(w__8806 ,w__8612 ,w__8758);
  and g__9529(w__8805 ,w__8608 ,w__8755);
  and g__9530(w__8804 ,w__8590 ,w__8778);
  and g__9531(w__8803 ,w__8582 ,w__8784);
  or g__9532(w__8802 ,w__8576 ,w__8774);
  or g__9533(w__8800 ,w__8603 ,w__8762);
  and g__9534(w__8799 ,w__8587 ,w__8785);
  and g__9535(w__8797 ,w__8610 ,w__8756);
  and g__9536(w__8796 ,w__8619 ,w__8740);
  and g__9537(w__8795 ,w__8601 ,w__8746);
  and g__9538(w__8794 ,w__8570 ,w__8752);
  or g__9539(w__8788 ,w__8567 ,w__8616);
  or g__9540(w__8787 ,w__8568 ,w__8573);
  or g__9541(w__8786 ,w__8566 ,w__8674);
  or g__9542(w__8785 ,w__8565 ,w__8649);
  or g__9543(w__8784 ,w__8492 ,w__8583);
  or g__9544(w__8783 ,w__8670 ,w__8564);
  or g__9545(w__8782 ,w__8480 ,w__8668);
  or g__9546(w__8781 ,w__8563 ,w__8665);
  or g__9547(w__8780 ,w__8562 ,w__8662);
  or g__9548(w__8779 ,w__8560 ,w__8663);
  or g__9549(w__8778 ,w__7866 ,w__8660);
  and g__9550(w__8777 ,w__8681 ,w__8659);
  or g__9551(w__8776 ,w__8558 ,w__8656);
  or g__9552(w__8775 ,w__8557 ,w__8655);
  nor g__9553(w__8774 ,w__8579 ,w__7725);
  or g__9554(w__8773 ,w__8556 ,w__8650);
  or g__9555(w__8772 ,w__8494 ,w__8643);
  or g__9556(w__8771 ,w__7746 ,w__8647);
  or g__9557(w__8770 ,w__8555 ,w__8642);
  or g__9558(w__8769 ,w__8478 ,w__8639);
  or g__9559(w__8768 ,w__8483 ,w__8636);
  or g__9560(w__8767 ,w__8521 ,w__8679);
  nor g__9561(w__8766 ,w__8520 ,w__8680);
  or g__9562(w__8765 ,w__8553 ,w__8629);
  or g__9563(w__8764 ,w__8552 ,w__8628);
  or g__9564(w__8763 ,w__8475 ,w__8630);
  and g__9565(w__8762 ,w__8626 ,w__8657);
  or g__9566(w__8761 ,w__8550 ,w__8677);
  or g__9567(w__8760 ,w__8554 ,w__8645);
  or g__9568(w__8759 ,w__8471 ,w__8614);
  or g__9569(w__8758 ,w__8468 ,w__8609);
  or g__9570(w__8757 ,w__8606 ,w__8491);
  or g__9571(w__8756 ,w__8472 ,w__8607);
  or g__9572(w__8755 ,w__8569 ,w__8605);
  or g__9573(w__8754 ,w__8482 ,w__8602);
  or g__9574(w__8753 ,w__8487 ,w__8604);
  or g__9575(w__8752 ,w__8586 ,w__8493);
  or g__9576(w__8751 ,w__8551 ,w__8588);
  or g__9577(w__8750 ,w__8479 ,w__8598);
  and g__9578(w__8749 ,w__8580 ,w__7677);
  or g__9579(w__8748 ,w__8559 ,w__8596);
  nor g__9580(w__8747 ,w__8428 ,w__8621);
  or g__9581(w__8746 ,w__8561 ,w__8646);
  and g__9582(w__8745 ,w__8428 ,w__8621);
  or g__9583(w__8744 ,w__8490 ,w__8594);
  nor g__9584(w__8743 ,w__8469 ,w__8637);
  or g__9585(w__8742 ,w__8575 ,w__8484);
  or g__9586(w__8741 ,w__8481 ,w__8651);
  or g__9587(w__8740 ,w__7744 ,w__8615);
  xnor g__9588(w__13368 ,w__8495 ,w__8416);
  xnor g__9589(w__8739 ,w__8427 ,w__7727);
  xnor g__9590(w__8738 ,w__8461 ,w__7919);
  xnor g__9591(w__8737 ,w__8441 ,w__8420);
  xnor g__9592(w__8736 ,w__8506 ,w__7746);
  xnor g__9593(w__8729 ,w__8423 ,w__8490);
  xnor g__9594(w__8728 ,w__8540 ,w__7939);
  xnor g__9595(w__8727 ,w__8468 ,w__7913);
  xnor g__9596(w__8726 ,w__8568 ,w__7945);
  xnor g__9597(w__8725 ,w__7675 ,w__7915);
  xnor g__9598(w__8724 ,w__8510 ,w__8497);
  xnor g__9599(w__8723 ,w__8567 ,w__8174);
  xnor g__9600(w__8722 ,w__8179 ,w__8463);
  xnor g__9601(w__8721 ,w__8480 ,w__8177);
  xnor g__9602(w__8720 ,w__8555 ,w__8175);
  xnor g__9603(w__8719 ,w__8479 ,w__8178);
  xnor g__9604(w__8718 ,w__8487 ,w__8176);
  xnor g__9605(w__8717 ,w__8443 ,w__7941);
  xnor g__9606(w__8716 ,w__8505 ,w__8442);
  xnor g__9607(w__8715 ,w__8440 ,w__7917);
  xnor g__9608(w__8714 ,w__8438 ,w__7943);
  xnor g__9609(w__8713 ,w__8483 ,w__7914);
  xnor g__9610(w__8712 ,w__8465 ,w__8425);
  xnor g__9611(w__8711 ,w__8458 ,w__8433);
  xnor g__9612(w__8710 ,w__8525 ,w__8478);
  xnor g__9613(w__8709 ,w__8529 ,w__8471);
  xnor g__9614(w__8708 ,w__8553 ,w__8530);
  xnor g__9615(w__8707 ,w__8528 ,w__8494);
  xnor g__9616(w__8706 ,w__8562 ,w__8539);
  xnor g__9617(w__8705 ,w__8434 ,w__8436);
  xnor g__9618(w__8704 ,w__8426 ,w__8459);
  xnor g__9619(w__8703 ,w__8449 ,w__8445);
  xnor g__9620(w__8702 ,w__8561 ,w__7918);
  xnor g__9621(w__8701 ,w__8509 ,w__8513);
  xnor g__9622(w__8700 ,w__8429 ,w__8511);
  xnor g__9623(w__8699 ,w__8462 ,w__8446);
  xnor g__9624(w__8698 ,w__8448 ,w__8565);
  xnor g__9625(w__8697 ,w__8453 ,w__8523);
  xnor g__9626(w__8696 ,w__8532 ,w__8563);
  xnor g__9627(w__8695 ,w__8543 ,w__8545);
  xnor g__9628(w__8694 ,w__8566 ,w__8547);
  xnor g__9629(w__8693 ,w__8491 ,w__8541);
  xnor g__9630(w__8692 ,w__7923 ,w__8496);
  xnor g__9631(w__8691 ,w__8557 ,w__8536);
  xnor g__9632(w__8690 ,w__8455 ,w__8527);
  xnor g__9633(w__8689 ,w__8560 ,w__8512);
  xnor g__9634(w__8688 ,w__8531 ,w__8533);
  xnor g__9635(w__8687 ,w__8514 ,w__8516);
  xnor g__9636(w__8686 ,w__8507 ,w__8508);
  xnor g__9637(w__8685 ,w__8564 ,w__8546);
  xnor g__9638(w__8684 ,w__8515 ,w__8519);
  xnor g__9639(w__8683 ,w__8435 ,w__8492);
  xnor g__9640(w__8682 ,w__8452 ,w__8432);
  xnor g__9641(w__8735 ,w__8488 ,w__8410);
  xnor g__9642(w__8734 ,w__8404 ,w__8470);
  xnor g__9643(w__8733 ,w__8412 ,w__8466);
  xnor g__9644(w__8732 ,w__8414 ,w__8476);
  xnor g__9645(w__8731 ,w__8408 ,w__8473);
  xnor g__9646(w__8730 ,w__8406 ,w__8485);
  not g__9647(w__8679 ,w__8680);
  or g__9648(w__8678 ,w__7747 ,w__8528);
  and g__9649(w__8677 ,w__8523 ,w__8453);
  or g__9650(w__8676 ,w__7748 ,w__8547);
  or g__9651(w__8675 ,w__8529 ,w__8534);
  and g__9652(w__8674 ,w__7940 ,w__8547);
  or g__9653(w__8673 ,w__7757 ,w__8541);
  or g__9654(w__8672 ,w__7755 ,w__8546);
  or g__9655(w__8671 ,w__8539 ,w__8518);
  and g__9656(w__8670 ,w__7942 ,w__8546);
  or g__9657(w__8669 ,w__8177 ,w__8535);
  and g__9658(w__8668 ,w__8177 ,w__8535);
  or g__9659(w__8667 ,w__8532 ,w__8517);
  or g__9660(w__8666 ,w__8512 ,w__8549);
  and g__9661(w__8665 ,w__8532 ,w__8517);
  nor g__9662(w__8664 ,w__8545 ,w__8543);
  and g__9663(w__8663 ,w__8512 ,w__8549);
  and g__9664(w__8662 ,w__8539 ,w__8518);
  or g__9665(w__8661 ,w__7753 ,w__8540);
  and g__9666(w__8660 ,w__8445 ,w__8449);
  or g__9667(w__8659 ,w__8544 ,w__8542);
  or g__9668(w__8658 ,w__8538 ,w__8536);
  or g__9669(w__8657 ,w__8431 ,w__8451);
  and g__9670(w__8656 ,w__7939 ,w__8540);
  and g__9671(w__8655 ,w__8538 ,w__8536);
  or g__9672(w__8654 ,w__8527 ,w__8455);
  or g__9673(w__8653 ,w__8530 ,w__8524);
  or g__9674(w__8652 ,w__8533 ,w__8531);
  and g__9675(w__8651 ,w__8442 ,w__8505);
  and g__9676(w__8650 ,w__8527 ,w__8455);
  and g__9677(w__8649 ,w__8450 ,w__8448);
  or g__9678(w__8648 ,w__8523 ,w__8453);
  and g__9679(w__8647 ,w__8533 ,w__8531);
  and g__9680(w__8646 ,w__7752 ,w__8447);
  and g__9681(w__8645 ,w__8513 ,w__8509);
  or g__9682(w__8644 ,w__8175 ,w__8457);
  and g__9683(w__8643 ,w__7944 ,w__8528);
  and g__9684(w__8642 ,w__8175 ,w__8457);
  or g__9685(w__8641 ,w__8526 ,w__8525);
  or g__9686(w__8640 ,w__8511 ,w__8429);
  and g__9687(w__8639 ,w__8526 ,w__8525);
  or g__9688(w__8638 ,w__7751 ,w__8522);
  and g__9689(w__8637 ,w__8180 ,w__8463);
  and g__9690(w__8636 ,w__7914 ,w__8522);
  and g__9691(w__8635 ,w__8508 ,w__8507);
  or g__9692(w__8634 ,w__7679 ,w__8510);
  or g__9693(w__8633 ,w__8519 ,w__8515);
  or g__9694(w__8632 ,w__8516 ,w__8514);
  or g__9695(w__8631 ,w__8513 ,w__8509);
  and g__9696(w__8630 ,w__8516 ,w__8514);
  and g__9697(w__8629 ,w__8530 ,w__8524);
  and g__9698(w__8628 ,w__8519 ,w__8515);
  or g__9699(w__8627 ,w__8508 ,w__8507);
  and g__9700(w__8681 ,w__8409 ,w__8474);
  and g__9701(w__8680 ,w__8411 ,w__8489);
  not g__9702(w__8624 ,w__8625);
  not g__9703(w__8623 ,w__8622);
  not g__9704(w__8621 ,w__8620);
  or g__9705(w__8619 ,w__8499 ,w__8506);
  and g__9706(w__8618 ,w__7912 ,w__8427);
  or g__9707(w__8617 ,w__8174 ,w__8504);
  and g__9708(w__8616 ,w__8174 ,w__8504);
  and g__9709(w__8615 ,w__8499 ,w__8506);
  and g__9710(w__8614 ,w__8529 ,w__8534);
  or g__9711(w__8613 ,w__8176 ,w__8548);
  or g__9712(w__8612 ,w__7749 ,w__8437);
  nor g__9713(w__8611 ,w__7912 ,w__8427);
  or g__9714(w__8610 ,w__8459 ,w__8426);
  and g__9715(w__8609 ,w__7913 ,w__8437);
  or g__9716(w__8608 ,w__8433 ,w__8458);
  and g__9717(w__8607 ,w__8459 ,w__8426);
  and g__9718(w__8606 ,w__7921 ,w__8541);
  and g__9719(w__8605 ,w__8433 ,w__8458);
  and g__9720(w__8604 ,w__8176 ,w__8548);
  nor g__9721(w__8603 ,w__8432 ,w__8452);
  and g__9722(w__8602 ,w__8446 ,w__8462);
  or g__9723(w__8601 ,w__7918 ,w__8447);
  or g__9724(w__8600 ,w__8436 ,w__8434);
  or g__9725(w__8599 ,w__8178 ,w__8430);
  and g__9726(w__8598 ,w__8178 ,w__8430);
  and g__9727(w__8597 ,w__8441 ,w__8421);
  and g__9728(w__8596 ,w__8511 ,w__8429);
  nor g__9729(w__8595 ,w__8180 ,w__8463);
  and g__9730(w__8594 ,w__8456 ,w__8423);
  or g__9731(w__8593 ,w__8441 ,w__8421);
  or g__9732(w__8592 ,w__8424 ,w__8464);
  or g__9733(w__8591 ,w__8456 ,w__8423);
  or g__9734(w__8590 ,w__8445 ,w__8449);
  and g__9735(w__8589 ,w__7679 ,w__8510);
  and g__9736(w__8588 ,w__8436 ,w__8434);
  or g__9737(w__8587 ,w__8450 ,w__8448);
  nor g__9738(w__8586 ,w__7920 ,w__8461);
  nor g__9739(w__8585 ,w__8425 ,w__8465);
  or g__9740(w__8584 ,w__8442 ,w__8505);
  and g__9741(w__8583 ,w__8444 ,w__8435);
  or g__9742(w__8582 ,w__8444 ,w__8435);
  or g__9743(w__8581 ,w__8446 ,w__8462);
  or g__9744(w__8580 ,w__7916 ,w__8439);
  and g__9745(w__8579 ,w__7758 ,w__8443);
  or g__9746(w__8578 ,w__7754 ,w__8438);
  nor g__9747(w__8577 ,w__7917 ,w__8440);
  nor g__9748(w__8576 ,w__7758 ,w__8443);
  and g__9749(w__8575 ,w__7943 ,w__8438);
  or g__9750(w__8574 ,w__7756 ,w__7681);
  and g__9751(w__8573 ,w__7945 ,w__7681);
  or g__9752(w__8572 ,w__7750 ,w__7675);
  and g__9753(w__8571 ,w__7915 ,w__8418);
  or g__9754(w__8570 ,w__7919 ,w__8460);
  and g__9755(w__13304 ,w__8417 ,w__8495);
  and g__9756(w__8626 ,w__8415 ,w__8477);
  and g__9757(w__8625 ,w__8407 ,w__8486);
  and g__9758(w__8622 ,w__8413 ,w__8467);
  and g__9759(w__8620 ,w__8405 ,w__8470);
  not g__9760(w__8544 ,w__8545);
  not g__9761(w__8542 ,w__8543);
  not g__9762(w__8520 ,w__8521);
  not g__9763(w__8501 ,w__8502);
  not g__9764(w__8499 ,w__8500);
  not g__9765(w__8498 ,w__8497);
  or g__9766(w__8496 ,w__8187 ,w__8290);
  and g__9767(w__8569 ,w__8215 ,w__8319);
  and g__9768(w__8568 ,w__8238 ,w__8293);
  and g__9769(w__8567 ,w__8249 ,w__8332);
  and g__9770(w__8566 ,w__8126 ,w__8283);
  and g__9771(w__8565 ,w__8138 ,w__8296);
  and g__9772(w__8564 ,w__8237 ,w__8365);
  and g__9773(w__8563 ,w__8234 ,w__8366);
  and g__9774(w__8562 ,w__8233 ,w__8361);
  and g__9775(w__8561 ,w__8120 ,w__8271);
  and g__9776(w__8560 ,w__8231 ,w__8292);
  and g__9777(w__8559 ,w__8223 ,w__8347);
  and g__9778(w__8558 ,w__8225 ,w__8354);
  and g__9779(w__8557 ,w__8244 ,w__8352);
  and g__9780(w__8556 ,w__8220 ,w__8350);
  and g__9781(w__8555 ,w__8194 ,w__8345);
  and g__9782(w__8554 ,w__8229 ,w__8329);
  and g__9783(w__8553 ,w__8205 ,w__8402);
  and g__9784(w__8552 ,w__8209 ,w__8338);
  and g__9785(w__8551 ,w__8214 ,w__8311);
  and g__9786(w__8550 ,w__8164 ,w__8378);
  and g__9787(w__8549 ,w__8236 ,w__8364);
  and g__9788(w__8548 ,w__8157 ,w__8317);
  and g__9789(w__8547 ,w__8201 ,w__8376);
  or g__9790(w__8546 ,w__8183 ,w__8289);
  and g__9791(w__8545 ,w__8148 ,w__8359);
  and g__9792(w__8543 ,w__8150 ,w__8358);
  or g__9793(w__8541 ,w__8192 ,w__8286);
  and g__9794(w__8540 ,w__8227 ,w__8355);
  or g__9795(w__8539 ,w__8190 ,w__8288);
  and g__9796(w__8538 ,w__8242 ,w__8356);
  and g__9797(w__8537 ,w__8243 ,w__8373);
  and g__9798(w__8536 ,w__8226 ,w__8353);
  and g__9799(w__8535 ,w__8240 ,w__8372);
  and g__9800(w__8534 ,w__8206 ,w__8330);
  and g__9801(w__8533 ,w__8221 ,w__8297);
  and g__9802(w__8532 ,w__8135 ,w__8369);
  and g__9803(w__8531 ,w__8121 ,w__8279);
  or g__9804(w__8530 ,w__8185 ,w__8287);
  and g__9805(w__8529 ,w__8202 ,w__8331);
  and g__9806(w__8528 ,w__8130 ,w__8278);
  and g__9807(w__8527 ,w__8136 ,w__8351);
  and g__9808(w__8526 ,w__8213 ,w__8343);
  and g__9809(w__8525 ,w__8212 ,w__8342);
  and g__9810(w__8524 ,w__8128 ,w__8280);
  and g__9811(w__8523 ,w__8140 ,w__8315);
  and g__9812(w__8522 ,w__8151 ,w__8381);
  and g__9813(w__8521 ,w__8207 ,w__8389);
  and g__9814(w__8519 ,w__8154 ,w__8395);
  and g__9815(w__8518 ,w__8235 ,w__8367);
  and g__9816(w__8517 ,w__8210 ,w__8403);
  and g__9817(w__8516 ,w__8197 ,w__8377);
  and g__9818(w__8515 ,w__8204 ,w__8399);
  and g__9819(w__8514 ,w__8167 ,w__8268);
  or g__9820(w__8513 ,w__8181 ,w__8285);
  or g__9821(w__8512 ,w__8188 ,w__8284);
  and g__9822(w__8511 ,w__8166 ,w__8299);
  and g__9823(w__8510 ,w__8122 ,w__8282);
  and g__9824(w__8509 ,w__8195 ,w__8335);
  and g__9825(w__8508 ,w__8158 ,w__8328);
  and g__9826(w__8507 ,w__8196 ,w__8336);
  and g__9827(w__8506 ,w__8127 ,w__8275);
  and g__9828(w__8505 ,w__8153 ,w__8340);
  and g__9829(w__8504 ,w__8246 ,w__8334);
  and g__9830(w__8503 ,w__8241 ,w__8333);
  and g__9831(w__8502 ,w__8132 ,w__8281);
  and g__9832(w__8500 ,w__8218 ,w__8349);
  and g__9833(w__8497 ,w__8199 ,w__8337);
  not g__9834(w__8489 ,w__8488);
  not g__9835(w__8486 ,w__8485);
  not g__9836(w__8477 ,w__8476);
  not g__9837(w__8474 ,w__8473);
  not g__9838(w__8467 ,w__8466);
  not g__9839(w__8464 ,w__8465);
  not g__9840(w__8460 ,w__8461);
  not g__9841(w__8451 ,w__8452);
  not g__9842(w__8439 ,w__8440);
  not g__9843(w__8431 ,w__8432);
  not g__9844(w__8424 ,w__8425);
  not g__9845(w__8421 ,w__8420);
  not g__9846(w__8419 ,w__8418);
  or g__9847(w__13369 ,w__8261 ,w__8392);
  or g__9848(w__13370 ,w__8255 ,w__8368);
  or g__9849(w__13305 ,w__8247 ,w__8302);
  or g__9850(w__8495 ,w__8262 ,w__8384);
  and g__9851(w__8494 ,w__8216 ,w__8348);
  and g__9852(w__8493 ,w__8208 ,w__8312);
  and g__9853(w__8492 ,w__8265 ,w__8374);
  and g__9854(w__8491 ,w__8124 ,w__8277);
  and g__9855(w__8490 ,w__8145 ,w__8303);
  and g__9856(w__8488 ,w__8159 ,w__8394);
  and g__9857(w__8487 ,w__8252 ,w__8390);
  and g__9858(w__8485 ,w__8251 ,w__8383);
  and g__9859(w__8484 ,w__8134 ,w__8274);
  and g__9860(w__8483 ,w__8189 ,w__8387);
  and g__9861(w__8482 ,w__8123 ,w__8272);
  and g__9862(w__8481 ,w__8217 ,w__8380);
  and g__9863(w__8480 ,w__8263 ,w__8400);
  and g__9864(w__8479 ,w__8264 ,w__8388);
  and g__9865(w__8478 ,w__8259 ,w__8397);
  and g__9866(w__8476 ,w__8258 ,w__8396);
  and g__9867(w__8475 ,w__8260 ,w__8391);
  and g__9868(w__8473 ,w__8256 ,w__8398);
  and g__9869(w__8472 ,w__8254 ,w__8393);
  and g__9870(w__8471 ,w__8253 ,w__8401);
  or g__9871(w__8470 ,w__8228 ,w__8386);
  and g__9872(w__8469 ,w__8257 ,w__8385);
  and g__9873(w__8468 ,w__8125 ,w__8273);
  and g__9874(w__8466 ,w__8198 ,w__8325);
  and g__9875(w__8465 ,w__8203 ,w__8304);
  and g__9876(w__8463 ,w__8147 ,w__8306);
  and g__9877(w__8462 ,w__8211 ,w__8370);
  or g__9878(w__8461 ,w__7922 ,w__8382);
  and g__9879(w__8459 ,w__8219 ,w__8324);
  and g__9880(w__8458 ,w__8239 ,w__8360);
  and g__9881(w__8457 ,w__8165 ,w__8346);
  and g__9882(w__8456 ,w__8137 ,w__8357);
  and g__9883(w__8455 ,w__8160 ,w__8320);
  and g__9884(w__8454 ,w__8161 ,w__8318);
  and g__9885(w__8453 ,w__8245 ,w__8322);
  and g__9886(w__8452 ,w__8149 ,w__8321);
  and g__9887(w__8450 ,w__8146 ,w__8294);
  and g__9888(w__8449 ,w__8141 ,w__8375);
  and g__9889(w__8448 ,w__8131 ,w__8339);
  and g__9890(w__8447 ,w__8155 ,w__8298);
  and g__9891(w__8446 ,w__8144 ,w__8326);
  and g__9892(w__8445 ,w__8139 ,w__8295);
  and g__9893(w__8444 ,w__8224 ,w__8371);
  and g__9894(w__8443 ,w__8193 ,w__8379);
  and g__9895(w__8442 ,w__8182 ,w__8363);
  and g__9896(w__8441 ,w__8186 ,w__8344);
  and g__9897(w__8440 ,w__8191 ,w__8362);
  and g__9898(w__8438 ,w__8184 ,w__8301);
  and g__9899(w__8437 ,w__8163 ,w__8327);
  and g__9900(w__8436 ,w__8248 ,w__8314);
  and g__9901(w__8435 ,w__8133 ,w__8269);
  and g__9902(w__8434 ,w__8162 ,w__8313);
  and g__9903(w__8432 ,w__8156 ,w__8316);
  and g__9904(w__8430 ,w__8222 ,w__8309);
  and g__9905(w__8429 ,w__8200 ,w__8308);
  and g__9906(w__8428 ,w__8230 ,w__8307);
  or g__9907(w__8427 ,w__8187 ,w__8276);
  and g__9908(w__8426 ,w__8232 ,w__8323);
  and g__9909(w__8425 ,w__8250 ,w__8305);
  and g__9910(w__8423 ,w__8129 ,w__8270);
  and g__9911(w__8422 ,w__8142 ,w__8310);
  and g__9912(w__8420 ,w__8143 ,w__8341);
  and g__9913(w__8418 ,w__8152 ,w__8300);
  not g__9914(w__8417 ,w__8416);
  not g__9915(w__8415 ,w__8414);
  not g__9916(w__8413 ,w__8412);
  not g__9917(w__8411 ,w__8410);
  not g__9918(w__8409 ,w__8408);
  not g__9919(w__8407 ,w__8406);
  not g__9920(w__8405 ,w__8404);
  or g__9921(w__8403 ,w__8007 ,w__7593);
  or g__9922(w__8402 ,w__8021 ,w__7578);
  or g__9923(w__8401 ,w__7983 ,w__7552);
  or g__9924(w__8400 ,w__7971 ,w__7644);
  or g__9925(w__8399 ,w__8079 ,w__7575);
  or g__9926(w__8398 ,w__7976 ,w__7552);
  or g__9927(w__8397 ,w__7978 ,w__7619);
  or g__9928(w__8396 ,w__7972 ,w__7640);
  or g__9929(w__8395 ,w__7969 ,w__7635);
  or g__9930(w__8394 ,w__8004 ,w__7571);
  or g__9931(w__8393 ,w__7980 ,w__7641);
  nor g__9932(w__8392 ,w__7643 ,w__7973);
  or g__9933(w__8391 ,w__7974 ,w__7619);
  or g__9934(w__8390 ,w__7979 ,w__7620);
  or g__9935(w__8389 ,w__7975 ,w__7632);
  or g__9936(w__8388 ,w__7981 ,w__7643);
  or g__9937(w__8387 ,w__8030 ,w__7637);
  nor g__9938(w__8386 ,w__7641 ,w__7985);
  or g__9939(w__8385 ,w__7982 ,w__7671);
  nor g__9940(w__8384 ,w__7644 ,w__7984);
  or g__9941(w__8383 ,w__7977 ,w__7670);
  nor g__9942(w__8382 ,w__7640 ,w__7970);
  or g__9943(w__8381 ,w__8100 ,w__7584);
  or g__9944(w__8380 ,w__8056 ,w__7563);
  or g__9945(w__8379 ,w__8057 ,w__7611);
  or g__9946(w__8378 ,w__8102 ,w__7590);
  or g__9947(w__8377 ,w__8066 ,w__7587);
  or g__9948(w__8376 ,w__8031 ,w__7605);
  or g__9949(w__8375 ,w__7989 ,w__7634);
  or g__9950(w__8374 ,w__7994 ,w__7566);
  or g__9951(w__8373 ,w__8061 ,w__7610);
  or g__9952(w__8372 ,w__8083 ,w__7652);
  or g__9953(w__8371 ,w__8018 ,w__7646);
  or g__9954(w__8370 ,w__8072 ,w__7569);
  or g__9955(w__8369 ,w__8097 ,w__7608);
  nor g__9956(w__8368 ,w__7620 ,w__7947);
  or g__9957(w__8367 ,w__8078 ,w__7664);
  or g__9958(w__8366 ,w__8062 ,w__7604);
  or g__9959(w__8365 ,w__8026 ,w__7565);
  or g__9960(w__8364 ,w__7996 ,w__7649);
  or g__9961(w__8363 ,w__8088 ,w__7631);
  or g__9962(w__8362 ,w__8080 ,w__7560);
  or g__9963(w__8361 ,w__8073 ,w__7568);
  or g__9964(w__8360 ,w__8082 ,w__7587);
  or g__9965(w__8359 ,w__8103 ,w__7563);
  or g__9966(w__8358 ,w__8074 ,w__7589);
  or g__9967(w__8357 ,w__8006 ,w__7586);
  or g__9968(w__8356 ,w__7949 ,w__7562);
  or g__9969(w__8355 ,w__8070 ,w__7578);
  or g__9970(w__8354 ,w__8071 ,w__7607);
  or g__9971(w__8353 ,w__8075 ,w__7577);
  or g__9972(w__8352 ,w__8065 ,w__7661);
  or g__9973(w__8351 ,w__8101 ,w__7655);
  or g__9974(w__8350 ,w__8063 ,w__7586);
  or g__9975(w__8349 ,w__8060 ,w__7569);
  or g__9976(w__8348 ,w__8014 ,w__7577);
  or g__9977(w__8347 ,w__8012 ,w__7562);
  or g__9978(w__8346 ,w__8022 ,w__7559);
  or g__9979(w__8345 ,w__8024 ,w__7637);
  or g__9980(w__8344 ,w__7988 ,w__7604);
  or g__9981(w__8343 ,w__8067 ,w__7590);
  or g__9982(w__8342 ,w__8086 ,w__7649);
  or g__9983(w__8341 ,w__8064 ,w__7634);
  or g__9984(w__8340 ,w__8027 ,w__7575);
  or g__9985(w__8416 ,w__7907 ,w__8118);
  or g__9986(w__8414 ,w__7932 ,w__8115);
  or g__9987(w__8412 ,w__7900 ,w__8116);
  or g__9988(w__8410 ,w__7905 ,w__8114);
  or g__9989(w__8408 ,w__7903 ,w__8113);
  or g__9990(w__8406 ,w__7908 ,w__8119);
  or g__9991(w__8404 ,w__7897 ,w__8117);
  or g__9992(w__8339 ,w__8042 ,w__7595);
  or g__9993(w__8338 ,w__8003 ,w__7566);
  or g__9994(w__8337 ,w__8009 ,w__7610);
  or g__9995(w__8336 ,w__8019 ,w__7583);
  or g__9996(w__8335 ,w__8011 ,w__7574);
  or g__9997(w__8334 ,w__8089 ,w__7574);
  or g__9998(w__8333 ,w__8084 ,w__7560);
  or g__9999(w__8332 ,w__8032 ,w__7546);
  or g__10000(w__8331 ,w__8020 ,w__7568);
  or g__10001(w__8330 ,w__8092 ,w__7593);
  or g__10002(w__8329 ,w__7997 ,w__7646);
  or g__10003(w__8328 ,w__7950 ,w__7589);
  or g__10004(w__8327 ,w__8017 ,w__7653);
  or g__10005(w__8326 ,w__8068 ,w__7664);
  or g__10006(w__8325 ,w__8090 ,w__7572);
  or g__10007(w__8324 ,w__8037 ,w__7548);
  or g__10008(w__8323 ,w__7987 ,w__7607);
  or g__10009(w__8322 ,w__8095 ,w__7592);
  or g__10010(w__8321 ,w__8002 ,w__7546);
  or g__10011(w__8320 ,w__7986 ,w__7622);
  or g__10012(w__8319 ,w__8028 ,w__7592);
  or g__10013(w__8318 ,w__8010 ,w__7584);
  or g__10014(w__8317 ,w__7999 ,w__7655);
  or g__10015(w__8316 ,w__8016 ,w__7631);
  or g__10016(w__8315 ,w__7998 ,w__7548);
  or g__10017(w__8314 ,w__7946 ,w__7559);
  or g__10018(w__8313 ,w__8099 ,w__7623);
  or g__10019(w__8312 ,w__8000 ,w__7622);
  or g__10020(w__8311 ,w__7992 ,w__7661);
  or g__10021(w__8310 ,w__8059 ,w__7650);
  or g__10022(w__8309 ,w__8013 ,w__7572);
  or g__10023(w__8308 ,w__8069 ,w__7583);
  or g__10024(w__8307 ,w__8077 ,w__7540);
  or g__10025(w__8306 ,w__8008 ,w__7638);
  or g__10026(w__8305 ,w__8034 ,w__7540);
  or g__10027(w__8304 ,w__8098 ,w__7571);
  or g__10028(w__8303 ,w__7993 ,w__7544);
  nor g__10029(w__8302 ,w__7638 ,w__8039);
  or g__10030(w__8301 ,w__8023 ,w__7550);
  or g__10031(w__8300 ,w__8096 ,w__7550);
  or g__10032(w__8299 ,w__8025 ,w__7647);
  or g__10033(w__8298 ,w__8015 ,w__7565);
  or g__10034(w__8297 ,w__7991 ,w__7538);
  or g__10035(w__8296 ,w__7990 ,w__7652);
  or g__10036(w__8295 ,w__8105 ,w__7538);
  or g__10037(w__8294 ,w__8001 ,w__7544);
  or g__10038(w__8293 ,w__8005 ,w__7665);
  or g__10039(w__8292 ,w__7995 ,w__7662);
  nor g__10040(w__8290 ,w__7629 ,w__7599);
  nor g__10041(w__8289 ,w__7635 ,w__7884);
  nor g__10042(w__8288 ,w__7608 ,w__7887);
  nor g__10043(w__8287 ,w__7605 ,w__7885);
  nor g__10044(w__8286 ,w__7611 ,w__7872);
  nor g__10045(w__8285 ,w__7632 ,w__7886);
  nor g__10046(w__8284 ,w__7623 ,w__7888);
  or g__10047(w__8283 ,w__8094 ,w__7596);
  or g__10048(w__8282 ,w__8091 ,w__7601);
  or g__10049(w__8281 ,w__8085 ,w__7598);
  or g__10050(w__8280 ,w__8093 ,w__7595);
  or g__10051(w__8279 ,w__8081 ,w__7596);
  or g__10052(w__8278 ,w__8107 ,w__7536);
  or g__10053(w__8277 ,w__8058 ,w__7668);
  nor g__10054(w__8276 ,w__7602 ,w__8076);
  or g__10055(w__8275 ,w__8087 ,w__7601);
  or g__10056(w__8274 ,w__8104 ,w__7598);
  or g__10057(w__8273 ,w__8109 ,w__7602);
  or g__10058(w__8272 ,w__8110 ,w__7667);
  or g__10059(w__8271 ,w__8108 ,w__7667);
  or g__10060(w__8270 ,w__8111 ,w__7599);
  or g__10061(w__8269 ,w__8106 ,w__7536);
  or g__10062(w__8268 ,w__8029 ,w__7656);
  or g__10063(w__8265 ,w__8078 ,w__7796);
  or g__10064(w__8264 ,w__7626 ,w__7972);
  or g__10065(w__8263 ,w__7614 ,w__7977);
  nor g__10066(w__8262 ,w__7626 ,w__7982);
  nor g__10067(w__8261 ,w__7614 ,w__7984);
  or g__10068(w__8260 ,w__7613 ,w__7978);
  or g__10069(w__8259 ,w__7625 ,w__7976);
  or g__10070(w__8258 ,w__7616 ,w__7979);
  or g__10071(w__8257 ,w__7625 ,w__7985);
  or g__10072(w__8256 ,w__7613 ,w__7971);
  nor g__10073(w__8255 ,w__7617 ,w__7973);
  or g__10074(w__8254 ,w__7616 ,w__7983);
  or g__10075(w__8253 ,w__7617 ,w__7974);
  or g__10076(w__8252 ,w__7554 ,w__7980);
  or g__10077(w__8251 ,w__7554 ,w__7970);
  or g__10078(w__8250 ,w__8077 ,w__7835);
  or g__10079(w__8249 ,w__8004 ,w__7820);
  or g__10080(w__8248 ,w__7999 ,w__7784);
  nor g__10081(w__8247 ,w__8008 ,w__7827);
  or g__10082(w__8246 ,w__8029 ,w__7793);
  or g__10083(w__8245 ,w__8069 ,w__7838);
  or g__10084(w__8244 ,w__8007 ,w__7838);
  or g__10085(w__8243 ,w__8012 ,w__7805);
  or g__10086(w__8242 ,w__8103 ,w__7805);
  or g__10087(w__8241 ,w__8079 ,w__7793);
  or g__10088(w__8240 ,w__7990 ,w__7826);
  or g__10089(w__8239 ,w__8060 ,w__7808);
  or g__10090(w__8238 ,w__8009 ,w__7797);
  or g__10091(w__8237 ,w__8057 ,w__7800);
  or g__10092(w__8236 ,w__8031 ,w__7814);
  or g__10093(w__8235 ,w__8015 ,w__7796);
  or g__10094(w__8234 ,w__7998 ,w__7814);
  or g__10095(w__8233 ,w__7988 ,w__7809);
  or g__10096(w__8232 ,w__8089 ,w__7785);
  or g__10097(w__8231 ,w__8088 ,w__7836);
  or g__10098(w__8230 ,w__7992 ,w__7835);
  or g__10099(w__8229 ,w__8018 ,w__7760);
  nor g__10100(w__8228 ,w__7699 ,w__7981);
  or g__10101(w__8227 ,w__8096 ,w__7769);
  or g__10102(w__8226 ,w__8074 ,w__7769);
  or g__10103(w__8225 ,w__8027 ,w__7788);
  or g__10104(w__8224 ,w__8014 ,w__7761);
  or g__10105(w__8223 ,w__8105 ,w__7799);
  or g__10106(w__8222 ,w__8099 ,w__7821);
  or g__10107(w__8221 ,w__8056 ,w__7802);
  or g__10108(w__8220 ,w__8062 ,w__7812);
  or g__10109(w__8219 ,w__8020 ,w__7808);
  or g__10110(w__8218 ,w__7996 ,w__7811);
  or g__10111(w__8217 ,w__8068 ,w__7802);
  or g__10112(w__8216 ,w__8064 ,w__7764);
  or g__10113(w__8215 ,w__8100 ,w__7832);
  or g__10114(w__8214 ,w__8016 ,w__7963);
  or g__10115(w__8213 ,w__8075 ,w__7760);
  or g__10116(w__8212 ,w__8063 ,w__7817);
  or g__10117(w__8211 ,w__8059 ,w__7817);
  or g__10118(w__8210 ,w__8095 ,w__7832);
  or g__10119(w__8209 ,w__7991 ,w__7799);
  or g__10120(w__8208 ,w__8017 ,w__7824);
  or g__10121(w__8207 ,w__8065 ,w__7833);
  or g__10122(w__8206 ,w__8019 ,w__7836);
  or g__10123(w__8205 ,w__8023 ,w__7763);
  or g__10124(w__8204 ,w__8071 ,w__7784);
  or g__10125(w__8203 ,w__8013 ,w__7820);
  or g__10126(w__8202 ,w__8066 ,w__7811);
  or g__10127(w__8201 ,w__8072 ,w__7815);
  or g__10128(w__8200 ,w__8028 ,w__7839);
  or g__10129(w__8199 ,w__8026 ,w__7806);
  or g__10130(w__8198 ,w__8032 ,w__7823);
  or g__10131(w__8197 ,w__8086 ,w__7812);
  or g__10132(w__8196 ,w__7975 ,w__7729);
  or g__10133(w__8195 ,w__8080 ,w__7787);
  or g__10134(w__8194 ,w__7986 ,w__7830);
  or g__10135(w__8267 ,w__7952 ,w__7688);
  or g__10136(w__8266 ,in17[0] ,w__8041);
  not g__10137(w__8193 ,w__8192);
  not g__10138(w__8191 ,w__8190);
  not g__10139(w__8189 ,w__8188);
  not g__10140(w__8186 ,w__8185);
  not g__10141(w__8184 ,w__8183);
  not g__10142(w__8182 ,w__8181);
  not g__10143(w__8180 ,w__8179);
  or g__10144(w__8167 ,w__8022 ,w__7790);
  or g__10145(w__8166 ,w__7989 ,w__7766);
  or g__10146(w__8165 ,w__8101 ,w__7790);
  or g__10147(w__8164 ,w__8025 ,w__7766);
  or g__10148(w__8163 ,w__8030 ,w__7829);
  or g__10149(w__8162 ,w__8002 ,w__7823);
  or g__10150(w__8161 ,w__8092 ,w__7729);
  or g__10151(w__8160 ,w__8083 ,w__7826);
  or g__10152(w__8159 ,w__8024 ,w__7824);
  or g__10153(w__8158 ,w__8067 ,w__7763);
  or g__10154(w__8157 ,w__7987 ,w__7787);
  or g__10155(w__8156 ,w__8010 ,w__7839);
  or g__10156(w__8155 ,w__8005 ,w__7800);
  or g__10157(w__8154 ,w__8070 ,w__7770);
  or g__10158(w__8153 ,w__8011 ,w__7794);
  or g__10159(w__8152 ,w__7997 ,w__7764);
  or g__10160(w__8151 ,w__7995 ,w__7833);
  or g__10161(w__8150 ,w__8102 ,w__7767);
  or g__10162(w__8149 ,w__8090 ,w__7829);
  or g__10163(w__8148 ,w__8061 ,w__7803);
  or g__10164(w__8147 ,w__8098 ,w__7821);
  or g__10165(w__8146 ,w__7993 ,w__7788);
  or g__10166(w__8145 ,w__8084 ,w__7791);
  or g__10167(w__8144 ,w__7994 ,w__7797);
  or g__10168(w__8143 ,w__8021 ,w__7761);
  or g__10169(w__8142 ,w__8073 ,w__7818);
  or g__10170(w__8141 ,w__7969 ,w__7770);
  or g__10171(w__8140 ,w__8006 ,w__7809);
  or g__10172(w__8139 ,w__8003 ,w__7806);
  or g__10173(w__8138 ,w__8000 ,w__7827);
  or g__10174(w__8137 ,w__8082 ,w__7815);
  or g__10175(w__8136 ,w__8097 ,w__7785);
  or g__10176(w__8135 ,w__8001 ,w__7794);
  or g__10177(w__8134 ,w__7772 ,w__8091);
  or g__10178(w__8133 ,w__7781 ,w__8107);
  or g__10179(w__8132 ,w__7781 ,w__8058);
  or g__10180(w__8131 ,w__7773 ,w__8111);
  or g__10181(w__8130 ,w__7776 ,w__8108);
  or g__10182(w__8129 ,w__7772 ,w__8109);
  or g__10183(w__8128 ,w__7775 ,w__8104);
  or g__10184(w__8127 ,w__7778 ,w__8081);
  or g__10185(w__8126 ,w__7778 ,w__8110);
  or g__10186(w__8125 ,w__7775 ,w__8087);
  or g__10187(w__8124 ,w__7782 ,w__8076);
  or g__10188(w__8123 ,w__7776 ,w__8106);
  or g__10189(w__8122 ,w__7779 ,w__8085);
  or g__10190(w__8121 ,w__7773 ,w__8094);
  or g__10191(w__8120 ,w__7782 ,w__8093);
  or g__10192(w__8119 ,w__7659 ,w__8045);
  or g__10193(w__8118 ,w__7888 ,w__8048);
  or g__10194(w__8117 ,w__7886 ,w__8049);
  or g__10195(w__8116 ,w__7885 ,w__8047);
  or g__10196(w__8115 ,w__7887 ,w__8043);
  or g__10197(w__8114 ,w__7884 ,w__8044);
  or g__10198(w__8113 ,w__7872 ,w__8046);
  nor g__10199(w__8112 ,w__7830 ,w__7525);
  and g__10200(w__8192 ,in17[13] ,w__7691);
  and g__10201(w__8190 ,in17[7] ,w__7689);
  and g__10202(w__8188 ,in17[3] ,w__7682);
  and g__10203(w__8187 ,in17[15] ,w__7690);
  and g__10204(w__8185 ,in17[9] ,w__7693);
  and g__10205(w__8183 ,in17[11] ,w__7687);
  and g__10206(w__8181 ,in17[5] ,w__7683);
  and g__10207(w__8179 ,in16[0] ,w__7697);
  or g__10208(w__8178 ,w__7673 ,w__7791);
  or g__10209(w__8177 ,w__7673 ,w__7779);
  or g__10210(w__8176 ,w__7889 ,w__7818);
  or g__10211(w__8175 ,w__7672 ,w__7803);
  or g__10212(w__8174 ,w__7672 ,w__7767);
  or g__10213(w__8173 ,w__8040 ,w__7685);
  or g__10214(w__8172 ,w__8035 ,w__7694);
  or g__10215(w__8171 ,w__8033 ,w__7684);
  or g__10216(w__8170 ,w__7948 ,w__7696);
  or g__10217(w__8169 ,w__8036 ,w__7692);
  or g__10218(w__8168 ,w__7951 ,w__7686);
  not g__10219(w__8055 ,w__7689);
  not g__10220(w__8054 ,w__7694);
  not g__10221(w__8052 ,w__7688);
  not g__10222(w__8051 ,w__7690);
  nor g__10223(w__8049 ,w__7737 ,w__7935);
  nor g__10224(w__8048 ,w__7873 ,w__7898);
  nor g__10225(w__8047 ,w__7735 ,w__7904);
  nor g__10226(w__8046 ,w__7733 ,w__7937);
  nor g__10227(w__8045 ,w__7731 ,w__7899);
  nor g__10228(w__8044 ,w__7739 ,w__7924);
  nor g__10229(w__8043 ,w__7741 ,w__7929);
  or g__10230(w__8042 ,w__7920 ,w__7909);
  xnor g__10231(w__8040 ,in17[13] ,in17[12]);
  xnor g__10232(w__8039 ,in16[0] ,in17[3]);
  nor g__10233(w__8038 ,w__13308 ,w__7743);
  xnor g__10234(w__8037 ,in16[0] ,in17[9]);
  xnor g__10235(w__8036 ,in17[9] ,in17[8]);
  xnor g__10236(w__8035 ,in17[7] ,in17[6]);
  xnor g__10237(w__8034 ,in16[0] ,in17[5]);
  xnor g__10238(w__8033 ,in17[3] ,in17[2]);
  or g__10239(w__8111 ,w__7841 ,w__7928);
  or g__10240(w__8110 ,w__7916 ,w__7925);
  or g__10241(w__8109 ,w__7842 ,w__7938);
  or g__10242(w__8108 ,w__7852 ,w__7933);
  or g__10243(w__8107 ,w__7844 ,w__7930);
  or g__10244(w__8106 ,w__7851 ,w__7926);
  xnor g__10245(w__8105 ,in16[4] ,in17[13]);
  or g__10246(w__8104 ,w__7849 ,w__7901);
  xnor g__10247(w__8103 ,in16[1] ,in17[13]);
  xnor g__10248(w__8102 ,in16[4] ,in17[11]);
  xnor g__10249(w__8101 ,in16[6] ,in17[7]);
  xnor g__10250(w__8100 ,in16[13] ,in17[5]);
  xnor g__10251(w__8099 ,in16[4] ,in17[3]);
  xnor g__10252(w__8098 ,in16[2] ,in17[3]);
  xnor g__10253(w__8097 ,in16[7] ,in17[7]);
  xnor g__10254(w__8096 ,in16[9] ,in17[11]);
  xnor g__10255(w__8095 ,in16[10] ,in17[5]);
  or g__10256(w__8094 ,w__7843 ,w__7934);
  or g__10257(w__8093 ,w__7850 ,w__7902);
  xnor g__10258(w__8092 ,in16[5] ,in17[5]);
  or g__10259(w__8091 ,w__7848 ,w__7906);
  xnor g__10260(w__8090 ,in16[6] ,in17[3]);
  xnor g__10261(w__8089 ,in16[3] ,in17[7]);
  xnor g__10262(w__8088 ,in16[15] ,in17[5]);
  or g__10263(w__8087 ,w__7846 ,w__7927);
  xnor g__10264(w__8086 ,in16[3] ,in17[9]);
  or g__10265(w__8085 ,w__7845 ,w__7931);
  xnor g__10266(w__8084 ,in16[10] ,in17[7]);
  xnor g__10267(w__8083 ,in16[11] ,in17[3]);
  xnor g__10268(w__8082 ,in16[8] ,in17[9]);
  or g__10269(w__8081 ,w__7847 ,w__7936);
  xnor g__10270(w__8080 ,in16[15] ,in17[7]);
  xnor g__10271(w__8079 ,in16[11] ,in17[7]);
  xnor g__10272(w__8078 ,in16[10] ,in17[13]);
  xnor g__10273(w__8077 ,in16[1] ,in17[5]);
  xnor g__10274(w__8076 ,in16[15] ,in17[15]);
  xnor g__10275(w__8075 ,in16[2] ,in17[11]);
  xnor g__10276(w__8074 ,in16[3] ,in17[11]);
  xnor g__10277(w__8073 ,in16[14] ,in17[9]);
  xnor g__10278(w__8072 ,in16[12] ,in17[9]);
  xnor g__10279(w__8071 ,in16[12] ,in17[7]);
  xnor g__10280(w__8070 ,in16[8] ,in17[11]);
  xnor g__10281(w__8069 ,in16[11] ,in17[5]);
  xnor g__10282(w__8068 ,in16[8] ,in17[13]);
  xnor g__10283(w__8067 ,in16[1] ,in17[11]);
  xnor g__10284(w__8066 ,in16[2] ,in17[9]);
  xnor g__10285(w__8065 ,in16[8] ,in17[5]);
  xnor g__10286(w__8064 ,in16[13] ,in17[11]);
  xnor g__10287(w__8063 ,in16[4] ,in17[9]);
  xnor g__10288(w__8062 ,in16[5] ,in17[9]);
  xnor g__10289(w__8061 ,in16[2] ,in17[13]);
  xnor g__10290(w__8060 ,in16[9] ,in17[9]);
  xnor g__10291(w__8059 ,in16[13] ,in17[9]);
  or g__10292(w__8058 ,w__7727 ,w__7910);
  xnor g__10293(w__8057 ,in16[15] ,in17[13]);
  xnor g__10294(w__8056 ,in16[7] ,in17[13]);
  xnor g__10295(w__8053 ,w__7741 ,in17[6]);
  xnor g__10296(w__8050 ,w__7731 ,in17[14]);
  not g__10297(w__7968 ,w__7687);
  not g__10298(w__7967 ,w__7686);
  not g__10299(w__7965 ,w__7697);
  not g__10300(w__7963 ,w__7683);
  not g__10301(w__7962 ,w__7696);
  not g__10302(w__7961 ,w__7682);
  not g__10303(w__7960 ,w__7684);
  not g__10304(w__7958 ,w__7693);
  not g__10305(w__7957 ,w__7692);
  not g__10306(w__7955 ,w__7691);
  not g__10307(w__7954 ,w__7685);
  xnor g__10308(w__7952 ,in17[15] ,in17[14]);
  xnor g__10309(w__7951 ,in17[11] ,in17[10]);
  xnor g__10310(w__7950 ,in16[0] ,in17[11]);
  xnor g__10311(w__7949 ,in16[0] ,in17[13]);
  xnor g__10312(w__7948 ,in17[5] ,in17[4]);
  xnor g__10313(w__7947 ,in16[0] ,in17[1]);
  xnor g__10314(w__7946 ,in16[0] ,in17[7]);
  xnor g__10315(w__8032 ,in16[7] ,in17[3]);
  xnor g__10316(w__8031 ,in16[11] ,in17[9]);
  xnor g__10317(w__8030 ,in16[15] ,in17[3]);
  xnor g__10318(w__8029 ,in16[4] ,in17[7]);
  xnor g__10319(w__8028 ,in16[12] ,in17[5]);
  xnor g__10320(w__8027 ,in16[13] ,in17[7]);
  xnor g__10321(w__8026 ,in16[14] ,in17[13]);
  xnor g__10322(w__8025 ,in16[5] ,in17[11]);
  xnor g__10323(w__8024 ,in16[9] ,in17[3]);
  xnor g__10324(w__8023 ,in16[15] ,in17[11]);
  xnor g__10325(w__8022 ,in16[5] ,in17[7]);
  xnor g__10326(w__8021 ,in16[14] ,in17[11]);
  xnor g__10327(w__8020 ,in16[1] ,in17[9]);
  xnor g__10328(w__8019 ,in16[6] ,in17[5]);
  xnor g__10329(w__8018 ,in16[11] ,in17[11]);
  xnor g__10330(w__8017 ,in16[14] ,in17[3]);
  xnor g__10331(w__8016 ,in16[3] ,in17[5]);
  xnor g__10332(w__8015 ,in16[11] ,in17[13]);
  xnor g__10333(w__8014 ,in16[12] ,in17[11]);
  xnor g__10334(w__8013 ,in16[3] ,in17[3]);
  xnor g__10335(w__8012 ,in16[3] ,in17[13]);
  xnor g__10336(w__8011 ,in16[14] ,in17[7]);
  xnor g__10337(w__8010 ,in16[4] ,in17[5]);
  xnor g__10338(w__8009 ,in16[13] ,in17[13]);
  xnor g__10339(w__8008 ,in16[1] ,in17[3]);
  xnor g__10340(w__8007 ,in16[9] ,in17[5]);
  xnor g__10341(w__8006 ,in16[7] ,in17[9]);
  xnor g__10342(w__8005 ,in16[12] ,in17[13]);
  xnor g__10343(w__8004 ,in16[8] ,in17[3]);
  xnor g__10344(w__8003 ,in16[5] ,in17[13]);
  xnor g__10345(w__8002 ,in16[5] ,in17[3]);
  xnor g__10346(w__8001 ,in16[8] ,in17[7]);
  xnor g__10347(w__8000 ,in16[13] ,in17[3]);
  xnor g__10348(w__7999 ,in16[1] ,in17[7]);
  xnor g__10349(w__7998 ,in16[6] ,in17[9]);
  xnor g__10350(w__7997 ,in16[10] ,in17[11]);
  xnor g__10351(w__7996 ,in16[10] ,in17[9]);
  xnor g__10352(w__7995 ,in16[14] ,in17[5]);
  xnor g__10353(w__7994 ,in16[9] ,in17[13]);
  xnor g__10354(w__7993 ,in16[9] ,in17[7]);
  xnor g__10355(w__7992 ,in16[2] ,in17[5]);
  xnor g__10356(w__7991 ,in16[6] ,in17[13]);
  xnor g__10357(w__7990 ,in16[12] ,in17[3]);
  xnor g__10358(w__7989 ,in16[6] ,in17[11]);
  xnor g__10359(w__7988 ,in16[15] ,in17[9]);
  xnor g__10360(w__7987 ,in16[2] ,in17[7]);
  xnor g__10361(w__7986 ,in16[10] ,in17[3]);
  xnor g__10362(w__7985 ,in16[4] ,in17[1]);
  xnor g__10363(w__7984 ,in16[2] ,in17[1]);
  xnor g__10364(w__7983 ,in16[9] ,in17[1]);
  xnor g__10365(w__7982 ,in16[3] ,in17[1]);
  xnor g__10366(w__7981 ,in16[5] ,in17[1]);
  xnor g__10367(w__7980 ,in16[8] ,in17[1]);
  xnor g__10368(w__7979 ,in16[7] ,in17[1]);
  xnor g__10369(w__7978 ,in16[11] ,in17[1]);
  xnor g__10370(w__7977 ,in16[14] ,in17[1]);
  xnor g__10371(w__7976 ,in16[12] ,in17[1]);
  xnor g__10372(w__7975 ,in16[7] ,in17[5]);
  xnor g__10373(w__7974 ,in16[10] ,in17[1]);
  xnor g__10374(w__7973 ,in16[1] ,in17[1]);
  xnor g__10375(w__7972 ,in16[6] ,in17[1]);
  xnor g__10376(w__7971 ,in16[13] ,in17[1]);
  xnor g__10377(w__7970 ,in16[15] ,in17[1]);
  xnor g__10378(w__7969 ,in16[7] ,in17[11]);
  xnor g__10379(w__7966 ,w__7739 ,in17[10]);
  xnor g__10380(w__7964 ,w__7737 ,in17[4]);
  xnor g__10381(w__7959 ,w__7743 ,in17[2]);
  xnor g__10382(w__7956 ,w__7735 ,in17[8]);
  xnor g__10383(w__7953 ,w__7733 ,in17[12]);
  nor g__10384(w__7938 ,in16[2] ,in17[15]);
  nor g__10385(w__7937 ,in16[0] ,in17[12]);
  nor g__10386(w__7936 ,in16[4] ,in17[15]);
  nor g__10387(w__7935 ,in16[0] ,in17[4]);
  nor g__10388(w__7934 ,in16[5] ,in17[15]);
  nor g__10389(w__7933 ,in16[9] ,in17[15]);
  and g__10390(w__7932 ,in16[0] ,in17[6]);
  nor g__10391(w__7931 ,in16[13] ,in17[15]);
  nor g__10392(w__7930 ,in16[8] ,in17[15]);
  nor g__10393(w__7929 ,in16[0] ,in17[6]);
  nor g__10394(w__7928 ,in16[1] ,in17[15]);
  nor g__10395(w__7927 ,in16[3] ,in17[15]);
  nor g__10396(w__7926 ,in16[7] ,in17[15]);
  nor g__10397(w__7925 ,in16[6] ,in17[15]);
  nor g__10398(w__7924 ,in16[0] ,in17[10]);
  or g__10399(w__7923 ,w__7893 ,w__7556);
  or g__10400(w__7945 ,w__7895 ,w__7580);
  or g__10401(w__7944 ,w__7896 ,w__7658);
  or g__10402(w__7943 ,w__7878 ,w__7628);
  or g__10403(w__7942 ,w__7882 ,w__7557);
  or g__10404(w__7941 ,w__7891 ,w__7581);
  or g__10405(w__7940 ,w__7890 ,w__7542);
  or g__10406(w__7939 ,w__7881 ,w__7628);
  not g__10407(w__7919 ,w__7920);
  not g__10408(w__7916 ,w__7917);
  not g__10409(w__7911 ,w__7912);
  nor g__10410(w__7910 ,in16[14] ,in17[15]);
  nor g__10411(w__7909 ,in16[0] ,in17[15]);
  and g__10412(w__7908 ,in16[0] ,in17[14]);
  and g__10413(w__7907 ,in16[0] ,in17[2]);
  nor g__10414(w__7906 ,in16[12] ,in17[15]);
  and g__10415(w__7905 ,in16[0] ,in17[10]);
  nor g__10416(w__7904 ,in16[0] ,in17[8]);
  and g__10417(w__7903 ,in16[0] ,in17[12]);
  nor g__10418(w__7902 ,in16[10] ,in17[15]);
  nor g__10419(w__7901 ,in16[11] ,in17[15]);
  and g__10420(w__7900 ,in16[0] ,in17[8]);
  nor g__10421(w__7899 ,in16[0] ,in17[14]);
  nor g__10422(w__7898 ,in16[0] ,in17[2]);
  and g__10423(w__7897 ,in16[0] ,in17[4]);
  and g__10424(w__13308 ,in16[0] ,in17[0]);
  and g__10425(w__7922 ,in17[1] ,in17[0]);
  or g__10426(w__7921 ,w__7879 ,w__7556);
  and g__10427(w__7920 ,in16[0] ,in17[15]);
  or g__10428(w__7918 ,w__7877 ,w__7580);
  or g__10429(w__7917 ,w__7892 ,w__7658);
  or g__10430(w__7915 ,w__7883 ,w__7581);
  or g__10431(w__7914 ,w__7876 ,w__7557);
  or g__10432(w__7913 ,w__7894 ,w__7542);
  or g__10433(w__7912 ,w__7880 ,w__7629);
  not g__10434(w__7896 ,in16[7]);
  not g__10435(w__7895 ,in16[9]);
  not g__10436(w__7894 ,in16[1]);
  not g__10437(w__7893 ,in16[15]);
  not g__10438(w__7892 ,in16[6]);
  not g__10439(w__7891 ,in16[12]);
  not g__10440(w__7890 ,in16[4]);
  not g__10441(w__7889 ,in16[0]);
  not g__10442(w__7888 ,in17[3]);
  not g__10443(w__7887 ,in17[7]);
  not g__10444(w__7886 ,in17[5]);
  not g__10445(w__7885 ,in17[9]);
  not g__10446(w__7884 ,in17[11]);
  not g__10447(w__7883 ,in16[5]);
  not g__10448(w__7882 ,in16[11]);
  not g__10449(w__7881 ,in16[3]);
  not g__10450(w__7880 ,in16[14]);
  not g__10451(w__7879 ,in16[13]);
  not g__10452(w__7878 ,in16[10]);
  not g__10453(w__7877 ,in16[8]);
  not g__10454(w__7876 ,in16[2]);
  not g__10455(w__7875 ,in17[0]);
  not g__10456(w__7874 ,in17[15]);
  not g__10457(w__7873 ,in17[1]);
  not g__10458(w__7872 ,in17[13]);
  not g__10459(w__7526 ,w__7840);
  not g__10460(w__7840 ,w__7889);
  not g__10461(w__7839 ,w__7837);
  not g__10462(w__7838 ,w__7837);
  not g__10463(w__7837 ,w__7859);
  not g__10464(w__7836 ,w__7834);
  not g__10465(w__7835 ,w__7834);
  not g__10466(w__7834 ,w__7965);
  not g__10467(w__7833 ,w__7831);
  not g__10468(w__7832 ,w__7831);
  not g__10469(w__7831 ,w__7962);
  not g__10470(w__7830 ,w__7828);
  not g__10471(w__7829 ,w__7828);
  not g__10472(w__7828 ,w__7960);
  not g__10473(w__7827 ,w__7825);
  not g__10474(w__7826 ,w__7825);
  not g__10475(w__7825 ,w__7961);
  not g__10476(w__7824 ,w__7822);
  not g__10477(w__7823 ,w__7822);
  not g__10478(w__7822 ,w__7858);
  not g__10479(w__7821 ,w__7819);
  not g__10480(w__7820 ,w__7819);
  not g__10481(w__7819 ,w__7857);
  not g__10482(w__7818 ,w__7816);
  not g__10483(w__7817 ,w__7816);
  not g__10484(w__7816 ,w__7957);
  not g__10485(w__7815 ,w__7813);
  not g__10486(w__7814 ,w__7813);
  not g__10487(w__7813 ,w__7958);
  not g__10488(w__7812 ,w__7810);
  not g__10489(w__7811 ,w__7810);
  not g__10490(w__7810 ,w__7856);
  not g__10491(w__7809 ,w__7807);
  not g__10492(w__7808 ,w__7807);
  not g__10493(w__7807 ,w__7855);
  not g__10494(w__7806 ,w__7804);
  not g__10495(w__7805 ,w__7804);
  not g__10496(w__7804 ,w__7955);
  not g__10497(w__7803 ,w__7801);
  not g__10498(w__7802 ,w__7801);
  not g__10499(w__7801 ,w__7954);
  not g__10500(w__7800 ,w__7798);
  not g__10501(w__7799 ,w__7798);
  not g__10502(w__7798 ,w__7854);
  not g__10503(w__7797 ,w__7795);
  not g__10504(w__7796 ,w__7795);
  not g__10505(w__7795 ,w__7853);
  not g__10506(w__7794 ,w__7792);
  not g__10507(w__7793 ,w__7792);
  not g__10508(w__7792 ,w__8055);
  not g__10509(w__7791 ,w__7789);
  not g__10510(w__7790 ,w__7789);
  not g__10511(w__7789 ,w__8054);
  not g__10512(w__7788 ,w__7786);
  not g__10513(w__7787 ,w__7786);
  not g__10514(w__7786 ,w__7865);
  not g__10515(w__7785 ,w__7783);
  not g__10516(w__7784 ,w__7783);
  not g__10517(w__7783 ,w__7864);
  not g__10518(w__7782 ,w__7780);
  not g__10519(w__7781 ,w__7780);
  not g__10520(w__7780 ,w__8052);
  not g__10521(w__7779 ,w__7777);
  not g__10522(w__7778 ,w__7777);
  not g__10523(w__7777 ,w__8051);
  not g__10524(w__7776 ,w__7774);
  not g__10525(w__7775 ,w__7774);
  not g__10526(w__7774 ,w__7863);
  not g__10527(w__7773 ,w__7771);
  not g__10528(w__7772 ,w__7771);
  not g__10529(w__7771 ,w__7862);
  not g__10530(w__7770 ,w__7768);
  not g__10531(w__7769 ,w__7768);
  not g__10532(w__7768 ,w__7968);
  not g__10533(w__7767 ,w__7765);
  not g__10534(w__7766 ,w__7765);
  not g__10535(w__7765 ,w__7967);
  not g__10536(w__7764 ,w__7762);
  not g__10537(w__7763 ,w__7762);
  not g__10538(w__7762 ,w__7861);
  not g__10539(w__7761 ,w__7759);
  not g__10540(w__7760 ,w__7759);
  not g__10541(w__7759 ,w__7860);
  not g__10542(w__7758 ,w__7848);
  not g__10543(w__7848 ,w__7941);
  not g__10544(w__7757 ,w__7845);
  not g__10545(w__7845 ,w__7921);
  not g__10546(w__7756 ,w__7852);
  not g__10547(w__7852 ,w__7945);
  not g__10548(w__7755 ,w__7849);
  not g__10549(w__7849 ,w__7942);
  not g__10550(w__7754 ,w__7850);
  not g__10551(w__7850 ,w__7943);
  not g__10552(w__7753 ,w__7846);
  not g__10553(w__7846 ,w__7939);
  not g__10554(w__7752 ,w__7844);
  not g__10555(w__7844 ,w__7918);
  not g__10556(w__7751 ,w__7842);
  not g__10557(w__7842 ,w__7914);
  not g__10558(w__7750 ,w__7843);
  not g__10559(w__7843 ,w__7915);
  not g__10560(w__7749 ,w__7841);
  not g__10561(w__7841 ,w__7913);
  not g__10562(w__7748 ,w__7847);
  not g__10563(w__7847 ,w__7940);
  not g__10564(w__7747 ,w__7851);
  not g__10565(w__7851 ,w__7944);
  not g__10566(w__7746 ,w__7745);
  not g__10567(w__7745 ,w__8500);
  not g__10568(w__7744 ,w__7866);
  not g__10569(w__7866 ,w__8503);
  not g__10570(w__7743 ,w__7742);
  not g__10571(w__7742 ,w__7873);
  not g__10572(w__7741 ,w__7740);
  not g__10573(w__7740 ,w__7886);
  not g__10574(w__7739 ,w__7738);
  not g__10575(w__7738 ,w__7885);
  not g__10576(w__7737 ,w__7736);
  not g__10577(w__7736 ,w__7888);
  not g__10578(w__7735 ,w__7734);
  not g__10579(w__7734 ,w__7887);
  not g__10580(w__7733 ,w__7732);
  not g__10581(w__7732 ,w__7884);
  not g__10582(w__7731 ,w__7730);
  not g__10583(w__7730 ,w__7872);
  not g__10584(w__7729 ,w__7728);
  not g__10585(w__7728 ,w__7963);
  buf g__10586(w__13306 ,w__8112);
  buf g__10587(w__13307 ,w__8038);
  not g__10588(w__7727 ,w__7726);
  not g__10589(w__7726 ,w__7911);
  not g__10590(w__7725 ,w__7724);
  not g__10591(w__7724 ,w__8501);
  not g__10592(w__7723 ,w__7868);
  not g__10593(w__7868 ,w__8857);
  not g__10594(w__7722 ,w__7869);
  not g__10595(w__7869 ,w__8873);
  not g__10596(w__7721 ,w__7870);
  not g__10597(w__7870 ,w__9113);
  not g__10598(w__7720 ,w__7867);
  not g__10599(w__7867 ,w__8856);
  not g__10600(w__7719 ,w__7871);
  not g__10601(w__7871 ,w__9114);
  not g__10602(w__7718 ,w__7717);
  not g__10603(w__7717 ,w__8266);
  not g__10604(w__7716 ,w__7715);
  not g__10605(w__7715 ,w__8173);
  not g__10606(w__7714 ,w__7713);
  not g__10607(w__7713 ,w__8172);
  not g__10608(w__7712 ,w__7711);
  not g__10609(w__7711 ,w__8169);
  not g__10610(w__7710 ,w__7709);
  not g__10611(w__7709 ,w__8168);
  not g__10612(w__7708 ,w__7707);
  not g__10613(w__7707 ,w__8171);
  not g__10614(w__7706 ,w__7705);
  not g__10615(w__7705 ,w__8170);
  not g__10616(w__7704 ,w__7703);
  not g__10617(w__7703 ,w__7874);
  not g__10618(w__7702 ,w__7701);
  not g__10619(w__7701 ,w__8267);
  not g__10620(w__7700 ,w__7698);
  not g__10621(w__7699 ,w__7698);
  not g__10622(w__7698 ,w__7875);
  not g__10623(w__7697 ,w__7695);
  not g__10624(w__7696 ,w__7695);
  not g__10625(w__7695 ,w__7964);
  not g__10626(w__7694 ,w__7864);
  not g__10627(w__7864 ,w__8053);
  not g__10628(w__7693 ,w__7856);
  not g__10629(w__7856 ,w__7956);
  not g__10630(w__7692 ,w__7855);
  not g__10631(w__7855 ,w__7956);
  not g__10632(w__7691 ,w__7854);
  not g__10633(w__7854 ,w__7953);
  not g__10634(w__7690 ,w__7862);
  not g__10635(w__7862 ,w__8050);
  not g__10636(w__7689 ,w__7865);
  not g__10637(w__7865 ,w__8053);
  not g__10638(w__7688 ,w__7863);
  not g__10639(w__7863 ,w__8050);
  not g__10640(w__7687 ,w__7861);
  not g__10641(w__7861 ,w__7966);
  not g__10642(w__7686 ,w__7860);
  not g__10643(w__7860 ,w__7966);
  not g__10644(w__7685 ,w__7853);
  not g__10645(w__7853 ,w__7953);
  not g__10646(w__7684 ,w__7857);
  not g__10647(w__7857 ,w__7959);
  not g__10648(w__7683 ,w__7859);
  not g__10649(w__7859 ,w__7964);
  not g__10650(w__7682 ,w__7858);
  not g__10651(w__7858 ,w__7959);
  not g__10652(w__7681 ,w__7680);
  not g__10653(w__7680 ,w__8420);
  not g__10654(w__7679 ,w__7678);
  not g__10655(w__7678 ,w__8497);
  not g__10656(w__7677 ,w__7676);
  not g__10657(w__7676 ,w__8422);
  not g__10658(w__7675 ,w__7674);
  not g__10659(w__7674 ,w__8418);
  not g__10660(w__7525 ,w__7534);
  not g__10661(w__7673 ,w__7534);
  not g__10662(w__7534 ,w__7526);
  not g__10663(w__7672 ,w__7840);
  not g__10664(w__7671 ,w__7669);
  not g__10665(w__7670 ,w__7669);
  not g__10666(w__7669 ,w__8266);
  not g__10667(w__7668 ,w__7666);
  not g__10668(w__7667 ,w__7666);
  not g__10669(w__7666 ,w__8267);
  not g__10670(w__7665 ,w__7663);
  not g__10671(w__7664 ,w__7663);
  not g__10672(w__7663 ,w__8173);
  not g__10673(w__7662 ,w__7660);
  not g__10674(w__7661 ,w__7660);
  not g__10675(w__7660 ,w__8170);
  not g__10676(w__7659 ,w__7657);
  not g__10677(w__7658 ,w__7657);
  not g__10678(w__7657 ,w__7874);
  not g__10679(w__7656 ,w__7654);
  not g__10680(w__7655 ,w__7654);
  not g__10681(w__7654 ,w__8172);
  not g__10682(w__7653 ,w__7651);
  not g__10683(w__7652 ,w__7651);
  not g__10684(w__7651 ,w__8171);
  not g__10685(w__7650 ,w__7648);
  not g__10686(w__7649 ,w__7648);
  not g__10687(w__7648 ,w__8169);
  not g__10688(w__7647 ,w__7645);
  not g__10689(w__7646 ,w__7645);
  not g__10690(w__7645 ,w__8168);
  not g__10691(w__7644 ,w__7642);
  not g__10692(w__7643 ,w__7642);
  not g__10693(w__7642 ,w__8266);
  not g__10694(w__7641 ,w__7639);
  not g__10695(w__7640 ,w__7639);
  not g__10696(w__7639 ,w__7718);
  not g__10697(w__7638 ,w__7636);
  not g__10698(w__7637 ,w__7636);
  not g__10699(w__7636 ,w__7708);
  not g__10700(w__7635 ,w__7633);
  not g__10701(w__7634 ,w__7633);
  not g__10702(w__7633 ,w__7710);
  not g__10703(w__7632 ,w__7630);
  not g__10704(w__7631 ,w__7630);
  not g__10705(w__7630 ,w__7706);
  not g__10706(w__7629 ,w__7627);
  not g__10707(w__7628 ,w__7627);
  not g__10708(w__7627 ,w__7704);
  not g__10709(w__7626 ,w__7624);
  not g__10710(w__7625 ,w__7624);
  not g__10711(w__7624 ,w__7700);
  not g__10712(w__7623 ,w__7621);
  not g__10713(w__7622 ,w__7621);
  not g__10714(w__7621 ,w__8171);
  not g__10715(w__7620 ,w__7618);
  not g__10716(w__7619 ,w__7618);
  not g__10717(w__7618 ,w__7718);
  not g__10718(w__7617 ,w__7615);
  not g__10719(w__7616 ,w__7615);
  not g__10720(w__7615 ,w__7875);
  not g__10721(w__7614 ,w__7612);
  not g__10722(w__7613 ,w__7612);
  not g__10723(w__7612 ,w__7875);
  not g__10724(w__7611 ,w__7609);
  not g__10725(w__7610 ,w__7609);
  not g__10726(w__7609 ,w__7716);
  not g__10727(w__7608 ,w__7606);
  not g__10728(w__7607 ,w__7606);
  not g__10729(w__7606 ,w__7714);
  not g__10730(w__7605 ,w__7603);
  not g__10731(w__7604 ,w__7603);
  not g__10732(w__7603 ,w__7712);
  not g__10733(w__7602 ,w__7600);
  not g__10734(w__7601 ,w__7600);
  not g__10735(w__7600 ,w__8267);
  not g__10736(w__7599 ,w__7597);
  not g__10737(w__7598 ,w__7597);
  not g__10738(w__7597 ,w__7702);
  not g__10739(w__7596 ,w__7594);
  not g__10740(w__7595 ,w__7594);
  not g__10741(w__7594 ,w__7702);
  not g__10742(w__7593 ,w__7591);
  not g__10743(w__7592 ,w__7591);
  not g__10744(w__7591 ,w__8170);
  not g__10745(w__7590 ,w__7588);
  not g__10746(w__7589 ,w__7588);
  not g__10747(w__7588 ,w__7710);
  not g__10748(w__7587 ,w__7585);
  not g__10749(w__7586 ,w__7585);
  not g__10750(w__7585 ,w__8169);
  not g__10751(w__7584 ,w__7582);
  not g__10752(w__7583 ,w__7582);
  not g__10753(w__7582 ,w__7706);
  not g__10754(w__7581 ,w__7579);
  not g__10755(w__7580 ,w__7579);
  not g__10756(w__7579 ,w__7704);
  not g__10757(w__7578 ,w__7576);
  not g__10758(w__7577 ,w__7576);
  not g__10759(w__7576 ,w__8168);
  not g__10760(w__7575 ,w__7573);
  not g__10761(w__7574 ,w__7573);
  not g__10762(w__7573 ,w__8172);
  not g__10763(w__7572 ,w__7570);
  not g__10764(w__7571 ,w__7570);
  not g__10765(w__7570 ,w__7708);
  not g__10766(w__7569 ,w__7567);
  not g__10767(w__7568 ,w__7567);
  not g__10768(w__7567 ,w__7712);
  not g__10769(w__7566 ,w__7564);
  not g__10770(w__7565 ,w__7564);
  not g__10771(w__7564 ,w__7716);
  not g__10772(w__7563 ,w__7561);
  not g__10773(w__7562 ,w__7561);
  not g__10774(w__7561 ,w__8173);
  not g__10775(w__7560 ,w__7558);
  not g__10776(w__7559 ,w__7558);
  not g__10777(w__7558 ,w__7714);
  not g__10778(w__7557 ,w__7555);
  not g__10779(w__7556 ,w__7555);
  not g__10780(w__7555 ,w__7874);
  not g__10781(w__7554 ,w__7553);
  not g__10782(w__7553 ,w__7699);
  not g__10783(w__7552 ,w__7551);
  not g__10784(w__7551 ,w__7670);
  not g__10785(w__7550 ,w__7549);
  not g__10786(w__7549 ,w__7647);
  not g__10787(w__7548 ,w__7547);
  not g__10788(w__7547 ,w__7650);
  not g__10789(w__7546 ,w__7545);
  not g__10790(w__7545 ,w__7653);
  not g__10791(w__7544 ,w__7543);
  not g__10792(w__7543 ,w__7656);
  not g__10793(w__7542 ,w__7541);
  not g__10794(w__7541 ,w__7659);
  not g__10795(w__7540 ,w__7539);
  not g__10796(w__7539 ,w__7662);
  not g__10797(w__7538 ,w__7537);
  not g__10798(w__7537 ,w__7665);
  not g__10799(w__7536 ,w__7535);
  not g__10800(w__7535 ,w__7668);
  xor g__10801(w__7533 ,w__9115 ,w__9210);
  xor g__10802(w__13283 ,w__9091 ,w__9180);
  xor g__10803(w__7532 ,w__9073 ,w__9094);
  xor g__10804(w__7531 ,w__8732 ,w__8810);
  xor g__10805(w__7530 ,w__8726 ,w__7680);
  xor g__10806(w__7529 ,w__8836 ,w__7678);
  xor g__10807(w__7528 ,w__8715 ,w__7676);
  xor g__10808(w__7527 ,w__8823 ,w__7674);
  xnor g__10809(w__13224 ,w__10907 ,w__10942);
  xnor g__10810(w__13225 ,w__10910 ,w__9242);
  xnor g__10811(w__13227 ,w__10920 ,w__10934);
  xnor g__10812(w__13226 ,w__10916 ,w__10933);
  xnor g__10813(w__13223 ,w__10900 ,w__10935);
  or g__10814(w__13163 ,w__10905 ,w__10941);
  or g__10815(w__13162 ,w__10928 ,w__10940);
  or g__10816(w__13159 ,w__10923 ,w__10937);
  or g__10817(w__13158 ,w__10932 ,w__10939);
  or g__10818(w__13160 ,w__10921 ,w__10938);
  or g__10819(w__13161 ,w__10930 ,w__10936);
  xnor g__10820(w__13222 ,w__10886 ,w__10914);
  xnor g__10821(w__13228 ,w__10917 ,w__10913);
  xnor g__10822(w__13221 ,w__10888 ,w__10912);
  xnor g__10823(w__10942 ,w__10802 ,w__10918);
  and g__10824(w__10941 ,w__10894 ,w__10917);
  and g__10825(w__10940 ,w__10927 ,w__10920);
  or g__10826(w__13156 ,w__10902 ,w__10922);
  and g__10827(w__10939 ,w__10900 ,w__10924);
  nor g__10828(w__10938 ,w__10931 ,w__10919);
  or g__10829(w__13164 ,w__10884 ,w__10925);
  or g__10830(w__13157 ,w__10904 ,w__10926);
  and g__10831(w__10937 ,w__10915 ,w__10918);
  xnor g__10832(w__13229 ,w__10899 ,w__10891);
  xnor g__10833(w__13220 ,w__10887 ,w__10890);
  xnor g__10834(w__13230 ,w__10805 ,w__10892);
  nor g__10835(w__10936 ,w__10929 ,w__10916);
  xnor g__10836(w__10935 ,w__10896 ,w__10822);
  xnor g__10837(w__10934 ,w__10909 ,w__10823);
  xnor g__10838(w__10933 ,w__10897 ,w__10911);
  nor g__10839(w__10932 ,w__9430 ,w__10896);
  and g__10840(w__10931 ,w__10824 ,w__10910);
  nor g__10841(w__10930 ,w__10898 ,w__10911);
  and g__10842(w__10929 ,w__10898 ,w__10911);
  nor g__10843(w__10928 ,w__9428 ,w__10909);
  or g__10844(w__10927 ,w__9580 ,w__10908);
  nor g__10845(w__10926 ,w__10886 ,w__10903);
  and g__10846(w__10925 ,w__10883 ,w__10899);
  or g__10847(w__10924 ,w__9579 ,w__10895);
  nor g__10848(w__10923 ,w__10802 ,w__10907);
  nor g__10849(w__10922 ,w__10888 ,w__10901);
  nor g__10850(w__10921 ,w__10824 ,w__10910);
  or g__10851(w__10915 ,w__10801 ,w__10906);
  or g__10852(w__13219 ,w__10877 ,w__10893);
  xnor g__10853(w__13231 ,w__10831 ,w__9241);
  xnor g__10854(w__13233 ,w__10741 ,w__10861);
  xnor g__10855(w__13154 ,w__10809 ,w__10862);
  xnor g__10856(w__10914 ,w__10773 ,w__10868);
  xnor g__10857(w__10913 ,w__10871 ,w__10826);
  xnor g__10858(w__10912 ,w__10763 ,w__10872);
  xnor g__10859(w__10920 ,w__10808 ,w__10864);
  xnor g__10860(w__10919 ,w__10857 ,w__10860);
  xnor g__10861(w__10918 ,w__10834 ,w__10863);
  xnor g__10862(w__10917 ,w__10806 ,w__10858);
  xnor g__10863(w__10916 ,w__10830 ,w__10859);
  not g__10864(w__10908 ,w__10909);
  not g__10865(w__10906 ,w__10907);
  nor g__10866(w__10905 ,w__10826 ,w__10871);
  nor g__10867(w__10904 ,w__10773 ,w__10869);
  and g__10868(w__10903 ,w__10773 ,w__10869);
  or g__10869(w__13165 ,w__10848 ,w__10882);
  nor g__10870(w__10902 ,w__10763 ,w__10873);
  or g__10871(w__13166 ,w__10846 ,w__10881);
  or g__10872(w__13168 ,w__10842 ,w__10880);
  or g__10873(w__13218 ,w__10840 ,w__10878);
  and g__10874(w__10901 ,w__10763 ,w__10873);
  and g__10875(w__10911 ,w__10854 ,w__10874);
  and g__10876(w__10910 ,w__10837 ,w__10875);
  and g__10877(w__10909 ,w__10852 ,w__10885);
  and g__10878(w__10907 ,w__10843 ,w__10879);
  not g__10879(w__10898 ,w__10897);
  not g__10880(w__10895 ,w__10896);
  or g__10881(w__10894 ,w__10825 ,w__10870);
  nor g__10882(w__10893 ,w__10887 ,w__10876);
  or g__10883(w__13217 ,w__10836 ,w__10865);
  xnor g__10884(w__13232 ,w__10833 ,w__10814);
  or g__10885(w__13167 ,w__10794 ,w__10867);
  xnor g__10886(w__10892 ,w__10777 ,w__10829);
  xnor g__10887(w__10891 ,w__10821 ,w__10819);
  xnor g__10888(w__10890 ,w__10758 ,w__10827);
  xnor g__10889(w__10889 ,w__10832 ,w__10717);
  or g__10890(w__10900 ,w__10849 ,w__10866);
  xnor g__10891(w__10899 ,w__10760 ,w__10812);
  xnor g__10892(w__10897 ,w__10640 ,w__10811);
  xnor g__10893(w__10896 ,w__10807 ,w__10813);
  or g__10894(w__10885 ,w__10806 ,w__10850);
  nor g__10895(w__10884 ,w__10819 ,w__10821);
  or g__10896(w__10883 ,w__10818 ,w__10820);
  and g__10897(w__10882 ,w__10847 ,w__10829);
  nor g__10898(w__10881 ,w__10856 ,w__10831);
  and g__10899(w__10880 ,w__10741 ,w__10841);
  or g__10900(w__13169 ,w__10743 ,w__10839);
  or g__10901(w__10879 ,w__10857 ,w__10838);
  nor g__10902(w__10878 ,w__10815 ,w__10832);
  nor g__10903(w__10877 ,w__10758 ,w__10828);
  and g__10904(w__10876 ,w__10758 ,w__10828);
  or g__10905(w__10875 ,w__10830 ,w__10855);
  or g__10906(w__10874 ,w__10808 ,w__10853);
  and g__10907(w__10888 ,w__10735 ,w__10844);
  and g__10908(w__10887 ,w__10670 ,w__10817);
  and g__10909(w__10886 ,w__10798 ,w__10851);
  not g__10910(w__10873 ,w__10872);
  not g__10911(w__10870 ,w__10871);
  not g__10912(w__10869 ,w__10868);
  nor g__10913(w__10867 ,w__10795 ,w__10833);
  nor g__10914(w__10866 ,w__10845 ,w__10834);
  nor g__10915(w__10865 ,w__10809 ,w__10835);
  xnor g__10916(w__13234 ,w__10789 ,w__10769);
  xnor g__10917(w__13153 ,w__10738 ,w__10767);
  xnor g__10918(w__10864 ,w__10643 ,w__10775);
  xnor g__10919(w__10863 ,w__10762 ,w__10786);
  xnor g__10920(w__10862 ,w__10543 ,w__10784);
  xnor g__10921(w__10861 ,w__10781 ,w__10582);
  xnor g__10922(w__10860 ,w__10783 ,w__10757);
  xnor g__10923(w__10859 ,w__10772 ,w__10513);
  xnor g__10924(w__10858 ,w__10712 ,w__10779);
  xnor g__10925(w__10872 ,w__10788 ,w__10727);
  and g__10926(w__10871 ,w__10770 ,w__10816);
  xnor g__10927(w__10868 ,w__10810 ,w__10768);
  and g__10928(w__10856 ,w__10782 ,w__10803);
  and g__10929(w__10855 ,w__10513 ,w__10772);
  or g__10930(w__10854 ,w__10642 ,w__10775);
  nor g__10931(w__10853 ,w__10643 ,w__10774);
  or g__10932(w__10852 ,w__10712 ,w__10778);
  or g__10933(w__10851 ,w__10796 ,w__10807);
  nor g__10934(w__10850 ,w__10711 ,w__10779);
  nor g__10935(w__10849 ,w__10762 ,w__10787);
  nor g__10936(w__10848 ,w__10805 ,w__10777);
  or g__10937(w__10847 ,w__10804 ,w__10776);
  nor g__10938(w__10846 ,w__10782 ,w__10803);
  and g__10939(w__10845 ,w__10762 ,w__10787);
  or g__10940(w__10844 ,w__10745 ,w__10810);
  or g__10941(w__10843 ,w__10757 ,w__10783);
  nor g__10942(w__10842 ,w__9431 ,w__10781);
  or g__10943(w__10841 ,w__9578 ,w__10780);
  nor g__10944(w__10840 ,w__10717 ,w__10800);
  and g__10945(w__10839 ,w__10744 ,w__10789);
  and g__10946(w__10838 ,w__10757 ,w__10783);
  or g__10947(w__13215 ,w__10749 ,w__10791);
  or g__10948(w__13216 ,w__10752 ,w__10790);
  or g__10949(w__10837 ,w__10513 ,w__10772);
  nor g__10950(w__10836 ,w__10543 ,w__10785);
  and g__10951(w__10835 ,w__10543 ,w__10785);
  and g__10952(w__10857 ,w__10660 ,w__10799);
  not g__10953(w__10828 ,w__10827);
  not g__10954(w__10826 ,w__10825);
  not g__10955(w__10820 ,w__10821);
  not g__10956(w__10818 ,w__10819);
  xnor g__10957(w__13151 ,w__10511 ,w__10733);
  xnor g__10958(w__13235 ,w__10739 ,w__10726);
  or g__10959(w__10817 ,w__10704 ,w__10788);
  or g__10960(w__10816 ,w__10740 ,w__10771);
  and g__10961(w__10815 ,w__10717 ,w__10800);
  or g__10962(w__13170 ,w__10663 ,w__10797);
  xnor g__10963(w__13236 ,w__10635 ,w__10724);
  xnor g__10964(w__13152 ,w__10716 ,w__10730);
  xnor g__10965(w__10814 ,w__10674 ,w__10764);
  xnor g__10966(w__10813 ,w__10761 ,w__10673);
  xnor g__10967(w__10812 ,w__10548 ,w__10740);
  xnor g__10968(w__10811 ,w__10766 ,w__10576);
  xnor g__10969(w__10834 ,w__10541 ,w__10722);
  xnor g__10970(w__10833 ,w__10645 ,w__10723);
  xnor g__10971(w__10832 ,w__9239 ,w__10725);
  xnor g__10972(w__10831 ,w__10678 ,w__10732);
  and g__10973(w__10830 ,w__10669 ,w__10792);
  xnor g__10974(w__10829 ,w__10765 ,w__10731);
  xnor g__10975(w__10827 ,w__10679 ,w__10729);
  xnor g__10976(w__10825 ,w__10579 ,w__10728);
  xnor g__10977(w__10824 ,w__10505 ,w__10721);
  xnor g__10978(w__10823 ,w__10737 ,w__10718);
  xnor g__10979(w__10822 ,w__10580 ,w__10719);
  xnor g__10980(w__10821 ,w__10574 ,w__10720);
  and g__10981(w__10819 ,w__10698 ,w__10793);
  not g__10982(w__10804 ,w__10805);
  not g__10983(w__10801 ,w__10802);
  or g__10984(w__10799 ,w__10659 ,w__10766);
  or g__10985(w__10798 ,w__10673 ,w__10761);
  nor g__10986(w__10797 ,w__10662 ,w__10739);
  and g__10987(w__10796 ,w__10673 ,w__10761);
  and g__10988(w__10795 ,w__10675 ,w__10764);
  nor g__10989(w__10794 ,w__10675 ,w__10764);
  or g__10990(w__10793 ,w__10765 ,w__10695);
  or g__10991(w__10792 ,w__10667 ,w__10737);
  and g__10992(w__10791 ,w__10644 ,w__10751);
  and g__10993(w__10790 ,w__10738 ,w__10747);
  and g__10994(w__10810 ,w__10710 ,w__10754);
  and g__10995(w__10809 ,w__10683 ,w__10734);
  and g__10996(w__10808 ,w__10709 ,w__10755);
  and g__10997(w__10807 ,w__10665 ,w__10748);
  and g__10998(w__10806 ,w__10703 ,w__10753);
  and g__10999(w__10805 ,w__10694 ,w__10746);
  and g__11000(w__10803 ,w__10690 ,w__10756);
  and g__11001(w__10802 ,w__10688 ,w__10742);
  and g__11002(w__10800 ,w__10708 ,w__10750);
  not g__11003(w__10787 ,w__10786);
  not g__11004(w__10785 ,w__10784);
  not g__11005(w__10780 ,w__10781);
  not g__11006(w__10778 ,w__10779);
  not g__11007(w__10776 ,w__10777);
  not g__11008(w__10774 ,w__10775);
  xnor g__11009(w__13237 ,w__10591 ,w__9240);
  or g__11010(w__13171 ,w__10681 ,w__10736);
  nor g__11011(w__10771 ,w__10548 ,w__10759);
  or g__11012(w__10770 ,w__10547 ,w__10760);
  xnor g__11013(w__10769 ,w__10714 ,w__10565);
  xnor g__11014(w__10768 ,w__9237 ,w__10672);
  xnor g__11015(w__10767 ,w__10677 ,w__10566);
  xnor g__11016(w__10789 ,w__10598 ,w__10652);
  xnor g__11017(w__10788 ,w__10593 ,w__10649);
  xnor g__11018(w__10786 ,w__10550 ,w__9236);
  xnor g__11019(w__10784 ,w__10594 ,w__9238);
  xnor g__11020(w__10783 ,w__10587 ,w__10648);
  xnor g__11021(w__10782 ,w__10552 ,w__10646);
  xnor g__11022(w__10781 ,w__10592 ,w__10647);
  xnor g__11023(w__10779 ,w__10526 ,w__10654);
  xnor g__11024(w__10777 ,w__10599 ,w__10655);
  xnor g__11025(w__10775 ,w__10503 ,w__10651);
  xnor g__11026(w__10773 ,w__10584 ,w__10653);
  xnor g__11027(w__10772 ,w__10585 ,w__10650);
  not g__11028(w__10759 ,w__10760);
  or g__11029(w__10756 ,w__10645 ,w__10689);
  or g__11030(w__10755 ,w__10590 ,w__10707);
  or g__11031(w__10754 ,w__10589 ,w__10706);
  or g__11032(w__10753 ,w__10588 ,w__10701);
  nor g__11033(w__10752 ,w__9432 ,w__10677);
  or g__11034(w__10751 ,w__10537 ,w__10715);
  or g__11035(w__10750 ,w__10700 ,w__10680);
  nor g__11036(w__10749 ,w__10538 ,w__10716);
  or g__11037(w__13214 ,w__10600 ,w__10668);
  or g__11038(w__10748 ,w__10595 ,w__10664);
  or g__11039(w__10747 ,w__9577 ,w__10676);
  or g__11040(w__10746 ,w__10678 ,w__10692);
  or g__11041(w__13172 ,w__10608 ,w__10693);
  nor g__11042(w__10745 ,w__9237 ,w__10671);
  or g__11043(w__10744 ,w__9576 ,w__10713);
  nor g__11044(w__10743 ,w__9429 ,w__10714);
  or g__11045(w__10742 ,w__10586 ,w__10686);
  and g__11046(w__10766 ,w__10609 ,w__10696);
  and g__11047(w__10765 ,w__10627 ,w__10697);
  and g__11048(w__10764 ,w__10619 ,w__10687);
  and g__11049(w__10763 ,w__10623 ,w__10682);
  and g__11050(w__10762 ,w__10624 ,w__10691);
  and g__11051(w__10761 ,w__10632 ,w__10702);
  and g__11052(w__10760 ,w__10631 ,w__10699);
  and g__11053(w__10758 ,w__10616 ,w__10656);
  and g__11054(w__10757 ,w__10615 ,w__10684);
  or g__11055(w__13173 ,w__10456 ,w__10657);
  nor g__11056(w__10736 ,w__10597 ,w__10685);
  or g__11057(w__10735 ,w__10641 ,w__10672);
  xnor g__11058(w__13238 ,w__10596 ,w__10499);
  or g__11059(w__10734 ,w__9239 ,w__10705);
  xnor g__11060(w__10733 ,w__10583 ,w__10211);
  xnor g__11061(w__10732 ,w__10568 ,w__10569);
  xnor g__11062(w__10731 ,w__10571 ,w__10638);
  xnor g__11063(w__10730 ,w__10538 ,w__10644);
  xnor g__11064(w__10729 ,w__10572 ,w__10546);
  xnor g__11065(w__10728 ,w__10558 ,w__10590);
  xnor g__11066(w__10727 ,w__10518 ,w__10562);
  xnor g__11067(w__10726 ,w__10509 ,w__10564);
  xnor g__11068(w__10725 ,w__10560 ,w__10504);
  xnor g__11069(w__10724 ,w__10597 ,w__10521);
  xnor g__11070(w__10723 ,w__10567 ,w__10563);
  xnor g__11071(w__10722 ,w__10581 ,w__10595);
  xnor g__11072(w__10721 ,w__10577 ,w__10586);
  xnor g__11073(w__10720 ,w__10588 ,w__10534);
  xnor g__11074(w__10719 ,w__10589 ,w__10540);
  xnor g__11075(w__10718 ,w__10573 ,w__10559);
  or g__11076(w__10741 ,w__10614 ,w__10658);
  xnor g__11077(w__10740 ,w__10549 ,w__10556);
  xnor g__11078(w__10739 ,w__10524 ,w__10555);
  or g__11079(w__10738 ,w__10630 ,w__10661);
  and g__11080(w__10737 ,w__10602 ,w__10666);
  not g__11081(w__10715 ,w__10716);
  not g__11082(w__10713 ,w__10714);
  not g__11083(w__10711 ,w__10712);
  or g__11084(w__13213 ,w__10327 ,w__10605);
  or g__11085(w__10710 ,w__10540 ,w__10580);
  or g__11086(w__10709 ,w__10557 ,w__10579);
  or g__11087(w__10708 ,w__10546 ,w__10572);
  nor g__11088(w__10707 ,w__10558 ,w__10578);
  and g__11089(w__10706 ,w__10540 ,w__10580);
  and g__11090(w__10705 ,w__10504 ,w__10560);
  nor g__11091(w__10704 ,w__10518 ,w__10561);
  or g__11092(w__10703 ,w__10534 ,w__10574);
  or g__11093(w__10702 ,w__10550 ,w__10629);
  and g__11094(w__10701 ,w__10534 ,w__10574);
  and g__11095(w__10700 ,w__10546 ,w__10572);
  or g__11096(w__10699 ,w__10599 ,w__10628);
  or g__11097(w__10698 ,w__10571 ,w__10637);
  or g__11098(w__10697 ,w__10552 ,w__10626);
  or g__11099(w__10696 ,w__10522 ,w__10606);
  nor g__11100(w__10695 ,w__10570 ,w__10638);
  or g__11101(w__10694 ,w__10569 ,w__10568);
  nor g__11102(w__10693 ,w__10607 ,w__10591);
  and g__11103(w__10692 ,w__10569 ,w__10568);
  or g__11104(w__10691 ,w__10622 ,w__10587);
  or g__11105(w__10690 ,w__10563 ,w__10567);
  and g__11106(w__10689 ,w__10563 ,w__10567);
  or g__11107(w__10688 ,w__10505 ,w__10577);
  or g__11108(w__10687 ,w__10618 ,w__10592);
  and g__11109(w__10686 ,w__10505 ,w__10577);
  and g__11110(w__10685 ,w__10521 ,w__10636);
  or g__11111(w__10684 ,w__10611 ,w__10585);
  or g__11112(w__10683 ,w__10504 ,w__10560);
  or g__11113(w__10682 ,w__10610 ,w__10584);
  nor g__11114(w__10681 ,w__10521 ,w__10636);
  and g__11115(w__10717 ,w__10302 ,w__10625);
  and g__11116(w__10716 ,w__10343 ,w__10617);
  and g__11117(w__10714 ,w__10500 ,w__10612);
  and g__11118(w__10712 ,w__10527 ,w__10633);
  not g__11119(w__10680 ,w__10679);
  not g__11120(w__10676 ,w__10677);
  not g__11121(w__10675 ,w__10674);
  not g__11122(w__10671 ,w__10672);
  xnor g__11123(w__13150 ,w__10554 ,w__10448);
  or g__11124(w__10670 ,w__10517 ,w__10562);
  or g__11125(w__10669 ,w__10559 ,w__10573);
  nor g__11126(w__10668 ,w__10620 ,w__10583);
  and g__11127(w__10667 ,w__10559 ,w__10573);
  or g__11128(w__10666 ,w__10526 ,w__10613);
  or g__11129(w__10665 ,w__10541 ,w__10581);
  and g__11130(w__10664 ,w__10541 ,w__10581);
  nor g__11131(w__10663 ,w__10510 ,w__10564);
  and g__11132(w__10662 ,w__10510 ,w__10564);
  nor g__11133(w__10661 ,w__10621 ,w__10594);
  or g__11134(w__10660 ,w__10576 ,w__10639);
  nor g__11135(w__10659 ,w__10575 ,w__10640);
  nor g__11136(w__10658 ,w__10634 ,w__10598);
  nor g__11137(w__10657 ,w__10454 ,w__10596);
  or g__11138(w__10656 ,w__10604 ,w__10593);
  xnor g__11139(w__10655 ,w__10542 ,w__10544);
  xnor g__11140(w__10654 ,w__10334 ,w__10508);
  xnor g__11141(w__10653 ,w__10516 ,w__10533);
  xnor g__11142(w__10652 ,w__10331 ,w__10506);
  xnor g__11143(w__10651 ,w__10522 ,w__10520);
  xnor g__11144(w__10650 ,w__10514 ,w__10515);
  xnor g__11145(w__10649 ,w__10512 ,w__10131);
  xnor g__11146(w__10648 ,w__10535 ,w__10536);
  xnor g__11147(w__10647 ,w__10530 ,w__10531);
  xnor g__11148(w__10646 ,w__10539 ,w__10440);
  xnor g__11149(w__10679 ,w__10553 ,w__10446);
  and g__11150(w__10678 ,w__10476 ,w__10601);
  xnor g__11151(w__10677 ,w__10523 ,w__10433);
  xnor g__11152(w__10674 ,w__10551 ,w__10498);
  xnor g__11153(w__10673 ,w__10525 ,w__10434);
  and g__11154(w__10672 ,w__10281 ,w__10603);
  not g__11155(w__10642 ,w__10643);
  not g__11156(w__10641 ,w__9237);
  not g__11157(w__10639 ,w__10640);
  not g__11158(w__10637 ,w__10638);
  not g__11159(w__10636 ,w__10635);
  and g__11160(w__10634 ,w__10332 ,w__10506);
  or g__11161(w__10633 ,w__10528 ,w__10549);
  or g__11162(w__10632 ,w__10128 ,w__10532);
  or g__11163(w__10631 ,w__10544 ,w__10542);
  nor g__11164(w__10630 ,w__10207 ,w__10545);
  and g__11165(w__10629 ,w__10128 ,w__10532);
  and g__11166(w__10628 ,w__10544 ,w__10542);
  or g__11167(w__10627 ,w__10440 ,w__10539);
  and g__11168(w__10626 ,w__10440 ,w__10539);
  or g__11169(w__10625 ,w__10306 ,w__10553);
  or g__11170(w__10624 ,w__10536 ,w__10535);
  or g__11171(w__10623 ,w__10533 ,w__10516);
  and g__11172(w__10622 ,w__10536 ,w__10535);
  and g__11173(w__10621 ,w__10207 ,w__10545);
  nor g__11174(w__10620 ,w__10210 ,w__10511);
  or g__11175(w__10619 ,w__10531 ,w__10530);
  and g__11176(w__10618 ,w__10531 ,w__10530);
  or g__11177(w__10617 ,w__10298 ,w__10523);
  or g__11178(w__10616 ,w__10131 ,w__10512);
  or g__11179(w__10615 ,w__10515 ,w__10514);
  nor g__11180(w__10614 ,w__10332 ,w__10506);
  nor g__11181(w__10613 ,w__10334 ,w__10507);
  or g__11182(w__10612 ,w__10524 ,w__10501);
  and g__11183(w__10611 ,w__10515 ,w__10514);
  and g__11184(w__10610 ,w__10533 ,w__10516);
  or g__11185(w__10609 ,w__10503 ,w__10520);
  nor g__11186(w__10608 ,w__10441 ,w__10519);
  and g__11187(w__10607 ,w__10441 ,w__10519);
  or g__11188(w__13174 ,w__10294 ,w__10502);
  and g__11189(w__10606 ,w__10503 ,w__10520);
  nor g__11190(w__10605 ,w__10320 ,w__10554);
  and g__11191(w__10604 ,w__9386 ,w__10512);
  or g__11192(w__10603 ,w__10280 ,w__10525);
  or g__11193(w__10602 ,w__10333 ,w__10508);
  or g__11194(w__10601 ,w__10475 ,w__10551);
  and g__11195(w__10600 ,w__9434 ,w__10511);
  and g__11196(w__10645 ,w__10336 ,w__10529);
  xnor g__11197(w__10644 ,w__10426 ,w__10211);
  xnor g__11198(w__10643 ,w__10412 ,w__9453);
  xnor g__11199(w__10640 ,w__10445 ,w__10212);
  xnor g__11200(w__10638 ,w__10390 ,w__10404);
  xnor g__11201(w__10635 ,w__10335 ,w__10391);
  not g__11202(w__10578 ,w__10579);
  not g__11203(w__10575 ,w__10576);
  not g__11204(w__10570 ,w__10571);
  not g__11205(w__10561 ,w__10562);
  not g__11206(w__10557 ,w__10558);
  xnor g__11207(w__13240 ,w__10178 ,w__10431);
  xnor g__11208(w__13149 ,w__10401 ,w__9620);
  xnor g__11209(w__13239 ,w__10443 ,w__10421);
  xnor g__11210(w__10556 ,w__10439 ,w__10246);
  xnor g__11211(w__10555 ,w__10442 ,w__10163);
  xnor g__11212(w__10599 ,w__10244 ,w__10430);
  xnor g__11213(w__10598 ,w__10213 ,w__10432);
  xnor g__11214(w__10597 ,w__10257 ,w__10427);
  xnor g__11215(w__10596 ,w__10139 ,w__10428);
  xnor g__11216(w__10595 ,w__10403 ,w__9649);
  xnor g__11217(w__10594 ,w__10193 ,w__10423);
  xnor g__11218(w__10593 ,w__10416 ,w__9653);
  xnor g__11219(w__10592 ,w__10184 ,w__10396);
  xnor g__11220(w__10591 ,w__10260 ,w__10414);
  xnor g__11221(w__10590 ,w__10268 ,w__10409);
  xnor g__11222(w__10589 ,w__10191 ,w__10408);
  xnor g__11223(w__10588 ,w__10259 ,w__10406);
  xnor g__11224(w__10587 ,w__10258 ,w__10398);
  xnor g__11225(w__10586 ,w__10267 ,w__10437);
  xnor g__11226(w__10585 ,w__10261 ,w__10393);
  xnor g__11227(w__10584 ,w__10153 ,w__10392);
  xnor g__11228(w__10583 ,w__10402 ,w__9630);
  xnor g__11229(w__10582 ,w__10444 ,w__10395);
  xnor g__11230(w__10581 ,w__10190 ,w__10425);
  xnor g__11231(w__10580 ,w__10263 ,w__10410);
  xnor g__11232(w__10579 ,w__10165 ,w__10438);
  xnor g__11233(w__10577 ,w__10397 ,w__10209);
  xnor g__11234(w__10576 ,w__10231 ,w__10422);
  xnor g__11235(w__10574 ,w__10159 ,w__10407);
  xnor g__11236(w__10573 ,w__10278 ,w__10420);
  xnor g__11237(w__10572 ,w__10156 ,w__10411);
  xnor g__11238(w__10571 ,w__10226 ,w__10405);
  xnor g__11239(w__10569 ,w__10247 ,w__10400);
  xnor g__11240(w__10568 ,w__10265 ,w__10399);
  xnor g__11241(w__10567 ,w__10235 ,w__10419);
  xnor g__11242(w__10566 ,w__10394 ,w__9651);
  xnor g__11243(w__10565 ,w__10243 ,w__10418);
  xnor g__11244(w__10564 ,w__10181 ,w__10413);
  xnor g__11245(w__10563 ,w__10166 ,w__10429);
  xnor g__11246(w__10562 ,w__10227 ,w__10415);
  xnor g__11247(w__10560 ,w__10233 ,w__10417);
  xnor g__11248(w__10559 ,w__10146 ,w__10436);
  xnor g__11249(w__10558 ,w__10202 ,w__10447);
  not g__11250(w__10547 ,w__10548);
  not g__11251(w__10537 ,w__10538);
  or g__11252(w__10529 ,w__10344 ,w__10444);
  and g__11253(w__10528 ,w__10246 ,w__10439);
  or g__11254(w__10527 ,w__10246 ,w__10439);
  and g__11255(w__10554 ,w__10382 ,w__10466);
  and g__11256(w__10553 ,w__10387 ,w__10481);
  and g__11257(w__10552 ,w__10350 ,w__10478);
  and g__11258(w__10551 ,w__10341 ,w__10472);
  and g__11259(w__10550 ,w__10370 ,w__10485);
  and g__11260(w__10549 ,w__10378 ,w__10491);
  or g__11261(w__10548 ,w__10373 ,w__10486);
  and g__11262(w__10546 ,w__10380 ,w__10489);
  and g__11263(w__10545 ,w__10362 ,w__10474);
  and g__11264(w__10544 ,w__10367 ,w__10484);
  and g__11265(w__10543 ,w__10283 ,w__10496);
  and g__11266(w__10542 ,w__10363 ,w__10482);
  and g__11267(w__10541 ,w__10361 ,w__10480);
  and g__11268(w__10540 ,w__10385 ,w__10495);
  and g__11269(w__10539 ,w__10353 ,w__10479);
  and g__11270(w__10538 ,w__10381 ,w__10492);
  and g__11271(w__10536 ,w__10347 ,w__10477);
  and g__11272(w__10535 ,w__10342 ,w__10473);
  and g__11273(w__10534 ,w__10376 ,w__10490);
  and g__11274(w__10533 ,w__10340 ,w__10469);
  and g__11275(w__10532 ,w__10375 ,w__10488);
  and g__11276(w__10531 ,w__10326 ,w__10497);
  and g__11277(w__10530 ,w__10384 ,w__10468);
  not g__11278(w__10517 ,w__10518);
  not g__11279(w__10510 ,w__10509);
  not g__11280(w__10507 ,w__10508);
  and g__11281(w__10502 ,w__10301 ,w__10443);
  or g__11282(w__13175 ,w__10304 ,w__10452);
  and g__11283(w__10501 ,w__10163 ,w__10442);
  or g__11284(w__10500 ,w__10163 ,w__10442);
  xnor g__11285(w__10499 ,w__10137 ,w__10329);
  xnor g__11286(w__10498 ,w__10230 ,w__10389);
  and g__11287(w__10526 ,w__10357 ,w__10470);
  and g__11288(w__10525 ,w__10293 ,w__10450);
  and g__11289(w__10524 ,w__10322 ,w__10462);
  and g__11290(w__10523 ,w__10287 ,w__10451);
  and g__11291(w__10522 ,w__10300 ,w__10453);
  and g__11292(w__10521 ,w__10309 ,w__10460);
  and g__11293(w__10520 ,w__10349 ,w__10457);
  and g__11294(w__10519 ,w__10308 ,w__10459);
  or g__11295(w__10518 ,w__10286 ,w__10458);
  and g__11296(w__10516 ,w__10290 ,w__10463);
  and g__11297(w__10515 ,w__10321 ,w__10467);
  and g__11298(w__10514 ,w__10317 ,w__10464);
  and g__11299(w__10513 ,w__10299 ,w__10487);
  and g__11300(w__10512 ,w__10291 ,w__10493);
  or g__11301(w__10511 ,w__10285 ,w__10483);
  or g__11302(w__10509 ,w__10312 ,w__10471);
  and g__11303(w__10508 ,w__10296 ,w__10494);
  and g__11304(w__10506 ,w__10319 ,w__10465);
  and g__11305(w__10505 ,w__10328 ,w__10449);
  and g__11306(w__10504 ,w__10310 ,w__10455);
  and g__11307(w__10503 ,w__10279 ,w__10461);
  or g__11308(w__10497 ,w__10276 ,w__10325);
  or g__11309(w__10496 ,w__10277 ,w__10282);
  or g__11310(w__10495 ,w__10275 ,w__10383);
  or g__11311(w__10494 ,w__10274 ,w__10358);
  or g__11312(w__10493 ,w__10201 ,w__10292);
  or g__11313(w__10492 ,w__10379 ,w__10273);
  or g__11314(w__10491 ,w__10189 ,w__10377);
  or g__11315(w__10490 ,w__10272 ,w__10374);
  or g__11316(w__10489 ,w__10271 ,w__10371);
  or g__11317(w__10488 ,w__10269 ,w__10372);
  or g__11318(w__10487 ,w__9575 ,w__10369);
  and g__11319(w__10486 ,w__10390 ,w__10368);
  or g__11320(w__10485 ,w__10267 ,w__10365);
  or g__11321(w__10484 ,w__10266 ,w__10364);
  nor g__11322(w__10483 ,w__10288 ,w__9434);
  or g__11323(w__10482 ,w__10265 ,w__10359);
  or g__11324(w__10481 ,w__10203 ,w__10352);
  or g__11325(w__10480 ,w__9455 ,w__10356);
  or g__11326(w__10479 ,w__10264 ,w__10351);
  or g__11327(w__10478 ,w__10187 ,w__10348);
  or g__11328(w__10477 ,w__10192 ,w__10345);
  or g__11329(w__10476 ,w__10230 ,w__10388);
  nor g__11330(w__10475 ,w__10229 ,w__10389);
  or g__11331(w__10474 ,w__10262 ,w__10338);
  or g__11332(w__10473 ,w__10261 ,w__10337);
  or g__11333(w__10472 ,w__10184 ,w__10339);
  and g__11334(w__10471 ,w__10335 ,w__10366);
  or g__11335(w__10470 ,w__10259 ,w__10386);
  or g__11336(w__10469 ,w__10263 ,w__10354);
  or g__11337(w__10468 ,w__10180 ,w__10323);
  or g__11338(w__10467 ,w__10177 ,w__10318);
  or g__11339(w__10466 ,w__10315 ,w__10200);
  or g__11340(w__10465 ,w__10181 ,w__10316);
  or g__11341(w__10464 ,w__10278 ,w__10314);
  or g__11342(w__10463 ,w__10191 ,w__10311);
  or g__11343(w__10462 ,w__10196 ,w__10313);
  or g__11344(w__10461 ,w__10295 ,w__10202);
  or g__11345(w__10460 ,w__10260 ,w__10297);
  or g__11346(w__10459 ,w__10188 ,w__10307);
  and g__11347(w__10458 ,w__10289 ,w__9386);
  or g__11348(w__10457 ,w__10268 ,w__10305);
  nor g__11349(w__10456 ,w__10137 ,w__10330);
  or g__11350(w__10455 ,w__10270 ,w__10355);
  and g__11351(w__10454 ,w__10137 ,w__10330);
  or g__11352(w__10453 ,w__10199 ,w__10303);
  nor g__11353(w__10452 ,w__10178 ,w__10346);
  or g__11354(w__10451 ,w__10284 ,w__10193);
  or g__11355(w__10450 ,w__10190 ,w__10360);
  or g__11356(w__10449 ,w__9453 ,w__10324);
  xnor g__11357(w__13241 ,w__10204 ,w__10125);
  xnor g__11358(w__10448 ,w__10136 ,w__9436);
  xnor g__11359(w__10447 ,w__10170 ,w__9628);
  xnor g__11360(w__10446 ,w__10150 ,w__10129);
  xnor g__11361(w__10445 ,w__10215 ,w__9455);
  xnor g__11362(w__10438 ,w__10132 ,w__10199);
  xnor g__11363(w__10437 ,w__10249 ,w__9648);
  xnor g__11364(w__10436 ,w__10177 ,w__9622);
  xnor g__11365(w__10435 ,w__10277 ,w__9654);
  xnor g__11366(w__10434 ,w__9384 ,w__9624);
  xnor g__11367(w__10433 ,w__10219 ,w__10206);
  xnor g__11368(w__10432 ,w__10276 ,w__9883);
  xnor g__11369(w__10431 ,w__9888 ,w__10172);
  xnor g__11370(w__10430 ,w__10189 ,w__9886);
  xnor g__11371(w__10429 ,w__10264 ,w__9884);
  xnor g__11372(w__10428 ,w__10188 ,w__9887);
  xnor g__11373(w__10427 ,w__10196 ,w__9885);
  xnor g__11374(w__10426 ,w__10152 ,w__9650);
  xnor g__11375(w__10425 ,w__10214 ,w__10151);
  xnor g__11376(w__10424 ,w__10149 ,w__9626);
  xnor g__11377(w__10423 ,w__10147 ,w__9652);
  xnor g__11378(w__10422 ,w__10192 ,w__9623);
  xnor g__11379(w__10421 ,w__10174 ,w__10134);
  xnor g__11380(w__10420 ,w__10167 ,w__10142);
  xnor g__11381(w__10419 ,w__10234 ,w__10187);
  xnor g__11382(w__10418 ,w__10238 ,w__10180);
  xnor g__11383(w__10417 ,w__10262 ,w__10239);
  xnor g__11384(w__10416 ,w__10237 ,w__10203);
  xnor g__11385(w__10415 ,w__10271 ,w__10248);
  xnor g__11386(w__10414 ,w__10143 ,w__10145);
  xnor g__11387(w__10413 ,w__10135 ,w__10168);
  xnor g__11388(w__10412 ,w__10158 ,w__10154);
  xnor g__11389(w__10411 ,w__10270 ,w__9627);
  xnor g__11390(w__10410 ,w__10218 ,w__10222);
  xnor g__11391(w__10409 ,w__10138 ,w__10220);
  xnor g__11392(w__10408 ,w__10171 ,w__10155);
  xnor g__11393(w__10407 ,w__10157 ,w__10274);
  xnor g__11394(w__10406 ,w__10162 ,w__10232);
  xnor g__11395(w__10405 ,w__10241 ,w__10272);
  xnor g__11396(w__10404 ,w__10252 ,w__10254);
  xnor g__11397(w__10403 ,w__10275 ,w__10256);
  xnor g__11398(w__10402 ,w__10200 ,w__10250);
  xnor g__11399(w__10401 ,w__9632 ,w__10205);
  xnor g__11400(w__10400 ,w__10266 ,w__10245);
  xnor g__11401(w__10399 ,w__10164 ,w__10236);
  xnor g__11402(w__10398 ,w__10269 ,w__10221);
  xnor g__11403(w__10397 ,w__10240 ,w__10242);
  xnor g__11404(w__10396 ,w__10223 ,w__10225);
  xnor g__11405(w__10395 ,w__10216 ,w__10217);
  xnor g__11406(w__10394 ,w__10273 ,w__10255);
  xnor g__11407(w__10393 ,w__10224 ,w__10228);
  xnor g__11408(w__10392 ,w__10144 ,w__10201);
  xnor g__11409(w__10391 ,w__10161 ,w__10141);
  xnor g__11410(w__10444 ,w__10197 ,w__10119);
  xnor g__11411(w__10443 ,w__10113 ,w__10179);
  xnor g__11412(w__10442 ,w__10121 ,w__10175);
  xnor g__11413(w__10441 ,w__10123 ,w__10185);
  xnor g__11414(w__10440 ,w__10117 ,w__10182);
  xnor g__11415(w__10439 ,w__10115 ,w__10194);
  not g__11416(w__10388 ,w__10389);
  or g__11417(w__10387 ,w__9456 ,w__10237);
  and g__11418(w__10386 ,w__10232 ,w__10162);
  or g__11419(w__10385 ,w__9457 ,w__10256);
  or g__11420(w__10384 ,w__10238 ,w__10243);
  and g__11421(w__10383 ,w__9649 ,w__10256);
  or g__11422(w__10382 ,w__9466 ,w__10250);
  or g__11423(w__10381 ,w__9464 ,w__10255);
  or g__11424(w__10380 ,w__10248 ,w__10227);
  and g__11425(w__10379 ,w__9651 ,w__10255);
  or g__11426(w__10378 ,w__9886 ,w__10244);
  and g__11427(w__10377 ,w__9886 ,w__10244);
  or g__11428(w__10376 ,w__10241 ,w__10226);
  or g__11429(w__10375 ,w__10221 ,w__10258);
  and g__11430(w__10374 ,w__10241 ,w__10226);
  nor g__11431(w__10373 ,w__10254 ,w__10252);
  and g__11432(w__10372 ,w__10221 ,w__10258);
  and g__11433(w__10371 ,w__10248 ,w__10227);
  or g__11434(w__10370 ,w__9462 ,w__10249);
  and g__11435(w__10369 ,w__10154 ,w__10158);
  or g__11436(w__10368 ,w__10253 ,w__10251);
  or g__11437(w__10367 ,w__10247 ,w__10245);
  or g__11438(w__10366 ,w__10140 ,w__10160);
  and g__11439(w__10365 ,w__9648 ,w__10249);
  and g__11440(w__10364 ,w__10247 ,w__10245);
  or g__11441(w__10363 ,w__10236 ,w__10164);
  or g__11442(w__10362 ,w__10239 ,w__10233);
  or g__11443(w__10361 ,w__10242 ,w__10240);
  and g__11444(w__10360 ,w__10151 ,w__10214);
  and g__11445(w__10359 ,w__10236 ,w__10164);
  and g__11446(w__10358 ,w__10159 ,w__10157);
  or g__11447(w__10357 ,w__10232 ,w__10162);
  and g__11448(w__10356 ,w__10242 ,w__10240);
  and g__11449(w__10355 ,w__9461 ,w__10156);
  and g__11450(w__10354 ,w__10222 ,w__10218);
  or g__11451(w__10353 ,w__9884 ,w__10166);
  and g__11452(w__10352 ,w__9653 ,w__10237);
  and g__11453(w__10351 ,w__9884 ,w__10166);
  or g__11454(w__10350 ,w__10235 ,w__10234);
  or g__11455(w__10349 ,w__10220 ,w__10138);
  and g__11456(w__10348 ,w__10235 ,w__10234);
  or g__11457(w__10347 ,w__9460 ,w__10231);
  and g__11458(w__10346 ,w__9889 ,w__10172);
  and g__11459(w__10345 ,w__9623 ,w__10231);
  and g__11460(w__10344 ,w__10217 ,w__10216);
  or g__11461(w__10343 ,w__9388 ,w__10219);
  or g__11462(w__10342 ,w__10228 ,w__10224);
  or g__11463(w__10341 ,w__10225 ,w__10223);
  or g__11464(w__10340 ,w__10222 ,w__10218);
  and g__11465(w__10339 ,w__10225 ,w__10223);
  and g__11466(w__10338 ,w__10239 ,w__10233);
  and g__11467(w__10337 ,w__10228 ,w__10224);
  or g__11468(w__10336 ,w__10217 ,w__10216);
  and g__11469(w__10390 ,w__10118 ,w__10183);
  and g__11470(w__10389 ,w__10120 ,w__10198);
  not g__11471(w__10333 ,w__10334);
  not g__11472(w__10332 ,w__10331);
  not g__11473(w__10330 ,w__10329);
  or g__11474(w__10328 ,w__10208 ,w__10215);
  and g__11475(w__10327 ,w__9621 ,w__10136);
  or g__11476(w__10326 ,w__9883 ,w__10213);
  and g__11477(w__10325 ,w__9883 ,w__10213);
  and g__11478(w__10324 ,w__10208 ,w__10215);
  and g__11479(w__10323 ,w__10238 ,w__10243);
  or g__11480(w__10322 ,w__9885 ,w__10257);
  or g__11481(w__10321 ,w__9458 ,w__10146);
  nor g__11482(w__10320 ,w__9621 ,w__10136);
  or g__11483(w__10319 ,w__10168 ,w__10135);
  and g__11484(w__10318 ,w__9622 ,w__10146);
  or g__11485(w__10317 ,w__10142 ,w__10167);
  and g__11486(w__10316 ,w__10168 ,w__10135);
  and g__11487(w__10315 ,w__9630 ,w__10250);
  and g__11488(w__10314 ,w__10142 ,w__10167);
  and g__11489(w__10313 ,w__9885 ,w__10257);
  nor g__11490(w__10312 ,w__10141 ,w__10161);
  and g__11491(w__10311 ,w__10155 ,w__10171);
  or g__11492(w__10310 ,w__9627 ,w__10156);
  or g__11493(w__10309 ,w__10145 ,w__10143);
  or g__11494(w__10308 ,w__9887 ,w__10139);
  and g__11495(w__10307 ,w__9887 ,w__10139);
  and g__11496(w__10306 ,w__10150 ,w__10130);
  and g__11497(w__10305 ,w__10220 ,w__10138);
  nor g__11498(w__10304 ,w__9889 ,w__10172);
  and g__11499(w__10303 ,w__10165 ,w__10132);
  or g__11500(w__10302 ,w__10150 ,w__10130);
  or g__11501(w__10301 ,w__10133 ,w__10173);
  or g__11502(w__10300 ,w__10165 ,w__10132);
  or g__11503(w__10299 ,w__10154 ,w__10158);
  and g__11504(w__10298 ,w__9388 ,w__10219);
  and g__11505(w__10297 ,w__10145 ,w__10143);
  or g__11506(w__10296 ,w__10159 ,w__10157);
  nor g__11507(w__10295 ,w__9629 ,w__10170);
  nor g__11508(w__10294 ,w__10134 ,w__10174);
  or g__11509(w__10293 ,w__10151 ,w__10214);
  and g__11510(w__10292 ,w__10153 ,w__10144);
  or g__11511(w__10291 ,w__10153 ,w__10144);
  or g__11512(w__10290 ,w__10155 ,w__10171);
  or g__11513(w__10289 ,w__9625 ,w__10148);
  and g__11514(w__10288 ,w__9467 ,w__10152);
  or g__11515(w__10287 ,w__9463 ,w__10147);
  nor g__11516(w__10286 ,w__9626 ,w__10149);
  nor g__11517(w__10285 ,w__9467 ,w__10152);
  and g__11518(w__10284 ,w__9652 ,w__10147);
  or g__11519(w__10283 ,w__9465 ,w__9390);
  and g__11520(w__10282 ,w__9654 ,w__9390);
  or g__11521(w__10281 ,w__9459 ,w__9384);
  and g__11522(w__10280 ,w__9624 ,w__10127);
  or g__11523(w__10279 ,w__9628 ,w__10169);
  and g__11524(w__13176 ,w__10126 ,w__10204);
  and g__11525(w__10335 ,w__10124 ,w__10186);
  and g__11526(w__10334 ,w__10116 ,w__10195);
  and g__11527(w__10331 ,w__10122 ,w__10176);
  and g__11528(w__10329 ,w__10114 ,w__10179);
  not g__11529(w__10253 ,w__10254);
  not g__11530(w__10251 ,w__10252);
  not g__11531(w__10229 ,w__10230);
  not g__11532(w__10210 ,w__10211);
  not g__11533(w__10208 ,w__10209);
  not g__11534(w__10207 ,w__10206);
  or g__11535(w__10205 ,w__9896 ,w__9999);
  and g__11536(w__10278 ,w__9924 ,w__10028);
  and g__11537(w__10277 ,w__9947 ,w__10002);
  and g__11538(w__10276 ,w__9958 ,w__10041);
  and g__11539(w__10275 ,w__9835 ,w__9992);
  and g__11540(w__10274 ,w__9847 ,w__10005);
  and g__11541(w__10273 ,w__9946 ,w__10074);
  and g__11542(w__10272 ,w__9943 ,w__10075);
  and g__11543(w__10271 ,w__9942 ,w__10070);
  and g__11544(w__10270 ,w__9829 ,w__9980);
  and g__11545(w__10269 ,w__9940 ,w__10001);
  and g__11546(w__10268 ,w__9932 ,w__10056);
  and g__11547(w__10267 ,w__9934 ,w__10063);
  and g__11548(w__10266 ,w__9953 ,w__10061);
  and g__11549(w__10265 ,w__9929 ,w__10059);
  and g__11550(w__10264 ,w__9903 ,w__10054);
  and g__11551(w__10263 ,w__9938 ,w__10038);
  and g__11552(w__10262 ,w__9914 ,w__10111);
  and g__11553(w__10261 ,w__9918 ,w__10047);
  and g__11554(w__10260 ,w__9923 ,w__10020);
  and g__11555(w__10259 ,w__9873 ,w__10087);
  and g__11556(w__10258 ,w__9945 ,w__10073);
  and g__11557(w__10257 ,w__9866 ,w__10026);
  and g__11558(w__10256 ,w__9910 ,w__10085);
  or g__11559(w__10255 ,w__9892 ,w__9998);
  and g__11560(w__10254 ,w__9857 ,w__10068);
  and g__11561(w__10252 ,w__9859 ,w__10067);
  or g__11562(w__10250 ,w__9901 ,w__9995);
  and g__11563(w__10249 ,w__9936 ,w__10064);
  or g__11564(w__10248 ,w__9899 ,w__9997);
  and g__11565(w__10247 ,w__9951 ,w__10065);
  and g__11566(w__10246 ,w__9952 ,w__10082);
  and g__11567(w__10245 ,w__9935 ,w__10062);
  and g__11568(w__10244 ,w__9949 ,w__10081);
  and g__11569(w__10243 ,w__9915 ,w__10039);
  and g__11570(w__10242 ,w__9930 ,w__10006);
  and g__11571(w__10241 ,w__9844 ,w__10078);
  and g__11572(w__10240 ,w__9830 ,w__9988);
  or g__11573(w__10239 ,w__9894 ,w__9996);
  and g__11574(w__10238 ,w__9911 ,w__10040);
  and g__11575(w__10237 ,w__9839 ,w__9987);
  and g__11576(w__10236 ,w__9845 ,w__10060);
  and g__11577(w__10235 ,w__9922 ,w__10052);
  and g__11578(w__10234 ,w__9921 ,w__10051);
  and g__11579(w__10233 ,w__9837 ,w__9989);
  and g__11580(w__10232 ,w__9849 ,w__10024);
  and g__11581(w__10231 ,w__9860 ,w__10090);
  and g__11582(w__10230 ,w__9916 ,w__10098);
  and g__11583(w__10228 ,w__9863 ,w__10104);
  and g__11584(w__10227 ,w__9944 ,w__10076);
  and g__11585(w__10226 ,w__9919 ,w__10112);
  and g__11586(w__10225 ,w__9906 ,w__10086);
  and g__11587(w__10224 ,w__9913 ,w__10108);
  and g__11588(w__10223 ,w__9876 ,w__9977);
  or g__11589(w__10222 ,w__9890 ,w__9994);
  or g__11590(w__10221 ,w__9897 ,w__9993);
  and g__11591(w__10220 ,w__9875 ,w__10008);
  and g__11592(w__10219 ,w__9831 ,w__9991);
  and g__11593(w__10218 ,w__9904 ,w__10044);
  and g__11594(w__10217 ,w__9867 ,w__10037);
  and g__11595(w__10216 ,w__9905 ,w__10045);
  and g__11596(w__10215 ,w__9836 ,w__9984);
  and g__11597(w__10214 ,w__9862 ,w__10049);
  and g__11598(w__10213 ,w__9955 ,w__10043);
  and g__11599(w__10212 ,w__9950 ,w__10042);
  and g__11600(w__10211 ,w__9841 ,w__9990);
  and g__11601(w__10209 ,w__9927 ,w__10058);
  and g__11602(w__10206 ,w__9908 ,w__10046);
  not g__11603(w__10198 ,w__10197);
  not g__11604(w__10195 ,w__10194);
  not g__11605(w__10186 ,w__10185);
  not g__11606(w__10183 ,w__10182);
  not g__11607(w__10176 ,w__10175);
  not g__11608(w__10173 ,w__10174);
  not g__11609(w__10169 ,w__10170);
  not g__11610(w__10160 ,w__10161);
  not g__11611(w__10148 ,w__10149);
  not g__11612(w__10140 ,w__10141);
  not g__11613(w__10133 ,w__10134);
  not g__11614(w__10130 ,w__10129);
  not g__11615(w__10128 ,w__10127);
  or g__11616(w__13242 ,w__9970 ,w__10101);
  or g__11617(w__13243 ,w__9964 ,w__10077);
  or g__11618(w__13177 ,w__9956 ,w__10011);
  or g__11619(w__10204 ,w__9971 ,w__10093);
  and g__11620(w__10203 ,w__9925 ,w__10057);
  and g__11621(w__10202 ,w__9917 ,w__10021);
  and g__11622(w__10201 ,w__9974 ,w__10083);
  and g__11623(w__10200 ,w__9833 ,w__9986);
  and g__11624(w__10199 ,w__9854 ,w__10012);
  and g__11625(w__10197 ,w__9868 ,w__10103);
  and g__11626(w__10196 ,w__9961 ,w__10099);
  and g__11627(w__10194 ,w__9960 ,w__10092);
  and g__11628(w__10193 ,w__9843 ,w__9983);
  and g__11629(w__10192 ,w__9898 ,w__10096);
  and g__11630(w__10191 ,w__9832 ,w__9981);
  and g__11631(w__10190 ,w__9926 ,w__10089);
  and g__11632(w__10189 ,w__9972 ,w__10109);
  and g__11633(w__10188 ,w__9973 ,w__10097);
  and g__11634(w__10187 ,w__9968 ,w__10106);
  and g__11635(w__10185 ,w__9967 ,w__10105);
  and g__11636(w__10184 ,w__9969 ,w__10100);
  and g__11637(w__10182 ,w__9965 ,w__10107);
  and g__11638(w__10181 ,w__9963 ,w__10102);
  and g__11639(w__10180 ,w__9962 ,w__10110);
  or g__11640(w__10179 ,w__9937 ,w__10095);
  and g__11641(w__10178 ,w__9966 ,w__10094);
  and g__11642(w__10177 ,w__9834 ,w__9982);
  and g__11643(w__10175 ,w__9907 ,w__10034);
  and g__11644(w__10174 ,w__9912 ,w__10013);
  and g__11645(w__10172 ,w__9856 ,w__10015);
  and g__11646(w__10171 ,w__9920 ,w__10079);
  or g__11647(w__10170 ,w__9631 ,w__10091);
  and g__11648(w__10168 ,w__9928 ,w__10033);
  and g__11649(w__10167 ,w__9948 ,w__10069);
  and g__11650(w__10166 ,w__9874 ,w__10055);
  and g__11651(w__10165 ,w__9846 ,w__10066);
  and g__11652(w__10164 ,w__9869 ,w__10029);
  and g__11653(w__10163 ,w__9870 ,w__10027);
  and g__11654(w__10162 ,w__9954 ,w__10031);
  and g__11655(w__10161 ,w__9858 ,w__10030);
  and g__11656(w__10159 ,w__9855 ,w__10003);
  and g__11657(w__10158 ,w__9850 ,w__10084);
  and g__11658(w__10157 ,w__9840 ,w__10048);
  and g__11659(w__10156 ,w__9864 ,w__10007);
  and g__11660(w__10155 ,w__9853 ,w__10035);
  and g__11661(w__10154 ,w__9848 ,w__10004);
  and g__11662(w__10153 ,w__9933 ,w__10080);
  and g__11663(w__10152 ,w__9902 ,w__10088);
  and g__11664(w__10151 ,w__9891 ,w__10072);
  and g__11665(w__10150 ,w__9895 ,w__10053);
  and g__11666(w__10149 ,w__9900 ,w__10071);
  and g__11667(w__10147 ,w__9893 ,w__10010);
  and g__11668(w__10146 ,w__9872 ,w__10036);
  and g__11669(w__10145 ,w__9957 ,w__10023);
  and g__11670(w__10144 ,w__9842 ,w__9978);
  and g__11671(w__10143 ,w__9871 ,w__10022);
  and g__11672(w__10141 ,w__9865 ,w__10025);
  and g__11673(w__10139 ,w__9931 ,w__10018);
  and g__11674(w__10138 ,w__9909 ,w__10017);
  and g__11675(w__10137 ,w__9939 ,w__10016);
  or g__11676(w__10136 ,w__9896 ,w__9985);
  and g__11677(w__10135 ,w__9941 ,w__10032);
  and g__11678(w__10134 ,w__9959 ,w__10014);
  and g__11679(w__10132 ,w__9838 ,w__9979);
  and g__11680(w__10131 ,w__9851 ,w__10019);
  and g__11681(w__10129 ,w__9852 ,w__10050);
  and g__11682(w__10127 ,w__9861 ,w__10009);
  not g__11683(w__10126 ,w__10125);
  not g__11684(w__10124 ,w__10123);
  not g__11685(w__10122 ,w__10121);
  not g__11686(w__10120 ,w__10119);
  not g__11687(w__10118 ,w__10117);
  not g__11688(w__10116 ,w__10115);
  not g__11689(w__10114 ,w__10113);
  or g__11690(w__10112 ,w__9716 ,w__9302);
  or g__11691(w__10111 ,w__9730 ,w__9287);
  or g__11692(w__10110 ,w__9692 ,w__9261);
  or g__11693(w__10109 ,w__9680 ,w__9353);
  or g__11694(w__10108 ,w__9788 ,w__9284);
  or g__11695(w__10107 ,w__9685 ,w__9261);
  or g__11696(w__10106 ,w__9687 ,w__9328);
  or g__11697(w__10105 ,w__9681 ,w__9349);
  or g__11698(w__10104 ,w__9678 ,w__9344);
  or g__11699(w__10103 ,w__9713 ,w__9280);
  or g__11700(w__10102 ,w__9689 ,w__9350);
  nor g__11701(w__10101 ,w__9352 ,w__9682);
  or g__11702(w__10100 ,w__9683 ,w__9328);
  or g__11703(w__10099 ,w__9688 ,w__9329);
  or g__11704(w__10098 ,w__9684 ,w__9341);
  or g__11705(w__10097 ,w__9690 ,w__9352);
  or g__11706(w__10096 ,w__9739 ,w__9346);
  nor g__11707(w__10095 ,w__9350 ,w__9694);
  or g__11708(w__10094 ,w__9691 ,w__9380);
  nor g__11709(w__10093 ,w__9353 ,w__9693);
  or g__11710(w__10092 ,w__9686 ,w__9379);
  nor g__11711(w__10091 ,w__9349 ,w__9679);
  or g__11712(w__10090 ,w__9809 ,w__9293);
  or g__11713(w__10089 ,w__9765 ,w__9272);
  or g__11714(w__10088 ,w__9766 ,w__9320);
  or g__11715(w__10087 ,w__9811 ,w__9299);
  or g__11716(w__10086 ,w__9775 ,w__9296);
  or g__11717(w__10085 ,w__9740 ,w__9314);
  or g__11718(w__10084 ,w__9698 ,w__9343);
  or g__11719(w__10083 ,w__9703 ,w__9275);
  or g__11720(w__10082 ,w__9770 ,w__9319);
  or g__11721(w__10081 ,w__9792 ,w__9361);
  or g__11722(w__10080 ,w__9727 ,w__9355);
  or g__11723(w__10079 ,w__9781 ,w__9278);
  or g__11724(w__10078 ,w__9806 ,w__9317);
  nor g__11725(w__10077 ,w__9329 ,w__9656);
  or g__11726(w__10076 ,w__9787 ,w__9373);
  or g__11727(w__10075 ,w__9771 ,w__9313);
  or g__11728(w__10074 ,w__9735 ,w__9274);
  or g__11729(w__10073 ,w__9705 ,w__9358);
  or g__11730(w__10072 ,w__9797 ,w__9340);
  or g__11731(w__10071 ,w__9789 ,w__9269);
  or g__11732(w__10070 ,w__9782 ,w__9277);
  or g__11733(w__10069 ,w__9791 ,w__9296);
  or g__11734(w__10068 ,w__9812 ,w__9272);
  or g__11735(w__10067 ,w__9783 ,w__9298);
  or g__11736(w__10066 ,w__9715 ,w__9295);
  or g__11737(w__10065 ,w__9658 ,w__9271);
  or g__11738(w__10064 ,w__9779 ,w__9287);
  or g__11739(w__10063 ,w__9780 ,w__9316);
  or g__11740(w__10062 ,w__9784 ,w__9286);
  or g__11741(w__10061 ,w__9774 ,w__9370);
  or g__11742(w__10060 ,w__9810 ,w__9364);
  or g__11743(w__10059 ,w__9772 ,w__9295);
  or g__11744(w__10058 ,w__9769 ,w__9278);
  or g__11745(w__10057 ,w__9723 ,w__9286);
  or g__11746(w__10056 ,w__9721 ,w__9271);
  or g__11747(w__10055 ,w__9731 ,w__9268);
  or g__11748(w__10054 ,w__9733 ,w__9346);
  or g__11749(w__10053 ,w__9697 ,w__9313);
  or g__11750(w__10052 ,w__9776 ,w__9299);
  or g__11751(w__10051 ,w__9795 ,w__9358);
  or g__11752(w__10050 ,w__9773 ,w__9343);
  or g__11753(w__10049 ,w__9736 ,w__9284);
  or g__11754(w__10125 ,w__9616 ,w__9827);
  or g__11755(w__10123 ,w__9641 ,w__9824);
  or g__11756(w__10121 ,w__9609 ,w__9825);
  or g__11757(w__10119 ,w__9614 ,w__9823);
  or g__11758(w__10117 ,w__9612 ,w__9822);
  or g__11759(w__10115 ,w__9617 ,w__9828);
  or g__11760(w__10113 ,w__9606 ,w__9826);
  or g__11761(w__10048 ,w__9751 ,w__9304);
  or g__11762(w__10047 ,w__9712 ,w__9275);
  or g__11763(w__10046 ,w__9718 ,w__9319);
  or g__11764(w__10045 ,w__9728 ,w__9292);
  or g__11765(w__10044 ,w__9720 ,w__9283);
  or g__11766(w__10043 ,w__9798 ,w__9283);
  or g__11767(w__10042 ,w__9793 ,w__9269);
  or g__11768(w__10041 ,w__9741 ,w__9255);
  or g__11769(w__10040 ,w__9729 ,w__9277);
  or g__11770(w__10039 ,w__9801 ,w__9302);
  or g__11771(w__10038 ,w__9706 ,w__9355);
  or g__11772(w__10037 ,w__9659 ,w__9298);
  or g__11773(w__10036 ,w__9726 ,w__9362);
  or g__11774(w__10035 ,w__9777 ,w__9373);
  or g__11775(w__10034 ,w__9799 ,w__9281);
  or g__11776(w__10033 ,w__9746 ,w__9257);
  or g__11777(w__10032 ,w__9696 ,w__9316);
  or g__11778(w__10031 ,w__9804 ,w__9301);
  or g__11779(w__10030 ,w__9711 ,w__9255);
  or g__11780(w__10029 ,w__9695 ,w__9331);
  or g__11781(w__10028 ,w__9737 ,w__9301);
  or g__11782(w__10027 ,w__9719 ,w__9293);
  or g__11783(w__10026 ,w__9708 ,w__9364);
  or g__11784(w__10025 ,w__9725 ,w__9340);
  or g__11785(w__10024 ,w__9707 ,w__9257);
  or g__11786(w__10023 ,w__9655 ,w__9268);
  or g__11787(w__10022 ,w__9808 ,w__9332);
  or g__11788(w__10021 ,w__9709 ,w__9331);
  or g__11789(w__10020 ,w__9701 ,w__9370);
  or g__11790(w__10019 ,w__9768 ,w__9359);
  or g__11791(w__10018 ,w__9722 ,w__9281);
  or g__11792(w__10017 ,w__9778 ,w__9292);
  or g__11793(w__10016 ,w__9786 ,w__9249);
  or g__11794(w__10015 ,w__9717 ,w__9347);
  or g__11795(w__10014 ,w__9743 ,w__9249);
  or g__11796(w__10013 ,w__9807 ,w__9280);
  or g__11797(w__10012 ,w__9702 ,w__9253);
  nor g__11798(w__10011 ,w__9347 ,w__9748);
  or g__11799(w__10010 ,w__9732 ,w__9259);
  or g__11800(w__10009 ,w__9805 ,w__9259);
  or g__11801(w__10008 ,w__9734 ,w__9356);
  or g__11802(w__10007 ,w__9724 ,w__9274);
  or g__11803(w__10006 ,w__9700 ,w__9247);
  or g__11804(w__10005 ,w__9699 ,w__9361);
  or g__11805(w__10004 ,w__9814 ,w__9247);
  or g__11806(w__10003 ,w__9710 ,w__9253);
  or g__11807(w__10002 ,w__9714 ,w__9374);
  or g__11808(w__10001 ,w__9704 ,w__9371);
  nor g__11809(w__9999 ,w__9338 ,w__9308);
  nor g__11810(w__9998 ,w__9344 ,w__9593);
  nor g__11811(w__9997 ,w__9317 ,w__9596);
  nor g__11812(w__9996 ,w__9314 ,w__9594);
  nor g__11813(w__9995 ,w__9320 ,w__9581);
  nor g__11814(w__9994 ,w__9341 ,w__9595);
  nor g__11815(w__9993 ,w__9332 ,w__9597);
  or g__11816(w__9992 ,w__9803 ,w__9305);
  or g__11817(w__9991 ,w__9800 ,w__9310);
  or g__11818(w__9990 ,w__9794 ,w__9307);
  or g__11819(w__9989 ,w__9802 ,w__9304);
  or g__11820(w__9988 ,w__9790 ,w__9305);
  or g__11821(w__9987 ,w__9816 ,w__9245);
  or g__11822(w__9986 ,w__9767 ,w__9377);
  nor g__11823(w__9985 ,w__9311 ,w__9785);
  or g__11824(w__9984 ,w__9796 ,w__9310);
  or g__11825(w__9983 ,w__9813 ,w__9307);
  or g__11826(w__9982 ,w__9818 ,w__9311);
  or g__11827(w__9981 ,w__9819 ,w__9376);
  or g__11828(w__9980 ,w__9817 ,w__9376);
  or g__11829(w__9979 ,w__9820 ,w__9308);
  or g__11830(w__9978 ,w__9815 ,w__9245);
  or g__11831(w__9977 ,w__9738 ,w__9365);
  or g__11832(w__9974 ,w__9787 ,w__9505);
  or g__11833(w__9973 ,w__9335 ,w__9681);
  or g__11834(w__9972 ,w__9323 ,w__9686);
  nor g__11835(w__9971 ,w__9335 ,w__9691);
  nor g__11836(w__9970 ,w__9323 ,w__9693);
  or g__11837(w__9969 ,w__9322 ,w__9687);
  or g__11838(w__9968 ,w__9334 ,w__9685);
  or g__11839(w__9967 ,w__9325 ,w__9688);
  or g__11840(w__9966 ,w__9334 ,w__9694);
  or g__11841(w__9965 ,w__9322 ,w__9680);
  nor g__11842(w__9964 ,w__9326 ,w__9682);
  or g__11843(w__9963 ,w__9325 ,w__9692);
  or g__11844(w__9962 ,w__9326 ,w__9683);
  or g__11845(w__9961 ,w__9263 ,w__9689);
  or g__11846(w__9960 ,w__9263 ,w__9679);
  or g__11847(w__9959 ,w__9786 ,w__9544);
  or g__11848(w__9958 ,w__9713 ,w__9529);
  or g__11849(w__9957 ,w__9708 ,w__9493);
  nor g__11850(w__9956 ,w__9717 ,w__9536);
  or g__11851(w__9955 ,w__9738 ,w__9502);
  or g__11852(w__9954 ,w__9778 ,w__9547);
  or g__11853(w__9953 ,w__9716 ,w__9547);
  or g__11854(w__9952 ,w__9721 ,w__9514);
  or g__11855(w__9951 ,w__9812 ,w__9514);
  or g__11856(w__9950 ,w__9788 ,w__9502);
  or g__11857(w__9949 ,w__9699 ,w__9535);
  or g__11858(w__9948 ,w__9769 ,w__9517);
  or g__11859(w__9947 ,w__9718 ,w__9506);
  or g__11860(w__9946 ,w__9766 ,w__9509);
  or g__11861(w__9945 ,w__9740 ,w__9523);
  or g__11862(w__9944 ,w__9724 ,w__9505);
  or g__11863(w__9943 ,w__9707 ,w__9523);
  or g__11864(w__9942 ,w__9697 ,w__9518);
  or g__11865(w__9941 ,w__9798 ,w__9494);
  or g__11866(w__9940 ,w__9797 ,w__9545);
  or g__11867(w__9939 ,w__9701 ,w__9544);
  or g__11868(w__9938 ,w__9727 ,w__9469);
  nor g__11869(w__9937 ,w__9408 ,w__9690);
  or g__11870(w__9936 ,w__9805 ,w__9478);
  or g__11871(w__9935 ,w__9783 ,w__9478);
  or g__11872(w__9934 ,w__9736 ,w__9497);
  or g__11873(w__9933 ,w__9723 ,w__9470);
  or g__11874(w__9932 ,w__9814 ,w__9508);
  or g__11875(w__9931 ,w__9808 ,w__9530);
  or g__11876(w__9930 ,w__9765 ,w__9511);
  or g__11877(w__9929 ,w__9771 ,w__9521);
  or g__11878(w__9928 ,w__9729 ,w__9517);
  or g__11879(w__9927 ,w__9705 ,w__9520);
  or g__11880(w__9926 ,w__9777 ,w__9511);
  or g__11881(w__9925 ,w__9773 ,w__9473);
  or g__11882(w__9924 ,w__9809 ,w__9541);
  or g__11883(w__9923 ,w__9725 ,w__9672);
  or g__11884(w__9922 ,w__9784 ,w__9469);
  or g__11885(w__9921 ,w__9772 ,w__9526);
  or g__11886(w__9920 ,w__9768 ,w__9526);
  or g__11887(w__9919 ,w__9804 ,w__9541);
  or g__11888(w__9918 ,w__9700 ,w__9508);
  or g__11889(w__9917 ,w__9726 ,w__9533);
  or g__11890(w__9916 ,w__9774 ,w__9542);
  or g__11891(w__9915 ,w__9728 ,w__9545);
  or g__11892(w__9914 ,w__9732 ,w__9472);
  or g__11893(w__9913 ,w__9780 ,w__9493);
  or g__11894(w__9912 ,w__9722 ,w__9529);
  or g__11895(w__9911 ,w__9775 ,w__9520);
  or g__11896(w__9910 ,w__9781 ,w__9524);
  or g__11897(w__9909 ,w__9737 ,w__9548);
  or g__11898(w__9908 ,w__9735 ,w__9515);
  or g__11899(w__9907 ,w__9741 ,w__9532);
  or g__11900(w__9906 ,w__9795 ,w__9521);
  or g__11901(w__9905 ,w__9684 ,w__9438);
  or g__11902(w__9904 ,w__9789 ,w__9496);
  or g__11903(w__9903 ,w__9695 ,w__9539);
  or g__11904(w__9976 ,w__9661 ,w__9397);
  or g__11905(w__9975 ,in21[0] ,w__9750);
  not g__11906(w__9902 ,w__9901);
  not g__11907(w__9900 ,w__9899);
  not g__11908(w__9898 ,w__9897);
  not g__11909(w__9895 ,w__9894);
  not g__11910(w__9893 ,w__9892);
  not g__11911(w__9891 ,w__9890);
  not g__11912(w__9889 ,w__9888);
  or g__11913(w__9876 ,w__9731 ,w__9499);
  or g__11914(w__9875 ,w__9698 ,w__9475);
  or g__11915(w__9874 ,w__9810 ,w__9499);
  or g__11916(w__9873 ,w__9734 ,w__9475);
  or g__11917(w__9872 ,w__9739 ,w__9538);
  or g__11918(w__9871 ,w__9711 ,w__9532);
  or g__11919(w__9870 ,w__9801 ,w__9438);
  or g__11920(w__9869 ,w__9792 ,w__9535);
  or g__11921(w__9868 ,w__9733 ,w__9533);
  or g__11922(w__9867 ,w__9776 ,w__9472);
  or g__11923(w__9866 ,w__9696 ,w__9496);
  or g__11924(w__9865 ,w__9719 ,w__9548);
  or g__11925(w__9864 ,w__9714 ,w__9509);
  or g__11926(w__9863 ,w__9779 ,w__9479);
  or g__11927(w__9862 ,w__9720 ,w__9503);
  or g__11928(w__9861 ,w__9706 ,w__9473);
  or g__11929(w__9860 ,w__9704 ,w__9542);
  or g__11930(w__9859 ,w__9811 ,w__9476);
  or g__11931(w__9858 ,w__9799 ,w__9538);
  or g__11932(w__9857 ,w__9770 ,w__9512);
  or g__11933(w__9856 ,w__9807 ,w__9530);
  or g__11934(w__9855 ,w__9702 ,w__9497);
  or g__11935(w__9854 ,w__9793 ,w__9500);
  or g__11936(w__9853 ,w__9703 ,w__9506);
  or g__11937(w__9852 ,w__9730 ,w__9470);
  or g__11938(w__9851 ,w__9782 ,w__9527);
  or g__11939(w__9850 ,w__9678 ,w__9479);
  or g__11940(w__9849 ,w__9715 ,w__9518);
  or g__11941(w__9848 ,w__9712 ,w__9515);
  or g__11942(w__9847 ,w__9709 ,w__9536);
  or g__11943(w__9846 ,w__9791 ,w__9524);
  or g__11944(w__9845 ,w__9806 ,w__9494);
  or g__11945(w__9844 ,w__9710 ,w__9503);
  or g__11946(w__9843 ,w__9481 ,w__9800);
  or g__11947(w__9842 ,w__9490 ,w__9816);
  or g__11948(w__9841 ,w__9490 ,w__9767);
  or g__11949(w__9840 ,w__9482 ,w__9820);
  or g__11950(w__9839 ,w__9485 ,w__9817);
  or g__11951(w__9838 ,w__9481 ,w__9818);
  or g__11952(w__9837 ,w__9484 ,w__9813);
  or g__11953(w__9836 ,w__9487 ,w__9790);
  or g__11954(w__9835 ,w__9487 ,w__9819);
  or g__11955(w__9834 ,w__9484 ,w__9796);
  or g__11956(w__9833 ,w__9491 ,w__9785);
  or g__11957(w__9832 ,w__9485 ,w__9815);
  or g__11958(w__9831 ,w__9488 ,w__9794);
  or g__11959(w__9830 ,w__9482 ,w__9803);
  or g__11960(w__9829 ,w__9491 ,w__9802);
  or g__11961(w__9828 ,w__9368 ,w__9754);
  or g__11962(w__9827 ,w__9597 ,w__9757);
  or g__11963(w__9826 ,w__9595 ,w__9758);
  or g__11964(w__9825 ,w__9594 ,w__9756);
  or g__11965(w__9824 ,w__9596 ,w__9752);
  or g__11966(w__9823 ,w__9593 ,w__9753);
  or g__11967(w__9822 ,w__9581 ,w__9755);
  nor g__11968(w__9821 ,w__9539 ,w__9234);
  and g__11969(w__9901 ,in21[13] ,w__9400);
  and g__11970(w__9899 ,in21[7] ,w__9398);
  and g__11971(w__9897 ,in21[3] ,w__9391);
  and g__11972(w__9896 ,in21[15] ,w__9399);
  and g__11973(w__9894 ,in21[9] ,w__9402);
  and g__11974(w__9892 ,in21[11] ,w__9396);
  and g__11975(w__9890 ,in21[5] ,w__9392);
  and g__11976(w__9888 ,in20[0] ,w__9406);
  or g__11977(w__9887 ,w__9382 ,w__9500);
  or g__11978(w__9886 ,w__9382 ,w__9488);
  or g__11979(w__9885 ,w__9598 ,w__9527);
  or g__11980(w__9884 ,w__9381 ,w__9512);
  or g__11981(w__9883 ,w__9381 ,w__9476);
  or g__11982(w__9882 ,w__9749 ,w__9394);
  or g__11983(w__9881 ,w__9744 ,w__9403);
  or g__11984(w__9880 ,w__9742 ,w__9393);
  or g__11985(w__9879 ,w__9657 ,w__9405);
  or g__11986(w__9878 ,w__9745 ,w__9401);
  or g__11987(w__9877 ,w__9660 ,w__9395);
  not g__11988(w__9764 ,w__9398);
  not g__11989(w__9763 ,w__9403);
  not g__11990(w__9761 ,w__9397);
  not g__11991(w__9760 ,w__9399);
  nor g__11992(w__9758 ,w__9446 ,w__9644);
  nor g__11993(w__9757 ,w__9582 ,w__9607);
  nor g__11994(w__9756 ,w__9444 ,w__9613);
  nor g__11995(w__9755 ,w__9442 ,w__9646);
  nor g__11996(w__9754 ,w__9440 ,w__9608);
  nor g__11997(w__9753 ,w__9448 ,w__9633);
  nor g__11998(w__9752 ,w__9450 ,w__9638);
  or g__11999(w__9751 ,w__9629 ,w__9618);
  xnor g__12000(w__9749 ,in21[13] ,in21[12]);
  xnor g__12001(w__9748 ,in20[0] ,in21[3]);
  nor g__12002(w__9747 ,w__13180 ,w__9452);
  xnor g__12003(w__9746 ,in20[0] ,in21[9]);
  xnor g__12004(w__9745 ,in21[9] ,in21[8]);
  xnor g__12005(w__9744 ,in21[7] ,in21[6]);
  xnor g__12006(w__9743 ,in20[0] ,in21[5]);
  xnor g__12007(w__9742 ,in21[3] ,in21[2]);
  or g__12008(w__9820 ,w__9550 ,w__9637);
  or g__12009(w__9819 ,w__9625 ,w__9634);
  or g__12010(w__9818 ,w__9551 ,w__9647);
  or g__12011(w__9817 ,w__9561 ,w__9642);
  or g__12012(w__9816 ,w__9553 ,w__9639);
  or g__12013(w__9815 ,w__9560 ,w__9635);
  xnor g__12014(w__9814 ,in20[4] ,in21[13]);
  or g__12015(w__9813 ,w__9558 ,w__9610);
  xnor g__12016(w__9812 ,in20[1] ,in21[13]);
  xnor g__12017(w__9811 ,in20[4] ,in21[11]);
  xnor g__12018(w__9810 ,in20[6] ,in21[7]);
  xnor g__12019(w__9809 ,in20[13] ,in21[5]);
  xnor g__12020(w__9808 ,in20[4] ,in21[3]);
  xnor g__12021(w__9807 ,in20[2] ,in21[3]);
  xnor g__12022(w__9806 ,in20[7] ,in21[7]);
  xnor g__12023(w__9805 ,in20[9] ,in21[11]);
  xnor g__12024(w__9804 ,in20[10] ,in21[5]);
  or g__12025(w__9803 ,w__9552 ,w__9643);
  or g__12026(w__9802 ,w__9559 ,w__9611);
  xnor g__12027(w__9801 ,in20[5] ,in21[5]);
  or g__12028(w__9800 ,w__9557 ,w__9615);
  xnor g__12029(w__9799 ,in20[6] ,in21[3]);
  xnor g__12030(w__9798 ,in20[3] ,in21[7]);
  xnor g__12031(w__9797 ,in20[15] ,in21[5]);
  or g__12032(w__9796 ,w__9555 ,w__9636);
  xnor g__12033(w__9795 ,in20[3] ,in21[9]);
  or g__12034(w__9794 ,w__9554 ,w__9640);
  xnor g__12035(w__9793 ,in20[10] ,in21[7]);
  xnor g__12036(w__9792 ,in20[11] ,in21[3]);
  xnor g__12037(w__9791 ,in20[8] ,in21[9]);
  or g__12038(w__9790 ,w__9556 ,w__9645);
  xnor g__12039(w__9789 ,in20[15] ,in21[7]);
  xnor g__12040(w__9788 ,in20[11] ,in21[7]);
  xnor g__12041(w__9787 ,in20[10] ,in21[13]);
  xnor g__12042(w__9786 ,in20[1] ,in21[5]);
  xnor g__12043(w__9785 ,in20[15] ,in21[15]);
  xnor g__12044(w__9784 ,in20[2] ,in21[11]);
  xnor g__12045(w__9783 ,in20[3] ,in21[11]);
  xnor g__12046(w__9782 ,in20[14] ,in21[9]);
  xnor g__12047(w__9781 ,in20[12] ,in21[9]);
  xnor g__12048(w__9780 ,in20[12] ,in21[7]);
  xnor g__12049(w__9779 ,in20[8] ,in21[11]);
  xnor g__12050(w__9778 ,in20[11] ,in21[5]);
  xnor g__12051(w__9777 ,in20[8] ,in21[13]);
  xnor g__12052(w__9776 ,in20[1] ,in21[11]);
  xnor g__12053(w__9775 ,in20[2] ,in21[9]);
  xnor g__12054(w__9774 ,in20[8] ,in21[5]);
  xnor g__12055(w__9773 ,in20[13] ,in21[11]);
  xnor g__12056(w__9772 ,in20[4] ,in21[9]);
  xnor g__12057(w__9771 ,in20[5] ,in21[9]);
  xnor g__12058(w__9770 ,in20[2] ,in21[13]);
  xnor g__12059(w__9769 ,in20[9] ,in21[9]);
  xnor g__12060(w__9768 ,in20[13] ,in21[9]);
  or g__12061(w__9767 ,w__9436 ,w__9619);
  xnor g__12062(w__9766 ,in20[15] ,in21[13]);
  xnor g__12063(w__9765 ,in20[7] ,in21[13]);
  xnor g__12064(w__9762 ,w__9450 ,in21[6]);
  xnor g__12065(w__9759 ,w__9440 ,in21[14]);
  not g__12066(w__9677 ,w__9396);
  not g__12067(w__9676 ,w__9395);
  not g__12068(w__9674 ,w__9406);
  not g__12069(w__9672 ,w__9392);
  not g__12070(w__9671 ,w__9405);
  not g__12071(w__9670 ,w__9391);
  not g__12072(w__9669 ,w__9393);
  not g__12073(w__9667 ,w__9402);
  not g__12074(w__9666 ,w__9401);
  not g__12075(w__9664 ,w__9400);
  not g__12076(w__9663 ,w__9394);
  xnor g__12077(w__9661 ,in21[15] ,in21[14]);
  xnor g__12078(w__9660 ,in21[11] ,in21[10]);
  xnor g__12079(w__9659 ,in20[0] ,in21[11]);
  xnor g__12080(w__9658 ,in20[0] ,in21[13]);
  xnor g__12081(w__9657 ,in21[5] ,in21[4]);
  xnor g__12082(w__9656 ,in20[0] ,in21[1]);
  xnor g__12083(w__9655 ,in20[0] ,in21[7]);
  xnor g__12084(w__9741 ,in20[7] ,in21[3]);
  xnor g__12085(w__9740 ,in20[11] ,in21[9]);
  xnor g__12086(w__9739 ,in20[15] ,in21[3]);
  xnor g__12087(w__9738 ,in20[4] ,in21[7]);
  xnor g__12088(w__9737 ,in20[12] ,in21[5]);
  xnor g__12089(w__9736 ,in20[13] ,in21[7]);
  xnor g__12090(w__9735 ,in20[14] ,in21[13]);
  xnor g__12091(w__9734 ,in20[5] ,in21[11]);
  xnor g__12092(w__9733 ,in20[9] ,in21[3]);
  xnor g__12093(w__9732 ,in20[15] ,in21[11]);
  xnor g__12094(w__9731 ,in20[5] ,in21[7]);
  xnor g__12095(w__9730 ,in20[14] ,in21[11]);
  xnor g__12096(w__9729 ,in20[1] ,in21[9]);
  xnor g__12097(w__9728 ,in20[6] ,in21[5]);
  xnor g__12098(w__9727 ,in20[11] ,in21[11]);
  xnor g__12099(w__9726 ,in20[14] ,in21[3]);
  xnor g__12100(w__9725 ,in20[3] ,in21[5]);
  xnor g__12101(w__9724 ,in20[11] ,in21[13]);
  xnor g__12102(w__9723 ,in20[12] ,in21[11]);
  xnor g__12103(w__9722 ,in20[3] ,in21[3]);
  xnor g__12104(w__9721 ,in20[3] ,in21[13]);
  xnor g__12105(w__9720 ,in20[14] ,in21[7]);
  xnor g__12106(w__9719 ,in20[4] ,in21[5]);
  xnor g__12107(w__9718 ,in20[13] ,in21[13]);
  xnor g__12108(w__9717 ,in20[1] ,in21[3]);
  xnor g__12109(w__9716 ,in20[9] ,in21[5]);
  xnor g__12110(w__9715 ,in20[7] ,in21[9]);
  xnor g__12111(w__9714 ,in20[12] ,in21[13]);
  xnor g__12112(w__9713 ,in20[8] ,in21[3]);
  xnor g__12113(w__9712 ,in20[5] ,in21[13]);
  xnor g__12114(w__9711 ,in20[5] ,in21[3]);
  xnor g__12115(w__9710 ,in20[8] ,in21[7]);
  xnor g__12116(w__9709 ,in20[13] ,in21[3]);
  xnor g__12117(w__9708 ,in20[1] ,in21[7]);
  xnor g__12118(w__9707 ,in20[6] ,in21[9]);
  xnor g__12119(w__9706 ,in20[10] ,in21[11]);
  xnor g__12120(w__9705 ,in20[10] ,in21[9]);
  xnor g__12121(w__9704 ,in20[14] ,in21[5]);
  xnor g__12122(w__9703 ,in20[9] ,in21[13]);
  xnor g__12123(w__9702 ,in20[9] ,in21[7]);
  xnor g__12124(w__9701 ,in20[2] ,in21[5]);
  xnor g__12125(w__9700 ,in20[6] ,in21[13]);
  xnor g__12126(w__9699 ,in20[12] ,in21[3]);
  xnor g__12127(w__9698 ,in20[6] ,in21[11]);
  xnor g__12128(w__9697 ,in20[15] ,in21[9]);
  xnor g__12129(w__9696 ,in20[2] ,in21[7]);
  xnor g__12130(w__9695 ,in20[10] ,in21[3]);
  xnor g__12131(w__9694 ,in20[4] ,in21[1]);
  xnor g__12132(w__9693 ,in20[2] ,in21[1]);
  xnor g__12133(w__9692 ,in20[9] ,in21[1]);
  xnor g__12134(w__9691 ,in20[3] ,in21[1]);
  xnor g__12135(w__9690 ,in20[5] ,in21[1]);
  xnor g__12136(w__9689 ,in20[8] ,in21[1]);
  xnor g__12137(w__9688 ,in20[7] ,in21[1]);
  xnor g__12138(w__9687 ,in20[11] ,in21[1]);
  xnor g__12139(w__9686 ,in20[14] ,in21[1]);
  xnor g__12140(w__9685 ,in20[12] ,in21[1]);
  xnor g__12141(w__9684 ,in20[7] ,in21[5]);
  xnor g__12142(w__9683 ,in20[10] ,in21[1]);
  xnor g__12143(w__9682 ,in20[1] ,in21[1]);
  xnor g__12144(w__9681 ,in20[6] ,in21[1]);
  xnor g__12145(w__9680 ,in20[13] ,in21[1]);
  xnor g__12146(w__9679 ,in20[15] ,in21[1]);
  xnor g__12147(w__9678 ,in20[7] ,in21[11]);
  xnor g__12148(w__9675 ,w__9448 ,in21[10]);
  xnor g__12149(w__9673 ,w__9446 ,in21[4]);
  xnor g__12150(w__9668 ,w__9452 ,in21[2]);
  xnor g__12151(w__9665 ,w__9444 ,in21[8]);
  xnor g__12152(w__9662 ,w__9442 ,in21[12]);
  nor g__12153(w__9647 ,in20[2] ,in21[15]);
  nor g__12154(w__9646 ,in20[0] ,in21[12]);
  nor g__12155(w__9645 ,in20[4] ,in21[15]);
  nor g__12156(w__9644 ,in20[0] ,in21[4]);
  nor g__12157(w__9643 ,in20[5] ,in21[15]);
  nor g__12158(w__9642 ,in20[9] ,in21[15]);
  and g__12159(w__9641 ,in20[0] ,in21[6]);
  nor g__12160(w__9640 ,in20[13] ,in21[15]);
  nor g__12161(w__9639 ,in20[8] ,in21[15]);
  nor g__12162(w__9638 ,in20[0] ,in21[6]);
  nor g__12163(w__9637 ,in20[1] ,in21[15]);
  nor g__12164(w__9636 ,in20[3] ,in21[15]);
  nor g__12165(w__9635 ,in20[7] ,in21[15]);
  nor g__12166(w__9634 ,in20[6] ,in21[15]);
  nor g__12167(w__9633 ,in20[0] ,in21[10]);
  or g__12168(w__9632 ,w__9602 ,w__9265);
  or g__12169(w__9654 ,w__9604 ,w__9289);
  or g__12170(w__9653 ,w__9605 ,w__9367);
  or g__12171(w__9652 ,w__9587 ,w__9337);
  or g__12172(w__9651 ,w__9591 ,w__9266);
  or g__12173(w__9650 ,w__9600 ,w__9290);
  or g__12174(w__9649 ,w__9599 ,w__9251);
  or g__12175(w__9648 ,w__9590 ,w__9337);
  not g__12176(w__9628 ,w__9629);
  not g__12177(w__9625 ,w__9626);
  not g__12178(w__9620 ,w__9621);
  nor g__12179(w__9619 ,in20[14] ,in21[15]);
  nor g__12180(w__9618 ,in20[0] ,in21[15]);
  and g__12181(w__9617 ,in20[0] ,in21[14]);
  and g__12182(w__9616 ,in20[0] ,in21[2]);
  nor g__12183(w__9615 ,in20[12] ,in21[15]);
  and g__12184(w__9614 ,in20[0] ,in21[10]);
  nor g__12185(w__9613 ,in20[0] ,in21[8]);
  and g__12186(w__9612 ,in20[0] ,in21[12]);
  nor g__12187(w__9611 ,in20[10] ,in21[15]);
  nor g__12188(w__9610 ,in20[11] ,in21[15]);
  and g__12189(w__9609 ,in20[0] ,in21[8]);
  nor g__12190(w__9608 ,in20[0] ,in21[14]);
  nor g__12191(w__9607 ,in20[0] ,in21[2]);
  and g__12192(w__9606 ,in20[0] ,in21[4]);
  and g__12193(w__13180 ,in20[0] ,in21[0]);
  and g__12194(w__9631 ,in21[1] ,in21[0]);
  or g__12195(w__9630 ,w__9588 ,w__9265);
  and g__12196(w__9629 ,in20[0] ,in21[15]);
  or g__12197(w__9627 ,w__9586 ,w__9289);
  or g__12198(w__9626 ,w__9601 ,w__9367);
  or g__12199(w__9624 ,w__9592 ,w__9290);
  or g__12200(w__9623 ,w__9585 ,w__9266);
  or g__12201(w__9622 ,w__9603 ,w__9251);
  or g__12202(w__9621 ,w__9589 ,w__9338);
  not g__12203(w__9605 ,in20[7]);
  not g__12204(w__9604 ,in20[9]);
  not g__12205(w__9603 ,in20[1]);
  not g__12206(w__9602 ,in20[15]);
  not g__12207(w__9601 ,in20[6]);
  not g__12208(w__9600 ,in20[12]);
  not g__12209(w__9599 ,in20[4]);
  not g__12210(w__9598 ,in20[0]);
  not g__12211(w__9597 ,in21[3]);
  not g__12212(w__9596 ,in21[7]);
  not g__12213(w__9595 ,in21[5]);
  not g__12214(w__9594 ,in21[9]);
  not g__12215(w__9593 ,in21[11]);
  not g__12216(w__9592 ,in20[5]);
  not g__12217(w__9591 ,in20[11]);
  not g__12218(w__9590 ,in20[3]);
  not g__12219(w__9589 ,in20[14]);
  not g__12220(w__9588 ,in20[13]);
  not g__12221(w__9587 ,in20[10]);
  not g__12222(w__9586 ,in20[8]);
  not g__12223(w__9585 ,in20[2]);
  not g__12224(w__9584 ,in21[0]);
  not g__12225(w__9583 ,in21[15]);
  not g__12226(w__9582 ,in21[1]);
  not g__12227(w__9581 ,in21[13]);
  not g__12228(w__9235 ,w__9549);
  not g__12229(w__9549 ,w__9598);
  not g__12230(w__9548 ,w__9546);
  not g__12231(w__9547 ,w__9546);
  not g__12232(w__9546 ,w__9568);
  not g__12233(w__9545 ,w__9543);
  not g__12234(w__9544 ,w__9543);
  not g__12235(w__9543 ,w__9674);
  not g__12236(w__9542 ,w__9540);
  not g__12237(w__9541 ,w__9540);
  not g__12238(w__9540 ,w__9671);
  not g__12239(w__9539 ,w__9537);
  not g__12240(w__9538 ,w__9537);
  not g__12241(w__9537 ,w__9669);
  not g__12242(w__9536 ,w__9534);
  not g__12243(w__9535 ,w__9534);
  not g__12244(w__9534 ,w__9670);
  not g__12245(w__9533 ,w__9531);
  not g__12246(w__9532 ,w__9531);
  not g__12247(w__9531 ,w__9567);
  not g__12248(w__9530 ,w__9528);
  not g__12249(w__9529 ,w__9528);
  not g__12250(w__9528 ,w__9566);
  not g__12251(w__9527 ,w__9525);
  not g__12252(w__9526 ,w__9525);
  not g__12253(w__9525 ,w__9666);
  not g__12254(w__9524 ,w__9522);
  not g__12255(w__9523 ,w__9522);
  not g__12256(w__9522 ,w__9667);
  not g__12257(w__9521 ,w__9519);
  not g__12258(w__9520 ,w__9519);
  not g__12259(w__9519 ,w__9565);
  not g__12260(w__9518 ,w__9516);
  not g__12261(w__9517 ,w__9516);
  not g__12262(w__9516 ,w__9564);
  not g__12263(w__9515 ,w__9513);
  not g__12264(w__9514 ,w__9513);
  not g__12265(w__9513 ,w__9664);
  not g__12266(w__9512 ,w__9510);
  not g__12267(w__9511 ,w__9510);
  not g__12268(w__9510 ,w__9663);
  not g__12269(w__9509 ,w__9507);
  not g__12270(w__9508 ,w__9507);
  not g__12271(w__9507 ,w__9563);
  not g__12272(w__9506 ,w__9504);
  not g__12273(w__9505 ,w__9504);
  not g__12274(w__9504 ,w__9562);
  not g__12275(w__9503 ,w__9501);
  not g__12276(w__9502 ,w__9501);
  not g__12277(w__9501 ,w__9764);
  not g__12278(w__9500 ,w__9498);
  not g__12279(w__9499 ,w__9498);
  not g__12280(w__9498 ,w__9763);
  not g__12281(w__9497 ,w__9495);
  not g__12282(w__9496 ,w__9495);
  not g__12283(w__9495 ,w__9574);
  not g__12284(w__9494 ,w__9492);
  not g__12285(w__9493 ,w__9492);
  not g__12286(w__9492 ,w__9573);
  not g__12287(w__9491 ,w__9489);
  not g__12288(w__9490 ,w__9489);
  not g__12289(w__9489 ,w__9761);
  not g__12290(w__9488 ,w__9486);
  not g__12291(w__9487 ,w__9486);
  not g__12292(w__9486 ,w__9760);
  not g__12293(w__9485 ,w__9483);
  not g__12294(w__9484 ,w__9483);
  not g__12295(w__9483 ,w__9572);
  not g__12296(w__9482 ,w__9480);
  not g__12297(w__9481 ,w__9480);
  not g__12298(w__9480 ,w__9571);
  not g__12299(w__9479 ,w__9477);
  not g__12300(w__9478 ,w__9477);
  not g__12301(w__9477 ,w__9677);
  not g__12302(w__9476 ,w__9474);
  not g__12303(w__9475 ,w__9474);
  not g__12304(w__9474 ,w__9676);
  not g__12305(w__9473 ,w__9471);
  not g__12306(w__9472 ,w__9471);
  not g__12307(w__9471 ,w__9570);
  not g__12308(w__9470 ,w__9468);
  not g__12309(w__9469 ,w__9468);
  not g__12310(w__9468 ,w__9569);
  not g__12311(w__9467 ,w__9557);
  not g__12312(w__9557 ,w__9650);
  not g__12313(w__9466 ,w__9554);
  not g__12314(w__9554 ,w__9630);
  not g__12315(w__9465 ,w__9561);
  not g__12316(w__9561 ,w__9654);
  not g__12317(w__9464 ,w__9558);
  not g__12318(w__9558 ,w__9651);
  not g__12319(w__9463 ,w__9559);
  not g__12320(w__9559 ,w__9652);
  not g__12321(w__9462 ,w__9555);
  not g__12322(w__9555 ,w__9648);
  not g__12323(w__9461 ,w__9553);
  not g__12324(w__9553 ,w__9627);
  not g__12325(w__9460 ,w__9551);
  not g__12326(w__9551 ,w__9623);
  not g__12327(w__9459 ,w__9552);
  not g__12328(w__9552 ,w__9624);
  not g__12329(w__9458 ,w__9550);
  not g__12330(w__9550 ,w__9622);
  not g__12331(w__9457 ,w__9556);
  not g__12332(w__9556 ,w__9649);
  not g__12333(w__9456 ,w__9560);
  not g__12334(w__9560 ,w__9653);
  not g__12335(w__9455 ,w__9454);
  not g__12336(w__9454 ,w__10209);
  not g__12337(w__9453 ,w__9575);
  not g__12338(w__9575 ,w__10212);
  not g__12339(w__9452 ,w__9451);
  not g__12340(w__9451 ,w__9582);
  not g__12341(w__9450 ,w__9449);
  not g__12342(w__9449 ,w__9595);
  not g__12343(w__9448 ,w__9447);
  not g__12344(w__9447 ,w__9594);
  not g__12345(w__9446 ,w__9445);
  not g__12346(w__9445 ,w__9597);
  not g__12347(w__9444 ,w__9443);
  not g__12348(w__9443 ,w__9596);
  not g__12349(w__9442 ,w__9441);
  not g__12350(w__9441 ,w__9593);
  not g__12351(w__9440 ,w__9439);
  not g__12352(w__9439 ,w__9581);
  not g__12353(w__9438 ,w__9437);
  not g__12354(w__9437 ,w__9672);
  buf g__12355(w__13178 ,w__9821);
  buf g__12356(w__13179 ,w__9747);
  not g__12357(w__9436 ,w__9435);
  not g__12358(w__9435 ,w__9620);
  not g__12359(w__9434 ,w__9433);
  not g__12360(w__9433 ,w__10210);
  not g__12361(w__9432 ,w__9577);
  not g__12362(w__9577 ,w__10566);
  not g__12363(w__9431 ,w__9578);
  not g__12364(w__9578 ,w__10582);
  not g__12365(w__9430 ,w__9579);
  not g__12366(w__9579 ,w__10822);
  not g__12367(w__9429 ,w__9576);
  not g__12368(w__9576 ,w__10565);
  not g__12369(w__9428 ,w__9580);
  not g__12370(w__9580 ,w__10823);
  not g__12371(w__9427 ,w__9426);
  not g__12372(w__9426 ,w__9975);
  not g__12373(w__9425 ,w__9424);
  not g__12374(w__9424 ,w__9882);
  not g__12375(w__9423 ,w__9422);
  not g__12376(w__9422 ,w__9881);
  not g__12377(w__9421 ,w__9420);
  not g__12378(w__9420 ,w__9878);
  not g__12379(w__9419 ,w__9418);
  not g__12380(w__9418 ,w__9877);
  not g__12381(w__9417 ,w__9416);
  not g__12382(w__9416 ,w__9880);
  not g__12383(w__9415 ,w__9414);
  not g__12384(w__9414 ,w__9879);
  not g__12385(w__9413 ,w__9412);
  not g__12386(w__9412 ,w__9583);
  not g__12387(w__9411 ,w__9410);
  not g__12388(w__9410 ,w__9976);
  not g__12389(w__9409 ,w__9407);
  not g__12390(w__9408 ,w__9407);
  not g__12391(w__9407 ,w__9584);
  not g__12392(w__9406 ,w__9404);
  not g__12393(w__9405 ,w__9404);
  not g__12394(w__9404 ,w__9673);
  not g__12395(w__9403 ,w__9573);
  not g__12396(w__9573 ,w__9762);
  not g__12397(w__9402 ,w__9565);
  not g__12398(w__9565 ,w__9665);
  not g__12399(w__9401 ,w__9564);
  not g__12400(w__9564 ,w__9665);
  not g__12401(w__9400 ,w__9563);
  not g__12402(w__9563 ,w__9662);
  not g__12403(w__9399 ,w__9571);
  not g__12404(w__9571 ,w__9759);
  not g__12405(w__9398 ,w__9574);
  not g__12406(w__9574 ,w__9762);
  not g__12407(w__9397 ,w__9572);
  not g__12408(w__9572 ,w__9759);
  not g__12409(w__9396 ,w__9570);
  not g__12410(w__9570 ,w__9675);
  not g__12411(w__9395 ,w__9569);
  not g__12412(w__9569 ,w__9675);
  not g__12413(w__9394 ,w__9562);
  not g__12414(w__9562 ,w__9662);
  not g__12415(w__9393 ,w__9566);
  not g__12416(w__9566 ,w__9668);
  not g__12417(w__9392 ,w__9568);
  not g__12418(w__9568 ,w__9673);
  not g__12419(w__9391 ,w__9567);
  not g__12420(w__9567 ,w__9668);
  not g__12421(w__9390 ,w__9389);
  not g__12422(w__9389 ,w__10129);
  not g__12423(w__9388 ,w__9387);
  not g__12424(w__9387 ,w__10206);
  not g__12425(w__9386 ,w__9385);
  not g__12426(w__9385 ,w__10131);
  not g__12427(w__9384 ,w__9383);
  not g__12428(w__9383 ,w__10127);
  not g__12429(w__9234 ,w__9243);
  not g__12430(w__9382 ,w__9243);
  not g__12431(w__9243 ,w__9235);
  not g__12432(w__9381 ,w__9549);
  not g__12433(w__9380 ,w__9378);
  not g__12434(w__9379 ,w__9378);
  not g__12435(w__9378 ,w__9975);
  not g__12436(w__9377 ,w__9375);
  not g__12437(w__9376 ,w__9375);
  not g__12438(w__9375 ,w__9976);
  not g__12439(w__9374 ,w__9372);
  not g__12440(w__9373 ,w__9372);
  not g__12441(w__9372 ,w__9882);
  not g__12442(w__9371 ,w__9369);
  not g__12443(w__9370 ,w__9369);
  not g__12444(w__9369 ,w__9879);
  not g__12445(w__9368 ,w__9366);
  not g__12446(w__9367 ,w__9366);
  not g__12447(w__9366 ,w__9583);
  not g__12448(w__9365 ,w__9363);
  not g__12449(w__9364 ,w__9363);
  not g__12450(w__9363 ,w__9881);
  not g__12451(w__9362 ,w__9360);
  not g__12452(w__9361 ,w__9360);
  not g__12453(w__9360 ,w__9880);
  not g__12454(w__9359 ,w__9357);
  not g__12455(w__9358 ,w__9357);
  not g__12456(w__9357 ,w__9878);
  not g__12457(w__9356 ,w__9354);
  not g__12458(w__9355 ,w__9354);
  not g__12459(w__9354 ,w__9877);
  not g__12460(w__9353 ,w__9351);
  not g__12461(w__9352 ,w__9351);
  not g__12462(w__9351 ,w__9975);
  not g__12463(w__9350 ,w__9348);
  not g__12464(w__9349 ,w__9348);
  not g__12465(w__9348 ,w__9427);
  not g__12466(w__9347 ,w__9345);
  not g__12467(w__9346 ,w__9345);
  not g__12468(w__9345 ,w__9417);
  not g__12469(w__9344 ,w__9342);
  not g__12470(w__9343 ,w__9342);
  not g__12471(w__9342 ,w__9419);
  not g__12472(w__9341 ,w__9339);
  not g__12473(w__9340 ,w__9339);
  not g__12474(w__9339 ,w__9415);
  not g__12475(w__9338 ,w__9336);
  not g__12476(w__9337 ,w__9336);
  not g__12477(w__9336 ,w__9413);
  not g__12478(w__9335 ,w__9333);
  not g__12479(w__9334 ,w__9333);
  not g__12480(w__9333 ,w__9409);
  not g__12481(w__9332 ,w__9330);
  not g__12482(w__9331 ,w__9330);
  not g__12483(w__9330 ,w__9880);
  not g__12484(w__9329 ,w__9327);
  not g__12485(w__9328 ,w__9327);
  not g__12486(w__9327 ,w__9427);
  not g__12487(w__9326 ,w__9324);
  not g__12488(w__9325 ,w__9324);
  not g__12489(w__9324 ,w__9584);
  not g__12490(w__9323 ,w__9321);
  not g__12491(w__9322 ,w__9321);
  not g__12492(w__9321 ,w__9584);
  not g__12493(w__9320 ,w__9318);
  not g__12494(w__9319 ,w__9318);
  not g__12495(w__9318 ,w__9425);
  not g__12496(w__9317 ,w__9315);
  not g__12497(w__9316 ,w__9315);
  not g__12498(w__9315 ,w__9423);
  not g__12499(w__9314 ,w__9312);
  not g__12500(w__9313 ,w__9312);
  not g__12501(w__9312 ,w__9421);
  not g__12502(w__9311 ,w__9309);
  not g__12503(w__9310 ,w__9309);
  not g__12504(w__9309 ,w__9976);
  not g__12505(w__9308 ,w__9306);
  not g__12506(w__9307 ,w__9306);
  not g__12507(w__9306 ,w__9411);
  not g__12508(w__9305 ,w__9303);
  not g__12509(w__9304 ,w__9303);
  not g__12510(w__9303 ,w__9411);
  not g__12511(w__9302 ,w__9300);
  not g__12512(w__9301 ,w__9300);
  not g__12513(w__9300 ,w__9879);
  not g__12514(w__9299 ,w__9297);
  not g__12515(w__9298 ,w__9297);
  not g__12516(w__9297 ,w__9419);
  not g__12517(w__9296 ,w__9294);
  not g__12518(w__9295 ,w__9294);
  not g__12519(w__9294 ,w__9878);
  not g__12520(w__9293 ,w__9291);
  not g__12521(w__9292 ,w__9291);
  not g__12522(w__9291 ,w__9415);
  not g__12523(w__9290 ,w__9288);
  not g__12524(w__9289 ,w__9288);
  not g__12525(w__9288 ,w__9413);
  not g__12526(w__9287 ,w__9285);
  not g__12527(w__9286 ,w__9285);
  not g__12528(w__9285 ,w__9877);
  not g__12529(w__9284 ,w__9282);
  not g__12530(w__9283 ,w__9282);
  not g__12531(w__9282 ,w__9881);
  not g__12532(w__9281 ,w__9279);
  not g__12533(w__9280 ,w__9279);
  not g__12534(w__9279 ,w__9417);
  not g__12535(w__9278 ,w__9276);
  not g__12536(w__9277 ,w__9276);
  not g__12537(w__9276 ,w__9421);
  not g__12538(w__9275 ,w__9273);
  not g__12539(w__9274 ,w__9273);
  not g__12540(w__9273 ,w__9425);
  not g__12541(w__9272 ,w__9270);
  not g__12542(w__9271 ,w__9270);
  not g__12543(w__9270 ,w__9882);
  not g__12544(w__9269 ,w__9267);
  not g__12545(w__9268 ,w__9267);
  not g__12546(w__9267 ,w__9423);
  not g__12547(w__9266 ,w__9264);
  not g__12548(w__9265 ,w__9264);
  not g__12549(w__9264 ,w__9583);
  not g__12550(w__9263 ,w__9262);
  not g__12551(w__9262 ,w__9408);
  not g__12552(w__9261 ,w__9260);
  not g__12553(w__9260 ,w__9379);
  not g__12554(w__9259 ,w__9258);
  not g__12555(w__9258 ,w__9356);
  not g__12556(w__9257 ,w__9256);
  not g__12557(w__9256 ,w__9359);
  not g__12558(w__9255 ,w__9254);
  not g__12559(w__9254 ,w__9362);
  not g__12560(w__9253 ,w__9252);
  not g__12561(w__9252 ,w__9365);
  not g__12562(w__9251 ,w__9250);
  not g__12563(w__9250 ,w__9368);
  not g__12564(w__9249 ,w__9248);
  not g__12565(w__9248 ,w__9371);
  not g__12566(w__9247 ,w__9246);
  not g__12567(w__9246 ,w__9374);
  not g__12568(w__9245 ,w__9244);
  not g__12569(w__9244 ,w__9377);
  xor g__12570(w__9242 ,w__10824 ,w__10919);
  xor g__12571(w__13155 ,w__10800 ,w__10889);
  xor g__12572(w__9241 ,w__10782 ,w__10803);
  xor g__12573(w__9240 ,w__10441 ,w__10519);
  xor g__12574(w__9239 ,w__10435 ,w__9389);
  xor g__12575(w__9238 ,w__10545 ,w__9387);
  xor g__12576(w__9237 ,w__10424 ,w__9385);
  xor g__12577(w__9236 ,w__10532 ,w__9383);
  xnor g__12578(w__13096 ,w__12616 ,w__12651);
  xnor g__12579(w__13097 ,w__12619 ,w__10951);
  xnor g__12580(w__13099 ,w__12629 ,w__12643);
  xnor g__12581(w__13098 ,w__12625 ,w__12642);
  xnor g__12582(w__13095 ,w__12609 ,w__12644);
  or g__12583(w__13044 ,w__12614 ,w__12650);
  or g__12584(w__13043 ,w__12637 ,w__12649);
  or g__12585(w__13040 ,w__12632 ,w__12646);
  or g__12586(w__13039 ,w__12641 ,w__12648);
  or g__12587(w__13041 ,w__12630 ,w__12647);
  or g__12588(w__13042 ,w__12639 ,w__12645);
  xnor g__12589(w__13094 ,w__12595 ,w__12623);
  xnor g__12590(w__13100 ,w__12626 ,w__12622);
  xnor g__12591(w__13093 ,w__12597 ,w__12621);
  xnor g__12592(w__12651 ,w__12511 ,w__12627);
  and g__12593(w__12650 ,w__12603 ,w__12626);
  and g__12594(w__12649 ,w__12636 ,w__12629);
  or g__12595(w__13037 ,w__12611 ,w__12631);
  and g__12596(w__12648 ,w__12609 ,w__12633);
  nor g__12597(w__12647 ,w__12640 ,w__12628);
  or g__12598(w__13045 ,w__12593 ,w__12634);
  or g__12599(w__13038 ,w__12613 ,w__12635);
  and g__12600(w__12646 ,w__12624 ,w__12627);
  xnor g__12601(w__13101 ,w__12608 ,w__12600);
  xnor g__12602(w__13092 ,w__12596 ,w__12599);
  xnor g__12603(w__13102 ,w__12514 ,w__12601);
  nor g__12604(w__12645 ,w__12638 ,w__12625);
  xnor g__12605(w__12644 ,w__12605 ,w__12531);
  xnor g__12606(w__12643 ,w__12618 ,w__12532);
  xnor g__12607(w__12642 ,w__12606 ,w__12620);
  nor g__12608(w__12641 ,w__11139 ,w__12605);
  and g__12609(w__12640 ,w__12533 ,w__12619);
  nor g__12610(w__12639 ,w__12607 ,w__12620);
  and g__12611(w__12638 ,w__12607 ,w__12620);
  nor g__12612(w__12637 ,w__11137 ,w__12618);
  or g__12613(w__12636 ,w__11289 ,w__12617);
  nor g__12614(w__12635 ,w__12595 ,w__12612);
  and g__12615(w__12634 ,w__12592 ,w__12608);
  or g__12616(w__12633 ,w__11288 ,w__12604);
  nor g__12617(w__12632 ,w__12511 ,w__12616);
  nor g__12618(w__12631 ,w__12597 ,w__12610);
  nor g__12619(w__12630 ,w__12533 ,w__12619);
  or g__12620(w__12624 ,w__12510 ,w__12615);
  or g__12621(w__13091 ,w__12586 ,w__12602);
  xnor g__12622(w__13103 ,w__12540 ,w__10950);
  xnor g__12623(w__13105 ,w__12450 ,w__12570);
  xnor g__12624(w__13035 ,w__12518 ,w__12571);
  xnor g__12625(w__12623 ,w__12482 ,w__12577);
  xnor g__12626(w__12622 ,w__12580 ,w__12535);
  xnor g__12627(w__12621 ,w__12472 ,w__12581);
  xnor g__12628(w__12629 ,w__12517 ,w__12573);
  xnor g__12629(w__12628 ,w__12566 ,w__12569);
  xnor g__12630(w__12627 ,w__12543 ,w__12572);
  xnor g__12631(w__12626 ,w__12515 ,w__12567);
  xnor g__12632(w__12625 ,w__12539 ,w__12568);
  not g__12633(w__12617 ,w__12618);
  not g__12634(w__12615 ,w__12616);
  nor g__12635(w__12614 ,w__12535 ,w__12580);
  nor g__12636(w__12613 ,w__12482 ,w__12578);
  and g__12637(w__12612 ,w__12482 ,w__12578);
  or g__12638(w__13046 ,w__12557 ,w__12591);
  nor g__12639(w__12611 ,w__12472 ,w__12582);
  or g__12640(w__13047 ,w__12555 ,w__12590);
  or g__12641(w__13049 ,w__12551 ,w__12589);
  or g__12642(w__13090 ,w__12549 ,w__12587);
  and g__12643(w__12610 ,w__12472 ,w__12582);
  and g__12644(w__12620 ,w__12563 ,w__12583);
  and g__12645(w__12619 ,w__12546 ,w__12584);
  and g__12646(w__12618 ,w__12561 ,w__12594);
  and g__12647(w__12616 ,w__12552 ,w__12588);
  not g__12648(w__12607 ,w__12606);
  not g__12649(w__12604 ,w__12605);
  or g__12650(w__12603 ,w__12534 ,w__12579);
  nor g__12651(w__12602 ,w__12596 ,w__12585);
  or g__12652(w__13089 ,w__12545 ,w__12574);
  xnor g__12653(w__13104 ,w__12542 ,w__12523);
  or g__12654(w__13048 ,w__12503 ,w__12576);
  xnor g__12655(w__12601 ,w__12486 ,w__12538);
  xnor g__12656(w__12600 ,w__12530 ,w__12528);
  xnor g__12657(w__12599 ,w__12467 ,w__12536);
  xnor g__12658(w__12598 ,w__12541 ,w__12426);
  or g__12659(w__12609 ,w__12558 ,w__12575);
  xnor g__12660(w__12608 ,w__12469 ,w__12521);
  xnor g__12661(w__12606 ,w__12349 ,w__12520);
  xnor g__12662(w__12605 ,w__12516 ,w__12522);
  or g__12663(w__12594 ,w__12515 ,w__12559);
  nor g__12664(w__12593 ,w__12528 ,w__12530);
  or g__12665(w__12592 ,w__12527 ,w__12529);
  and g__12666(w__12591 ,w__12556 ,w__12538);
  nor g__12667(w__12590 ,w__12565 ,w__12540);
  and g__12668(w__12589 ,w__12450 ,w__12550);
  or g__12669(w__13050 ,w__12452 ,w__12548);
  or g__12670(w__12588 ,w__12566 ,w__12547);
  nor g__12671(w__12587 ,w__12524 ,w__12541);
  nor g__12672(w__12586 ,w__12467 ,w__12537);
  and g__12673(w__12585 ,w__12467 ,w__12537);
  or g__12674(w__12584 ,w__12539 ,w__12564);
  or g__12675(w__12583 ,w__12517 ,w__12562);
  and g__12676(w__12597 ,w__12444 ,w__12553);
  and g__12677(w__12596 ,w__12379 ,w__12526);
  and g__12678(w__12595 ,w__12507 ,w__12560);
  not g__12679(w__12582 ,w__12581);
  not g__12680(w__12579 ,w__12580);
  not g__12681(w__12578 ,w__12577);
  nor g__12682(w__12576 ,w__12504 ,w__12542);
  nor g__12683(w__12575 ,w__12554 ,w__12543);
  nor g__12684(w__12574 ,w__12518 ,w__12544);
  xnor g__12685(w__13106 ,w__12498 ,w__12478);
  xnor g__12686(w__13034 ,w__12447 ,w__12476);
  xnor g__12687(w__12573 ,w__12352 ,w__12484);
  xnor g__12688(w__12572 ,w__12471 ,w__12495);
  xnor g__12689(w__12571 ,w__12252 ,w__12493);
  xnor g__12690(w__12570 ,w__12490 ,w__12291);
  xnor g__12691(w__12569 ,w__12492 ,w__12466);
  xnor g__12692(w__12568 ,w__12481 ,w__12222);
  xnor g__12693(w__12567 ,w__12421 ,w__12488);
  xnor g__12694(w__12581 ,w__12497 ,w__12436);
  and g__12695(w__12580 ,w__12479 ,w__12525);
  xnor g__12696(w__12577 ,w__12519 ,w__12477);
  and g__12697(w__12565 ,w__12491 ,w__12512);
  and g__12698(w__12564 ,w__12222 ,w__12481);
  or g__12699(w__12563 ,w__12351 ,w__12484);
  nor g__12700(w__12562 ,w__12352 ,w__12483);
  or g__12701(w__12561 ,w__12421 ,w__12487);
  or g__12702(w__12560 ,w__12505 ,w__12516);
  nor g__12703(w__12559 ,w__12420 ,w__12488);
  nor g__12704(w__12558 ,w__12471 ,w__12496);
  nor g__12705(w__12557 ,w__12514 ,w__12486);
  or g__12706(w__12556 ,w__12513 ,w__12485);
  nor g__12707(w__12555 ,w__12491 ,w__12512);
  and g__12708(w__12554 ,w__12471 ,w__12496);
  or g__12709(w__12553 ,w__12454 ,w__12519);
  or g__12710(w__12552 ,w__12466 ,w__12492);
  nor g__12711(w__12551 ,w__11140 ,w__12490);
  or g__12712(w__12550 ,w__11287 ,w__12489);
  nor g__12713(w__12549 ,w__12426 ,w__12509);
  and g__12714(w__12548 ,w__12453 ,w__12498);
  and g__12715(w__12547 ,w__12466 ,w__12492);
  or g__12716(w__13087 ,w__12458 ,w__12500);
  or g__12717(w__13088 ,w__12461 ,w__12499);
  or g__12718(w__12546 ,w__12222 ,w__12481);
  nor g__12719(w__12545 ,w__12252 ,w__12494);
  and g__12720(w__12544 ,w__12252 ,w__12494);
  and g__12721(w__12566 ,w__12369 ,w__12508);
  not g__12722(w__12537 ,w__12536);
  not g__12723(w__12535 ,w__12534);
  not g__12724(w__12529 ,w__12530);
  not g__12725(w__12527 ,w__12528);
  xnor g__12726(w__13032 ,w__12220 ,w__12442);
  xnor g__12727(w__13107 ,w__12448 ,w__12435);
  or g__12728(w__12526 ,w__12413 ,w__12497);
  or g__12729(w__12525 ,w__12449 ,w__12480);
  and g__12730(w__12524 ,w__12426 ,w__12509);
  or g__12731(w__13051 ,w__12372 ,w__12506);
  xnor g__12732(w__13108 ,w__12344 ,w__12433);
  xnor g__12733(w__13033 ,w__12425 ,w__12439);
  xnor g__12734(w__12523 ,w__12383 ,w__12473);
  xnor g__12735(w__12522 ,w__12470 ,w__12382);
  xnor g__12736(w__12521 ,w__12257 ,w__12449);
  xnor g__12737(w__12520 ,w__12475 ,w__12285);
  xnor g__12738(w__12543 ,w__12250 ,w__12431);
  xnor g__12739(w__12542 ,w__12354 ,w__12432);
  xnor g__12740(w__12541 ,w__10948 ,w__12434);
  xnor g__12741(w__12540 ,w__12387 ,w__12441);
  and g__12742(w__12539 ,w__12378 ,w__12501);
  xnor g__12743(w__12538 ,w__12474 ,w__12440);
  xnor g__12744(w__12536 ,w__12388 ,w__12438);
  xnor g__12745(w__12534 ,w__12288 ,w__12437);
  xnor g__12746(w__12533 ,w__12214 ,w__12430);
  xnor g__12747(w__12532 ,w__12446 ,w__12427);
  xnor g__12748(w__12531 ,w__12289 ,w__12428);
  xnor g__12749(w__12530 ,w__12283 ,w__12429);
  and g__12750(w__12528 ,w__12407 ,w__12502);
  not g__12751(w__12513 ,w__12514);
  not g__12752(w__12510 ,w__12511);
  or g__12753(w__12508 ,w__12368 ,w__12475);
  or g__12754(w__12507 ,w__12382 ,w__12470);
  nor g__12755(w__12506 ,w__12371 ,w__12448);
  and g__12756(w__12505 ,w__12382 ,w__12470);
  and g__12757(w__12504 ,w__12384 ,w__12473);
  nor g__12758(w__12503 ,w__12384 ,w__12473);
  or g__12759(w__12502 ,w__12474 ,w__12404);
  or g__12760(w__12501 ,w__12376 ,w__12446);
  and g__12761(w__12500 ,w__12353 ,w__12460);
  and g__12762(w__12499 ,w__12447 ,w__12456);
  and g__12763(w__12519 ,w__12419 ,w__12463);
  and g__12764(w__12518 ,w__12392 ,w__12443);
  and g__12765(w__12517 ,w__12418 ,w__12464);
  and g__12766(w__12516 ,w__12374 ,w__12457);
  and g__12767(w__12515 ,w__12412 ,w__12462);
  and g__12768(w__12514 ,w__12403 ,w__12455);
  and g__12769(w__12512 ,w__12399 ,w__12465);
  and g__12770(w__12511 ,w__12397 ,w__12451);
  and g__12771(w__12509 ,w__12417 ,w__12459);
  not g__12772(w__12496 ,w__12495);
  not g__12773(w__12494 ,w__12493);
  not g__12774(w__12489 ,w__12490);
  not g__12775(w__12487 ,w__12488);
  not g__12776(w__12485 ,w__12486);
  not g__12777(w__12483 ,w__12484);
  xnor g__12778(w__13109 ,w__12300 ,w__10949);
  or g__12779(w__13052 ,w__12390 ,w__12445);
  nor g__12780(w__12480 ,w__12257 ,w__12468);
  or g__12781(w__12479 ,w__12256 ,w__12469);
  xnor g__12782(w__12478 ,w__12423 ,w__12274);
  xnor g__12783(w__12477 ,w__10946 ,w__12381);
  xnor g__12784(w__12476 ,w__12386 ,w__12275);
  xnor g__12785(w__12498 ,w__12307 ,w__12361);
  xnor g__12786(w__12497 ,w__12302 ,w__12358);
  xnor g__12787(w__12495 ,w__12259 ,w__10945);
  xnor g__12788(w__12493 ,w__12303 ,w__10947);
  xnor g__12789(w__12492 ,w__12296 ,w__12357);
  xnor g__12790(w__12491 ,w__12261 ,w__12355);
  xnor g__12791(w__12490 ,w__12301 ,w__12356);
  xnor g__12792(w__12488 ,w__12235 ,w__12363);
  xnor g__12793(w__12486 ,w__12308 ,w__12364);
  xnor g__12794(w__12484 ,w__12212 ,w__12360);
  xnor g__12795(w__12482 ,w__12293 ,w__12362);
  xnor g__12796(w__12481 ,w__12294 ,w__12359);
  not g__12797(w__12468 ,w__12469);
  or g__12798(w__12465 ,w__12354 ,w__12398);
  or g__12799(w__12464 ,w__12299 ,w__12416);
  or g__12800(w__12463 ,w__12298 ,w__12415);
  or g__12801(w__12462 ,w__12297 ,w__12410);
  nor g__12802(w__12461 ,w__11141 ,w__12386);
  or g__12803(w__12460 ,w__12246 ,w__12424);
  or g__12804(w__12459 ,w__12409 ,w__12389);
  nor g__12805(w__12458 ,w__12247 ,w__12425);
  or g__12806(w__13086 ,w__12309 ,w__12377);
  or g__12807(w__12457 ,w__12304 ,w__12373);
  or g__12808(w__12456 ,w__11286 ,w__12385);
  or g__12809(w__12455 ,w__12387 ,w__12401);
  or g__12810(w__13053 ,w__12317 ,w__12402);
  nor g__12811(w__12454 ,w__10946 ,w__12380);
  or g__12812(w__12453 ,w__11285 ,w__12422);
  nor g__12813(w__12452 ,w__11138 ,w__12423);
  or g__12814(w__12451 ,w__12295 ,w__12395);
  and g__12815(w__12475 ,w__12318 ,w__12405);
  and g__12816(w__12474 ,w__12336 ,w__12406);
  and g__12817(w__12473 ,w__12328 ,w__12396);
  and g__12818(w__12472 ,w__12332 ,w__12391);
  and g__12819(w__12471 ,w__12333 ,w__12400);
  and g__12820(w__12470 ,w__12341 ,w__12411);
  and g__12821(w__12469 ,w__12340 ,w__12408);
  and g__12822(w__12467 ,w__12325 ,w__12365);
  and g__12823(w__12466 ,w__12324 ,w__12393);
  or g__12824(w__13054 ,w__12165 ,w__12366);
  nor g__12825(w__12445 ,w__12306 ,w__12394);
  or g__12826(w__12444 ,w__12350 ,w__12381);
  xnor g__12827(w__13110 ,w__12305 ,w__12208);
  or g__12828(w__12443 ,w__10948 ,w__12414);
  xnor g__12829(w__12442 ,w__12292 ,w__11920);
  xnor g__12830(w__12441 ,w__12277 ,w__12278);
  xnor g__12831(w__12440 ,w__12280 ,w__12347);
  xnor g__12832(w__12439 ,w__12247 ,w__12353);
  xnor g__12833(w__12438 ,w__12281 ,w__12255);
  xnor g__12834(w__12437 ,w__12267 ,w__12299);
  xnor g__12835(w__12436 ,w__12227 ,w__12271);
  xnor g__12836(w__12435 ,w__12218 ,w__12273);
  xnor g__12837(w__12434 ,w__12269 ,w__12213);
  xnor g__12838(w__12433 ,w__12306 ,w__12230);
  xnor g__12839(w__12432 ,w__12276 ,w__12272);
  xnor g__12840(w__12431 ,w__12290 ,w__12304);
  xnor g__12841(w__12430 ,w__12286 ,w__12295);
  xnor g__12842(w__12429 ,w__12297 ,w__12243);
  xnor g__12843(w__12428 ,w__12298 ,w__12249);
  xnor g__12844(w__12427 ,w__12282 ,w__12268);
  or g__12845(w__12450 ,w__12323 ,w__12367);
  xnor g__12846(w__12449 ,w__12258 ,w__12265);
  xnor g__12847(w__12448 ,w__12233 ,w__12264);
  or g__12848(w__12447 ,w__12339 ,w__12370);
  and g__12849(w__12446 ,w__12311 ,w__12375);
  not g__12850(w__12424 ,w__12425);
  not g__12851(w__12422 ,w__12423);
  not g__12852(w__12420 ,w__12421);
  or g__12853(w__13085 ,w__12036 ,w__12314);
  or g__12854(w__12419 ,w__12249 ,w__12289);
  or g__12855(w__12418 ,w__12266 ,w__12288);
  or g__12856(w__12417 ,w__12255 ,w__12281);
  nor g__12857(w__12416 ,w__12267 ,w__12287);
  and g__12858(w__12415 ,w__12249 ,w__12289);
  and g__12859(w__12414 ,w__12213 ,w__12269);
  nor g__12860(w__12413 ,w__12227 ,w__12270);
  or g__12861(w__12412 ,w__12243 ,w__12283);
  or g__12862(w__12411 ,w__12259 ,w__12338);
  and g__12863(w__12410 ,w__12243 ,w__12283);
  and g__12864(w__12409 ,w__12255 ,w__12281);
  or g__12865(w__12408 ,w__12308 ,w__12337);
  or g__12866(w__12407 ,w__12280 ,w__12346);
  or g__12867(w__12406 ,w__12261 ,w__12335);
  or g__12868(w__12405 ,w__12231 ,w__12315);
  nor g__12869(w__12404 ,w__12279 ,w__12347);
  or g__12870(w__12403 ,w__12278 ,w__12277);
  nor g__12871(w__12402 ,w__12316 ,w__12300);
  and g__12872(w__12401 ,w__12278 ,w__12277);
  or g__12873(w__12400 ,w__12331 ,w__12296);
  or g__12874(w__12399 ,w__12272 ,w__12276);
  and g__12875(w__12398 ,w__12272 ,w__12276);
  or g__12876(w__12397 ,w__12214 ,w__12286);
  or g__12877(w__12396 ,w__12327 ,w__12301);
  and g__12878(w__12395 ,w__12214 ,w__12286);
  and g__12879(w__12394 ,w__12230 ,w__12345);
  or g__12880(w__12393 ,w__12320 ,w__12294);
  or g__12881(w__12392 ,w__12213 ,w__12269);
  or g__12882(w__12391 ,w__12319 ,w__12293);
  nor g__12883(w__12390 ,w__12230 ,w__12345);
  and g__12884(w__12426 ,w__12011 ,w__12334);
  and g__12885(w__12425 ,w__12052 ,w__12326);
  and g__12886(w__12423 ,w__12209 ,w__12321);
  and g__12887(w__12421 ,w__12236 ,w__12342);
  not g__12888(w__12389 ,w__12388);
  not g__12889(w__12385 ,w__12386);
  not g__12890(w__12384 ,w__12383);
  not g__12891(w__12380 ,w__12381);
  xnor g__12892(w__13031 ,w__12263 ,w__12157);
  or g__12893(w__12379 ,w__12226 ,w__12271);
  or g__12894(w__12378 ,w__12268 ,w__12282);
  nor g__12895(w__12377 ,w__12329 ,w__12292);
  and g__12896(w__12376 ,w__12268 ,w__12282);
  or g__12897(w__12375 ,w__12235 ,w__12322);
  or g__12898(w__12374 ,w__12250 ,w__12290);
  and g__12899(w__12373 ,w__12250 ,w__12290);
  nor g__12900(w__12372 ,w__12219 ,w__12273);
  and g__12901(w__12371 ,w__12219 ,w__12273);
  nor g__12902(w__12370 ,w__12330 ,w__12303);
  or g__12903(w__12369 ,w__12285 ,w__12348);
  nor g__12904(w__12368 ,w__12284 ,w__12349);
  nor g__12905(w__12367 ,w__12343 ,w__12307);
  nor g__12906(w__12366 ,w__12163 ,w__12305);
  or g__12907(w__12365 ,w__12313 ,w__12302);
  xnor g__12908(w__12364 ,w__12251 ,w__12253);
  xnor g__12909(w__12363 ,w__12043 ,w__12217);
  xnor g__12910(w__12362 ,w__12225 ,w__12242);
  xnor g__12911(w__12361 ,w__12040 ,w__12215);
  xnor g__12912(w__12360 ,w__12231 ,w__12229);
  xnor g__12913(w__12359 ,w__12223 ,w__12224);
  xnor g__12914(w__12358 ,w__12221 ,w__11840);
  xnor g__12915(w__12357 ,w__12244 ,w__12245);
  xnor g__12916(w__12356 ,w__12239 ,w__12240);
  xnor g__12917(w__12355 ,w__12248 ,w__12149);
  xnor g__12918(w__12388 ,w__12262 ,w__12155);
  and g__12919(w__12387 ,w__12185 ,w__12310);
  xnor g__12920(w__12386 ,w__12232 ,w__12142);
  xnor g__12921(w__12383 ,w__12260 ,w__12207);
  xnor g__12922(w__12382 ,w__12234 ,w__12143);
  and g__12923(w__12381 ,w__11990 ,w__12312);
  not g__12924(w__12351 ,w__12352);
  not g__12925(w__12350 ,w__10946);
  not g__12926(w__12348 ,w__12349);
  not g__12927(w__12346 ,w__12347);
  not g__12928(w__12345 ,w__12344);
  and g__12929(w__12343 ,w__12041 ,w__12215);
  or g__12930(w__12342 ,w__12237 ,w__12258);
  or g__12931(w__12341 ,w__11837 ,w__12241);
  or g__12932(w__12340 ,w__12253 ,w__12251);
  nor g__12933(w__12339 ,w__11916 ,w__12254);
  and g__12934(w__12338 ,w__11837 ,w__12241);
  and g__12935(w__12337 ,w__12253 ,w__12251);
  or g__12936(w__12336 ,w__12149 ,w__12248);
  and g__12937(w__12335 ,w__12149 ,w__12248);
  or g__12938(w__12334 ,w__12015 ,w__12262);
  or g__12939(w__12333 ,w__12245 ,w__12244);
  or g__12940(w__12332 ,w__12242 ,w__12225);
  and g__12941(w__12331 ,w__12245 ,w__12244);
  and g__12942(w__12330 ,w__11916 ,w__12254);
  nor g__12943(w__12329 ,w__11919 ,w__12220);
  or g__12944(w__12328 ,w__12240 ,w__12239);
  and g__12945(w__12327 ,w__12240 ,w__12239);
  or g__12946(w__12326 ,w__12007 ,w__12232);
  or g__12947(w__12325 ,w__11840 ,w__12221);
  or g__12948(w__12324 ,w__12224 ,w__12223);
  nor g__12949(w__12323 ,w__12041 ,w__12215);
  nor g__12950(w__12322 ,w__12043 ,w__12216);
  or g__12951(w__12321 ,w__12233 ,w__12210);
  and g__12952(w__12320 ,w__12224 ,w__12223);
  and g__12953(w__12319 ,w__12242 ,w__12225);
  or g__12954(w__12318 ,w__12212 ,w__12229);
  nor g__12955(w__12317 ,w__12150 ,w__12228);
  and g__12956(w__12316 ,w__12150 ,w__12228);
  or g__12957(w__13055 ,w__12003 ,w__12211);
  and g__12958(w__12315 ,w__12212 ,w__12229);
  nor g__12959(w__12314 ,w__12029 ,w__12263);
  and g__12960(w__12313 ,w__11095 ,w__12221);
  or g__12961(w__12312 ,w__11989 ,w__12234);
  or g__12962(w__12311 ,w__12042 ,w__12217);
  or g__12963(w__12310 ,w__12184 ,w__12260);
  and g__12964(w__12309 ,w__11143 ,w__12220);
  and g__12965(w__12354 ,w__12045 ,w__12238);
  xnor g__12966(w__12353 ,w__12135 ,w__11920);
  xnor g__12967(w__12352 ,w__12121 ,w__11162);
  xnor g__12968(w__12349 ,w__12154 ,w__11921);
  xnor g__12969(w__12347 ,w__12099 ,w__12113);
  xnor g__12970(w__12344 ,w__12044 ,w__12100);
  not g__12971(w__12287 ,w__12288);
  not g__12972(w__12284 ,w__12285);
  not g__12973(w__12279 ,w__12280);
  not g__12974(w__12270 ,w__12271);
  not g__12975(w__12266 ,w__12267);
  xnor g__12976(w__13112 ,w__11887 ,w__12140);
  xnor g__12977(w__13030 ,w__12110 ,w__11329);
  xnor g__12978(w__13111 ,w__12152 ,w__12130);
  xnor g__12979(w__12265 ,w__12148 ,w__11955);
  xnor g__12980(w__12264 ,w__12151 ,w__11872);
  xnor g__12981(w__12308 ,w__11953 ,w__12139);
  xnor g__12982(w__12307 ,w__11922 ,w__12141);
  xnor g__12983(w__12306 ,w__11966 ,w__12136);
  xnor g__12984(w__12305 ,w__11848 ,w__12137);
  xnor g__12985(w__12304 ,w__12112 ,w__11358);
  xnor g__12986(w__12303 ,w__11902 ,w__12132);
  xnor g__12987(w__12302 ,w__12125 ,w__11362);
  xnor g__12988(w__12301 ,w__11893 ,w__12105);
  xnor g__12989(w__12300 ,w__11969 ,w__12123);
  xnor g__12990(w__12299 ,w__11977 ,w__12118);
  xnor g__12991(w__12298 ,w__11900 ,w__12117);
  xnor g__12992(w__12297 ,w__11968 ,w__12115);
  xnor g__12993(w__12296 ,w__11967 ,w__12107);
  xnor g__12994(w__12295 ,w__11976 ,w__12146);
  xnor g__12995(w__12294 ,w__11970 ,w__12102);
  xnor g__12996(w__12293 ,w__11862 ,w__12101);
  xnor g__12997(w__12292 ,w__12111 ,w__11339);
  xnor g__12998(w__12291 ,w__12153 ,w__12104);
  xnor g__12999(w__12290 ,w__11899 ,w__12134);
  xnor g__13000(w__12289 ,w__11972 ,w__12119);
  xnor g__13001(w__12288 ,w__11874 ,w__12147);
  xnor g__13002(w__12286 ,w__12106 ,w__11918);
  xnor g__13003(w__12285 ,w__11940 ,w__12131);
  xnor g__13004(w__12283 ,w__11868 ,w__12116);
  xnor g__13005(w__12282 ,w__11987 ,w__12129);
  xnor g__13006(w__12281 ,w__11865 ,w__12120);
  xnor g__13007(w__12280 ,w__11935 ,w__12114);
  xnor g__13008(w__12278 ,w__11956 ,w__12109);
  xnor g__13009(w__12277 ,w__11974 ,w__12108);
  xnor g__13010(w__12276 ,w__11944 ,w__12128);
  xnor g__13011(w__12275 ,w__12103 ,w__11360);
  xnor g__13012(w__12274 ,w__11952 ,w__12127);
  xnor g__13013(w__12273 ,w__11890 ,w__12122);
  xnor g__13014(w__12272 ,w__11875 ,w__12138);
  xnor g__13015(w__12271 ,w__11936 ,w__12124);
  xnor g__13016(w__12269 ,w__11942 ,w__12126);
  xnor g__13017(w__12268 ,w__11855 ,w__12145);
  xnor g__13018(w__12267 ,w__11911 ,w__12156);
  not g__13019(w__12256 ,w__12257);
  not g__13020(w__12246 ,w__12247);
  or g__13021(w__12238 ,w__12053 ,w__12153);
  and g__13022(w__12237 ,w__11955 ,w__12148);
  or g__13023(w__12236 ,w__11955 ,w__12148);
  and g__13024(w__12263 ,w__12091 ,w__12175);
  and g__13025(w__12262 ,w__12096 ,w__12190);
  and g__13026(w__12261 ,w__12059 ,w__12187);
  and g__13027(w__12260 ,w__12050 ,w__12181);
  and g__13028(w__12259 ,w__12079 ,w__12194);
  and g__13029(w__12258 ,w__12087 ,w__12200);
  or g__13030(w__12257 ,w__12082 ,w__12195);
  and g__13031(w__12255 ,w__12089 ,w__12198);
  and g__13032(w__12254 ,w__12071 ,w__12183);
  and g__13033(w__12253 ,w__12076 ,w__12193);
  and g__13034(w__12252 ,w__11992 ,w__12205);
  and g__13035(w__12251 ,w__12072 ,w__12191);
  and g__13036(w__12250 ,w__12070 ,w__12189);
  and g__13037(w__12249 ,w__12094 ,w__12204);
  and g__13038(w__12248 ,w__12062 ,w__12188);
  and g__13039(w__12247 ,w__12090 ,w__12201);
  and g__13040(w__12245 ,w__12056 ,w__12186);
  and g__13041(w__12244 ,w__12051 ,w__12182);
  and g__13042(w__12243 ,w__12085 ,w__12199);
  and g__13043(w__12242 ,w__12049 ,w__12178);
  and g__13044(w__12241 ,w__12084 ,w__12197);
  and g__13045(w__12240 ,w__12035 ,w__12206);
  and g__13046(w__12239 ,w__12093 ,w__12177);
  not g__13047(w__12226 ,w__12227);
  not g__13048(w__12219 ,w__12218);
  not g__13049(w__12216 ,w__12217);
  and g__13050(w__12211 ,w__12010 ,w__12152);
  or g__13051(w__13056 ,w__12013 ,w__12161);
  and g__13052(w__12210 ,w__11872 ,w__12151);
  or g__13053(w__12209 ,w__11872 ,w__12151);
  xnor g__13054(w__12208 ,w__11846 ,w__12038);
  xnor g__13055(w__12207 ,w__11939 ,w__12098);
  and g__13056(w__12235 ,w__12066 ,w__12179);
  and g__13057(w__12234 ,w__12002 ,w__12159);
  and g__13058(w__12233 ,w__12031 ,w__12171);
  and g__13059(w__12232 ,w__11996 ,w__12160);
  and g__13060(w__12231 ,w__12009 ,w__12162);
  and g__13061(w__12230 ,w__12018 ,w__12169);
  and g__13062(w__12229 ,w__12058 ,w__12166);
  and g__13063(w__12228 ,w__12017 ,w__12168);
  or g__13064(w__12227 ,w__11995 ,w__12167);
  and g__13065(w__12225 ,w__11999 ,w__12172);
  and g__13066(w__12224 ,w__12030 ,w__12176);
  and g__13067(w__12223 ,w__12026 ,w__12173);
  and g__13068(w__12222 ,w__12008 ,w__12196);
  and g__13069(w__12221 ,w__12000 ,w__12202);
  or g__13070(w__12220 ,w__11994 ,w__12192);
  or g__13071(w__12218 ,w__12021 ,w__12180);
  and g__13072(w__12217 ,w__12005 ,w__12203);
  and g__13073(w__12215 ,w__12028 ,w__12174);
  and g__13074(w__12214 ,w__12037 ,w__12158);
  and g__13075(w__12213 ,w__12019 ,w__12164);
  and g__13076(w__12212 ,w__11988 ,w__12170);
  or g__13077(w__12206 ,w__11985 ,w__12034);
  or g__13078(w__12205 ,w__11986 ,w__11991);
  or g__13079(w__12204 ,w__11984 ,w__12092);
  or g__13080(w__12203 ,w__11983 ,w__12067);
  or g__13081(w__12202 ,w__11910 ,w__12001);
  or g__13082(w__12201 ,w__12088 ,w__11982);
  or g__13083(w__12200 ,w__11898 ,w__12086);
  or g__13084(w__12199 ,w__11981 ,w__12083);
  or g__13085(w__12198 ,w__11980 ,w__12080);
  or g__13086(w__12197 ,w__11978 ,w__12081);
  or g__13087(w__12196 ,w__11284 ,w__12078);
  and g__13088(w__12195 ,w__12099 ,w__12077);
  or g__13089(w__12194 ,w__11976 ,w__12074);
  or g__13090(w__12193 ,w__11975 ,w__12073);
  nor g__13091(w__12192 ,w__11997 ,w__11143);
  or g__13092(w__12191 ,w__11974 ,w__12068);
  or g__13093(w__12190 ,w__11912 ,w__12061);
  or g__13094(w__12189 ,w__11164 ,w__12065);
  or g__13095(w__12188 ,w__11973 ,w__12060);
  or g__13096(w__12187 ,w__11896 ,w__12057);
  or g__13097(w__12186 ,w__11901 ,w__12054);
  or g__13098(w__12185 ,w__11939 ,w__12097);
  nor g__13099(w__12184 ,w__11938 ,w__12098);
  or g__13100(w__12183 ,w__11971 ,w__12047);
  or g__13101(w__12182 ,w__11970 ,w__12046);
  or g__13102(w__12181 ,w__11893 ,w__12048);
  and g__13103(w__12180 ,w__12044 ,w__12075);
  or g__13104(w__12179 ,w__11968 ,w__12095);
  or g__13105(w__12178 ,w__11972 ,w__12063);
  or g__13106(w__12177 ,w__11889 ,w__12032);
  or g__13107(w__12176 ,w__11886 ,w__12027);
  or g__13108(w__12175 ,w__12024 ,w__11909);
  or g__13109(w__12174 ,w__11890 ,w__12025);
  or g__13110(w__12173 ,w__11987 ,w__12023);
  or g__13111(w__12172 ,w__11900 ,w__12020);
  or g__13112(w__12171 ,w__11905 ,w__12022);
  or g__13113(w__12170 ,w__12004 ,w__11911);
  or g__13114(w__12169 ,w__11969 ,w__12006);
  or g__13115(w__12168 ,w__11897 ,w__12016);
  and g__13116(w__12167 ,w__11998 ,w__11095);
  or g__13117(w__12166 ,w__11977 ,w__12014);
  nor g__13118(w__12165 ,w__11846 ,w__12039);
  or g__13119(w__12164 ,w__11979 ,w__12064);
  and g__13120(w__12163 ,w__11846 ,w__12039);
  or g__13121(w__12162 ,w__11908 ,w__12012);
  nor g__13122(w__12161 ,w__11887 ,w__12055);
  or g__13123(w__12160 ,w__11993 ,w__11902);
  or g__13124(w__12159 ,w__11899 ,w__12069);
  or g__13125(w__12158 ,w__11162 ,w__12033);
  xnor g__13126(w__13113 ,w__11913 ,w__11834);
  xnor g__13127(w__12157 ,w__11845 ,w__11145);
  xnor g__13128(w__12156 ,w__11879 ,w__11337);
  xnor g__13129(w__12155 ,w__11859 ,w__11838);
  xnor g__13130(w__12154 ,w__11924 ,w__11164);
  xnor g__13131(w__12147 ,w__11841 ,w__11908);
  xnor g__13132(w__12146 ,w__11958 ,w__11357);
  xnor g__13133(w__12145 ,w__11886 ,w__11331);
  xnor g__13134(w__12144 ,w__11986 ,w__11363);
  xnor g__13135(w__12143 ,w__11093 ,w__11333);
  xnor g__13136(w__12142 ,w__11928 ,w__11915);
  xnor g__13137(w__12141 ,w__11985 ,w__11592);
  xnor g__13138(w__12140 ,w__11597 ,w__11881);
  xnor g__13139(w__12139 ,w__11898 ,w__11595);
  xnor g__13140(w__12138 ,w__11973 ,w__11593);
  xnor g__13141(w__12137 ,w__11897 ,w__11596);
  xnor g__13142(w__12136 ,w__11905 ,w__11594);
  xnor g__13143(w__12135 ,w__11861 ,w__11359);
  xnor g__13144(w__12134 ,w__11923 ,w__11860);
  xnor g__13145(w__12133 ,w__11858 ,w__11335);
  xnor g__13146(w__12132 ,w__11856 ,w__11361);
  xnor g__13147(w__12131 ,w__11901 ,w__11332);
  xnor g__13148(w__12130 ,w__11883 ,w__11843);
  xnor g__13149(w__12129 ,w__11876 ,w__11851);
  xnor g__13150(w__12128 ,w__11943 ,w__11896);
  xnor g__13151(w__12127 ,w__11947 ,w__11889);
  xnor g__13152(w__12126 ,w__11971 ,w__11948);
  xnor g__13153(w__12125 ,w__11946 ,w__11912);
  xnor g__13154(w__12124 ,w__11980 ,w__11957);
  xnor g__13155(w__12123 ,w__11852 ,w__11854);
  xnor g__13156(w__12122 ,w__11844 ,w__11877);
  xnor g__13157(w__12121 ,w__11867 ,w__11863);
  xnor g__13158(w__12120 ,w__11979 ,w__11336);
  xnor g__13159(w__12119 ,w__11927 ,w__11931);
  xnor g__13160(w__12118 ,w__11847 ,w__11929);
  xnor g__13161(w__12117 ,w__11880 ,w__11864);
  xnor g__13162(w__12116 ,w__11866 ,w__11983);
  xnor g__13163(w__12115 ,w__11871 ,w__11941);
  xnor g__13164(w__12114 ,w__11950 ,w__11981);
  xnor g__13165(w__12113 ,w__11961 ,w__11963);
  xnor g__13166(w__12112 ,w__11984 ,w__11965);
  xnor g__13167(w__12111 ,w__11909 ,w__11959);
  xnor g__13168(w__12110 ,w__11341 ,w__11914);
  xnor g__13169(w__12109 ,w__11975 ,w__11954);
  xnor g__13170(w__12108 ,w__11873 ,w__11945);
  xnor g__13171(w__12107 ,w__11978 ,w__11930);
  xnor g__13172(w__12106 ,w__11949 ,w__11951);
  xnor g__13173(w__12105 ,w__11932 ,w__11934);
  xnor g__13174(w__12104 ,w__11925 ,w__11926);
  xnor g__13175(w__12103 ,w__11982 ,w__11964);
  xnor g__13176(w__12102 ,w__11933 ,w__11937);
  xnor g__13177(w__12101 ,w__11853 ,w__11910);
  xnor g__13178(w__12100 ,w__11870 ,w__11850);
  xnor g__13179(w__12153 ,w__11906 ,w__11828);
  xnor g__13180(w__12152 ,w__11822 ,w__11888);
  xnor g__13181(w__12151 ,w__11830 ,w__11884);
  xnor g__13182(w__12150 ,w__11832 ,w__11894);
  xnor g__13183(w__12149 ,w__11826 ,w__11891);
  xnor g__13184(w__12148 ,w__11824 ,w__11903);
  not g__13185(w__12097 ,w__12098);
  or g__13186(w__12096 ,w__11165 ,w__11946);
  and g__13187(w__12095 ,w__11941 ,w__11871);
  or g__13188(w__12094 ,w__11166 ,w__11965);
  or g__13189(w__12093 ,w__11947 ,w__11952);
  and g__13190(w__12092 ,w__11358 ,w__11965);
  or g__13191(w__12091 ,w__11175 ,w__11959);
  or g__13192(w__12090 ,w__11173 ,w__11964);
  or g__13193(w__12089 ,w__11957 ,w__11936);
  and g__13194(w__12088 ,w__11360 ,w__11964);
  or g__13195(w__12087 ,w__11595 ,w__11953);
  and g__13196(w__12086 ,w__11595 ,w__11953);
  or g__13197(w__12085 ,w__11950 ,w__11935);
  or g__13198(w__12084 ,w__11930 ,w__11967);
  and g__13199(w__12083 ,w__11950 ,w__11935);
  nor g__13200(w__12082 ,w__11963 ,w__11961);
  and g__13201(w__12081 ,w__11930 ,w__11967);
  and g__13202(w__12080 ,w__11957 ,w__11936);
  or g__13203(w__12079 ,w__11171 ,w__11958);
  and g__13204(w__12078 ,w__11863 ,w__11867);
  or g__13205(w__12077 ,w__11962 ,w__11960);
  or g__13206(w__12076 ,w__11956 ,w__11954);
  or g__13207(w__12075 ,w__11849 ,w__11869);
  and g__13208(w__12074 ,w__11357 ,w__11958);
  and g__13209(w__12073 ,w__11956 ,w__11954);
  or g__13210(w__12072 ,w__11945 ,w__11873);
  or g__13211(w__12071 ,w__11948 ,w__11942);
  or g__13212(w__12070 ,w__11951 ,w__11949);
  and g__13213(w__12069 ,w__11860 ,w__11923);
  and g__13214(w__12068 ,w__11945 ,w__11873);
  and g__13215(w__12067 ,w__11868 ,w__11866);
  or g__13216(w__12066 ,w__11941 ,w__11871);
  and g__13217(w__12065 ,w__11951 ,w__11949);
  and g__13218(w__12064 ,w__11170 ,w__11865);
  and g__13219(w__12063 ,w__11931 ,w__11927);
  or g__13220(w__12062 ,w__11593 ,w__11875);
  and g__13221(w__12061 ,w__11362 ,w__11946);
  and g__13222(w__12060 ,w__11593 ,w__11875);
  or g__13223(w__12059 ,w__11944 ,w__11943);
  or g__13224(w__12058 ,w__11929 ,w__11847);
  and g__13225(w__12057 ,w__11944 ,w__11943);
  or g__13226(w__12056 ,w__11169 ,w__11940);
  and g__13227(w__12055 ,w__11598 ,w__11881);
  and g__13228(w__12054 ,w__11332 ,w__11940);
  and g__13229(w__12053 ,w__11926 ,w__11925);
  or g__13230(w__12052 ,w__11097 ,w__11928);
  or g__13231(w__12051 ,w__11937 ,w__11933);
  or g__13232(w__12050 ,w__11934 ,w__11932);
  or g__13233(w__12049 ,w__11931 ,w__11927);
  and g__13234(w__12048 ,w__11934 ,w__11932);
  and g__13235(w__12047 ,w__11948 ,w__11942);
  and g__13236(w__12046 ,w__11937 ,w__11933);
  or g__13237(w__12045 ,w__11926 ,w__11925);
  and g__13238(w__12099 ,w__11827 ,w__11892);
  and g__13239(w__12098 ,w__11829 ,w__11907);
  not g__13240(w__12042 ,w__12043);
  not g__13241(w__12041 ,w__12040);
  not g__13242(w__12039 ,w__12038);
  or g__13243(w__12037 ,w__11917 ,w__11924);
  and g__13244(w__12036 ,w__11330 ,w__11845);
  or g__13245(w__12035 ,w__11592 ,w__11922);
  and g__13246(w__12034 ,w__11592 ,w__11922);
  and g__13247(w__12033 ,w__11917 ,w__11924);
  and g__13248(w__12032 ,w__11947 ,w__11952);
  or g__13249(w__12031 ,w__11594 ,w__11966);
  or g__13250(w__12030 ,w__11167 ,w__11855);
  nor g__13251(w__12029 ,w__11330 ,w__11845);
  or g__13252(w__12028 ,w__11877 ,w__11844);
  and g__13253(w__12027 ,w__11331 ,w__11855);
  or g__13254(w__12026 ,w__11851 ,w__11876);
  and g__13255(w__12025 ,w__11877 ,w__11844);
  and g__13256(w__12024 ,w__11339 ,w__11959);
  and g__13257(w__12023 ,w__11851 ,w__11876);
  and g__13258(w__12022 ,w__11594 ,w__11966);
  nor g__13259(w__12021 ,w__11850 ,w__11870);
  and g__13260(w__12020 ,w__11864 ,w__11880);
  or g__13261(w__12019 ,w__11336 ,w__11865);
  or g__13262(w__12018 ,w__11854 ,w__11852);
  or g__13263(w__12017 ,w__11596 ,w__11848);
  and g__13264(w__12016 ,w__11596 ,w__11848);
  and g__13265(w__12015 ,w__11859 ,w__11839);
  and g__13266(w__12014 ,w__11929 ,w__11847);
  nor g__13267(w__12013 ,w__11598 ,w__11881);
  and g__13268(w__12012 ,w__11874 ,w__11841);
  or g__13269(w__12011 ,w__11859 ,w__11839);
  or g__13270(w__12010 ,w__11842 ,w__11882);
  or g__13271(w__12009 ,w__11874 ,w__11841);
  or g__13272(w__12008 ,w__11863 ,w__11867);
  and g__13273(w__12007 ,w__11097 ,w__11928);
  and g__13274(w__12006 ,w__11854 ,w__11852);
  or g__13275(w__12005 ,w__11868 ,w__11866);
  nor g__13276(w__12004 ,w__11338 ,w__11879);
  nor g__13277(w__12003 ,w__11843 ,w__11883);
  or g__13278(w__12002 ,w__11860 ,w__11923);
  and g__13279(w__12001 ,w__11862 ,w__11853);
  or g__13280(w__12000 ,w__11862 ,w__11853);
  or g__13281(w__11999 ,w__11864 ,w__11880);
  or g__13282(w__11998 ,w__11334 ,w__11857);
  and g__13283(w__11997 ,w__11176 ,w__11861);
  or g__13284(w__11996 ,w__11172 ,w__11856);
  nor g__13285(w__11995 ,w__11335 ,w__11858);
  nor g__13286(w__11994 ,w__11176 ,w__11861);
  and g__13287(w__11993 ,w__11361 ,w__11856);
  or g__13288(w__11992 ,w__11174 ,w__11099);
  and g__13289(w__11991 ,w__11363 ,w__11099);
  or g__13290(w__11990 ,w__11168 ,w__11093);
  and g__13291(w__11989 ,w__11333 ,w__11836);
  or g__13292(w__11988 ,w__11337 ,w__11878);
  and g__13293(w__13057 ,w__11835 ,w__11913);
  and g__13294(w__12044 ,w__11833 ,w__11895);
  and g__13295(w__12043 ,w__11825 ,w__11904);
  and g__13296(w__12040 ,w__11831 ,w__11885);
  and g__13297(w__12038 ,w__11823 ,w__11888);
  not g__13298(w__11962 ,w__11963);
  not g__13299(w__11960 ,w__11961);
  not g__13300(w__11938 ,w__11939);
  not g__13301(w__11919 ,w__11920);
  not g__13302(w__11917 ,w__11918);
  not g__13303(w__11916 ,w__11915);
  or g__13304(w__11914 ,w__11605 ,w__11708);
  and g__13305(w__11987 ,w__11633 ,w__11737);
  and g__13306(w__11986 ,w__11656 ,w__11711);
  and g__13307(w__11985 ,w__11667 ,w__11750);
  and g__13308(w__11984 ,w__11544 ,w__11701);
  and g__13309(w__11983 ,w__11556 ,w__11714);
  and g__13310(w__11982 ,w__11655 ,w__11783);
  and g__13311(w__11981 ,w__11652 ,w__11784);
  and g__13312(w__11980 ,w__11651 ,w__11779);
  and g__13313(w__11979 ,w__11538 ,w__11689);
  and g__13314(w__11978 ,w__11649 ,w__11710);
  and g__13315(w__11977 ,w__11641 ,w__11765);
  and g__13316(w__11976 ,w__11643 ,w__11772);
  and g__13317(w__11975 ,w__11662 ,w__11770);
  and g__13318(w__11974 ,w__11638 ,w__11768);
  and g__13319(w__11973 ,w__11612 ,w__11763);
  and g__13320(w__11972 ,w__11647 ,w__11747);
  and g__13321(w__11971 ,w__11623 ,w__11820);
  and g__13322(w__11970 ,w__11627 ,w__11756);
  and g__13323(w__11969 ,w__11632 ,w__11729);
  and g__13324(w__11968 ,w__11582 ,w__11796);
  and g__13325(w__11967 ,w__11654 ,w__11782);
  and g__13326(w__11966 ,w__11575 ,w__11735);
  and g__13327(w__11965 ,w__11619 ,w__11794);
  or g__13328(w__11964 ,w__11601 ,w__11707);
  and g__13329(w__11963 ,w__11566 ,w__11777);
  and g__13330(w__11961 ,w__11568 ,w__11776);
  or g__13331(w__11959 ,w__11610 ,w__11704);
  and g__13332(w__11958 ,w__11645 ,w__11773);
  or g__13333(w__11957 ,w__11608 ,w__11706);
  and g__13334(w__11956 ,w__11660 ,w__11774);
  and g__13335(w__11955 ,w__11661 ,w__11791);
  and g__13336(w__11954 ,w__11644 ,w__11771);
  and g__13337(w__11953 ,w__11658 ,w__11790);
  and g__13338(w__11952 ,w__11624 ,w__11748);
  and g__13339(w__11951 ,w__11639 ,w__11715);
  and g__13340(w__11950 ,w__11553 ,w__11787);
  and g__13341(w__11949 ,w__11539 ,w__11697);
  or g__13342(w__11948 ,w__11603 ,w__11705);
  and g__13343(w__11947 ,w__11620 ,w__11749);
  and g__13344(w__11946 ,w__11548 ,w__11696);
  and g__13345(w__11945 ,w__11554 ,w__11769);
  and g__13346(w__11944 ,w__11631 ,w__11761);
  and g__13347(w__11943 ,w__11630 ,w__11760);
  and g__13348(w__11942 ,w__11546 ,w__11698);
  and g__13349(w__11941 ,w__11558 ,w__11733);
  and g__13350(w__11940 ,w__11569 ,w__11799);
  and g__13351(w__11939 ,w__11625 ,w__11807);
  and g__13352(w__11937 ,w__11572 ,w__11813);
  and g__13353(w__11936 ,w__11653 ,w__11785);
  and g__13354(w__11935 ,w__11628 ,w__11821);
  and g__13355(w__11934 ,w__11615 ,w__11795);
  and g__13356(w__11933 ,w__11622 ,w__11817);
  and g__13357(w__11932 ,w__11585 ,w__11686);
  or g__13358(w__11931 ,w__11599 ,w__11703);
  or g__13359(w__11930 ,w__11606 ,w__11702);
  and g__13360(w__11929 ,w__11584 ,w__11717);
  and g__13361(w__11928 ,w__11540 ,w__11700);
  and g__13362(w__11927 ,w__11613 ,w__11753);
  and g__13363(w__11926 ,w__11576 ,w__11746);
  and g__13364(w__11925 ,w__11614 ,w__11754);
  and g__13365(w__11924 ,w__11545 ,w__11693);
  and g__13366(w__11923 ,w__11571 ,w__11758);
  and g__13367(w__11922 ,w__11664 ,w__11752);
  and g__13368(w__11921 ,w__11659 ,w__11751);
  and g__13369(w__11920 ,w__11550 ,w__11699);
  and g__13370(w__11918 ,w__11636 ,w__11767);
  and g__13371(w__11915 ,w__11617 ,w__11755);
  not g__13372(w__11907 ,w__11906);
  not g__13373(w__11904 ,w__11903);
  not g__13374(w__11895 ,w__11894);
  not g__13375(w__11892 ,w__11891);
  not g__13376(w__11885 ,w__11884);
  not g__13377(w__11882 ,w__11883);
  not g__13378(w__11878 ,w__11879);
  not g__13379(w__11869 ,w__11870);
  not g__13380(w__11857 ,w__11858);
  not g__13381(w__11849 ,w__11850);
  not g__13382(w__11842 ,w__11843);
  not g__13383(w__11839 ,w__11838);
  not g__13384(w__11837 ,w__11836);
  or g__13385(w__13114 ,w__11679 ,w__11810);
  or g__13386(w__13115 ,w__11673 ,w__11786);
  or g__13387(w__13058 ,w__11665 ,w__11720);
  or g__13388(w__11913 ,w__11680 ,w__11802);
  and g__13389(w__11912 ,w__11634 ,w__11766);
  and g__13390(w__11911 ,w__11626 ,w__11730);
  and g__13391(w__11910 ,w__11683 ,w__11792);
  and g__13392(w__11909 ,w__11542 ,w__11695);
  and g__13393(w__11908 ,w__11563 ,w__11721);
  and g__13394(w__11906 ,w__11577 ,w__11812);
  and g__13395(w__11905 ,w__11670 ,w__11808);
  and g__13396(w__11903 ,w__11669 ,w__11801);
  and g__13397(w__11902 ,w__11552 ,w__11692);
  and g__13398(w__11901 ,w__11607 ,w__11805);
  and g__13399(w__11900 ,w__11541 ,w__11690);
  and g__13400(w__11899 ,w__11635 ,w__11798);
  and g__13401(w__11898 ,w__11681 ,w__11818);
  and g__13402(w__11897 ,w__11682 ,w__11806);
  and g__13403(w__11896 ,w__11677 ,w__11815);
  and g__13404(w__11894 ,w__11676 ,w__11814);
  and g__13405(w__11893 ,w__11678 ,w__11809);
  and g__13406(w__11891 ,w__11674 ,w__11816);
  and g__13407(w__11890 ,w__11672 ,w__11811);
  and g__13408(w__11889 ,w__11671 ,w__11819);
  or g__13409(w__11888 ,w__11646 ,w__11804);
  and g__13410(w__11887 ,w__11675 ,w__11803);
  and g__13411(w__11886 ,w__11543 ,w__11691);
  and g__13412(w__11884 ,w__11616 ,w__11743);
  and g__13413(w__11883 ,w__11621 ,w__11722);
  and g__13414(w__11881 ,w__11565 ,w__11724);
  and g__13415(w__11880 ,w__11629 ,w__11788);
  or g__13416(w__11879 ,w__11340 ,w__11800);
  and g__13417(w__11877 ,w__11637 ,w__11742);
  and g__13418(w__11876 ,w__11657 ,w__11778);
  and g__13419(w__11875 ,w__11583 ,w__11764);
  and g__13420(w__11874 ,w__11555 ,w__11775);
  and g__13421(w__11873 ,w__11578 ,w__11738);
  and g__13422(w__11872 ,w__11579 ,w__11736);
  and g__13423(w__11871 ,w__11663 ,w__11740);
  and g__13424(w__11870 ,w__11567 ,w__11739);
  and g__13425(w__11868 ,w__11564 ,w__11712);
  and g__13426(w__11867 ,w__11559 ,w__11793);
  and g__13427(w__11866 ,w__11549 ,w__11757);
  and g__13428(w__11865 ,w__11573 ,w__11716);
  and g__13429(w__11864 ,w__11562 ,w__11744);
  and g__13430(w__11863 ,w__11557 ,w__11713);
  and g__13431(w__11862 ,w__11642 ,w__11789);
  and g__13432(w__11861 ,w__11611 ,w__11797);
  and g__13433(w__11860 ,w__11600 ,w__11781);
  and g__13434(w__11859 ,w__11604 ,w__11762);
  and g__13435(w__11858 ,w__11609 ,w__11780);
  and g__13436(w__11856 ,w__11602 ,w__11719);
  and g__13437(w__11855 ,w__11581 ,w__11745);
  and g__13438(w__11854 ,w__11666 ,w__11732);
  and g__13439(w__11853 ,w__11551 ,w__11687);
  and g__13440(w__11852 ,w__11580 ,w__11731);
  and g__13441(w__11850 ,w__11574 ,w__11734);
  and g__13442(w__11848 ,w__11640 ,w__11727);
  and g__13443(w__11847 ,w__11618 ,w__11726);
  and g__13444(w__11846 ,w__11648 ,w__11725);
  or g__13445(w__11845 ,w__11605 ,w__11694);
  and g__13446(w__11844 ,w__11650 ,w__11741);
  and g__13447(w__11843 ,w__11668 ,w__11723);
  and g__13448(w__11841 ,w__11547 ,w__11688);
  and g__13449(w__11840 ,w__11560 ,w__11728);
  and g__13450(w__11838 ,w__11561 ,w__11759);
  and g__13451(w__11836 ,w__11570 ,w__11718);
  not g__13452(w__11835 ,w__11834);
  not g__13453(w__11833 ,w__11832);
  not g__13454(w__11831 ,w__11830);
  not g__13455(w__11829 ,w__11828);
  not g__13456(w__11827 ,w__11826);
  not g__13457(w__11825 ,w__11824);
  not g__13458(w__11823 ,w__11822);
  or g__13459(w__11821 ,w__11425 ,w__11011);
  or g__13460(w__11820 ,w__11439 ,w__10996);
  or g__13461(w__11819 ,w__11401 ,w__10970);
  or g__13462(w__11818 ,w__11389 ,w__11062);
  or g__13463(w__11817 ,w__11497 ,w__10993);
  or g__13464(w__11816 ,w__11394 ,w__10970);
  or g__13465(w__11815 ,w__11396 ,w__11037);
  or g__13466(w__11814 ,w__11390 ,w__11058);
  or g__13467(w__11813 ,w__11387 ,w__11053);
  or g__13468(w__11812 ,w__11422 ,w__10989);
  or g__13469(w__11811 ,w__11398 ,w__11059);
  nor g__13470(w__11810 ,w__11061 ,w__11391);
  or g__13471(w__11809 ,w__11392 ,w__11037);
  or g__13472(w__11808 ,w__11397 ,w__11038);
  or g__13473(w__11807 ,w__11393 ,w__11050);
  or g__13474(w__11806 ,w__11399 ,w__11061);
  or g__13475(w__11805 ,w__11448 ,w__11055);
  nor g__13476(w__11804 ,w__11059 ,w__11403);
  or g__13477(w__11803 ,w__11400 ,w__11089);
  nor g__13478(w__11802 ,w__11062 ,w__11402);
  or g__13479(w__11801 ,w__11395 ,w__11088);
  nor g__13480(w__11800 ,w__11058 ,w__11388);
  or g__13481(w__11799 ,w__11518 ,w__11002);
  or g__13482(w__11798 ,w__11474 ,w__10981);
  or g__13483(w__11797 ,w__11475 ,w__11029);
  or g__13484(w__11796 ,w__11520 ,w__11008);
  or g__13485(w__11795 ,w__11484 ,w__11005);
  or g__13486(w__11794 ,w__11449 ,w__11023);
  or g__13487(w__11793 ,w__11407 ,w__11052);
  or g__13488(w__11792 ,w__11412 ,w__10984);
  or g__13489(w__11791 ,w__11479 ,w__11028);
  or g__13490(w__11790 ,w__11501 ,w__11070);
  or g__13491(w__11789 ,w__11436 ,w__11064);
  or g__13492(w__11788 ,w__11490 ,w__10987);
  or g__13493(w__11787 ,w__11515 ,w__11026);
  nor g__13494(w__11786 ,w__11038 ,w__11365);
  or g__13495(w__11785 ,w__11496 ,w__11082);
  or g__13496(w__11784 ,w__11480 ,w__11022);
  or g__13497(w__11783 ,w__11444 ,w__10983);
  or g__13498(w__11782 ,w__11414 ,w__11067);
  or g__13499(w__11781 ,w__11506 ,w__11049);
  or g__13500(w__11780 ,w__11498 ,w__10978);
  or g__13501(w__11779 ,w__11491 ,w__10986);
  or g__13502(w__11778 ,w__11500 ,w__11005);
  or g__13503(w__11777 ,w__11521 ,w__10981);
  or g__13504(w__11776 ,w__11492 ,w__11007);
  or g__13505(w__11775 ,w__11424 ,w__11004);
  or g__13506(w__11774 ,w__11367 ,w__10980);
  or g__13507(w__11773 ,w__11488 ,w__10996);
  or g__13508(w__11772 ,w__11489 ,w__11025);
  or g__13509(w__11771 ,w__11493 ,w__10995);
  or g__13510(w__11770 ,w__11483 ,w__11079);
  or g__13511(w__11769 ,w__11519 ,w__11073);
  or g__13512(w__11768 ,w__11481 ,w__11004);
  or g__13513(w__11767 ,w__11478 ,w__10987);
  or g__13514(w__11766 ,w__11432 ,w__10995);
  or g__13515(w__11765 ,w__11430 ,w__10980);
  or g__13516(w__11764 ,w__11440 ,w__10977);
  or g__13517(w__11763 ,w__11442 ,w__11055);
  or g__13518(w__11762 ,w__11406 ,w__11022);
  or g__13519(w__11761 ,w__11485 ,w__11008);
  or g__13520(w__11760 ,w__11504 ,w__11067);
  or g__13521(w__11759 ,w__11482 ,w__11052);
  or g__13522(w__11758 ,w__11445 ,w__10993);
  or g__13523(w__11834 ,w__11325 ,w__11536);
  or g__13524(w__11832 ,w__11350 ,w__11533);
  or g__13525(w__11830 ,w__11318 ,w__11534);
  or g__13526(w__11828 ,w__11323 ,w__11532);
  or g__13527(w__11826 ,w__11321 ,w__11531);
  or g__13528(w__11824 ,w__11326 ,w__11537);
  or g__13529(w__11822 ,w__11315 ,w__11535);
  or g__13530(w__11757 ,w__11460 ,w__11013);
  or g__13531(w__11756 ,w__11421 ,w__10984);
  or g__13532(w__11755 ,w__11427 ,w__11028);
  or g__13533(w__11754 ,w__11437 ,w__11001);
  or g__13534(w__11753 ,w__11429 ,w__10992);
  or g__13535(w__11752 ,w__11507 ,w__10992);
  or g__13536(w__11751 ,w__11502 ,w__10978);
  or g__13537(w__11750 ,w__11450 ,w__10964);
  or g__13538(w__11749 ,w__11438 ,w__10986);
  or g__13539(w__11748 ,w__11510 ,w__11011);
  or g__13540(w__11747 ,w__11415 ,w__11064);
  or g__13541(w__11746 ,w__11368 ,w__11007);
  or g__13542(w__11745 ,w__11435 ,w__11071);
  or g__13543(w__11744 ,w__11486 ,w__11082);
  or g__13544(w__11743 ,w__11508 ,w__10990);
  or g__13545(w__11742 ,w__11455 ,w__10966);
  or g__13546(w__11741 ,w__11405 ,w__11025);
  or g__13547(w__11740 ,w__11513 ,w__11010);
  or g__13548(w__11739 ,w__11420 ,w__10964);
  or g__13549(w__11738 ,w__11404 ,w__11040);
  or g__13550(w__11737 ,w__11446 ,w__11010);
  or g__13551(w__11736 ,w__11428 ,w__11002);
  or g__13552(w__11735 ,w__11417 ,w__11073);
  or g__13553(w__11734 ,w__11434 ,w__11049);
  or g__13554(w__11733 ,w__11416 ,w__10966);
  or g__13555(w__11732 ,w__11364 ,w__10977);
  or g__13556(w__11731 ,w__11517 ,w__11041);
  or g__13557(w__11730 ,w__11418 ,w__11040);
  or g__13558(w__11729 ,w__11410 ,w__11079);
  or g__13559(w__11728 ,w__11477 ,w__11068);
  or g__13560(w__11727 ,w__11431 ,w__10990);
  or g__13561(w__11726 ,w__11487 ,w__11001);
  or g__13562(w__11725 ,w__11495 ,w__10958);
  or g__13563(w__11724 ,w__11426 ,w__11056);
  or g__13564(w__11723 ,w__11452 ,w__10958);
  or g__13565(w__11722 ,w__11516 ,w__10989);
  or g__13566(w__11721 ,w__11411 ,w__10962);
  nor g__13567(w__11720 ,w__11056 ,w__11457);
  or g__13568(w__11719 ,w__11441 ,w__10968);
  or g__13569(w__11718 ,w__11514 ,w__10968);
  or g__13570(w__11717 ,w__11443 ,w__11065);
  or g__13571(w__11716 ,w__11433 ,w__10983);
  or g__13572(w__11715 ,w__11409 ,w__10956);
  or g__13573(w__11714 ,w__11408 ,w__11070);
  or g__13574(w__11713 ,w__11523 ,w__10956);
  or g__13575(w__11712 ,w__11419 ,w__10962);
  or g__13576(w__11711 ,w__11423 ,w__11083);
  or g__13577(w__11710 ,w__11413 ,w__11080);
  nor g__13578(w__11708 ,w__11047 ,w__11017);
  nor g__13579(w__11707 ,w__11053 ,w__11302);
  nor g__13580(w__11706 ,w__11026 ,w__11305);
  nor g__13581(w__11705 ,w__11023 ,w__11303);
  nor g__13582(w__11704 ,w__11029 ,w__11290);
  nor g__13583(w__11703 ,w__11050 ,w__11304);
  nor g__13584(w__11702 ,w__11041 ,w__11306);
  or g__13585(w__11701 ,w__11512 ,w__11014);
  or g__13586(w__11700 ,w__11509 ,w__11019);
  or g__13587(w__11699 ,w__11503 ,w__11016);
  or g__13588(w__11698 ,w__11511 ,w__11013);
  or g__13589(w__11697 ,w__11499 ,w__11014);
  or g__13590(w__11696 ,w__11525 ,w__10954);
  or g__13591(w__11695 ,w__11476 ,w__11086);
  nor g__13592(w__11694 ,w__11020 ,w__11494);
  or g__13593(w__11693 ,w__11505 ,w__11019);
  or g__13594(w__11692 ,w__11522 ,w__11016);
  or g__13595(w__11691 ,w__11527 ,w__11020);
  or g__13596(w__11690 ,w__11528 ,w__11085);
  or g__13597(w__11689 ,w__11526 ,w__11085);
  or g__13598(w__11688 ,w__11529 ,w__11017);
  or g__13599(w__11687 ,w__11524 ,w__10954);
  or g__13600(w__11686 ,w__11447 ,w__11074);
  or g__13601(w__11683 ,w__11496 ,w__11214);
  or g__13602(w__11682 ,w__11044 ,w__11390);
  or g__13603(w__11681 ,w__11032 ,w__11395);
  nor g__13604(w__11680 ,w__11044 ,w__11400);
  nor g__13605(w__11679 ,w__11032 ,w__11402);
  or g__13606(w__11678 ,w__11031 ,w__11396);
  or g__13607(w__11677 ,w__11043 ,w__11394);
  or g__13608(w__11676 ,w__11034 ,w__11397);
  or g__13609(w__11675 ,w__11043 ,w__11403);
  or g__13610(w__11674 ,w__11031 ,w__11389);
  nor g__13611(w__11673 ,w__11035 ,w__11391);
  or g__13612(w__11672 ,w__11034 ,w__11401);
  or g__13613(w__11671 ,w__11035 ,w__11392);
  or g__13614(w__11670 ,w__10972 ,w__11398);
  or g__13615(w__11669 ,w__10972 ,w__11388);
  or g__13616(w__11668 ,w__11495 ,w__11253);
  or g__13617(w__11667 ,w__11422 ,w__11238);
  or g__13618(w__11666 ,w__11417 ,w__11202);
  nor g__13619(w__11665 ,w__11426 ,w__11245);
  or g__13620(w__11664 ,w__11447 ,w__11211);
  or g__13621(w__11663 ,w__11487 ,w__11256);
  or g__13622(w__11662 ,w__11425 ,w__11256);
  or g__13623(w__11661 ,w__11430 ,w__11223);
  or g__13624(w__11660 ,w__11521 ,w__11223);
  or g__13625(w__11659 ,w__11497 ,w__11211);
  or g__13626(w__11658 ,w__11408 ,w__11244);
  or g__13627(w__11657 ,w__11478 ,w__11226);
  or g__13628(w__11656 ,w__11427 ,w__11215);
  or g__13629(w__11655 ,w__11475 ,w__11218);
  or g__13630(w__11654 ,w__11449 ,w__11232);
  or g__13631(w__11653 ,w__11433 ,w__11214);
  or g__13632(w__11652 ,w__11416 ,w__11232);
  or g__13633(w__11651 ,w__11406 ,w__11227);
  or g__13634(w__11650 ,w__11507 ,w__11203);
  or g__13635(w__11649 ,w__11506 ,w__11254);
  or g__13636(w__11648 ,w__11410 ,w__11253);
  or g__13637(w__11647 ,w__11436 ,w__11178);
  nor g__13638(w__11646 ,w__11117 ,w__11399);
  or g__13639(w__11645 ,w__11514 ,w__11187);
  or g__13640(w__11644 ,w__11492 ,w__11187);
  or g__13641(w__11643 ,w__11445 ,w__11206);
  or g__13642(w__11642 ,w__11432 ,w__11179);
  or g__13643(w__11641 ,w__11523 ,w__11217);
  or g__13644(w__11640 ,w__11517 ,w__11239);
  or g__13645(w__11639 ,w__11474 ,w__11220);
  or g__13646(w__11638 ,w__11480 ,w__11230);
  or g__13647(w__11637 ,w__11438 ,w__11226);
  or g__13648(w__11636 ,w__11414 ,w__11229);
  or g__13649(w__11635 ,w__11486 ,w__11220);
  or g__13650(w__11634 ,w__11482 ,w__11182);
  or g__13651(w__11633 ,w__11518 ,w__11250);
  or g__13652(w__11632 ,w__11434 ,w__11381);
  or g__13653(w__11631 ,w__11493 ,w__11178);
  or g__13654(w__11630 ,w__11481 ,w__11235);
  or g__13655(w__11629 ,w__11477 ,w__11235);
  or g__13656(w__11628 ,w__11513 ,w__11250);
  or g__13657(w__11627 ,w__11409 ,w__11217);
  or g__13658(w__11626 ,w__11435 ,w__11242);
  or g__13659(w__11625 ,w__11483 ,w__11251);
  or g__13660(w__11624 ,w__11437 ,w__11254);
  or g__13661(w__11623 ,w__11441 ,w__11181);
  or g__13662(w__11622 ,w__11489 ,w__11202);
  or g__13663(w__11621 ,w__11431 ,w__11238);
  or g__13664(w__11620 ,w__11484 ,w__11229);
  or g__13665(w__11619 ,w__11490 ,w__11233);
  or g__13666(w__11618 ,w__11446 ,w__11257);
  or g__13667(w__11617 ,w__11444 ,w__11224);
  or g__13668(w__11616 ,w__11450 ,w__11241);
  or g__13669(w__11615 ,w__11504 ,w__11230);
  or g__13670(w__11614 ,w__11393 ,w__11147);
  or g__13671(w__11613 ,w__11498 ,w__11205);
  or g__13672(w__11612 ,w__11404 ,w__11248);
  or g__13673(w__11685 ,w__11370 ,w__11106);
  or g__13674(w__11684 ,in25[0] ,w__11459);
  not g__13675(w__11611 ,w__11610);
  not g__13676(w__11609 ,w__11608);
  not g__13677(w__11607 ,w__11606);
  not g__13678(w__11604 ,w__11603);
  not g__13679(w__11602 ,w__11601);
  not g__13680(w__11600 ,w__11599);
  not g__13681(w__11598 ,w__11597);
  or g__13682(w__11585 ,w__11440 ,w__11208);
  or g__13683(w__11584 ,w__11407 ,w__11184);
  or g__13684(w__11583 ,w__11519 ,w__11208);
  or g__13685(w__11582 ,w__11443 ,w__11184);
  or g__13686(w__11581 ,w__11448 ,w__11247);
  or g__13687(w__11580 ,w__11420 ,w__11241);
  or g__13688(w__11579 ,w__11510 ,w__11147);
  or g__13689(w__11578 ,w__11501 ,w__11244);
  or g__13690(w__11577 ,w__11442 ,w__11242);
  or g__13691(w__11576 ,w__11485 ,w__11181);
  or g__13692(w__11575 ,w__11405 ,w__11205);
  or g__13693(w__11574 ,w__11428 ,w__11257);
  or g__13694(w__11573 ,w__11423 ,w__11218);
  or g__13695(w__11572 ,w__11488 ,w__11188);
  or g__13696(w__11571 ,w__11429 ,w__11212);
  or g__13697(w__11570 ,w__11415 ,w__11182);
  or g__13698(w__11569 ,w__11413 ,w__11251);
  or g__13699(w__11568 ,w__11520 ,w__11185);
  or g__13700(w__11567 ,w__11508 ,w__11247);
  or g__13701(w__11566 ,w__11479 ,w__11221);
  or g__13702(w__11565 ,w__11516 ,w__11239);
  or g__13703(w__11564 ,w__11411 ,w__11206);
  or g__13704(w__11563 ,w__11502 ,w__11209);
  or g__13705(w__11562 ,w__11412 ,w__11215);
  or g__13706(w__11561 ,w__11439 ,w__11179);
  or g__13707(w__11560 ,w__11491 ,w__11236);
  or g__13708(w__11559 ,w__11387 ,w__11188);
  or g__13709(w__11558 ,w__11424 ,w__11227);
  or g__13710(w__11557 ,w__11421 ,w__11224);
  or g__13711(w__11556 ,w__11418 ,w__11245);
  or g__13712(w__11555 ,w__11500 ,w__11233);
  or g__13713(w__11554 ,w__11515 ,w__11203);
  or g__13714(w__11553 ,w__11419 ,w__11212);
  or g__13715(w__11552 ,w__11190 ,w__11509);
  or g__13716(w__11551 ,w__11199 ,w__11525);
  or g__13717(w__11550 ,w__11199 ,w__11476);
  or g__13718(w__11549 ,w__11191 ,w__11529);
  or g__13719(w__11548 ,w__11194 ,w__11526);
  or g__13720(w__11547 ,w__11190 ,w__11527);
  or g__13721(w__11546 ,w__11193 ,w__11522);
  or g__13722(w__11545 ,w__11196 ,w__11499);
  or g__13723(w__11544 ,w__11196 ,w__11528);
  or g__13724(w__11543 ,w__11193 ,w__11505);
  or g__13725(w__11542 ,w__11200 ,w__11494);
  or g__13726(w__11541 ,w__11194 ,w__11524);
  or g__13727(w__11540 ,w__11197 ,w__11503);
  or g__13728(w__11539 ,w__11191 ,w__11512);
  or g__13729(w__11538 ,w__11200 ,w__11511);
  or g__13730(w__11537 ,w__11077 ,w__11463);
  or g__13731(w__11536 ,w__11306 ,w__11466);
  or g__13732(w__11535 ,w__11304 ,w__11467);
  or g__13733(w__11534 ,w__11303 ,w__11465);
  or g__13734(w__11533 ,w__11305 ,w__11461);
  or g__13735(w__11532 ,w__11302 ,w__11462);
  or g__13736(w__11531 ,w__11290 ,w__11464);
  nor g__13737(w__11530 ,w__11248 ,w__10943);
  and g__13738(w__11610 ,in25[13] ,w__11109);
  and g__13739(w__11608 ,in25[7] ,w__11107);
  and g__13740(w__11606 ,in25[3] ,w__11100);
  and g__13741(w__11605 ,in25[15] ,w__11108);
  and g__13742(w__11603 ,in25[9] ,w__11111);
  and g__13743(w__11601 ,in25[11] ,w__11105);
  and g__13744(w__11599 ,in25[5] ,w__11101);
  and g__13745(w__11597 ,in24[0] ,w__11115);
  or g__13746(w__11596 ,w__11091 ,w__11209);
  or g__13747(w__11595 ,w__11091 ,w__11197);
  or g__13748(w__11594 ,w__11307 ,w__11236);
  or g__13749(w__11593 ,w__11090 ,w__11221);
  or g__13750(w__11592 ,w__11090 ,w__11185);
  or g__13751(w__11591 ,w__11458 ,w__11103);
  or g__13752(w__11590 ,w__11453 ,w__11112);
  or g__13753(w__11589 ,w__11451 ,w__11102);
  or g__13754(w__11588 ,w__11366 ,w__11114);
  or g__13755(w__11587 ,w__11454 ,w__11110);
  or g__13756(w__11586 ,w__11369 ,w__11104);
  not g__13757(w__11473 ,w__11107);
  not g__13758(w__11472 ,w__11112);
  not g__13759(w__11470 ,w__11106);
  not g__13760(w__11469 ,w__11108);
  nor g__13761(w__11467 ,w__11155 ,w__11353);
  nor g__13762(w__11466 ,w__11291 ,w__11316);
  nor g__13763(w__11465 ,w__11153 ,w__11322);
  nor g__13764(w__11464 ,w__11151 ,w__11355);
  nor g__13765(w__11463 ,w__11149 ,w__11317);
  nor g__13766(w__11462 ,w__11157 ,w__11342);
  nor g__13767(w__11461 ,w__11159 ,w__11347);
  or g__13768(w__11460 ,w__11338 ,w__11327);
  xnor g__13769(w__11458 ,in25[13] ,in25[12]);
  xnor g__13770(w__11457 ,in24[0] ,in25[3]);
  nor g__13771(w__11456 ,w__13061 ,w__11161);
  xnor g__13772(w__11455 ,in24[0] ,in25[9]);
  xnor g__13773(w__11454 ,in25[9] ,in25[8]);
  xnor g__13774(w__11453 ,in25[7] ,in25[6]);
  xnor g__13775(w__11452 ,in24[0] ,in25[5]);
  xnor g__13776(w__11451 ,in25[3] ,in25[2]);
  or g__13777(w__11529 ,w__11259 ,w__11346);
  or g__13778(w__11528 ,w__11334 ,w__11343);
  or g__13779(w__11527 ,w__11260 ,w__11356);
  or g__13780(w__11526 ,w__11270 ,w__11351);
  or g__13781(w__11525 ,w__11262 ,w__11348);
  or g__13782(w__11524 ,w__11269 ,w__11344);
  xnor g__13783(w__11523 ,in24[4] ,in25[13]);
  or g__13784(w__11522 ,w__11267 ,w__11319);
  xnor g__13785(w__11521 ,in24[1] ,in25[13]);
  xnor g__13786(w__11520 ,in24[4] ,in25[11]);
  xnor g__13787(w__11519 ,in24[6] ,in25[7]);
  xnor g__13788(w__11518 ,in24[13] ,in25[5]);
  xnor g__13789(w__11517 ,in24[4] ,in25[3]);
  xnor g__13790(w__11516 ,in24[2] ,in25[3]);
  xnor g__13791(w__11515 ,in24[7] ,in25[7]);
  xnor g__13792(w__11514 ,in24[9] ,in25[11]);
  xnor g__13793(w__11513 ,in24[10] ,in25[5]);
  or g__13794(w__11512 ,w__11261 ,w__11352);
  or g__13795(w__11511 ,w__11268 ,w__11320);
  xnor g__13796(w__11510 ,in24[5] ,in25[5]);
  or g__13797(w__11509 ,w__11266 ,w__11324);
  xnor g__13798(w__11508 ,in24[6] ,in25[3]);
  xnor g__13799(w__11507 ,in24[3] ,in25[7]);
  xnor g__13800(w__11506 ,in24[15] ,in25[5]);
  or g__13801(w__11505 ,w__11264 ,w__11345);
  xnor g__13802(w__11504 ,in24[3] ,in25[9]);
  or g__13803(w__11503 ,w__11263 ,w__11349);
  xnor g__13804(w__11502 ,in24[10] ,in25[7]);
  xnor g__13805(w__11501 ,in24[11] ,in25[3]);
  xnor g__13806(w__11500 ,in24[8] ,in25[9]);
  or g__13807(w__11499 ,w__11265 ,w__11354);
  xnor g__13808(w__11498 ,in24[15] ,in25[7]);
  xnor g__13809(w__11497 ,in24[11] ,in25[7]);
  xnor g__13810(w__11496 ,in24[10] ,in25[13]);
  xnor g__13811(w__11495 ,in24[1] ,in25[5]);
  xnor g__13812(w__11494 ,in24[15] ,in25[15]);
  xnor g__13813(w__11493 ,in24[2] ,in25[11]);
  xnor g__13814(w__11492 ,in24[3] ,in25[11]);
  xnor g__13815(w__11491 ,in24[14] ,in25[9]);
  xnor g__13816(w__11490 ,in24[12] ,in25[9]);
  xnor g__13817(w__11489 ,in24[12] ,in25[7]);
  xnor g__13818(w__11488 ,in24[8] ,in25[11]);
  xnor g__13819(w__11487 ,in24[11] ,in25[5]);
  xnor g__13820(w__11486 ,in24[8] ,in25[13]);
  xnor g__13821(w__11485 ,in24[1] ,in25[11]);
  xnor g__13822(w__11484 ,in24[2] ,in25[9]);
  xnor g__13823(w__11483 ,in24[8] ,in25[5]);
  xnor g__13824(w__11482 ,in24[13] ,in25[11]);
  xnor g__13825(w__11481 ,in24[4] ,in25[9]);
  xnor g__13826(w__11480 ,in24[5] ,in25[9]);
  xnor g__13827(w__11479 ,in24[2] ,in25[13]);
  xnor g__13828(w__11478 ,in24[9] ,in25[9]);
  xnor g__13829(w__11477 ,in24[13] ,in25[9]);
  or g__13830(w__11476 ,w__11145 ,w__11328);
  xnor g__13831(w__11475 ,in24[15] ,in25[13]);
  xnor g__13832(w__11474 ,in24[7] ,in25[13]);
  xnor g__13833(w__11471 ,w__11159 ,in25[6]);
  xnor g__13834(w__11468 ,w__11149 ,in25[14]);
  not g__13835(w__11386 ,w__11105);
  not g__13836(w__11385 ,w__11104);
  not g__13837(w__11383 ,w__11115);
  not g__13838(w__11381 ,w__11101);
  not g__13839(w__11380 ,w__11114);
  not g__13840(w__11379 ,w__11100);
  not g__13841(w__11378 ,w__11102);
  not g__13842(w__11376 ,w__11111);
  not g__13843(w__11375 ,w__11110);
  not g__13844(w__11373 ,w__11109);
  not g__13845(w__11372 ,w__11103);
  xnor g__13846(w__11370 ,in25[15] ,in25[14]);
  xnor g__13847(w__11369 ,in25[11] ,in25[10]);
  xnor g__13848(w__11368 ,in24[0] ,in25[11]);
  xnor g__13849(w__11367 ,in24[0] ,in25[13]);
  xnor g__13850(w__11366 ,in25[5] ,in25[4]);
  xnor g__13851(w__11365 ,in24[0] ,in25[1]);
  xnor g__13852(w__11364 ,in24[0] ,in25[7]);
  xnor g__13853(w__11450 ,in24[7] ,in25[3]);
  xnor g__13854(w__11449 ,in24[11] ,in25[9]);
  xnor g__13855(w__11448 ,in24[15] ,in25[3]);
  xnor g__13856(w__11447 ,in24[4] ,in25[7]);
  xnor g__13857(w__11446 ,in24[12] ,in25[5]);
  xnor g__13858(w__11445 ,in24[13] ,in25[7]);
  xnor g__13859(w__11444 ,in24[14] ,in25[13]);
  xnor g__13860(w__11443 ,in24[5] ,in25[11]);
  xnor g__13861(w__11442 ,in24[9] ,in25[3]);
  xnor g__13862(w__11441 ,in24[15] ,in25[11]);
  xnor g__13863(w__11440 ,in24[5] ,in25[7]);
  xnor g__13864(w__11439 ,in24[14] ,in25[11]);
  xnor g__13865(w__11438 ,in24[1] ,in25[9]);
  xnor g__13866(w__11437 ,in24[6] ,in25[5]);
  xnor g__13867(w__11436 ,in24[11] ,in25[11]);
  xnor g__13868(w__11435 ,in24[14] ,in25[3]);
  xnor g__13869(w__11434 ,in24[3] ,in25[5]);
  xnor g__13870(w__11433 ,in24[11] ,in25[13]);
  xnor g__13871(w__11432 ,in24[12] ,in25[11]);
  xnor g__13872(w__11431 ,in24[3] ,in25[3]);
  xnor g__13873(w__11430 ,in24[3] ,in25[13]);
  xnor g__13874(w__11429 ,in24[14] ,in25[7]);
  xnor g__13875(w__11428 ,in24[4] ,in25[5]);
  xnor g__13876(w__11427 ,in24[13] ,in25[13]);
  xnor g__13877(w__11426 ,in24[1] ,in25[3]);
  xnor g__13878(w__11425 ,in24[9] ,in25[5]);
  xnor g__13879(w__11424 ,in24[7] ,in25[9]);
  xnor g__13880(w__11423 ,in24[12] ,in25[13]);
  xnor g__13881(w__11422 ,in24[8] ,in25[3]);
  xnor g__13882(w__11421 ,in24[5] ,in25[13]);
  xnor g__13883(w__11420 ,in24[5] ,in25[3]);
  xnor g__13884(w__11419 ,in24[8] ,in25[7]);
  xnor g__13885(w__11418 ,in24[13] ,in25[3]);
  xnor g__13886(w__11417 ,in24[1] ,in25[7]);
  xnor g__13887(w__11416 ,in24[6] ,in25[9]);
  xnor g__13888(w__11415 ,in24[10] ,in25[11]);
  xnor g__13889(w__11414 ,in24[10] ,in25[9]);
  xnor g__13890(w__11413 ,in24[14] ,in25[5]);
  xnor g__13891(w__11412 ,in24[9] ,in25[13]);
  xnor g__13892(w__11411 ,in24[9] ,in25[7]);
  xnor g__13893(w__11410 ,in24[2] ,in25[5]);
  xnor g__13894(w__11409 ,in24[6] ,in25[13]);
  xnor g__13895(w__11408 ,in24[12] ,in25[3]);
  xnor g__13896(w__11407 ,in24[6] ,in25[11]);
  xnor g__13897(w__11406 ,in24[15] ,in25[9]);
  xnor g__13898(w__11405 ,in24[2] ,in25[7]);
  xnor g__13899(w__11404 ,in24[10] ,in25[3]);
  xnor g__13900(w__11403 ,in24[4] ,in25[1]);
  xnor g__13901(w__11402 ,in24[2] ,in25[1]);
  xnor g__13902(w__11401 ,in24[9] ,in25[1]);
  xnor g__13903(w__11400 ,in24[3] ,in25[1]);
  xnor g__13904(w__11399 ,in24[5] ,in25[1]);
  xnor g__13905(w__11398 ,in24[8] ,in25[1]);
  xnor g__13906(w__11397 ,in24[7] ,in25[1]);
  xnor g__13907(w__11396 ,in24[11] ,in25[1]);
  xnor g__13908(w__11395 ,in24[14] ,in25[1]);
  xnor g__13909(w__11394 ,in24[12] ,in25[1]);
  xnor g__13910(w__11393 ,in24[7] ,in25[5]);
  xnor g__13911(w__11392 ,in24[10] ,in25[1]);
  xnor g__13912(w__11391 ,in24[1] ,in25[1]);
  xnor g__13913(w__11390 ,in24[6] ,in25[1]);
  xnor g__13914(w__11389 ,in24[13] ,in25[1]);
  xnor g__13915(w__11388 ,in24[15] ,in25[1]);
  xnor g__13916(w__11387 ,in24[7] ,in25[11]);
  xnor g__13917(w__11384 ,w__11157 ,in25[10]);
  xnor g__13918(w__11382 ,w__11155 ,in25[4]);
  xnor g__13919(w__11377 ,w__11161 ,in25[2]);
  xnor g__13920(w__11374 ,w__11153 ,in25[8]);
  xnor g__13921(w__11371 ,w__11151 ,in25[12]);
  nor g__13922(w__11356 ,in24[2] ,in25[15]);
  nor g__13923(w__11355 ,in24[0] ,in25[12]);
  nor g__13924(w__11354 ,in24[4] ,in25[15]);
  nor g__13925(w__11353 ,in24[0] ,in25[4]);
  nor g__13926(w__11352 ,in24[5] ,in25[15]);
  nor g__13927(w__11351 ,in24[9] ,in25[15]);
  and g__13928(w__11350 ,in24[0] ,in25[6]);
  nor g__13929(w__11349 ,in24[13] ,in25[15]);
  nor g__13930(w__11348 ,in24[8] ,in25[15]);
  nor g__13931(w__11347 ,in24[0] ,in25[6]);
  nor g__13932(w__11346 ,in24[1] ,in25[15]);
  nor g__13933(w__11345 ,in24[3] ,in25[15]);
  nor g__13934(w__11344 ,in24[7] ,in25[15]);
  nor g__13935(w__11343 ,in24[6] ,in25[15]);
  nor g__13936(w__11342 ,in24[0] ,in25[10]);
  or g__13937(w__11341 ,w__11311 ,w__10974);
  or g__13938(w__11363 ,w__11313 ,w__10998);
  or g__13939(w__11362 ,w__11314 ,w__11076);
  or g__13940(w__11361 ,w__11296 ,w__11046);
  or g__13941(w__11360 ,w__11300 ,w__10975);
  or g__13942(w__11359 ,w__11309 ,w__10999);
  or g__13943(w__11358 ,w__11308 ,w__10960);
  or g__13944(w__11357 ,w__11299 ,w__11046);
  not g__13945(w__11337 ,w__11338);
  not g__13946(w__11334 ,w__11335);
  not g__13947(w__11329 ,w__11330);
  nor g__13948(w__11328 ,in24[14] ,in25[15]);
  nor g__13949(w__11327 ,in24[0] ,in25[15]);
  and g__13950(w__11326 ,in24[0] ,in25[14]);
  and g__13951(w__11325 ,in24[0] ,in25[2]);
  nor g__13952(w__11324 ,in24[12] ,in25[15]);
  and g__13953(w__11323 ,in24[0] ,in25[10]);
  nor g__13954(w__11322 ,in24[0] ,in25[8]);
  and g__13955(w__11321 ,in24[0] ,in25[12]);
  nor g__13956(w__11320 ,in24[10] ,in25[15]);
  nor g__13957(w__11319 ,in24[11] ,in25[15]);
  and g__13958(w__11318 ,in24[0] ,in25[8]);
  nor g__13959(w__11317 ,in24[0] ,in25[14]);
  nor g__13960(w__11316 ,in24[0] ,in25[2]);
  and g__13961(w__11315 ,in24[0] ,in25[4]);
  and g__13962(w__13061 ,in24[0] ,in25[0]);
  and g__13963(w__11340 ,in25[1] ,in25[0]);
  or g__13964(w__11339 ,w__11297 ,w__10974);
  and g__13965(w__11338 ,in24[0] ,in25[15]);
  or g__13966(w__11336 ,w__11295 ,w__10998);
  or g__13967(w__11335 ,w__11310 ,w__11076);
  or g__13968(w__11333 ,w__11301 ,w__10999);
  or g__13969(w__11332 ,w__11294 ,w__10975);
  or g__13970(w__11331 ,w__11312 ,w__10960);
  or g__13971(w__11330 ,w__11298 ,w__11047);
  not g__13972(w__11314 ,in24[7]);
  not g__13973(w__11313 ,in24[9]);
  not g__13974(w__11312 ,in24[1]);
  not g__13975(w__11311 ,in24[15]);
  not g__13976(w__11310 ,in24[6]);
  not g__13977(w__11309 ,in24[12]);
  not g__13978(w__11308 ,in24[4]);
  not g__13979(w__11307 ,in24[0]);
  not g__13980(w__11306 ,in25[3]);
  not g__13981(w__11305 ,in25[7]);
  not g__13982(w__11304 ,in25[5]);
  not g__13983(w__11303 ,in25[9]);
  not g__13984(w__11302 ,in25[11]);
  not g__13985(w__11301 ,in24[5]);
  not g__13986(w__11300 ,in24[11]);
  not g__13987(w__11299 ,in24[3]);
  not g__13988(w__11298 ,in24[14]);
  not g__13989(w__11297 ,in24[13]);
  not g__13990(w__11296 ,in24[10]);
  not g__13991(w__11295 ,in24[8]);
  not g__13992(w__11294 ,in24[2]);
  not g__13993(w__11293 ,in25[0]);
  not g__13994(w__11292 ,in25[15]);
  not g__13995(w__11291 ,in25[1]);
  not g__13996(w__11290 ,in25[13]);
  not g__13997(w__10944 ,w__11258);
  not g__13998(w__11258 ,w__11307);
  not g__13999(w__11257 ,w__11255);
  not g__14000(w__11256 ,w__11255);
  not g__14001(w__11255 ,w__11277);
  not g__14002(w__11254 ,w__11252);
  not g__14003(w__11253 ,w__11252);
  not g__14004(w__11252 ,w__11383);
  not g__14005(w__11251 ,w__11249);
  not g__14006(w__11250 ,w__11249);
  not g__14007(w__11249 ,w__11380);
  not g__14008(w__11248 ,w__11246);
  not g__14009(w__11247 ,w__11246);
  not g__14010(w__11246 ,w__11378);
  not g__14011(w__11245 ,w__11243);
  not g__14012(w__11244 ,w__11243);
  not g__14013(w__11243 ,w__11379);
  not g__14014(w__11242 ,w__11240);
  not g__14015(w__11241 ,w__11240);
  not g__14016(w__11240 ,w__11276);
  not g__14017(w__11239 ,w__11237);
  not g__14018(w__11238 ,w__11237);
  not g__14019(w__11237 ,w__11275);
  not g__14020(w__11236 ,w__11234);
  not g__14021(w__11235 ,w__11234);
  not g__14022(w__11234 ,w__11375);
  not g__14023(w__11233 ,w__11231);
  not g__14024(w__11232 ,w__11231);
  not g__14025(w__11231 ,w__11376);
  not g__14026(w__11230 ,w__11228);
  not g__14027(w__11229 ,w__11228);
  not g__14028(w__11228 ,w__11274);
  not g__14029(w__11227 ,w__11225);
  not g__14030(w__11226 ,w__11225);
  not g__14031(w__11225 ,w__11273);
  not g__14032(w__11224 ,w__11222);
  not g__14033(w__11223 ,w__11222);
  not g__14034(w__11222 ,w__11373);
  not g__14035(w__11221 ,w__11219);
  not g__14036(w__11220 ,w__11219);
  not g__14037(w__11219 ,w__11372);
  not g__14038(w__11218 ,w__11216);
  not g__14039(w__11217 ,w__11216);
  not g__14040(w__11216 ,w__11272);
  not g__14041(w__11215 ,w__11213);
  not g__14042(w__11214 ,w__11213);
  not g__14043(w__11213 ,w__11271);
  not g__14044(w__11212 ,w__11210);
  not g__14045(w__11211 ,w__11210);
  not g__14046(w__11210 ,w__11473);
  not g__14047(w__11209 ,w__11207);
  not g__14048(w__11208 ,w__11207);
  not g__14049(w__11207 ,w__11472);
  not g__14050(w__11206 ,w__11204);
  not g__14051(w__11205 ,w__11204);
  not g__14052(w__11204 ,w__11283);
  not g__14053(w__11203 ,w__11201);
  not g__14054(w__11202 ,w__11201);
  not g__14055(w__11201 ,w__11282);
  not g__14056(w__11200 ,w__11198);
  not g__14057(w__11199 ,w__11198);
  not g__14058(w__11198 ,w__11470);
  not g__14059(w__11197 ,w__11195);
  not g__14060(w__11196 ,w__11195);
  not g__14061(w__11195 ,w__11469);
  not g__14062(w__11194 ,w__11192);
  not g__14063(w__11193 ,w__11192);
  not g__14064(w__11192 ,w__11281);
  not g__14065(w__11191 ,w__11189);
  not g__14066(w__11190 ,w__11189);
  not g__14067(w__11189 ,w__11280);
  not g__14068(w__11188 ,w__11186);
  not g__14069(w__11187 ,w__11186);
  not g__14070(w__11186 ,w__11386);
  not g__14071(w__11185 ,w__11183);
  not g__14072(w__11184 ,w__11183);
  not g__14073(w__11183 ,w__11385);
  not g__14074(w__11182 ,w__11180);
  not g__14075(w__11181 ,w__11180);
  not g__14076(w__11180 ,w__11279);
  not g__14077(w__11179 ,w__11177);
  not g__14078(w__11178 ,w__11177);
  not g__14079(w__11177 ,w__11278);
  not g__14080(w__11176 ,w__11266);
  not g__14081(w__11266 ,w__11359);
  not g__14082(w__11175 ,w__11263);
  not g__14083(w__11263 ,w__11339);
  not g__14084(w__11174 ,w__11270);
  not g__14085(w__11270 ,w__11363);
  not g__14086(w__11173 ,w__11267);
  not g__14087(w__11267 ,w__11360);
  not g__14088(w__11172 ,w__11268);
  not g__14089(w__11268 ,w__11361);
  not g__14090(w__11171 ,w__11264);
  not g__14091(w__11264 ,w__11357);
  not g__14092(w__11170 ,w__11262);
  not g__14093(w__11262 ,w__11336);
  not g__14094(w__11169 ,w__11260);
  not g__14095(w__11260 ,w__11332);
  not g__14096(w__11168 ,w__11261);
  not g__14097(w__11261 ,w__11333);
  not g__14098(w__11167 ,w__11259);
  not g__14099(w__11259 ,w__11331);
  not g__14100(w__11166 ,w__11265);
  not g__14101(w__11265 ,w__11358);
  not g__14102(w__11165 ,w__11269);
  not g__14103(w__11269 ,w__11362);
  not g__14104(w__11164 ,w__11163);
  not g__14105(w__11163 ,w__11918);
  not g__14106(w__11162 ,w__11284);
  not g__14107(w__11284 ,w__11921);
  not g__14108(w__11161 ,w__11160);
  not g__14109(w__11160 ,w__11291);
  not g__14110(w__11159 ,w__11158);
  not g__14111(w__11158 ,w__11304);
  not g__14112(w__11157 ,w__11156);
  not g__14113(w__11156 ,w__11303);
  not g__14114(w__11155 ,w__11154);
  not g__14115(w__11154 ,w__11306);
  not g__14116(w__11153 ,w__11152);
  not g__14117(w__11152 ,w__11305);
  not g__14118(w__11151 ,w__11150);
  not g__14119(w__11150 ,w__11302);
  not g__14120(w__11149 ,w__11148);
  not g__14121(w__11148 ,w__11290);
  not g__14122(w__11147 ,w__11146);
  not g__14123(w__11146 ,w__11381);
  buf g__14124(w__13059 ,w__11530);
  buf g__14125(w__13060 ,w__11456);
  not g__14126(w__11145 ,w__11144);
  not g__14127(w__11144 ,w__11329);
  not g__14128(w__11143 ,w__11142);
  not g__14129(w__11142 ,w__11919);
  not g__14130(w__11141 ,w__11286);
  not g__14131(w__11286 ,w__12275);
  not g__14132(w__11140 ,w__11287);
  not g__14133(w__11287 ,w__12291);
  not g__14134(w__11139 ,w__11288);
  not g__14135(w__11288 ,w__12531);
  not g__14136(w__11138 ,w__11285);
  not g__14137(w__11285 ,w__12274);
  not g__14138(w__11137 ,w__11289);
  not g__14139(w__11289 ,w__12532);
  not g__14140(w__11136 ,w__11135);
  not g__14141(w__11135 ,w__11684);
  not g__14142(w__11134 ,w__11133);
  not g__14143(w__11133 ,w__11591);
  not g__14144(w__11132 ,w__11131);
  not g__14145(w__11131 ,w__11590);
  not g__14146(w__11130 ,w__11129);
  not g__14147(w__11129 ,w__11587);
  not g__14148(w__11128 ,w__11127);
  not g__14149(w__11127 ,w__11586);
  not g__14150(w__11126 ,w__11125);
  not g__14151(w__11125 ,w__11589);
  not g__14152(w__11124 ,w__11123);
  not g__14153(w__11123 ,w__11588);
  not g__14154(w__11122 ,w__11121);
  not g__14155(w__11121 ,w__11292);
  not g__14156(w__11120 ,w__11119);
  not g__14157(w__11119 ,w__11685);
  not g__14158(w__11118 ,w__11116);
  not g__14159(w__11117 ,w__11116);
  not g__14160(w__11116 ,w__11293);
  not g__14161(w__11115 ,w__11113);
  not g__14162(w__11114 ,w__11113);
  not g__14163(w__11113 ,w__11382);
  not g__14164(w__11112 ,w__11282);
  not g__14165(w__11282 ,w__11471);
  not g__14166(w__11111 ,w__11274);
  not g__14167(w__11274 ,w__11374);
  not g__14168(w__11110 ,w__11273);
  not g__14169(w__11273 ,w__11374);
  not g__14170(w__11109 ,w__11272);
  not g__14171(w__11272 ,w__11371);
  not g__14172(w__11108 ,w__11280);
  not g__14173(w__11280 ,w__11468);
  not g__14174(w__11107 ,w__11283);
  not g__14175(w__11283 ,w__11471);
  not g__14176(w__11106 ,w__11281);
  not g__14177(w__11281 ,w__11468);
  not g__14178(w__11105 ,w__11279);
  not g__14179(w__11279 ,w__11384);
  not g__14180(w__11104 ,w__11278);
  not g__14181(w__11278 ,w__11384);
  not g__14182(w__11103 ,w__11271);
  not g__14183(w__11271 ,w__11371);
  not g__14184(w__11102 ,w__11275);
  not g__14185(w__11275 ,w__11377);
  not g__14186(w__11101 ,w__11277);
  not g__14187(w__11277 ,w__11382);
  not g__14188(w__11100 ,w__11276);
  not g__14189(w__11276 ,w__11377);
  not g__14190(w__11099 ,w__11098);
  not g__14191(w__11098 ,w__11838);
  not g__14192(w__11097 ,w__11096);
  not g__14193(w__11096 ,w__11915);
  not g__14194(w__11095 ,w__11094);
  not g__14195(w__11094 ,w__11840);
  not g__14196(w__11093 ,w__11092);
  not g__14197(w__11092 ,w__11836);
  not g__14198(w__10943 ,w__10952);
  not g__14199(w__11091 ,w__10952);
  not g__14200(w__10952 ,w__10944);
  not g__14201(w__11090 ,w__11258);
  not g__14202(w__11089 ,w__11087);
  not g__14203(w__11088 ,w__11087);
  not g__14204(w__11087 ,w__11684);
  not g__14205(w__11086 ,w__11084);
  not g__14206(w__11085 ,w__11084);
  not g__14207(w__11084 ,w__11685);
  not g__14208(w__11083 ,w__11081);
  not g__14209(w__11082 ,w__11081);
  not g__14210(w__11081 ,w__11591);
  not g__14211(w__11080 ,w__11078);
  not g__14212(w__11079 ,w__11078);
  not g__14213(w__11078 ,w__11588);
  not g__14214(w__11077 ,w__11075);
  not g__14215(w__11076 ,w__11075);
  not g__14216(w__11075 ,w__11292);
  not g__14217(w__11074 ,w__11072);
  not g__14218(w__11073 ,w__11072);
  not g__14219(w__11072 ,w__11590);
  not g__14220(w__11071 ,w__11069);
  not g__14221(w__11070 ,w__11069);
  not g__14222(w__11069 ,w__11589);
  not g__14223(w__11068 ,w__11066);
  not g__14224(w__11067 ,w__11066);
  not g__14225(w__11066 ,w__11587);
  not g__14226(w__11065 ,w__11063);
  not g__14227(w__11064 ,w__11063);
  not g__14228(w__11063 ,w__11586);
  not g__14229(w__11062 ,w__11060);
  not g__14230(w__11061 ,w__11060);
  not g__14231(w__11060 ,w__11684);
  not g__14232(w__11059 ,w__11057);
  not g__14233(w__11058 ,w__11057);
  not g__14234(w__11057 ,w__11136);
  not g__14235(w__11056 ,w__11054);
  not g__14236(w__11055 ,w__11054);
  not g__14237(w__11054 ,w__11126);
  not g__14238(w__11053 ,w__11051);
  not g__14239(w__11052 ,w__11051);
  not g__14240(w__11051 ,w__11128);
  not g__14241(w__11050 ,w__11048);
  not g__14242(w__11049 ,w__11048);
  not g__14243(w__11048 ,w__11124);
  not g__14244(w__11047 ,w__11045);
  not g__14245(w__11046 ,w__11045);
  not g__14246(w__11045 ,w__11122);
  not g__14247(w__11044 ,w__11042);
  not g__14248(w__11043 ,w__11042);
  not g__14249(w__11042 ,w__11118);
  not g__14250(w__11041 ,w__11039);
  not g__14251(w__11040 ,w__11039);
  not g__14252(w__11039 ,w__11589);
  not g__14253(w__11038 ,w__11036);
  not g__14254(w__11037 ,w__11036);
  not g__14255(w__11036 ,w__11136);
  not g__14256(w__11035 ,w__11033);
  not g__14257(w__11034 ,w__11033);
  not g__14258(w__11033 ,w__11293);
  not g__14259(w__11032 ,w__11030);
  not g__14260(w__11031 ,w__11030);
  not g__14261(w__11030 ,w__11293);
  not g__14262(w__11029 ,w__11027);
  not g__14263(w__11028 ,w__11027);
  not g__14264(w__11027 ,w__11134);
  not g__14265(w__11026 ,w__11024);
  not g__14266(w__11025 ,w__11024);
  not g__14267(w__11024 ,w__11132);
  not g__14268(w__11023 ,w__11021);
  not g__14269(w__11022 ,w__11021);
  not g__14270(w__11021 ,w__11130);
  not g__14271(w__11020 ,w__11018);
  not g__14272(w__11019 ,w__11018);
  not g__14273(w__11018 ,w__11685);
  not g__14274(w__11017 ,w__11015);
  not g__14275(w__11016 ,w__11015);
  not g__14276(w__11015 ,w__11120);
  not g__14277(w__11014 ,w__11012);
  not g__14278(w__11013 ,w__11012);
  not g__14279(w__11012 ,w__11120);
  not g__14280(w__11011 ,w__11009);
  not g__14281(w__11010 ,w__11009);
  not g__14282(w__11009 ,w__11588);
  not g__14283(w__11008 ,w__11006);
  not g__14284(w__11007 ,w__11006);
  not g__14285(w__11006 ,w__11128);
  not g__14286(w__11005 ,w__11003);
  not g__14287(w__11004 ,w__11003);
  not g__14288(w__11003 ,w__11587);
  not g__14289(w__11002 ,w__11000);
  not g__14290(w__11001 ,w__11000);
  not g__14291(w__11000 ,w__11124);
  not g__14292(w__10999 ,w__10997);
  not g__14293(w__10998 ,w__10997);
  not g__14294(w__10997 ,w__11122);
  not g__14295(w__10996 ,w__10994);
  not g__14296(w__10995 ,w__10994);
  not g__14297(w__10994 ,w__11586);
  not g__14298(w__10993 ,w__10991);
  not g__14299(w__10992 ,w__10991);
  not g__14300(w__10991 ,w__11590);
  not g__14301(w__10990 ,w__10988);
  not g__14302(w__10989 ,w__10988);
  not g__14303(w__10988 ,w__11126);
  not g__14304(w__10987 ,w__10985);
  not g__14305(w__10986 ,w__10985);
  not g__14306(w__10985 ,w__11130);
  not g__14307(w__10984 ,w__10982);
  not g__14308(w__10983 ,w__10982);
  not g__14309(w__10982 ,w__11134);
  not g__14310(w__10981 ,w__10979);
  not g__14311(w__10980 ,w__10979);
  not g__14312(w__10979 ,w__11591);
  not g__14313(w__10978 ,w__10976);
  not g__14314(w__10977 ,w__10976);
  not g__14315(w__10976 ,w__11132);
  not g__14316(w__10975 ,w__10973);
  not g__14317(w__10974 ,w__10973);
  not g__14318(w__10973 ,w__11292);
  not g__14319(w__10972 ,w__10971);
  not g__14320(w__10971 ,w__11117);
  not g__14321(w__10970 ,w__10969);
  not g__14322(w__10969 ,w__11088);
  not g__14323(w__10968 ,w__10967);
  not g__14324(w__10967 ,w__11065);
  not g__14325(w__10966 ,w__10965);
  not g__14326(w__10965 ,w__11068);
  not g__14327(w__10964 ,w__10963);
  not g__14328(w__10963 ,w__11071);
  not g__14329(w__10962 ,w__10961);
  not g__14330(w__10961 ,w__11074);
  not g__14331(w__10960 ,w__10959);
  not g__14332(w__10959 ,w__11077);
  not g__14333(w__10958 ,w__10957);
  not g__14334(w__10957 ,w__11080);
  not g__14335(w__10956 ,w__10955);
  not g__14336(w__10955 ,w__11083);
  not g__14337(w__10954 ,w__10953);
  not g__14338(w__10953 ,w__11086);
  xor g__14339(w__10951 ,w__12533 ,w__12628);
  xor g__14340(w__13036 ,w__12509 ,w__12598);
  xor g__14341(w__10950 ,w__12491 ,w__12512);
  xor g__14342(w__10949 ,w__12150 ,w__12228);
  xor g__14343(w__10948 ,w__12144 ,w__11098);
  xor g__14344(w__10947 ,w__12254 ,w__11096);
  xor g__14345(w__10946 ,w__12133 ,w__11094);
  xor g__14346(w__10945 ,w__12241 ,w__11092);
  not g__14347(w__11459 ,in25[1]);
  not g__14348(w__9750 ,in21[1]);
  not g__14349(w__8041 ,in17[1]);
  not g__14350(w__6332 ,in13[1]);
  buf g__14351(w__6238 ,in12[0]);
  not g__14352(w__2914 ,in2[1]);
  not g__14353(w__4623 ,in9[1]);
  buf g__14354(w__11709 ,in25[1]);
  buf g__14355(w__10000 ,in21[1]);
  buf g__14356(w__8291 ,in17[1]);
  buf g__14357(w__4873 ,in9[1]);
  buf g__14358(w__865 ,in5[0]);
  buf g__14359(w__11851 ,w__11709);
  buf g__14360(w__10142 ,w__10000);
  buf g__14361(w__8433 ,w__8291);
  buf g__14362(w__5015 ,w__4873);
  buf g__14363(w__225 ,w__12746);
  not g__14364(w__1147 ,w__12809);
  not g__14365(w__364 ,w__12746);
  not g__14366(w__1499 ,w__1201);
  buf g__14367(w__714 ,w__519);
  buf g__14368(w__1371 ,w__1208);
  buf g__14369(w__1326 ,w__12778);
  not g__14370(w__1459 ,w__787);
  buf g__14371(w__1575 ,w__1069);
endmodule
