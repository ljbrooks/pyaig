module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, out1, out2, out3, out4, out5, out6);
  input [10:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12;
  output out1, out2, out3, out4, out5, out6;
  wire [10:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12;
  wire out1, out2, out3, out4, out5, out6;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__139, w__140, w__141, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__157, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__171, w__172, w__173, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__665, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__680;
  wire w__681, w__682, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__697, w__698, w__699, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__714, w__715, w__716, w__717, w__718, w__719, w__720;
  wire w__721, w__722, w__723, w__724, w__725, w__726, w__727, w__728;
  wire w__729, w__730, w__731, w__732, w__733, w__734, w__735, w__736;
  wire w__737, w__738, w__739, w__740, w__741, w__742, w__743, w__744;
  wire w__745, w__746, w__747, w__748, w__749, w__750, w__751, w__752;
  wire w__753, w__754, w__755, w__756, w__757, w__758, w__759, w__760;
  wire w__761, w__762, w__763, w__764, w__765, w__766, w__767, w__768;
  wire w__769, w__770, w__771, w__772, w__773, w__774, w__775, w__776;
  wire w__777, w__778, w__779, w__780, w__781, w__782, w__783, w__784;
  wire w__785, w__786, w__787, w__788, w__789, w__790, w__791, w__792;
  wire w__793, w__794, w__795, w__796, w__797, w__798, w__799, w__800;
  wire w__801, w__802, w__803, w__804, w__805, w__806, w__807, w__808;
  wire w__809, w__810, w__811, w__812, w__813, w__814, w__815, w__816;
  wire w__817, w__818, w__819, w__820, w__821, w__822, w__823, w__824;
  wire w__825, w__826, w__827, w__828, w__829, w__830, w__831, w__832;
  wire w__833, w__834, w__835, w__836, w__837, w__838, w__839, w__840;
  wire w__841, w__842, w__843, w__844, w__845, w__846, w__847, w__848;
  wire w__849, w__850, w__851, w__852, w__853, w__854, w__855, w__856;
  wire w__857, w__858, w__859, w__860, w__861, w__862, w__863, w__864;
  wire w__865, w__866, w__867, w__868, w__869, w__870, w__871, w__872;
  wire w__873, w__874, w__875, w__876, w__877, w__878, w__879, w__880;
  wire w__881, w__882, w__883, w__884, w__885, w__886, w__887, w__888;
  wire w__889, w__890, w__891, w__892, w__893, w__894, w__895, w__896;
  wire w__897, w__898, w__899, w__900, w__901, w__902, w__903, w__904;
  wire w__905, w__906, w__907, w__908, w__909, w__910, w__911, w__912;
  wire w__913, w__914, w__915, w__916, w__917, w__918, w__919, w__920;
  wire w__921, w__922, w__923, w__924, w__925, w__926, w__927, w__928;
  wire w__929, w__930, w__931, w__932, w__933, w__934, w__935, w__936;
  wire w__937, w__938, w__939, w__940, w__941, w__942, w__943, w__944;
  wire w__945, w__946, w__947, w__948, w__949, w__950, w__951, w__952;
  wire w__953, w__954, w__955, w__956, w__957, w__958, w__959, w__960;
  wire w__961, w__962, w__963, w__964, w__965, w__966, w__967, w__968;
  wire w__969, w__970, w__971, w__972, w__973, w__974, w__975, w__976;
  wire w__977, w__978, w__979, w__980, w__981, w__982, w__983, w__984;
  wire w__985, w__986, w__987, w__988, w__989, w__990, w__991, w__992;
  wire w__993, w__994, w__995, w__996, w__997, w__998, w__999, w__1000;
  wire w__1001, w__1002, w__1003, w__1004, w__1005, w__1006, w__1007, w__1008;
  wire w__1009, w__1010, w__1011, w__1012, w__1013, w__1014, w__1015, w__1016;
  wire w__1017, w__1018, w__1019, w__1020, w__1021, w__1022, w__1023, w__1024;
  wire w__1025, w__1026, w__1027, w__1028, w__1029, w__1030, w__1031, w__1032;
  wire w__1033, w__1034, w__1035, w__1036, w__1037, w__1038, w__1039, w__1040;
  wire w__1041, w__1042, w__1043, w__1044, w__1045, w__1046, w__1047, w__1048;
  wire w__1049, w__1050, w__1051, w__1052, w__1053, w__1054, w__1055, w__1056;
  wire w__1057, w__1058, w__1059, w__1060, w__1061, w__1062, w__1063, w__1064;
  wire w__1065, w__1066, w__1067, w__1068, w__1069, w__1070, w__1071, w__1072;
  wire w__1073, w__1074, w__1075, w__1076, w__1077, w__1078, w__1079, w__1080;
  wire w__1081, w__1082, w__1083, w__1084, w__1085, w__1086, w__1087, w__1088;
  wire w__1089, w__1090, w__1091, w__1092, w__1093, w__1094, w__1095, w__1096;
  wire w__1097, w__1098, w__1099, w__1100, w__1101, w__1102, w__1103, w__1104;
  wire w__1105, w__1106, w__1107, w__1108, w__1109, w__1110, w__1111, w__1112;
  wire w__1113, w__1114, w__1115, w__1116, w__1117, w__1118, w__1119, w__1120;
  wire w__1121, w__1122, w__1123, w__1124, w__1125, w__1126, w__1127, w__1128;
  wire w__1129, w__1130, w__1131, w__1132, w__1133, w__1134, w__1135, w__1136;
  wire w__1137, w__1138, w__1139, w__1140, w__1141, w__1142, w__1143, w__1144;
  wire w__1145, w__1146, w__1147, w__1148, w__1149, w__1150, w__1151, w__1152;
  wire w__1153, w__1154, w__1155, w__1156, w__1157, w__1158, w__1159, w__1160;
  wire w__1161, w__1162, w__1163, w__1164, w__1165, w__1166, w__1167, w__1168;
  wire w__1169, w__1170, w__1171, w__1172, w__1173, w__1174, w__1175, w__1176;
  wire w__1177, w__1178, w__1179, w__1180, w__1181, w__1182, w__1183, w__1184;
  wire w__1185, w__1186, w__1187, w__1188, w__1189, w__1190, w__1191, w__1192;
  wire w__1193, w__1194, w__1195, w__1196, w__1197, w__1198, w__1199, w__1200;
  wire w__1201, w__1202, w__1203, w__1204, w__1205, w__1206, w__1207, w__1208;
  wire w__1209, w__1210, w__1211, w__1212, w__1213, w__1214, w__1215, w__1216;
  wire w__1217, w__1218, w__1219, w__1220, w__1221, w__1222, w__1223, w__1224;
  wire w__1225, w__1226, w__1227, w__1228, w__1229, w__1230, w__1231, w__1232;
  wire w__1233, w__1234, w__1235, w__1236, w__1237, w__1238, w__1239, w__1240;
  wire w__1241, w__1242, w__1243, w__1244, w__1245, w__1246, w__1247, w__1248;
  wire w__1249, w__1250, w__1251, w__1252, w__1253, w__1254, w__1255, w__1256;
  wire w__1257, w__1258, w__1259, w__1260, w__1261, w__1262, w__1263, w__1264;
  wire w__1265, w__1266, w__1267, w__1268, w__1269, w__1270, w__1271, w__1272;
  wire w__1273, w__1274, w__1275, w__1276, w__1277, w__1278, w__1279, w__1280;
  wire w__1281, w__1282, w__1283, w__1284, w__1285, w__1286, w__1287, w__1288;
  wire w__1289, w__1290, w__1291, w__1292, w__1293, w__1294, w__1295, w__1296;
  wire w__1297, w__1298, w__1299, w__1300, w__1301, w__1302, w__1303, w__1304;
  wire w__1305, w__1306, w__1307, w__1308, w__1309, w__1310, w__1311, w__1312;
  wire w__1313, w__1314, w__1315, w__1316, w__1317, w__1318, w__1319, w__1320;
  wire w__1321, w__1322, w__1323, w__1324, w__1325, w__1326, w__1327, w__1328;
  wire w__1329, w__1330, w__1331, w__1332, w__1333, w__1334, w__1335, w__1336;
  wire w__1337, w__1338, w__1339, w__1340, w__1341, w__1342, w__1343, w__1344;
  wire w__1345, w__1346, w__1347, w__1348, w__1349, w__1350, w__1351, w__1352;
  wire w__1353, w__1354, w__1355, w__1356, w__1357, w__1358, w__1359, w__1360;
  wire w__1361, w__1362, w__1363, w__1364, w__1365, w__1366, w__1367, w__1368;
  wire w__1369, w__1370, w__1371, w__1372, w__1373, w__1374, w__1375, w__1376;
  wire w__1377, w__1378, w__1379, w__1380, w__1381, w__1382, w__1383, w__1384;
  wire w__1385, w__1386, w__1387, w__1388, w__1389, w__1390, w__1391, w__1392;
  wire w__1393, w__1394, w__1395, w__1396, w__1397, w__1398, w__1399, w__1400;
  wire w__1401, w__1402, w__1403, w__1404, w__1405, w__1406, w__1407, w__1408;
  wire w__1409, w__1410, w__1411, w__1412, w__1413, w__1414, w__1415, w__1416;
  wire w__1417, w__1418, w__1419, w__1420, w__1421, w__1422, w__1423, w__1424;
  wire w__1425, w__1426, w__1427, w__1428, w__1429, w__1430, w__1431, w__1432;
  wire w__1433, w__1434, w__1435, w__1436, w__1437, w__1438, w__1439, w__1440;
  wire w__1441, w__1442, w__1443, w__1444, w__1445, w__1446, w__1447, w__1448;
  wire w__1449, w__1450, w__1451, w__1452, w__1453, w__1454, w__1455, w__1456;
  wire w__1457, w__1458, w__1459, w__1460, w__1461, w__1462, w__1463, w__1464;
  wire w__1465, w__1466, w__1467, w__1468, w__1469, w__1470, w__1471, w__1472;
  wire w__1473, w__1474, w__1475, w__1476, w__1477, w__1478, w__1479, w__1480;
  wire w__1481, w__1482, w__1483, w__1484, w__1485, w__1486, w__1487, w__1488;
  wire w__1489, w__1490, w__1491, w__1492, w__1493, w__1494, w__1495, w__1496;
  wire w__1497, w__1498, w__1499, w__1500, w__1501, w__1502, w__1503, w__1504;
  wire w__1505, w__1506, w__1507, w__1508, w__1509, w__1510, w__1511, w__1512;
  wire w__1513, w__1514, w__1515, w__1516, w__1517, w__1518, w__1519, w__1520;
  wire w__1521, w__1522, w__1523, w__1524, w__1525, w__1526, w__1527, w__1528;
  wire w__1529, w__1530, w__1531, w__1532, w__1533, w__1534, w__1535, w__1536;
  wire w__1537, w__1538, w__1539, w__1540, w__1541, w__1542, w__1543, w__1544;
  wire w__1545, w__1546, w__1547, w__1548, w__1549, w__1550, w__1551, w__1552;
  wire w__1553, w__1554, w__1555, w__1556, w__1557, w__1558, w__1559, w__1560;
  wire w__1561, w__1562, w__1563, w__1564, w__1565, w__1566, w__1567, w__1568;
  wire w__1569, w__1570, w__1571, w__1572, w__1573, w__1574, w__1575, w__1576;
  wire w__1577, w__1578, w__1579, w__1580, w__1581, w__1582, w__1583, w__1584;
  wire w__1585, w__1586, w__1587, w__1588, w__1589, w__1590, w__1591, w__1592;
  wire w__1593, w__1594, w__1595, w__1596, w__1597, w__1598, w__1599, w__1600;
  wire w__1601, w__1602, w__1603, w__1604, w__1605, w__1606, w__1607, w__1608;
  wire w__1609, w__1610, w__1611, w__1612, w__1613, w__1614, w__1615, w__1616;
  wire w__1617, w__1618, w__1619, w__1620, w__1621, w__1622, w__1623, w__1624;
  wire w__1625, w__1626, w__1627, w__1628, w__1629, w__1630, w__1631, w__1632;
  wire w__1633, w__1634, w__1635, w__1636, w__1637, w__1638, w__1639, w__1640;
  wire w__1641, w__1642, w__1643, w__1644, w__1645, w__1646, w__1647, w__1648;
  wire w__1649, w__1650, w__1651, w__1652, w__1653, w__1654, w__1655, w__1656;
  wire w__1657, w__1658, w__1659, w__1660, w__1661, w__1662, w__1663, w__1664;
  wire w__1665, w__1666, w__1667, w__1668, w__1669, w__1670, w__1671, w__1672;
  wire w__1673, w__1674, w__1675, w__1676, w__1677, w__1678, w__1679, w__1680;
  wire w__1681, w__1682, w__1683, w__1684, w__1685, w__1686, w__1687, w__1688;
  wire w__1689, w__1690, w__1691, w__1692, w__1693, w__1694, w__1695, w__1696;
  wire w__1697, w__1698, w__1699, w__1700, w__1701, w__1702, w__1703, w__1704;
  wire w__1705, w__1706, w__1707, w__1708, w__1709, w__1710, w__1711, w__1712;
  wire w__1713, w__1714, w__1715, w__1716, w__1717, w__1718, w__1719, w__1720;
  wire w__1721, w__1722, w__1723, w__1724, w__1725, w__1726, w__1727, w__1728;
  wire w__1729, w__1730, w__1731, w__1732, w__1733, w__1734, w__1735, w__1736;
  wire w__1737, w__1738, w__1739, w__1740, w__1741, w__1742, w__1743, w__1744;
  wire w__1745, w__1746, w__1747, w__1748, w__1749, w__1750, w__1751, w__1752;
  wire w__1753, w__1754, w__1755, w__1756, w__1757, w__1758, w__1759, w__1760;
  wire w__1761, w__1762, w__1763, w__1764, w__1765, w__1766, w__1767, w__1768;
  wire w__1769, w__1770, w__1771, w__1772, w__1773, w__1774, w__1775, w__1776;
  wire w__1777, w__1778, w__1779, w__1780, w__1781, w__1782, w__1783, w__1784;
  wire w__1785, w__1786, w__1787, w__1788, w__1789, w__1790, w__1791, w__1792;
  wire w__1793, w__1794, w__1795, w__1796, w__1797, w__1798, w__1799, w__1800;
  wire w__1801, w__1802, w__1803, w__1804, w__1805, w__1806, w__1807, w__1808;
  wire w__1809, w__1810, w__1811, w__1812, w__1813, w__1814, w__1815, w__1816;
  wire w__1817, w__1818, w__1819, w__1820, w__1821, w__1822, w__1823, w__1824;
  wire w__1825, w__1826, w__1827, w__1828, w__1829, w__1830, w__1831, w__1832;
  wire w__1833, w__1834, w__1835, w__1836, w__1837, w__1838, w__1839, w__1840;
  wire w__1841, w__1842, w__1843, w__1844, w__1845, w__1846, w__1847, w__1848;
  wire w__1849, w__1850, w__1851, w__1852, w__1853, w__1854, w__1855, w__1856;
  wire w__1857, w__1858, w__1859, w__1860, w__1861, w__1862, w__1863, w__1864;
  wire w__1865, w__1866, w__1867, w__1868, w__1869, w__1870, w__1871, w__1872;
  wire w__1873, w__1874, w__1875, w__1876, w__1877, w__1878, w__1879, w__1880;
  wire w__1881, w__1882, w__1883, w__1884, w__1885, w__1886, w__1887, w__1888;
  wire w__1889, w__1890, w__1891, w__1892, w__1893, w__1894, w__1895, w__1896;
  wire w__1897, w__1898, w__1899, w__1900, w__1901, w__1902, w__1903, w__1904;
  wire w__1905, w__1906, w__1907, w__1908, w__1909, w__1910, w__1911, w__1912;
  wire w__1913, w__1914, w__1915, w__1916, w__1917, w__1918, w__1919, w__1920;
  wire w__1921, w__1922, w__1923, w__1924, w__1925, w__1926, w__1927, w__1928;
  wire w__1929, w__1930, w__1931, w__1932, w__1933, w__1934, w__1935, w__1936;
  wire w__1937, w__1938, w__1939, w__1940, w__1941, w__1942, w__1943, w__1944;
  wire w__1945, w__1946, w__1947, w__1948, w__1949, w__1950, w__1951, w__1952;
  wire w__1953, w__1954, w__1955, w__1956, w__1957, w__1958, w__1959, w__1960;
  wire w__1961, w__1962, w__1963, w__1964, w__1965, w__1966, w__1967, w__1968;
  wire w__1969, w__1970, w__1971, w__1972, w__1973, w__1974, w__1975, w__1976;
  wire w__1977, w__1978, w__1979, w__1980, w__1981, w__1982, w__1983, w__1984;
  wire w__1985, w__1986, w__1987, w__1988, w__1989, w__1990, w__1991, w__1992;
  wire w__1993, w__1994, w__1995, w__1996, w__1997, w__1998, w__1999, w__2000;
  wire w__2001, w__2002, w__2003, w__2004, w__2005, w__2006, w__2007, w__2008;
  wire w__2009, w__2010, w__2011, w__2012, w__2013, w__2014, w__2015, w__2016;
  wire w__2017, w__2018, w__2019, w__2020, w__2021, w__2022, w__2023, w__2024;
  wire w__2025, w__2026, w__2027, w__2028, w__2029, w__2030, w__2031, w__2032;
  wire w__2033, w__2034, w__2035, w__2036, w__2037, w__2038, w__2039, w__2040;
  wire w__2041, w__2042, w__2043, w__2044, w__2045, w__2046, w__2047, w__2048;
  wire w__2049, w__2050, w__2051, w__2052, w__2053, w__2054, w__2055, w__2056;
  wire w__2057, w__2058, w__2059, w__2060, w__2061, w__2062, w__2063, w__2064;
  wire w__2065, w__2066, w__2067, w__2068, w__2069, w__2070, w__2071, w__2072;
  wire w__2073, w__2074, w__2075, w__2076, w__2077, w__2078, w__2079, w__2080;
  wire w__2081, w__2082, w__2083, w__2084, w__2085, w__2086, w__2087, w__2088;
  wire w__2089, w__2090, w__2091, w__2092, w__2093, w__2094, w__2095, w__2096;
  wire w__2097, w__2098, w__2099, w__2100, w__2101, w__2102, w__2103, w__2104;
  wire w__2105, w__2106, w__2107, w__2108, w__2109, w__2110, w__2111, w__2112;
  wire w__2113, w__2114, w__2115, w__2116, w__2117, w__2118, w__2119, w__2120;
  wire w__2121, w__2122, w__2123, w__2124, w__2125, w__2126, w__2127, w__2128;
  wire w__2129, w__2130, w__2131, w__2132, w__2133, w__2134, w__2135, w__2136;
  wire w__2137, w__2138, w__2139, w__2140, w__2141, w__2142, w__2143, w__2144;
  wire w__2145, w__2146, w__2147, w__2148, w__2149, w__2150, w__2151, w__2152;
  wire w__2153, w__2154, w__2155, w__2156, w__2157, w__2158, w__2159, w__2160;
  wire w__2161, w__2162, w__2163, w__2164, w__2165, w__2166, w__2167, w__2168;
  wire w__2169, w__2170, w__2171, w__2172, w__2173, w__2174, w__2175, w__2176;
  wire w__2177, w__2178, w__2179, w__2180, w__2181, w__2182, w__2183, w__2184;
  wire w__2185, w__2186, w__2187, w__2188, w__2189, w__2190, w__2191, w__2192;
  wire w__2193, w__2194, w__2195, w__2196, w__2197, w__2198, w__2199, w__2200;
  wire w__2201, w__2202, w__2203, w__2204, w__2205, w__2206, w__2207, w__2208;
  wire w__2209, w__2210, w__2211, w__2212, w__2213, w__2214, w__2215, w__2216;
  wire w__2217, w__2218, w__2219, w__2220, w__2221, w__2222, w__2223, w__2224;
  wire w__2225, w__2226, w__2227, w__2228, w__2229, w__2230, w__2231, w__2232;
  wire w__2233, w__2234, w__2235, w__2236, w__2237, w__2238, w__2239, w__2240;
  wire w__2241, w__2242, w__2243, w__2244, w__2245, w__2246, w__2247, w__2248;
  wire w__2249, w__2250, w__2251, w__2252, w__2253, w__2254, w__2255, w__2256;
  wire w__2257, w__2258, w__2259, w__2260, w__2261, w__2262, w__2263, w__2264;
  wire w__2265, w__2266, w__2267, w__2268, w__2269, w__2270, w__2271, w__2272;
  wire w__2273, w__2274, w__2275, w__2276, w__2277, w__2278, w__2279, w__2280;
  wire w__2281, w__2282, w__2283, w__2284, w__2285, w__2286, w__2287, w__2288;
  wire w__2289, w__2290, w__2291, w__2292, w__2293, w__2294, w__2295, w__2296;
  wire w__2297, w__2298, w__2299, w__2300, w__2301, w__2302, w__2303, w__2304;
  wire w__2305, w__2306, w__2307, w__2308, w__2309, w__2310, w__2311, w__2312;
  wire w__2313, w__2314, w__2315, w__2316, w__2317, w__2318, w__2319, w__2320;
  wire w__2321, w__2322, w__2323, w__2324, w__2325, w__2326, w__2327, w__2328;
  wire w__2329, w__2330, w__2331, w__2332, w__2333, w__2334, w__2335, w__2336;
  wire w__2337, w__2338, w__2339, w__2340, w__2341, w__2342, w__2343, w__2344;
  wire w__2345, w__2346, w__2347, w__2348, w__2349, w__2350, w__2351, w__2352;
  wire w__2353, w__2354, w__2355, w__2356, w__2357, w__2358, w__2359, w__2360;
  wire w__2361, w__2362, w__2363, w__2364, w__2365, w__2366, w__2367, w__2368;
  wire w__2369, w__2370, w__2371, w__2372, w__2373, w__2374, w__2375, w__2376;
  wire w__2377, w__2378, w__2379, w__2380, w__2381, w__2382, w__2383, w__2384;
  wire w__2385, w__2386, w__2387, w__2388, w__2389, w__2390, w__2391, w__2392;
  wire w__2393, w__2394, w__2395, w__2396, w__2397, w__2398, w__2399, w__2400;
  wire w__2401, w__2402, w__2403, w__2404, w__2405, w__2406, w__2407, w__2408;
  wire w__2409, w__2410, w__2411, w__2412, w__2413, w__2414, w__2415, w__2416;
  wire w__2417, w__2418, w__2419, w__2420, w__2421, w__2422, w__2423, w__2424;
  wire w__2425, w__2426, w__2427, w__2428, w__2429, w__2430, w__2431, w__2432;
  wire w__2433, w__2434, w__2435, w__2436, w__2437, w__2438, w__2439, w__2440;
  wire w__2441, w__2442, w__2443, w__2444, w__2445, w__2446, w__2447, w__2448;
  wire w__2449, w__2450, w__2451, w__2452, w__2453, w__2454, w__2455, w__2456;
  wire w__2457, w__2458, w__2459, w__2460, w__2461, w__2462, w__2463, w__2464;
  wire w__2465, w__2466, w__2467, w__2468, w__2469, w__2470, w__2471, w__2472;
  wire w__2473, w__2474, w__2475, w__2476, w__2477, w__2478, w__2479, w__2480;
  wire w__2481, w__2482, w__2483, w__2484, w__2485, w__2486, w__2487, w__2488;
  wire w__2489, w__2490, w__2491, w__2492, w__2493, w__2494, w__2495, w__2496;
  wire w__2497, w__2498, w__2499, w__2500, w__2501, w__2502, w__2503, w__2504;
  wire w__2505, w__2506, w__2507, w__2508, w__2509, w__2510, w__2511, w__2512;
  wire w__2513, w__2514, w__2515, w__2516, w__2517, w__2518, w__2519, w__2520;
  wire w__2521, w__2522, w__2523, w__2524, w__2525, w__2526, w__2527, w__2528;
  wire w__2529, w__2530, w__2531, w__2532, w__2533, w__2534, w__2535, w__2536;
  wire w__2537, w__2538, w__2539, w__2540, w__2541, w__2542, w__2543, w__2544;
  wire w__2545, w__2546, w__2547, w__2548, w__2549, w__2550, w__2551, w__2552;
  wire w__2553, w__2554, w__2555, w__2556, w__2557, w__2558, w__2559, w__2560;
  wire w__2561, w__2562, w__2563, w__2564, w__2565, w__2566, w__2567, w__2568;
  wire w__2569, w__2570, w__2571, w__2572, w__2573, w__2574, w__2575, w__2576;
  wire w__2577, w__2578, w__2579, w__2580, w__2581, w__2582, w__2583, w__2584;
  wire w__2585, w__2586, w__2587, w__2588, w__2589, w__2590, w__2591, w__2592;
  wire w__2593, w__2594, w__2595, w__2596, w__2597, w__2598, w__2599, w__2600;
  wire w__2601, w__2602, w__2603, w__2604, w__2605, w__2606, w__2607, w__2608;
  wire w__2609, w__2610, w__2611, w__2612, w__2613, w__2614, w__2615, w__2616;
  wire w__2617, w__2618, w__2619, w__2620, w__2621, w__2622, w__2623, w__2624;
  wire w__2625, w__2626, w__2627, w__2628, w__2629, w__2630, w__2631, w__2632;
  wire w__2633, w__2634, w__2635, w__2636, w__2637, w__2638, w__2639, w__2640;
  wire w__2641, w__2642, w__2643, w__2644, w__2645, w__2646, w__2647, w__2648;
  wire w__2649, w__2650, w__2651, w__2652, w__2653, w__2654, w__2655, w__2656;
  wire w__2657, w__2658, w__2659, w__2660, w__2661, w__2662, w__2663, w__2664;
  wire w__2665, w__2666, w__2667, w__2668, w__2669, w__2670, w__2671, w__2672;
  wire w__2673, w__2674, w__2675, w__2676, w__2677, w__2678, w__2679, w__2680;
  wire w__2681, w__2682, w__2683, w__2684, w__2685, w__2686, w__2687, w__2688;
  wire w__2689, w__2690, w__2691, w__2692, w__2693, w__2694, w__2695, w__2696;
  wire w__2697, w__2698, w__2699, w__2700, w__2701, w__2702, w__2703, w__2704;
  wire w__2705, w__2706, w__2707, w__2708, w__2709, w__2710, w__2711, w__2712;
  wire w__2713, w__2714, w__2715, w__2716, w__2717, w__2718, w__2719, w__2720;
  wire w__2721, w__2722, w__2723, w__2724, w__2725, w__2726, w__2727, w__2728;
  wire w__2729, w__2730, w__2731, w__2732, w__2733, w__2734, w__2735, w__2736;
  wire w__2737, w__2738, w__2739, w__2740, w__2741, w__2742, w__2743, w__2744;
  wire w__2745, w__2746, w__2747, w__2748, w__2749, w__2750, w__2751, w__2752;
  wire w__2753, w__2754, w__2755, w__2756, w__2757, w__2758, w__2759, w__2760;
  wire w__2761, w__2762, w__2763, w__2764, w__2765, w__2766, w__2767, w__2768;
  wire w__2769, w__2770, w__2771, w__2772, w__2773, w__2774, w__2775, w__2776;
  wire w__2777, w__2778, w__2779, w__2780, w__2781, w__2782, w__2783, w__2784;
  wire w__2785, w__2786, w__2787, w__2788, w__2789, w__2790, w__2791, w__2792;
  wire w__2793, w__2794, w__2795, w__2796, w__2797, w__2798, w__2799, w__2800;
  wire w__2801, w__2802, w__2803, w__2804, w__2805, w__2806, w__2807, w__2808;
  wire w__2809, w__2810, w__2811, w__2812, w__2813, w__2814, w__2815, w__2816;
  wire w__2817, w__2818, w__2819, w__2820, w__2821, w__2822, w__2823, w__2824;
  wire w__2825, w__2826, w__2827, w__2828, w__2829, w__2830, w__2831, w__2832;
  wire w__2833, w__2834, w__2835, w__2836, w__2837, w__2838, w__2839, w__2840;
  wire w__2841, w__2842, w__2843, w__2844, w__2845, w__2846, w__2847, w__2848;
  wire w__2849, w__2850, w__2851, w__2852, w__2853, w__2854, w__2855, w__2856;
  wire w__2857, w__2858, w__2859, w__2860, w__2861, w__2862, w__2863, w__2864;
  wire w__2865, w__2866, w__2867, w__2868, w__2869, w__2870, w__2871, w__2872;
  wire w__2873, w__2874, w__2875, w__2876, w__2877, w__2878, w__2879, w__2880;
  wire w__2881, w__2882, w__2883, w__2884, w__2885, w__2886, w__2887, w__2888;
  wire w__2889, w__2890, w__2891, w__2892, w__2893, w__2894, w__2895, w__2896;
  wire w__2897, w__2898, w__2899, w__2900, w__2901, w__2902, w__2903, w__2904;
  wire w__2905, w__2906, w__2907, w__2908, w__2909, w__2910, w__2911, w__2912;
  wire w__2913, w__2914, w__2915, w__2916, w__2917, w__2918, w__2919, w__2920;
  wire w__2921, w__2922, w__2923, w__2924, w__2925, w__2926, w__2927, w__2928;
  wire w__2929, w__2930, w__2931, w__2932, w__2933, w__2934, w__2935, w__2936;
  wire w__2937, w__2938, w__2939, w__2940, w__2941, w__2942, w__2943, w__2944;
  wire w__2945, w__2946, w__2947, w__2948, w__2949, w__2950, w__2951, w__2952;
  wire w__2953, w__2954, w__2955, w__2956, w__2957, w__2958, w__2959, w__2960;
  wire w__2961, w__2962, w__2963, w__2964, w__2965, w__2966, w__2967, w__2968;
  wire w__2969, w__2970, w__2971, w__2972, w__2973, w__2974, w__2975, w__2976;
  wire w__2977, w__2978, w__2979, w__2980, w__2981, w__2982, w__2983, w__2984;
  wire w__2985, w__2986, w__2987, w__2988, w__2989, w__2990, w__2991, w__2992;
  wire w__2993, w__2994, w__2995, w__2996, w__2997, w__2998, w__2999, w__3000;
  wire w__3001, w__3002, w__3003, w__3004, w__3005, w__3006, w__3007, w__3008;
  wire w__3009, w__3010, w__3011, w__3012, w__3013, w__3014, w__3015, w__3016;
  wire w__3017, w__3018, w__3019, w__3020, w__3021, w__3022, w__3023, w__3024;
  wire w__3025, w__3026, w__3027, w__3028, w__3029, w__3030, w__3031, w__3032;
  wire w__3033, w__3034, w__3035, w__3036, w__3037, w__3038, w__3039, w__3040;
  wire w__3041, w__3042, w__3043, w__3044, w__3045, w__3046, w__3047, w__3048;
  wire w__3049, w__3050, w__3051, w__3052, w__3053, w__3054, w__3055, w__3056;
  wire w__3057, w__3058, w__3059, w__3060, w__3061, w__3062, w__3063, w__3064;
  wire w__3065, w__3066, w__3067, w__3068, w__3069, w__3070, w__3071, w__3072;
  wire w__3073, w__3074, w__3075, w__3076, w__3077, w__3078, w__3079, w__3080;
  wire w__3081, w__3082, w__3083, w__3084, w__3085, w__3086, w__3087, w__3088;
  wire w__3089, w__3090, w__3091, w__3092, w__3093, w__3094, w__3095, w__3096;
  wire w__3097, w__3098, w__3099, w__3100, w__3101, w__3102, w__3103, w__3104;
  wire w__3105, w__3106, w__3107, w__3108, w__3109, w__3110, w__3111, w__3112;
  wire w__3113, w__3114, w__3115, w__3116, w__3117, w__3118, w__3119, w__3120;
  wire w__3121, w__3122, w__3123, w__3124, w__3125, w__3126, w__3127, w__3128;
  wire w__3129, w__3130, w__3131, w__3132, w__3133, w__3134, w__3135, w__3136;
  wire w__3137, w__3138, w__3139, w__3140, w__3141, w__3142, w__3143, w__3144;
  wire w__3145, w__3146, w__3147, w__3148, w__3149, w__3150, w__3151, w__3152;
  wire w__3153, w__3154, w__3155, w__3156, w__3157, w__3158, w__3159, w__3160;
  wire w__3161, w__3162, w__3163, w__3164, w__3165, w__3166, w__3167, w__3168;
  wire w__3169, w__3170, w__3171, w__3172, w__3173, w__3174, w__3175, w__3176;
  wire w__3177, w__3178, w__3179, w__3180, w__3181, w__3182, w__3183, w__3184;
  wire w__3185, w__3186, w__3187, w__3188, w__3189, w__3190, w__3191, w__3192;
  wire w__3193, w__3194, w__3195, w__3196, w__3197, w__3198, w__3199, w__3200;
  wire w__3201, w__3202, w__3203, w__3204, w__3205, w__3206, w__3207, w__3208;
  wire w__3209, w__3210, w__3211, w__3212, w__3213, w__3214, w__3215, w__3216;
  wire w__3217, w__3218, w__3219, w__3220, w__3221, w__3222, w__3223, w__3224;
  wire w__3225, w__3226, w__3227, w__3228, w__3229, w__3230, w__3231, w__3232;
  wire w__3233, w__3234, w__3235, w__3236, w__3237, w__3238, w__3239, w__3240;
  wire w__3241, w__3242, w__3243, w__3244, w__3245, w__3246, w__3247, w__3248;
  wire w__3249, w__3250, w__3251, w__3252, w__3253, w__3254, w__3255, w__3256;
  wire w__3257, w__3258, w__3259, w__3260, w__3261, w__3262, w__3263, w__3264;
  wire w__3265, w__3266, w__3267, w__3268, w__3269, w__3270, w__3271, w__3272;
  wire w__3273, w__3274, w__3275, w__3276, w__3277, w__3278, w__3279, w__3280;
  wire w__3281, w__3282, w__3283, w__3284, w__3285, w__3286, w__3287, w__3288;
  wire w__3289, w__3290, w__3291, w__3292, w__3293, w__3294, w__3295, w__3296;
  wire w__3297, w__3298, w__3299, w__3300, w__3301, w__3302, w__3303, w__3304;
  wire w__3305, w__3306, w__3307, w__3308, w__3309, w__3310, w__3311, w__3312;
  wire w__3313, w__3314, w__3315, w__3316, w__3317, w__3318, w__3319, w__3320;
  wire w__3321, w__3322, w__3323, w__3324, w__3325, w__3326, w__3327, w__3328;
  wire w__3329, w__3330, w__3331, w__3332, w__3333, w__3334, w__3335, w__3336;
  wire w__3337, w__3338, w__3339, w__3340, w__3341, w__3342, w__3343, w__3344;
  wire w__3345, w__3346, w__3347, w__3348, w__3349, w__3350, w__3351, w__3352;
  wire w__3353, w__3354, w__3355, w__3356, w__3357, w__3358, w__3359, w__3360;
  wire w__3361, w__3362, w__3363, w__3364, w__3365, w__3366, w__3367, w__3368;
  wire w__3369, w__3370, w__3371, w__3372, w__3373, w__3374, w__3375, w__3376;
  wire w__3377, w__3378, w__3379, w__3380, w__3381, w__3382, w__3383, w__3384;
  wire w__3385, w__3386, w__3387, w__3388, w__3389, w__3390, w__3391, w__3392;
  wire w__3393, w__3394, w__3395, w__3396, w__3397, w__3398, w__3399, w__3400;
  wire w__3401, w__3402, w__3403, w__3404, w__3405, w__3406, w__3407, w__3408;
  wire w__3409, w__3410, w__3411, w__3412, w__3413, w__3414, w__3415, w__3416;
  wire w__3417, w__3418, w__3419, w__3420, w__3421, w__3422, w__3423, w__3424;
  wire w__3425, w__3426, w__3427, w__3428, w__3429, w__3430, w__3431, w__3432;
  wire w__3433, w__3434, w__3435, w__3436, w__3437, w__3438, w__3439, w__3440;
  wire w__3441, w__3442, w__3443, w__3444, w__3445, w__3446, w__3447, w__3448;
  wire w__3449, w__3450, w__3451, w__3452, w__3453, w__3454, w__3455, w__3456;
  wire w__3457, w__3458, w__3459, w__3460, w__3461, w__3462, w__3463, w__3464;
  wire w__3465, w__3466, w__3467, w__3468, w__3469, w__3470, w__3471, w__3472;
  wire w__3473, w__3474, w__3475, w__3476, w__3477, w__3478, w__3479, w__3480;
  wire w__3481, w__3482, w__3483, w__3484, w__3485, w__3486, w__3487, w__3488;
  wire w__3489, w__3490, w__3491, w__3492, w__3493, w__3494, w__3495, w__3496;
  wire w__3497, w__3498, w__3499, w__3500, w__3501, w__3502, w__3503, w__3504;
  wire w__3505, w__3506, w__3507, w__3508, w__3509, w__3510, w__3511, w__3512;
  wire w__3513, w__3514, w__3515, w__3516, w__3517, w__3518, w__3519, w__3520;
  wire w__3521, w__3522, w__3523, w__3524, w__3525, w__3526, w__3527, w__3528;
  wire w__3529, w__3530, w__3531, w__3532, w__3533, w__3534, w__3535, w__3536;
  wire w__3537, w__3538, w__3539, w__3540, w__3541, w__3542, w__3543, w__3544;
  wire w__3545, w__3546, w__3547, w__3548, w__3549, w__3550, w__3551, w__3552;
  wire w__3553, w__3554, w__3555, w__3556, w__3557, w__3558, w__3559, w__3560;
  wire w__3561, w__3562, w__3563, w__3564, w__3565, w__3566, w__3567, w__3568;
  wire w__3569, w__3570, w__3571, w__3572, w__3573, w__3574, w__3575, w__3576;
  wire w__3577, w__3578, w__3579, w__3580, w__3581, w__3582, w__3583, w__3584;
  wire w__3585, w__3586, w__3587, w__3588, w__3589, w__3590, w__3591, w__3592;
  wire w__3593, w__3594, w__3595, w__3596, w__3597, w__3598, w__3599, w__3600;
  wire w__3601, w__3602, w__3603, w__3604, w__3605, w__3606, w__3607, w__3608;
  wire w__3609, w__3610, w__3611, w__3612, w__3613, w__3614, w__3615, w__3616;
  wire w__3617, w__3618, w__3619, w__3620, w__3621, w__3622, w__3623, w__3624;
  wire w__3625, w__3626, w__3627, w__3628, w__3629, w__3630, w__3631, w__3632;
  wire w__3633, w__3634, w__3635, w__3636, w__3637, w__3638, w__3639, w__3640;
  wire w__3641, w__3642, w__3643, w__3644, w__3645, w__3646, w__3647, w__3648;
  wire w__3649, w__3650, w__3651, w__3652, w__3653, w__3654, w__3655, w__3656;
  wire w__3657, w__3658, w__3659, w__3660, w__3661, w__3662, w__3663, w__3664;
  wire w__3665, w__3666, w__3667, w__3668, w__3669, w__3670, w__3671, w__3672;
  wire w__3673, w__3674, w__3675, w__3676, w__3677, w__3678, w__3679, w__3680;
  wire w__3681, w__3682, w__3683, w__3684, w__3685, w__3686, w__3687, w__3688;
  wire w__3689, w__3690, w__3691, w__3692, w__3693, w__3694, w__3695, w__3696;
  wire w__3697, w__3698, w__3699, w__3700, w__3701, w__3702, w__3703, w__3704;
  wire w__3705, w__3706, w__3707, w__3708, w__3709, w__3710, w__3711, w__3712;
  wire w__3713, w__3714, w__3715, w__3716, w__3717, w__3718, w__3719, w__3720;
  wire w__3721, w__3722, w__3723, w__3724, w__3725, w__3726, w__3727, w__3728;
  wire w__3729, w__3730, w__3731, w__3732, w__3733, w__3734, w__3735, w__3736;
  wire w__3737, w__3738, w__3739, w__3740, w__3741, w__3742, w__3743, w__3744;
  wire w__3745, w__3746, w__3747, w__3748, w__3749, w__3750, w__3751, w__3752;
  wire w__3753, w__3754, w__3755, w__3756, w__3757, w__3758, w__3759, w__3760;
  wire w__3761, w__3762, w__3763, w__3764, w__3765, w__3766, w__3767, w__3768;
  wire w__3769, w__3770, w__3771, w__3772, w__3773, w__3774, w__3775, w__3776;
  wire w__3777, w__3778, w__3779, w__3780, w__3781, w__3782, w__3783, w__3784;
  wire w__3785, w__3786, w__3787, w__3788, w__3789, w__3790, w__3791, w__3792;
  wire w__3793, w__3794, w__3795, w__3796, w__3797, w__3798, w__3799, w__3800;
  wire w__3801, w__3802, w__3803, w__3804, w__3805, w__3806, w__3807, w__3808;
  wire w__3809, w__3810, w__3811, w__3812, w__3813, w__3814, w__3815, w__3816;
  wire w__3817, w__3818, w__3819, w__3820, w__3821, w__3822, w__3823, w__3824;
  wire w__3825, w__3826, w__3827, w__3828, w__3829, w__3830, w__3831, w__3832;
  wire w__3833, w__3834, w__3835, w__3836, w__3837, w__3838, w__3839, w__3840;
  wire w__3841, w__3842, w__3843, w__3844, w__3845, w__3846, w__3847, w__3848;
  wire w__3849, w__3850, w__3851, w__3852, w__3853, w__3854, w__3855, w__3856;
  wire w__3857, w__3858, w__3859, w__3860, w__3861, w__3862, w__3863, w__3864;
  wire w__3865, w__3866, w__3867, w__3868, w__3869, w__3870, w__3871, w__3872;
  wire w__3873, w__3874, w__3875, w__3876, w__3877, w__3878, w__3879, w__3880;
  wire w__3881, w__3882, w__3883, w__3884, w__3885, w__3886, w__3887, w__3888;
  wire w__3889, w__3890, w__3891, w__3892, w__3893, w__3894, w__3895, w__3896;
  wire w__3897, w__3898, w__3899, w__3900, w__3901, w__3902, w__3903, w__3904;
  wire w__3905, w__3906, w__3907, w__3908, w__3909, w__3910, w__3911, w__3912;
  wire w__3913, w__3914, w__3915, w__3916, w__3917, w__3918, w__3919, w__3920;
  wire w__3921, w__3922, w__3923, w__3924, w__3925, w__3926, w__3927, w__3928;
  wire w__3929, w__3930, w__3931, w__3932, w__3933, w__3934, w__3935, w__3936;
  wire w__3937, w__3938, w__3939, w__3940, w__3941, w__3942, w__3943, w__3944;
  wire w__3945, w__3946, w__3947, w__3948, w__3949, w__3950, w__3951, w__3952;
  wire w__3953, w__3954, w__3955, w__3956, w__3957, w__3958, w__3959, w__3960;
  wire w__3961, w__3962, w__3963, w__3964, w__3965, w__3966, w__3967, w__3968;
  wire w__3969, w__3970, w__3971, w__3972, w__3973, w__3974, w__3975, w__3976;
  wire w__3977, w__3978, w__3979, w__3980, w__3981, w__3982, w__3983, w__3984;
  wire w__3985, w__3986, w__3987, w__3988, w__3989, w__3990, w__3991, w__3992;
  wire w__3993, w__3994, w__3995, w__3996, w__3997, w__3998, w__3999, w__4000;
  wire w__4001, w__4002, w__4003, w__4004, w__4005, w__4006, w__4007, w__4008;
  wire w__4009, w__4010, w__4011, w__4012, w__4013, w__4014, w__4015, w__4016;
  wire w__4017, w__4018, w__4019, w__4020, w__4021, w__4022, w__4023, w__4024;
  wire w__4025, w__4026, w__4027, w__4028, w__4029, w__4030, w__4031, w__4032;
  wire w__4033, w__4034, w__4035, w__4036, w__4037, w__4038, w__4039, w__4040;
  wire w__4041, w__4042, w__4043, w__4044, w__4045, w__4046, w__4047, w__4048;
  wire w__4049, w__4050, w__4051, w__4052, w__4053, w__4054, w__4055, w__4056;
  wire w__4057, w__4058, w__4059, w__4060, w__4061, w__4062, w__4063, w__4064;
  wire w__4065, w__4066, w__4067, w__4068, w__4069, w__4070, w__4071, w__4072;
  wire w__4073, w__4074, w__4075, w__4076, w__4077, w__4078, w__4079, w__4080;
  wire w__4081, w__4082, w__4083, w__4084, w__4085, w__4086, w__4087, w__4088;
  wire w__4089, w__4090, w__4091, w__4092, w__4093, w__4094, w__4095, w__4096;
  wire w__4097, w__4098, w__4099, w__4100, w__4101, w__4102, w__4103, w__4104;
  wire w__4105, w__4106, w__4107, w__4108, w__4109, w__4110, w__4111, w__4112;
  wire w__4113, w__4114, w__4115, w__4116, w__4117, w__4118, w__4119, w__4120;
  wire w__4121, w__4122, w__4123, w__4124, w__4125, w__4126, w__4127, w__4128;
  wire w__4129, w__4130, w__4131, w__4132, w__4133, w__4134, w__4135, w__4136;
  wire w__4137, w__4138, w__4139, w__4140, w__4141, w__4142, w__4143, w__4144;
  wire w__4145, w__4146, w__4147, w__4148, w__4149, w__4150, w__4151, w__4152;
  wire w__4153, w__4154, w__4155, w__4156, w__4157, w__4158, w__4159, w__4160;
  wire w__4161, w__4162, w__4163, w__4164, w__4165, w__4166, w__4167, w__4168;
  wire w__4169, w__4170, w__4171, w__4172, w__4173, w__4174, w__4175, w__4176;
  wire w__4177, w__4178, w__4179, w__4180, w__4181, w__4182, w__4183, w__4184;
  wire w__4185, w__4186, w__4187, w__4188, w__4189, w__4190, w__4191, w__4192;
  wire w__4193, w__4194, w__4195, w__4196, w__4197, w__4198, w__4199, w__4200;
  wire w__4201, w__4202, w__4203, w__4204, w__4205, w__4206, w__4207, w__4208;
  wire w__4209, w__4210, w__4211, w__4212, w__4213, w__4214, w__4215, w__4216;
  wire w__4217, w__4218, w__4219, w__4220, w__4221, w__4222, w__4223, w__4224;
  wire w__4225, w__4226, w__4227, w__4228, w__4229, w__4230, w__4231, w__4232;
  wire w__4233, w__4234, w__4235, w__4236, w__4237, w__4238, w__4239, w__4240;
  wire w__4241, w__4242, w__4243, w__4244, w__4245, w__4246, w__4247, w__4248;
  wire w__4249, w__4250, w__4251, w__4252, w__4253, w__4254, w__4255, w__4256;
  wire w__4257, w__4258, w__4259, w__4260, w__4261, w__4262, w__4263, w__4264;
  wire w__4265, w__4266, w__4267, w__4268, w__4269, w__4270, w__4271, w__4272;
  wire w__4273, w__4274, w__4275, w__4276, w__4277, w__4278, w__4279, w__4280;
  wire w__4281, w__4282, w__4283, w__4284, w__4285, w__4286, w__4287, w__4288;
  wire w__4289, w__4290, w__4291, w__4292, w__4293, w__4294, w__4295, w__4296;
  wire w__4297, w__4298, w__4299, w__4300, w__4301, w__4302, w__4303, w__4304;
  wire w__4305, w__4306, w__4307, w__4308, w__4309, w__4310, w__4311, w__4312;
  wire w__4313, w__4314, w__4315, w__4316, w__4317, w__4318, w__4319, w__4320;
  wire w__4321, w__4322, w__4323, w__4324, w__4325, w__4326, w__4327, w__4328;
  wire w__4329, w__4330, w__4331, w__4332, w__4333, w__4334, w__4335, w__4336;
  wire w__4337, w__4338, w__4339, w__4340, w__4341, w__4342, w__4343, w__4344;
  wire w__4345, w__4346, w__4347, w__4348, w__4349, w__4350, w__4351, w__4352;
  wire w__4353, w__4354, w__4355, w__4356, w__4357, w__4358, w__4359, w__4360;
  wire w__4361, w__4362, w__4363, w__4364, w__4365, w__4366, w__4367, w__4368;
  wire w__4369, w__4370, w__4371, w__4372, w__4373, w__4374, w__4375, w__4376;
  wire w__4377, w__4378, w__4379, w__4380, w__4381, w__4382, w__4383, w__4384;
  wire w__4385, w__4386, w__4387, w__4388, w__4389, w__4390, w__4391, w__4392;
  wire w__4393, w__4394, w__4395, w__4396, w__4397, w__4398, w__4399, w__4400;
  wire w__4401, w__4402, w__4403, w__4404, w__4405, w__4406, w__4407, w__4408;
  wire w__4409, w__4410, w__4411, w__4412, w__4413, w__4414, w__4415, w__4416;
  wire w__4417, w__4418, w__4419, w__4420, w__4421, w__4422, w__4423, w__4424;
  wire w__4425, w__4426, w__4427, w__4428, w__4429, w__4430, w__4431, w__4432;
  wire w__4433, w__4434, w__4435, w__4436, w__4437, w__4438, w__4439, w__4440;
  wire w__4441, w__4442, w__4443, w__4444, w__4445, w__4446, w__4447, w__4448;
  wire w__4449, w__4450, w__4451, w__4452, w__4453, w__4454, w__4455, w__4456;
  wire w__4457, w__4458, w__4459, w__4460, w__4461, w__4462, w__4463, w__4464;
  wire w__4465, w__4466, w__4467, w__4468, w__4469, w__4470, w__4471, w__4472;
  wire w__4473, w__4474, w__4475, w__4476, w__4477, w__4478, w__4479, w__4480;
  wire w__4481, w__4482, w__4483, w__4484, w__4485, w__4486, w__4487, w__4488;
  wire w__4489, w__4490, w__4491, w__4492, w__4493, w__4494, w__4495, w__4496;
  wire w__4497, w__4498, w__4499, w__4500, w__4501, w__4502, w__4503, w__4504;
  wire w__4505, w__4506, w__4507, w__4508, w__4509, w__4510, w__4511, w__4512;
  wire w__4513, w__4514, w__4515, w__4516, w__4517, w__4518, w__4519, w__4520;
  wire w__4521, w__4522, w__4523, w__4524, w__4525, w__4526, w__4527, w__4528;
  wire w__4529, w__4530, w__4531, w__4532, w__4533, w__4534, w__4535, w__4536;
  wire w__4537, w__4538, w__4539, w__4540, w__4541, w__4542, w__4543, w__4544;
  wire w__4545, w__4546, w__4547, w__4548, w__4549, w__4550, w__4551, w__4552;
  wire w__4553, w__4554, w__4555, w__4556, w__4557, w__4558, w__4559, w__4560;
  wire w__4561, w__4562, w__4563, w__4564, w__4565, w__4566, w__4567, w__4568;
  wire w__4569, w__4570, w__4571, w__4572, w__4573, w__4574, w__4575, w__4576;
  wire w__4577, w__4578, w__4579, w__4580, w__4581, w__4582, w__4583, w__4584;
  wire w__4585, w__4586, w__4587, w__4588, w__4589, w__4590, w__4591, w__4592;
  wire w__4593, w__4594, w__4595, w__4596, w__4597, w__4598, w__4599, w__4600;
  wire w__4601, w__4602, w__4603, w__4604, w__4605, w__4606, w__4607, w__4608;
  wire w__4609, w__4610, w__4611, w__4612, w__4613, w__4614, w__4615, w__4616;
  wire w__4617, w__4618, w__4619, w__4620, w__4621, w__4622, w__4623, w__4624;
  wire w__4625, w__4626, w__4627, w__4628, w__4629, w__4630, w__4631, w__4632;
  wire w__4633, w__4634, w__4635, w__4636, w__4637, w__4638, w__4639, w__4640;
  wire w__4641, w__4642, w__4643, w__4644, w__4645, w__4646, w__4647, w__4648;
  wire w__4649, w__4650, w__4651, w__4652, w__4653, w__4654, w__4655, w__4656;
  wire w__4657, w__4658, w__4659, w__4660, w__4661, w__4662, w__4663, w__4664;
  wire w__4665, w__4666, w__4667, w__4668, w__4669, w__4670, w__4671, w__4672;
  wire w__4673, w__4674, w__4675, w__4676, w__4677, w__4678, w__4679, w__4680;
  wire w__4681, w__4682, w__4683, w__4684, w__4685, w__4686, w__4687, w__4688;
  wire w__4689, w__4690, w__4691, w__4692, w__4693, w__4694, w__4695, w__4696;
  wire w__4697, w__4698, w__4699, w__4700, w__4701, w__4702, w__4703, w__4704;
  wire w__4705, w__4706, w__4707, w__4708, w__4709, w__4710, w__4711, w__4712;
  wire w__4713, w__4714, w__4715, w__4716, w__4717, w__4718, w__4719, w__4720;
  wire w__4721, w__4722, w__4723, w__4724, w__4725, w__4726, w__4727, w__4728;
  wire w__4729, w__4730, w__4731, w__4732, w__4733, w__4734, w__4735, w__4736;
  wire w__4737, w__4738, w__4739, w__4740, w__4741, w__4742, w__4743, w__4744;
  wire w__4745, w__4746, w__4747, w__4748, w__4749, w__4750, w__4751, w__4752;
  wire w__4753, w__4754, w__4755, w__4756, w__4757, w__4758, w__4759, w__4760;
  wire w__4761, w__4762, w__4763, w__4764, w__4765, w__4766, w__4767, w__4768;
  wire w__4769, w__4770, w__4771, w__4772, w__4773, w__4774, w__4775, w__4776;
  wire w__4777, w__4778, w__4779, w__4780, w__4781, w__4782, w__4783, w__4784;
  wire w__4785, w__4786, w__4787, w__4788, w__4789, w__4790, w__4791, w__4792;
  wire w__4793, w__4794, w__4795, w__4796, w__4797, w__4798, w__4799, w__4800;
  wire w__4801, w__4802, w__4803, w__4804, w__4805, w__4806, w__4807, w__4808;
  wire w__4809, w__4810, w__4811, w__4812, w__4813, w__4814, w__4815, w__4816;
  wire w__4817, w__4818, w__4819, w__4820, w__4821, w__4822, w__4823, w__4824;
  wire w__4825, w__4826, w__4827, w__4828, w__4829, w__4830, w__4831, w__4832;
  wire w__4833, w__4834, w__4835, w__4836, w__4837, w__4838, w__4839, w__4840;
  wire w__4841, w__4842, w__4843, w__4844, w__4845, w__4846, w__4847, w__4848;
  wire w__4849, w__4850, w__4851, w__4852, w__4853, w__4854, w__4855, w__4856;
  wire w__4857, w__4858, w__4859, w__4860, w__4861, w__4862, w__4863, w__4864;
  wire w__4865, w__4866, w__4867, w__4868, w__4869, w__4870, w__4871, w__4872;
  wire w__4873, w__4874, w__4875, w__4876, w__4877, w__4878, w__4879, w__4880;
  wire w__4881, w__4882, w__4883, w__4884, w__4885, w__4886, w__4887, w__4888;
  wire w__4889, w__4890, w__4891, w__4892, w__4893, w__4894, w__4895, w__4896;
  wire w__4897, w__4898, w__4899, w__4900, w__4901, w__4902, w__4903, w__4904;
  wire w__4905, w__4906, w__4907, w__4908, w__4909, w__4910, w__4911, w__4912;
  wire w__4913, w__4914, w__4915, w__4916, w__4917, w__4918, w__4919, w__4920;
  wire w__4921, w__4922, w__4923, w__4924, w__4925, w__4926, w__4927, w__4928;
  wire w__4929, w__4930, w__4931, w__4932, w__4933, w__4934, w__4935, w__4936;
  wire w__4937, w__4938, w__4939, w__4940, w__4941, w__4942, w__4943, w__4944;
  wire w__4945, w__4946, w__4947, w__4948, w__4949, w__4950, w__4951, w__4952;
  wire w__4953, w__4954, w__4955, w__4956, w__4957, w__4958, w__4959, w__4960;
  wire w__4961, w__4962, w__4963, w__4964, w__4965, w__4966, w__4967, w__4968;
  wire w__4969, w__4970, w__4971, w__4972, w__4973, w__4974, w__4975, w__4976;
  wire w__4977, w__4978, w__4979, w__4980, w__4981, w__4982, w__4983, w__4984;
  wire w__4985, w__4986, w__4987, w__4988, w__4989, w__4990, w__4991, w__4992;
  wire w__4993, w__4994, w__4995, w__4996, w__4997, w__4998, w__4999, w__5000;
  wire w__5001, w__5002, w__5003, w__5004, w__5005, w__5006, w__5007, w__5008;
  wire w__5009, w__5010, w__5011, w__5012, w__5013, w__5014, w__5015, w__5016;
  wire w__5017, w__5018, w__5019, w__5020, w__5021, w__5022, w__5023, w__5024;
  wire w__5025, w__5026, w__5027, w__5028, w__5029, w__5030, w__5031, w__5032;
  wire w__5033, w__5034, w__5035, w__5036, w__5037, w__5038, w__5039, w__5040;
  wire w__5041, w__5042, w__5043, w__5044, w__5045, w__5046, w__5047, w__5048;
  wire w__5049, w__5050, w__5051, w__5052, w__5053, w__5054, w__5055, w__5056;
  wire w__5057, w__5058, w__5059, w__5060, w__5061, w__5062, w__5063, w__5064;
  wire w__5065, w__5066, w__5067, w__5068, w__5069, w__5070, w__5071, w__5072;
  wire w__5073, w__5074, w__5075, w__5076, w__5077, w__5078, w__5079, w__5080;
  wire w__5081, w__5082, w__5083, w__5084, w__5085, w__5086, w__5087, w__5088;
  wire w__5089, w__5090, w__5091, w__5092, w__5093, w__5094, w__5095, w__5096;
  wire w__5097, w__5098, w__5099, w__5100, w__5101, w__5102, w__5103, w__5104;
  wire w__5105, w__5106, w__5107, w__5108, w__5109, w__5110, w__5111, w__5112;
  wire w__5113, w__5114, w__5115, w__5116, w__5117, w__5118, w__5119, w__5120;
  wire w__5121, w__5122, w__5123, w__5124, w__5125, w__5126, w__5127, w__5128;
  wire w__5129, w__5130, w__5131, w__5132, w__5133, w__5134, w__5135, w__5136;
  wire w__5137, w__5138, w__5139, w__5140, w__5141, w__5142, w__5143, w__5144;
  wire w__5145, w__5146, w__5147, w__5148, w__5149, w__5150, w__5151, w__5152;
  wire w__5153, w__5154, w__5155, w__5156, w__5157, w__5158, w__5159, w__5160;
  wire w__5161, w__5162, w__5163, w__5164, w__5165, w__5166, w__5167, w__5168;
  wire w__5169, w__5170, w__5171, w__5172, w__5173, w__5174, w__5175, w__5176;
  wire w__5177, w__5178, w__5179, w__5180, w__5181, w__5182, w__5183, w__5184;
  wire w__5185, w__5186, w__5187, w__5188, w__5189, w__5190, w__5191, w__5192;
  wire w__5193, w__5194, w__5195, w__5196, w__5197, w__5198, w__5199, w__5200;
  wire w__5201, w__5202, w__5203, w__5204, w__5205, w__5206, w__5207, w__5208;
  wire w__5209, w__5210, w__5211, w__5212, w__5213, w__5214, w__5215, w__5216;
  wire w__5217, w__5218, w__5219, w__5220, w__5221, w__5222, w__5223, w__5224;
  wire w__5225, w__5226, w__5227, w__5228, w__5229, w__5230, w__5231, w__5232;
  wire w__5233, w__5234, w__5235, w__5236, w__5237, w__5238, w__5239, w__5240;
  wire w__5241, w__5242, w__5243, w__5244, w__5245, w__5246, w__5247, w__5248;
  wire w__5249, w__5250, w__5251, w__5252, w__5253, w__5254, w__5255, w__5256;
  wire w__5257, w__5258, w__5259, w__5260, w__5261, w__5262, w__5263, w__5264;
  wire w__5265, w__5266, w__5267, w__5268, w__5269, w__5270, w__5271, w__5272;
  wire w__5273, w__5274, w__5275, w__5276, w__5277, w__5278, w__5279, w__5280;
  wire w__5281, w__5282, w__5283, w__5284, w__5285, w__5286, w__5287, w__5288;
  wire w__5289, w__5290, w__5291, w__5292, w__5293, w__5294, w__5295, w__5296;
  wire w__5297, w__5298, w__5299, w__5300, w__5301, w__5302, w__5303, w__5304;
  wire w__5305, w__5306, w__5307, w__5308, w__5309, w__5310, w__5311, w__5312;
  wire w__5313, w__5314, w__5315, w__5316, w__5317, w__5318, w__5319, w__5320;
  wire w__5321, w__5322, w__5323, w__5324, w__5325, w__5326, w__5327, w__5328;
  wire w__5329, w__5330, w__5331, w__5332, w__5333, w__5334, w__5335, w__5336;
  wire w__5337, w__5338, w__5339, w__5340, w__5341, w__5342, w__5343, w__5344;
  wire w__5345, w__5346, w__5347, w__5348, w__5349, w__5350, w__5351, w__5352;
  wire w__5353, w__5354, w__5355, w__5356, w__5357, w__5358, w__5359, w__5360;
  wire w__5361, w__5362, w__5363, w__5364, w__5365, w__5366, w__5367, w__5368;
  wire w__5369, w__5370, w__5371, w__5372, w__5373, w__5374, w__5375, w__5376;
  wire w__5377, w__5378, w__5379, w__5380, w__5381, w__5382, w__5383, w__5384;
  wire w__5385, w__5386, w__5387, w__5388, w__5389, w__5390, w__5391, w__5392;
  wire w__5393, w__5394, w__5395, w__5396, w__5397, w__5398, w__5399, w__5400;
  wire w__5401, w__5402, w__5403, w__5404, w__5405, w__5406, w__5407, w__5408;
  wire w__5409, w__5410, w__5411, w__5412, w__5413, w__5414, w__5415, w__5416;
  wire w__5417, w__5418, w__5419, w__5420, w__5421, w__5422, w__5423, w__5424;
  wire w__5425, w__5426, w__5427, w__5428, w__5429, w__5430, w__5431, w__5432;
  wire w__5433, w__5434, w__5435, w__5436, w__5437, w__5438, w__5439, w__5440;
  wire w__5441, w__5442, w__5443, w__5444, w__5445, w__5446, w__5447, w__5448;
  wire w__5449, w__5450, w__5451, w__5452, w__5453, w__5454, w__5455, w__5456;
  wire w__5457, w__5458, w__5459, w__5460, w__5461, w__5462, w__5463, w__5464;
  wire w__5465, w__5466, w__5467, w__5468, w__5469, w__5470, w__5471, w__5472;
  wire w__5473, w__5474, w__5475, w__5476, w__5477, w__5478, w__5479, w__5480;
  wire w__5481, w__5482, w__5483, w__5484, w__5485, w__5486, w__5487, w__5488;
  wire w__5489, w__5490, w__5491, w__5492, w__5493, w__5494, w__5495, w__5496;
  wire w__5497, w__5498, w__5499, w__5500, w__5501, w__5502, w__5503, w__5504;
  wire w__5505, w__5506, w__5507, w__5508, w__5509, w__5510, w__5511, w__5512;
  wire w__5513, w__5514, w__5515, w__5516, w__5517, w__5518, w__5519, w__5520;
  wire w__5521, w__5522, w__5523, w__5524, w__5525, w__5526, w__5527, w__5528;
  wire w__5529, w__5530, w__5531, w__5532, w__5533, w__5534, w__5535, w__5536;
  wire w__5537, w__5538, w__5539, w__5540, w__5541, w__5542, w__5543, w__5544;
  wire w__5545, w__5546, w__5547, w__5548, w__5549, w__5550, w__5551, w__5552;
  wire w__5553, w__5554, w__5555, w__5556, w__5557, w__5558, w__5559, w__5560;
  wire w__5561, w__5562, w__5563, w__5564, w__5565, w__5566, w__5567, w__5568;
  wire w__5569, w__5570, w__5571, w__5572, w__5573, w__5574, w__5575, w__5576;
  wire w__5577, w__5578, w__5579, w__5580, w__5581, w__5582, w__5583, w__5584;
  wire w__5585, w__5586, w__5587, w__5588, w__5589, w__5590, w__5591, w__5592;
  wire w__5593, w__5594, w__5595, w__5596, w__5597, w__5598, w__5599, w__5600;
  wire w__5601, w__5602, w__5603, w__5604, w__5605, w__5606, w__5607, w__5608;
  wire w__5609, w__5610, w__5611, w__5612, w__5613, w__5614, w__5615, w__5616;
  wire w__5617, w__5618, w__5619, w__5620, w__5621, w__5622, w__5623, w__5624;
  wire w__5625, w__5626, w__5627, w__5628, w__5629, w__5630, w__5631, w__5632;
  wire w__5633, w__5634, w__5635, w__5636, w__5637, w__5638, w__5639, w__5640;
  wire w__5641, w__5642, w__5643, w__5644, w__5645, w__5646, w__5647, w__5648;
  wire w__5649, w__5650, w__5651, w__5652, w__5653, w__5654, w__5655, w__5656;
  wire w__5657, w__5658, w__5659, w__5660, w__5661, w__5662, w__5663, w__5664;
  wire w__5665, w__5666, w__5667, w__5668, w__5669, w__5670, w__5671, w__5672;
  wire w__5673, w__5674, w__5675, w__5676, w__5677, w__5678, w__5679, w__5680;
  wire w__5681, w__5682, w__5683, w__5684, w__5685, w__5686, w__5687, w__5688;
  wire w__5689, w__5690, w__5691, w__5692, w__5693, w__5694, w__5695, w__5696;
  wire w__5697, w__5698, w__5699, w__5700, w__5701, w__5702, w__5703, w__5704;
  wire w__5705, w__5706, w__5707, w__5708, w__5709, w__5710, w__5711, w__5712;
  wire w__5713, w__5714, w__5715, w__5716, w__5717, w__5718, w__5719, w__5720;
  wire w__5721, w__5722, w__5723, w__5724, w__5725, w__5726, w__5727, w__5728;
  wire w__5729, w__5730, w__5731, w__5732, w__5733, w__5734, w__5735, w__5736;
  wire w__5737, w__5738, w__5739, w__5740, w__5741, w__5742, w__5743, w__5744;
  wire w__5745, w__5746, w__5747, w__5748, w__5749, w__5750, w__5751, w__5752;
  wire w__5753, w__5754, w__5755, w__5756, w__5757, w__5758, w__5759, w__5760;
  wire w__5761, w__5762, w__5763, w__5764, w__5765, w__5766, w__5767, w__5768;
  wire w__5769, w__5770, w__5771, w__5772, w__5773, w__5774, w__5775, w__5776;
  wire w__5777, w__5778, w__5779, w__5780, w__5781, w__5782, w__5783, w__5784;
  wire w__5785, w__5786, w__5787, w__5788, w__5789, w__5790, w__5791, w__5792;
  wire w__5793, w__5794, w__5795, w__5796, w__5797, w__5798, w__5799, w__5800;
  wire w__5801, w__5802, w__5803, w__5804, w__5805, w__5806, w__5807, w__5808;
  wire w__5809, w__5810, w__5811, w__5812, w__5813, w__5814, w__5815, w__5816;
  wire w__5817, w__5818, w__5819, w__5820, w__5821, w__5822, w__5823, w__5824;
  wire w__5825, w__5826, w__5827, w__5828, w__5829, w__5830, w__5831, w__5832;
  wire w__5833, w__5834, w__5835, w__5836, w__5837, w__5838, w__5839, w__5840;
  wire w__5841, w__5842, w__5843, w__5844, w__5845, w__5846, w__5847, w__5848;
  wire w__5849, w__5850, w__5851, w__5852, w__5853, w__5854, w__5855, w__5856;
  wire w__5857, w__5858, w__5859, w__5860, w__5861, w__5862, w__5863, w__5864;
  wire w__5865, w__5866, w__5867, w__5868, w__5869, w__5870, w__5871, w__5872;
  wire w__5873, w__5874, w__5875, w__5876, w__5877, w__5878, w__5879, w__5880;
  wire w__5881, w__5882, w__5883, w__5884, w__5885, w__5886, w__5887, w__5888;
  wire w__5889, w__5890, w__5891, w__5892, w__5893, w__5894, w__5895, w__5896;
  wire w__5897, w__5898, w__5899, w__5900, w__5901, w__5902, w__5903, w__5904;
  wire w__5905, w__5906, w__5907, w__5908, w__5909, w__5910, w__5911, w__5912;
  wire w__5913, w__5914, w__5915, w__5916, w__5917, w__5918, w__5919, w__5920;
  wire w__5921, w__5922, w__5923, w__5924, w__5925, w__5926, w__5927, w__5928;
  wire w__5929, w__5930, w__5931, w__5932, w__5933, w__5934, w__5935, w__5936;
  wire w__5937, w__5938, w__5939, w__5940, w__5941, w__5942, w__5943, w__5944;
  wire w__5945, w__5946, w__5947, w__5948, w__5949, w__5950, w__5951, w__5952;
  wire w__5953, w__5954, w__5955, w__5956, w__5957, w__5958, w__5959, w__5960;
  wire w__5961, w__5962, w__5963, w__5964, w__5965, w__5966, w__5967, w__5968;
  wire w__5969, w__5970, w__5971, w__5972, w__5973, w__5974, w__5975, w__5976;
  wire w__5977, w__5978, w__5979, w__5980, w__5981, w__5982, w__5983, w__5984;
  wire w__5985, w__5986, w__5987, w__5988, w__5989, w__5990, w__5991, w__5992;
  wire w__5993, w__5994, w__5995, w__5996, w__5997, w__5998, w__5999, w__6000;
  wire w__6001, w__6002, w__6003, w__6004, w__6005, w__6006, w__6007, w__6008;
  wire w__6009, w__6010, w__6011, w__6012, w__6013, w__6014, w__6015, w__6016;
  wire w__6017, w__6018, w__6019, w__6020, w__6021, w__6022, w__6023, w__6024;
  wire w__6025, w__6026, w__6027, w__6028, w__6029, w__6030, w__6031, w__6032;
  wire w__6033, w__6034, w__6035, w__6036, w__6037, w__6038, w__6039, w__6040;
  wire w__6041, w__6042, w__6043, w__6044, w__6045, w__6046, w__6047, w__6048;
  wire w__6049, w__6050, w__6051, w__6052, w__6053, w__6054, w__6055, w__6056;
  wire w__6057, w__6058, w__6059, w__6060, w__6061, w__6062, w__6063, w__6064;
  wire w__6065, w__6066, w__6067, w__6068, w__6069, w__6070, w__6071, w__6072;
  wire w__6073, w__6074, w__6075, w__6076, w__6077, w__6078, w__6079, w__6080;
  wire w__6081, w__6082, w__6083, w__6084, w__6085, w__6086, w__6087, w__6088;
  wire w__6089, w__6090, w__6091, w__6092, w__6093, w__6094, w__6095, w__6096;
  wire w__6097, w__6098, w__6099, w__6100, w__6101, w__6102, w__6103, w__6104;
  wire w__6105, w__6106, w__6107, w__6108, w__6109, w__6110, w__6111, w__6112;
  wire w__6113, w__6114, w__6115, w__6116, w__6117, w__6118, w__6119, w__6120;
  wire w__6121, w__6122, w__6123, w__6124, w__6125, w__6126, w__6127, w__6128;
  wire w__6129, w__6130, w__6131, w__6132, w__6133, w__6134, w__6135, w__6136;
  wire w__6137, w__6138, w__6139, w__6140, w__6141, w__6142, w__6143, w__6144;
  wire w__6145, w__6146, w__6147, w__6148, w__6149, w__6150, w__6151, w__6152;
  wire w__6153, w__6154, w__6155, w__6156, w__6157, w__6158, w__6159, w__6160;
  wire w__6161, w__6162, w__6163, w__6164, w__6165, w__6166, w__6167, w__6168;
  wire w__6169, w__6170, w__6171, w__6172, w__6173, w__6174, w__6175, w__6176;
  wire w__6177, w__6178, w__6179, w__6180, w__6181, w__6182, w__6183, w__6184;
  wire w__6185, w__6186, w__6187, w__6188, w__6189, w__6190, w__6191, w__6192;
  wire w__6193, w__6194, w__6195, w__6196, w__6197, w__6198, w__6199, w__6200;
  wire w__6201, w__6202, w__6203, w__6204, w__6205, w__6206, w__6207, w__6208;
  wire w__6209, w__6210, w__6211, w__6212, w__6213, w__6214, w__6215, w__6216;
  wire w__6217, w__6218, w__6219, w__6220, w__6221, w__6222, w__6223, w__6224;
  wire w__6225, w__6226, w__6227, w__6228, w__6229, w__6230, w__6231, w__6232;
  wire w__6233, w__6234, w__6235, w__6236, w__6237, w__6238, w__6239, w__6240;
  wire w__6241, w__6242, w__6243, w__6244, w__6245, w__6246, w__6247, w__6248;
  wire w__6249, w__6250, w__6251, w__6252, w__6253, w__6254, w__6255, w__6256;
  wire w__6257, w__6258, w__6259, w__6260, w__6261, w__6262, w__6263, w__6264;
  wire w__6265, w__6266, w__6267, w__6268, w__6269, w__6270, w__6271, w__6272;
  wire w__6273, w__6274, w__6275, w__6276, w__6277, w__6278, w__6279, w__6280;
  wire w__6281, w__6282, w__6283, w__6284, w__6285, w__6286, w__6287, w__6288;
  wire w__6289, w__6290, w__6291, w__6292, w__6293, w__6294, w__6295, w__6296;
  wire w__6297, w__6298, w__6299, w__6300, w__6301, w__6302, w__6303, w__6304;
  wire w__6305, w__6306, w__6307, w__6308, w__6309, w__6310, w__6311, w__6312;
  wire w__6313, w__6314, w__6315, w__6316, w__6317, w__6318, w__6319, w__6320;
  wire w__6321, w__6322, w__6323, w__6324, w__6325, w__6326, w__6327, w__6328;
  wire w__6329, w__6330, w__6331, w__6332, w__6333, w__6334, w__6335, w__6336;
  wire w__6337, w__6338, w__6339, w__6340, w__6341, w__6342, w__6343, w__6344;
  wire w__6345, w__6346, w__6347, w__6348, w__6349, w__6350, w__6351, w__6352;
  wire w__6353, w__6354, w__6355, w__6356, w__6357, w__6358, w__6359, w__6360;
  wire w__6361, w__6362, w__6363, w__6364, w__6365, w__6366, w__6367, w__6368;
  wire w__6369, w__6370, w__6371, w__6372, w__6373, w__6374, w__6375, w__6376;
  wire w__6377, w__6378, w__6379, w__6380, w__6381, w__6382, w__6383, w__6384;
  wire w__6385, w__6386, w__6387, w__6388, w__6389, w__6390, w__6391, w__6392;
  wire w__6393, w__6394, w__6395, w__6396, w__6397, w__6398, w__6399, w__6400;
  wire w__6401, w__6402, w__6403, w__6404, w__6405, w__6406, w__6407, w__6408;
  wire w__6409, w__6410, w__6411, w__6412, w__6413, w__6414, w__6415, w__6416;
  wire w__6417, w__6418, w__6419, w__6420, w__6421, w__6422, w__6423, w__6424;
  wire w__6425, w__6426, w__6427, w__6428, w__6429, w__6430, w__6431, w__6432;
  wire w__6433, w__6434, w__6435, w__6436, w__6437, w__6438, w__6439, w__6440;
  wire w__6441, w__6442, w__6443, w__6444, w__6445, w__6446, w__6447, w__6448;
  wire w__6449, w__6450, w__6451, w__6452, w__6453, w__6454, w__6455, w__6456;
  wire w__6457, w__6458, w__6459, w__6460, w__6461, w__6462, w__6463, w__6464;
  wire w__6465, w__6466, w__6467, w__6468, w__6469, w__6470, w__6471, w__6472;
  wire w__6473, w__6474, w__6475, w__6476, w__6477, w__6478, w__6479, w__6480;
  wire w__6481, w__6482, w__6483, w__6484, w__6485, w__6486, w__6487, w__6488;
  wire w__6489, w__6490, w__6491, w__6492, w__6493, w__6494, w__6495, w__6496;
  wire w__6497, w__6498, w__6499, w__6500, w__6501, w__6502, w__6503, w__6504;
  wire w__6505, w__6506, w__6507, w__6508, w__6509, w__6510, w__6511, w__6512;
  wire w__6513, w__6514, w__6515, w__6516, w__6517, w__6518, w__6519, w__6520;
  wire w__6521, w__6522, w__6523, w__6524, w__6525, w__6526, w__6527, w__6528;
  wire w__6529, w__6530, w__6531, w__6532, w__6533, w__6534, w__6535, w__6536;
  wire w__6537, w__6538, w__6539, w__6540, w__6541, w__6542, w__6543, w__6544;
  wire w__6545, w__6546, w__6547, w__6548, w__6549, w__6550, w__6551, w__6552;
  wire w__6553, w__6554, w__6555, w__6556, w__6557, w__6558, w__6559, w__6560;
  wire w__6561, w__6562, w__6563, w__6564, w__6565, w__6566, w__6567, w__6568;
  wire w__6569, w__6570, w__6571, w__6572, w__6573, w__6574, w__6575, w__6576;
  wire w__6577, w__6578, w__6579, w__6580, w__6581, w__6582, w__6583, w__6584;
  wire w__6585, w__6586, w__6587, w__6588, w__6589, w__6590, w__6591, w__6592;
  wire w__6593, w__6594, w__6595, w__6596, w__6597, w__6598, w__6599, w__6600;
  wire w__6601, w__6602, w__6603, w__6604, w__6605, w__6606, w__6607, w__6608;
  wire w__6609, w__6610, w__6611, w__6612, w__6613, w__6614, w__6615, w__6616;
  wire w__6617, w__6618, w__6619, w__6620, w__6621, w__6622, w__6623, w__6624;
  wire w__6625, w__6626, w__6627, w__6628, w__6629, w__6630, w__6631, w__6632;
  wire w__6633, w__6634, w__6635, w__6636, w__6637, w__6638, w__6639, w__6640;
  wire w__6641, w__6642, w__6643, w__6644, w__6645, w__6646, w__6647, w__6648;
  wire w__6649, w__6650, w__6651, w__6652, w__6653, w__6654, w__6655, w__6656;
  wire w__6657, w__6658, w__6659, w__6660, w__6661, w__6662, w__6663, w__6664;
  wire w__6665, w__6666, w__6667, w__6668, w__6669, w__6670, w__6671, w__6672;
  wire w__6673, w__6674, w__6675, w__6676, w__6677, w__6678, w__6679, w__6680;
  wire w__6681, w__6682, w__6683, w__6684, w__6685, w__6686, w__6687, w__6688;
  wire w__6689, w__6690, w__6691, w__6692, w__6693, w__6694, w__6695, w__6696;
  wire w__6697, w__6698, w__6699, w__6700, w__6701, w__6702, w__6703, w__6704;
  wire w__6705, w__6706, w__6707, w__6708, w__6709, w__6710, w__6711, w__6712;
  wire w__6713, w__6714, w__6715, w__6716, w__6717, w__6718, w__6719, w__6720;
  wire w__6721, w__6722, w__6723, w__6724, w__6725, w__6726, w__6727, w__6728;
  wire w__6729, w__6730, w__6731, w__6732, w__6733, w__6734, w__6735, w__6736;
  wire w__6737, w__6738, w__6739, w__6740, w__6741, w__6742, w__6743, w__6744;
  wire w__6745, w__6746, w__6747, w__6748, w__6749, w__6750, w__6751, w__6752;
  wire w__6753, w__6754, w__6755, w__6756, w__6757, w__6758, w__6759, w__6760;
  wire w__6761, w__6762, w__6763, w__6764, w__6765, w__6766, w__6767, w__6768;
  wire w__6769, w__6770, w__6771, w__6772, w__6773, w__6774, w__6775, w__6776;
  wire w__6777, w__6778, w__6779, w__6780, w__6781, w__6782, w__6783, w__6784;
  wire w__6785, w__6786, w__6787, w__6788, w__6789, w__6790, w__6791, w__6792;
  wire w__6793, w__6794, w__6795, w__6796, w__6797, w__6798, w__6799, w__6800;
  wire w__6801, w__6802, w__6803, w__6804, w__6805, w__6806, w__6807, w__6808;
  wire w__6809, w__6810, w__6811, w__6812, w__6813, w__6814, w__6815, w__6816;
  wire w__6817, w__6818, w__6819, w__6820, w__6821, w__6822, w__6823, w__6824;
  wire w__6825, w__6826, w__6827, w__6828, w__6829, w__6830, w__6831, w__6832;
  wire w__6833, w__6834, w__6835, w__6836, w__6837, w__6838, w__6839, w__6840;
  wire w__6841, w__6842, w__6843, w__6844, w__6845, w__6846, w__6847, w__6848;
  wire w__6849, w__6850, w__6851, w__6852, w__6853, w__6854, w__6855, w__6856;
  wire w__6857, w__6858, w__6859, w__6860, w__6861, w__6862, w__6863, w__6864;
  wire w__6865, w__6866, w__6867, w__6868, w__6869, w__6870, w__6871, w__6872;
  wire w__6873, w__6874, w__6875, w__6876, w__6877, w__6878, w__6879, w__6880;
  wire w__6881, w__6882, w__6883, w__6884, w__6885, w__6886, w__6887, w__6888;
  wire w__6889, w__6890, w__6891, w__6892, w__6893, w__6894, w__6895, w__6896;
  wire w__6897, w__6898, w__6899, w__6900, w__6901, w__6902, w__6903, w__6904;
  wire w__6905, w__6906, w__6907, w__6908, w__6909, w__6910, w__6911, w__6912;
  wire w__6913, w__6914, w__6915, w__6916, w__6917, w__6918, w__6919, w__6920;
  wire w__6921, w__6922, w__6923, w__6924, w__6925, w__6926, w__6927, w__6928;
  wire w__6929, w__6930, w__6931, w__6932, w__6933, w__6934, w__6935, w__6936;
  wire w__6937, w__6938, w__6939, w__6940, w__6941, w__6942, w__6943, w__6944;
  wire w__6945, w__6946, w__6947, w__6948, w__6949, w__6950, w__6951, w__6952;
  wire w__6953, w__6954, w__6955, w__6956, w__6957, w__6958, w__6959, w__6960;
  wire w__6961, w__6962, w__6963, w__6964, w__6965, w__6966, w__6967, w__6968;
  wire w__6969, w__6970, w__6971, w__6972, w__6973, w__6974, w__6975, w__6976;
  wire w__6977, w__6978, w__6979, w__6980, w__6981, w__6982, w__6983, w__6984;
  wire w__6985, w__6986, w__6987, w__6988, w__6989, w__6990, w__6991, w__6992;
  wire w__6993, w__6994, w__6995, w__6996, w__6997, w__6998, w__6999, w__7000;
  wire w__7001, w__7002, w__7003, w__7004, w__7005, w__7006, w__7007, w__7008;
  wire w__7009, w__7010, w__7011, w__7012, w__7013, w__7014, w__7015, w__7016;
  wire w__7017, w__7018, w__7019, w__7020, w__7021, w__7022, w__7023, w__7024;
  wire w__7025, w__7026, w__7027, w__7028, w__7029, w__7030, w__7031, w__7032;
  wire w__7033, w__7034, w__7035, w__7036, w__7037, w__7038, w__7039, w__7040;
  wire w__7041, w__7042, w__7043, w__7044, w__7045, w__7046, w__7047, w__7048;
  wire w__7049, w__7050, w__7051, w__7052, w__7053, w__7054, w__7055, w__7056;
  wire w__7057, w__7058, w__7059, w__7060, w__7061, w__7062, w__7063, w__7064;
  wire w__7065, w__7066, w__7067, w__7068, w__7069, w__7070, w__7071, w__7072;
  wire w__7073, w__7074, w__7075, w__7076, w__7077, w__7078, w__7079, w__7080;
  wire w__7081, w__7082, w__7083, w__7084, w__7085, w__7086, w__7087, w__7088;
  wire w__7089, w__7090, w__7091, w__7092, w__7093, w__7094, w__7095, w__7096;
  wire w__7097, w__7098, w__7099, w__7100, w__7101, w__7102, w__7103, w__7104;
  wire w__7105, w__7106, w__7107, w__7108, w__7109, w__7110, w__7111, w__7112;
  wire w__7113, w__7114, w__7115, w__7116, w__7117, w__7118, w__7119, w__7120;
  wire w__7121, w__7122, w__7123, w__7124, w__7125, w__7126, w__7127, w__7128;
  wire w__7129, w__7130, w__7131, w__7132, w__7133, w__7134, w__7135, w__7136;
  wire w__7137, w__7138, w__7139, w__7140, w__7141, w__7142, w__7143, w__7144;
  wire w__7145, w__7146, w__7147, w__7148, w__7149, w__7150, w__7151, w__7152;
  wire w__7153, w__7154, w__7155, w__7156, w__7157, w__7158, w__7159, w__7160;
  wire w__7161, w__7162, w__7163, w__7164, w__7165, w__7166, w__7167, w__7168;
  wire w__7169, w__7170, w__7171, w__7172, w__7173, w__7174, w__7175, w__7176;
  wire w__7177, w__7178, w__7179, w__7180, w__7181, w__7182, w__7183, w__7184;
  wire w__7185, w__7186, w__7187, w__7188, w__7189, w__7190, w__7191, w__7192;
  wire w__7193, w__7194, w__7195, w__7196, w__7197, w__7198, w__7199, w__7200;
  wire w__7201, w__7202, w__7203, w__7204, w__7205, w__7206, w__7207, w__7208;
  wire w__7209, w__7210, w__7211, w__7212, w__7213, w__7214, w__7215, w__7216;
  wire w__7217, w__7218, w__7219, w__7220, w__7221, w__7222, w__7223, w__7224;
  wire w__7225, w__7226, w__7227, w__7228, w__7229, w__7230, w__7231, w__7232;
  wire w__7233, w__7234, w__7235, w__7236, w__7237, w__7238, w__7239, w__7240;
  wire w__7241, w__7242, w__7243, w__7244, w__7245, w__7246, w__7247, w__7248;
  wire w__7249, w__7250, w__7251, w__7252, w__7253, w__7254, w__7255, w__7256;
  wire w__7257, w__7258, w__7259, w__7260, w__7261, w__7262, w__7263, w__7264;
  wire w__7265, w__7266, w__7267, w__7268, w__7269, w__7270, w__7271, w__7272;
  wire w__7273, w__7274, w__7275, w__7276, w__7277, w__7278, w__7279, w__7280;
  wire w__7281, w__7282, w__7283, w__7284, w__7285, w__7286, w__7287, w__7288;
  wire w__7289, w__7290, w__7291, w__7292, w__7293, w__7294, w__7295, w__7296;
  wire w__7297, w__7298, w__7299, w__7300, w__7301, w__7302, w__7303, w__7304;
  wire w__7305, w__7306, w__7307, w__7308, w__7309, w__7310, w__7311, w__7312;
  wire w__7313, w__7314, w__7315, w__7316, w__7317, w__7318, w__7319, w__7320;
  wire w__7321, w__7322, w__7323, w__7324, w__7325, w__7326, w__7327, w__7328;
  wire w__7329, w__7330, w__7331, w__7332, w__7333, w__7334, w__7335, w__7336;
  wire w__7337, w__7338, w__7339, w__7340, w__7341, w__7342, w__7343, w__7344;
  wire w__7345, w__7346, w__7347, w__7348, w__7349, w__7350, w__7351, w__7352;
  wire w__7353, w__7354, w__7355, w__7356, w__7357, w__7358, w__7359, w__7360;
  wire w__7361, w__7362, w__7363, w__7364, w__7365, w__7366, w__7367, w__7368;
  wire w__7369, w__7370, w__7371, w__7372, w__7373, w__7374, w__7375, w__7376;
  wire w__7377, w__7378, w__7379, w__7380, w__7381, w__7382, w__7383, w__7384;
  wire w__7385, w__7386, w__7387, w__7388, w__7389, w__7390, w__7391, w__7392;
  wire w__7393, w__7394, w__7395, w__7396, w__7397, w__7398, w__7399, w__7400;
  wire w__7401, w__7402, w__7403, w__7404, w__7405, w__7406, w__7407, w__7408;
  wire w__7409, w__7410, w__7411, w__7412, w__7413, w__7414, w__7415, w__7416;
  wire w__7417, w__7418, w__7419, w__7420, w__7421, w__7422, w__7423, w__7424;
  wire w__7425, w__7426, w__7427, w__7428, w__7429, w__7430, w__7431, w__7432;
  wire w__7433, w__7434, w__7435, w__7436, w__7437, w__7438, w__7439, w__7440;
  wire w__7441, w__7442, w__7443, w__7444, w__7445, w__7446, w__7447, w__7448;
  wire w__7449, w__7450, w__7451, w__7452, w__7453, w__7454, w__7455, w__7456;
  wire w__7457, w__7458, w__7459, w__7460, w__7461, w__7462, w__7463, w__7464;
  wire w__7465, w__7466, w__7467, w__7468, w__7469, w__7470, w__7471, w__7472;
  wire w__7473, w__7474, w__7475, w__7476, w__7477, w__7478, w__7479, w__7480;
  wire w__7481, w__7482, w__7483, w__7484, w__7485, w__7486, w__7487, w__7488;
  wire w__7489, w__7490, w__7491, w__7492, w__7493, w__7494, w__7495, w__7496;
  wire w__7497, w__7498, w__7499, w__7500, w__7501, w__7502, w__7503, w__7504;
  wire w__7505, w__7506, w__7507, w__7508, w__7509, w__7510, w__7511, w__7512;
  wire w__7513, w__7514, w__7515, w__7516, w__7517, w__7518, w__7519, w__7520;
  wire w__7521, w__7522, w__7523, w__7524, w__7525, w__7526, w__7527, w__7528;
  wire w__7529, w__7530, w__7531, w__7532, w__7533, w__7534, w__7535, w__7536;
  wire w__7537, w__7538, w__7539, w__7540, w__7541, w__7542, w__7543, w__7544;
  wire w__7545, w__7546, w__7547, w__7548, w__7549, w__7550, w__7551, w__7552;
  wire w__7553, w__7554, w__7555, w__7556, w__7557, w__7558, w__7559, w__7560;
  wire w__7561, w__7562, w__7563, w__7564, w__7565, w__7566, w__7567, w__7568;
  wire w__7569, w__7570, w__7571, w__7572, w__7573, w__7574, w__7575, w__7576;
  wire w__7577, w__7578, w__7579, w__7580, w__7581, w__7582, w__7583, w__7584;
  wire w__7585, w__7586, w__7587, w__7588, w__7589, w__7590, w__7591, w__7592;
  wire w__7593, w__7594, w__7595, w__7596, w__7597, w__7598, w__7599, w__7600;
  wire w__7601, w__7602, w__7603, w__7604, w__7605, w__7606, w__7607, w__7608;
  wire w__7609, w__7610, w__7611, w__7612, w__7613, w__7614, w__7615, w__7616;
  wire w__7617, w__7618, w__7619, w__7620, w__7621, w__7622, w__7623, w__7624;
  wire w__7625, w__7626, w__7627, w__7628, w__7629, w__7630, w__7631, w__7632;
  wire w__7633, w__7634, w__7635, w__7636, w__7637, w__7638, w__7639, w__7640;
  wire w__7641, w__7642, w__7643, w__7644, w__7645, w__7646, w__7647, w__7648;
  wire w__7649, w__7650, w__7651, w__7652, w__7653, w__7654, w__7655, w__7656;
  wire w__7657, w__7658, w__7659, w__7660, w__7661, w__7662, w__7663, w__7664;
  wire w__7665, w__7666, w__7667, w__7668, w__7669, w__7670, w__7671, w__7672;
  wire w__7673, w__7674, w__7675, w__7676, w__7677, w__7678, w__7679, w__7680;
  wire w__7681, w__7682, w__7683, w__7684, w__7685, w__7686, w__7687, w__7688;
  wire w__7689, w__7690, w__7691, w__7692, w__7693, w__7694, w__7695, w__7696;
  wire w__7697, w__7698, w__7699, w__7700, w__7701, w__7702, w__7703, w__7704;
  wire w__7705, w__7706, w__7707, w__7708, w__7709, w__7710, w__7711, w__7712;
  wire w__7713, w__7714, w__7715, w__7716, w__7717, w__7718, w__7719, w__7720;
  wire w__7721, w__7722, w__7723, w__7724, w__7725, w__7726, w__7727, w__7728;
  wire w__7729, w__7730, w__7731, w__7732, w__7733, w__7734, w__7735, w__7736;
  wire w__7737, w__7738, w__7739, w__7740, w__7741, w__7742, w__7743, w__7744;
  wire w__7745, w__7746, w__7747, w__7748, w__7749, w__7750, w__7751, w__7752;
  wire w__7753, w__7754, w__7755, w__7756, w__7757, w__7758, w__7759, w__7760;
  wire w__7761, w__7762, w__7763, w__7764, w__7765, w__7766, w__7767, w__7768;
  wire w__7769, w__7770, w__7771, w__7772, w__7773, w__7774, w__7775, w__7776;
  wire w__7777, w__7778, w__7779, w__7780, w__7781, w__7782, w__7783, w__7784;
  wire w__7785, w__7786, w__7787, w__7788, w__7789, w__7790, w__7791, w__7792;
  wire w__7793, w__7794, w__7795, w__7796, w__7797, w__7798, w__7799, w__7800;
  wire w__7801, w__7802, w__7803, w__7804, w__7805, w__7806, w__7807, w__7808;
  wire w__7809, w__7810, w__7811, w__7812, w__7813, w__7814, w__7815, w__7816;
  wire w__7817, w__7818, w__7819, w__7820, w__7821, w__7822, w__7823, w__7824;
  wire w__7825, w__7826, w__7827, w__7828, w__7829, w__7830, w__7831, w__7832;
  wire w__7833, w__7834, w__7835, w__7836, w__7837, w__7838, w__7839, w__7840;
  wire w__7841, w__7842, w__7843, w__7844, w__7845, w__7846, w__7847, w__7848;
  wire w__7849, w__7850, w__7851, w__7852, w__7853, w__7854, w__7855, w__7856;
  wire w__7857, w__7858, w__7859, w__7860, w__7861, w__7862, w__7863, w__7864;
  wire w__7865, w__7866, w__7867, w__7868, w__7869, w__7870, w__7871, w__7872;
  wire w__7873, w__7874, w__7875, w__7876, w__7877, w__7878, w__7879, w__7880;
  wire w__7881, w__7882, w__7883, w__7884, w__7885, w__7886, w__7887, w__7888;
  wire w__7889, w__7890, w__7891, w__7892, w__7893, w__7894, w__7895, w__7896;
  wire w__7897, w__7898, w__7899, w__7900, w__7901, w__7902, w__7903, w__7904;
  wire w__7905, w__7906, w__7907, w__7908, w__7909, w__7910, w__7911, w__7912;
  wire w__7913, w__7914, w__7915, w__7916, w__7917, w__7918, w__7919, w__7920;
  wire w__7921, w__7922, w__7923, w__7924, w__7925, w__7926, w__7927, w__7928;
  wire w__7929, w__7930, w__7931, w__7932, w__7933, w__7934, w__7935, w__7936;
  wire w__7937, w__7938, w__7939, w__7940, w__7941, w__7942, w__7943, w__7944;
  wire w__7945, w__7946, w__7947, w__7948, w__7949, w__7950, w__7951, w__7952;
  wire w__7953, w__7954, w__7955, w__7956, w__7957, w__7958, w__7959, w__7960;
  wire w__7961, w__7962, w__7963, w__7964, w__7965, w__7966, w__7967, w__7968;
  wire w__7969, w__7970, w__7971, w__7972, w__7973, w__7974, w__7975, w__7976;
  wire w__7977, w__7978, w__7979, w__7980, w__7981, w__7982, w__7983, w__7984;
  wire w__7985, w__7986, w__7987, w__7988, w__7989, w__7990, w__7991, w__7992;
  wire w__7993, w__7994, w__7995, w__7996, w__7997, w__7998, w__7999, w__8000;
  wire w__8001, w__8002, w__8003, w__8004, w__8005, w__8006, w__8007, w__8008;
  wire w__8009, w__8010, w__8011, w__8012, w__8013, w__8014, w__8015, w__8016;
  wire w__8017, w__8018, w__8019, w__8020, w__8021, w__8022, w__8023, w__8024;
  wire w__8025, w__8026, w__8027, w__8028, w__8029, w__8030, w__8031, w__8032;
  wire w__8033, w__8034, w__8035, w__8036, w__8037, w__8038, w__8039, w__8040;
  wire w__8041, w__8042, w__8043, w__8044, w__8045, w__8046, w__8047, w__8048;
  wire w__8049, w__8050, w__8051, w__8052, w__8053, w__8054, w__8055, w__8056;
  wire w__8057, w__8058, w__8059, w__8060, w__8061, w__8062, w__8063, w__8064;
  wire w__8065, w__8066, w__8067, w__8068, w__8069, w__8070, w__8071, w__8072;
  wire w__8073, w__8074, w__8075, w__8076, w__8077, w__8078, w__8079, w__8080;
  wire w__8081, w__8082, w__8083, w__8084, w__8085, w__8086, w__8087, w__8088;
  wire w__8089, w__8090, w__8091, w__8092, w__8093, w__8094, w__8095, w__8096;
  wire w__8097, w__8098, w__8099, w__8100, w__8101, w__8102, w__8103, w__8104;
  wire w__8105, w__8106, w__8107, w__8108, w__8109, w__8110, w__8111, w__8112;
  wire w__8113, w__8114, w__8115, w__8116, w__8117, w__8118, w__8119, w__8120;
  wire w__8121, w__8122, w__8123, w__8124, w__8125, w__8126, w__8127, w__8128;
  wire w__8129, w__8130, w__8131, w__8132, w__8133, w__8134, w__8135, w__8136;
  wire w__8137, w__8138, w__8139, w__8140, w__8141, w__8142, w__8143, w__8144;
  wire w__8145, w__8146, w__8147, w__8148, w__8149, w__8150, w__8151, w__8152;
  wire w__8153, w__8154, w__8155, w__8156, w__8157, w__8158, w__8159, w__8160;
  wire w__8161, w__8162, w__8163, w__8164, w__8165, w__8166, w__8167, w__8168;
  wire w__8169, w__8170, w__8171, w__8172, w__8173, w__8174, w__8175, w__8176;
  wire w__8177, w__8178, w__8179, w__8180, w__8181, w__8182, w__8183, w__8184;
  wire w__8185, w__8186, w__8187, w__8188, w__8189, w__8190, w__8191, w__8192;
  wire w__8193, w__8194, w__8195, w__8196, w__8197, w__8198, w__8199, w__8200;
  wire w__8201, w__8202, w__8203, w__8204, w__8205, w__8206, w__8207, w__8208;
  wire w__8209, w__8210, w__8211, w__8212, w__8213, w__8214, w__8215, w__8216;
  wire w__8217, w__8218, w__8219, w__8220, w__8221, w__8222, w__8223, w__8224;
  wire w__8225, w__8226, w__8227, w__8228, w__8229, w__8230, w__8231, w__8232;
  wire w__8233, w__8234, w__8235, w__8236, w__8237, w__8238, w__8239, w__8240;
  wire w__8241, w__8242, w__8243, w__8244, w__8245, w__8246, w__8247, w__8248;
  wire w__8249, w__8250, w__8251, w__8252, w__8253, w__8254, w__8255, w__8256;
  wire w__8257, w__8258, w__8259, w__8260, w__8261, w__8262, w__8263, w__8264;
  wire w__8265, w__8266, w__8267, w__8268, w__8269, w__8270, w__8271, w__8272;
  wire w__8273, w__8274, w__8275, w__8276, w__8277, w__8278, w__8279, w__8280;
  wire w__8281, w__8282, w__8283, w__8284, w__8285, w__8286, w__8287, w__8288;
  wire w__8289, w__8290, w__8291, w__8292, w__8293, w__8294, w__8295, w__8296;
  wire w__8297, w__8298, w__8299, w__8300, w__8301, w__8302, w__8303, w__8304;
  wire w__8305, w__8306, w__8307, w__8308, w__8309, w__8310, w__8311, w__8312;
  wire w__8313, w__8314, w__8315, w__8316, w__8317, w__8318, w__8319, w__8320;
  wire w__8321, w__8322, w__8323, w__8324, w__8325, w__8326, w__8327, w__8328;
  wire w__8329, w__8330, w__8331, w__8332, w__8333, w__8334, w__8335, w__8336;
  wire w__8337, w__8338, w__8339, w__8340, w__8341, w__8342, w__8343, w__8344;
  wire w__8345, w__8346, w__8347, w__8348, w__8349, w__8350, w__8351, w__8352;
  wire w__8353, w__8354, w__8355, w__8356, w__8357, w__8358, w__8359, w__8360;
  wire w__8361, w__8362, w__8363, w__8364, w__8365, w__8366, w__8367, w__8368;
  wire w__8369, w__8370, w__8371, w__8372, w__8373, w__8374, w__8375, w__8376;
  wire w__8377, w__8378, w__8379, w__8380, w__8381, w__8382, w__8383, w__8384;
  wire w__8385, w__8386, w__8387, w__8388, w__8389, w__8390, w__8391, w__8392;
  wire w__8393, w__8394, w__8395, w__8396, w__8397, w__8398, w__8399, w__8400;
  wire w__8401, w__8402, w__8403, w__8404, w__8405, w__8406, w__8407, w__8408;
  wire w__8409, w__8410, w__8411, w__8412, w__8413, w__8414, w__8415, w__8416;
  wire w__8417, w__8418, w__8419, w__8420, w__8421, w__8422, w__8423, w__8424;
  wire w__8425, w__8426, w__8427, w__8428, w__8429, w__8430, w__8431, w__8432;
  wire w__8433, w__8434, w__8435, w__8436, w__8437, w__8438, w__8439, w__8440;
  wire w__8441, w__8442, w__8443, w__8444, w__8445, w__8446, w__8447, w__8448;
  wire w__8449, w__8450, w__8451, w__8452, w__8453, w__8454, w__8455, w__8456;
  wire w__8457, w__8458, w__8459, w__8460, w__8461, w__8462, w__8463, w__8464;
  wire w__8465, w__8466, w__8467, w__8468, w__8469, w__8470, w__8471, w__8472;
  wire w__8473, w__8474, w__8475, w__8476, w__8477, w__8478, w__8479, w__8480;
  wire w__8481, w__8482, w__8483, w__8484, w__8485, w__8486, w__8487, w__8488;
  wire w__8489, w__8490, w__8491, w__8492, w__8493, w__8494, w__8495, w__8496;
  wire w__8497, w__8498, w__8499, w__8500, w__8501, w__8502, w__8503, w__8504;
  wire w__8505, w__8506, w__8507, w__8508, w__8509, w__8510, w__8511, w__8512;
  wire w__8513, w__8514, w__8515, w__8516, w__8517, w__8518, w__8519, w__8520;
  wire w__8521, w__8522, w__8523, w__8524, w__8525, w__8526, w__8527, w__8528;
  wire w__8529, w__8530, w__8531, w__8532;
  or g__1(w__8532 ,w__831 ,w__1063);
  xnor g__2(w__8531 ,w__1062 ,w__848);
  and g__3(w__1063 ,w__830 ,w__1062);
  or g__4(w__1062 ,w__903 ,w__1061);
  xnor g__5(w__8530 ,w__1060 ,w__913);
  and g__6(w__1061 ,w__904 ,w__1060);
  or g__7(w__1060 ,w__954 ,w__1059);
  xnor g__8(w__8529 ,w__1058 ,w__966);
  and g__9(w__1059 ,w__961 ,w__1058);
  or g__10(w__1058 ,w__980 ,w__1057);
  xnor g__11(w__8528 ,w__1056 ,w__991);
  and g__12(w__1057 ,w__969 ,w__1056);
  or g__13(w__1056 ,w__994 ,w__1055);
  xnor g__14(w__8527 ,w__1054 ,w__1008);
  and g__15(w__1055 ,w__1003 ,w__1054);
  or g__16(w__1054 ,w__1026 ,w__1053);
  xnor g__17(w__8526 ,w__1052 ,w__1032);
  nor g__18(w__1053 ,w__1027 ,w__1052);
  and g__19(w__1052 ,w__1051 ,w__1028);
  or g__20(w__1051 ,w__1020 ,w__1050);
  and g__21(w__1050 ,w__1036 ,w__1049);
  or g__22(w__1049 ,w__1035 ,w__1048);
  and g__23(w__1048 ,w__1047 ,w__1037);
  or g__24(w__1047 ,w__1034 ,w__1046);
  and g__25(w__1046 ,w__1025 ,w__1045);
  or g__26(w__1045 ,w__1024 ,w__1044);
  and g__27(w__1044 ,w__1013 ,w__1043);
  or g__28(w__1043 ,w__1014 ,w__1042);
  and g__29(w__1042 ,w__998 ,w__1041);
  xnor g__30(w__8520 ,w__1040 ,w__1007);
  or g__31(w__1041 ,w__992 ,w__1040);
  and g__32(w__1040 ,w__970 ,w__1033);
  xnor g__33(w__1039 ,w__1021 ,w__1016);
  xnor g__34(w__1038 ,w__1022 ,w__1029);
  or g__35(w__1037 ,w__1016 ,w__1021);
  or g__36(w__1036 ,w__1029 ,w__1022);
  and g__37(w__1035 ,w__1029 ,w__1022);
  and g__38(w__1034 ,w__1016 ,w__1021);
  or g__39(w__1033 ,w__971 ,w__1023);
  xnor g__40(w__1032 ,w__1018 ,w__996);
  xnor g__41(w__1031 ,w__1012 ,w__1017);
  xnor g__42(w__1030 ,w__1005 ,w__1011);
  or g__43(w__1028 ,w__1017 ,w__1012);
  and g__44(w__1027 ,w__1018 ,w__997);
  nor g__45(w__1026 ,w__1018 ,w__997);
  or g__46(w__1025 ,w__1004 ,w__1010);
  nor g__47(w__1024 ,w__1005 ,w__1011);
  and g__48(w__1029 ,w__1002 ,w__1015);
  and g__49(w__1020 ,w__1017 ,w__1012);
  xnor g__50(w__8518 ,w__1006 ,w__967);
  xnor g__51(w__1019 ,w__995 ,w__986);
  and g__52(w__1023 ,w__941 ,w__1009);
  xnor g__53(w__1022 ,w__948 ,w__989);
  xnor g__54(w__1021 ,w__985 ,w__990);
  or g__55(w__1015 ,w__950 ,w__1001);
  and g__56(w__1014 ,w__986 ,w__995);
  or g__57(w__1013 ,w__986 ,w__995);
  and g__58(w__1018 ,w__956 ,w__999);
  and g__59(w__1017 ,w__982 ,w__993);
  and g__60(w__1016 ,w__981 ,w__1000);
  not g__61(w__1010 ,w__1011);
  or g__62(w__1009 ,w__955 ,w__1006);
  xnor g__63(w__8517 ,w__947 ,w__965);
  xnor g__64(w__1008 ,w__973 ,w__975);
  xnor g__65(w__1007 ,w__944 ,w__976);
  xnor g__66(w__1012 ,w__987 ,w__968);
  xnor g__67(w__1011 ,w__943 ,w__964);
  not g__68(w__1004 ,w__1005);
  or g__69(w__1003 ,w__974 ,w__972);
  or g__70(w__1002 ,w__916 ,w__985);
  and g__71(w__1001 ,w__916 ,w__985);
  or g__72(w__1000 ,w__938 ,w__979);
  or g__73(w__999 ,w__987 ,w__953);
  or g__74(w__998 ,w__944 ,w__977);
  and g__75(w__1006 ,w__960 ,w__984);
  or g__76(w__1005 ,w__929 ,w__978);
  not g__77(w__997 ,w__996);
  nor g__78(w__994 ,w__975 ,w__973);
  or g__79(w__993 ,w__948 ,w__983);
  and g__80(w__992 ,w__944 ,w__977);
  xnor g__81(w__991 ,w__963 ,w__917);
  xnor g__82(w__990 ,w__950 ,w__916);
  xnor g__83(w__989 ,w__946 ,w__890);
  xnor g__84(w__988 ,w__945 ,w__936);
  xnor g__85(w__996 ,w__937 ,w__939);
  xnor g__86(w__995 ,w__949 ,w__940);
  or g__87(w__984 ,w__959 ,w__947);
  and g__88(w__983 ,w__890 ,w__946);
  or g__89(w__982 ,w__890 ,w__946);
  or g__90(w__981 ,w__874 ,w__942);
  nor g__91(w__980 ,w__222 ,w__963);
  nor g__92(w__979 ,w__873 ,w__943);
  and g__93(w__978 ,w__926 ,w__949);
  and g__94(w__987 ,w__927 ,w__952);
  and g__95(w__986 ,w__898 ,w__951);
  and g__96(w__985 ,w__932 ,w__957);
  not g__97(w__977 ,w__976);
  not g__98(w__975 ,w__974);
  not g__99(w__972 ,w__973);
  and g__100(w__971 ,w__936 ,w__945);
  or g__101(w__970 ,w__936 ,w__945);
  or g__102(w__969 ,w__224 ,w__962);
  xnor g__103(w__968 ,w__924 ,w__905);
  xnor g__104(w__967 ,w__889 ,w__923);
  xnor g__105(w__966 ,w__919 ,w__858);
  xnor g__106(w__965 ,w__784 ,w__921);
  xnor g__107(w__964 ,w__938 ,w__874);
  xnor g__108(w__976 ,w__925 ,w__911);
  xnor g__109(w__974 ,w__908 ,w__912);
  and g__110(w__973 ,w__914 ,w__958);
  not g__111(w__963 ,w__962);
  or g__112(w__961 ,w__857 ,w__918);
  or g__113(w__960 ,w__783 ,w__921);
  nor g__114(w__959 ,w__784 ,w__920);
  or g__115(w__958 ,w__934 ,w__937);
  or g__116(w__957 ,w__798 ,w__931);
  or g__117(w__956 ,w__905 ,w__924);
  nor g__118(w__955 ,w__888 ,w__923);
  nor g__119(w__954 ,w__858 ,w__919);
  and g__120(w__953 ,w__905 ,w__924);
  or g__121(w__952 ,w__791 ,w__930);
  or g__122(w__951 ,w__902 ,w__925);
  or g__123(w__962 ,w__899 ,w__928);
  not g__124(w__942 ,w__943);
  xnor g__125(w__8516 ,w__909 ,w__882);
  or g__126(w__941 ,w__889 ,w__922);
  xnor g__127(w__940 ,w__856 ,w__907);
  xnor g__128(w__939 ,w__840 ,w__895);
  xnor g__129(w__950 ,w__910 ,w__880);
  xnor g__130(w__949 ,w__787 ,w__883);
  and g__131(w__948 ,w__852 ,w__935);
  and g__132(w__947 ,w__871 ,w__915);
  xnor g__133(w__946 ,w__893 ,w__885);
  xnor g__134(w__945 ,w__896 ,w__884);
  and g__135(w__944 ,w__867 ,w__933);
  xnor g__136(w__943 ,w__892 ,w__881);
  or g__137(w__935 ,w__872 ,w__910);
  nor g__138(w__934 ,w__839 ,w__895);
  or g__139(w__933 ,w__850 ,w__896);
  or g__140(w__932 ,w__820 ,w__891);
  nor g__141(w__931 ,w__819 ,w__892);
  and g__142(w__930 ,w__815 ,w__893);
  nor g__143(w__929 ,w__855 ,w__907);
  nor g__144(w__928 ,w__897 ,w__908);
  or g__145(w__927 ,w__815 ,w__893);
  or g__146(w__926 ,w__856 ,w__906);
  and g__147(w__938 ,w__863 ,w__901);
  and g__148(w__937 ,w__866 ,w__900);
  and g__149(w__936 ,w__854 ,w__887);
  not g__150(w__922 ,w__923);
  not g__151(w__920 ,w__921);
  not g__152(w__918 ,w__919);
  or g__153(w__915 ,w__870 ,w__909);
  or g__154(w__914 ,w__840 ,w__894);
  xnor g__155(w__8515 ,w__821 ,w__846);
  xnor g__156(w__913 ,w__878 ,w__771);
  xnor g__157(w__912 ,w__735 ,w__859);
  xnor g__158(w__911 ,w__876 ,w__814);
  xnor g__159(w__925 ,w__792 ,w__844);
  xnor g__160(w__924 ,w__818 ,w__842);
  xnor g__161(w__923 ,w__809 ,w__845);
  xnor g__162(w__921 ,w__719 ,w__841);
  and g__163(w__919 ,w__824 ,w__886);
  xnor g__164(w__917 ,w__879 ,w__843);
  xnor g__165(w__916 ,w__767 ,w__847);
  not g__166(w__906 ,w__907);
  or g__167(w__904 ,w__223 ,w__877);
  nor g__168(w__903 ,w__221 ,w__878);
  nor g__169(w__902 ,w__875 ,w__814);
  or g__170(w__901 ,w__793 ,w__861);
  or g__171(w__900 ,w__797 ,w__864);
  nor g__172(w__899 ,w__736 ,w__859);
  or g__173(w__898 ,w__876 ,w__813);
  and g__174(w__897 ,w__736 ,w__859);
  and g__175(w__910 ,w__837 ,w__868);
  and g__176(w__909 ,w__836 ,w__869);
  and g__177(w__908 ,w__823 ,w__865);
  and g__178(w__907 ,w__827 ,w__860);
  and g__179(w__905 ,w__838 ,w__862);
  not g__180(w__895 ,w__894);
  not g__181(w__891 ,w__892);
  not g__182(w__888 ,w__889);
  or g__183(w__887 ,w__790 ,w__853);
  or g__184(w__886 ,w__879 ,w__828);
  xnor g__185(w__885 ,w__815 ,w__791);
  xnor g__186(w__884 ,w__812 ,w__785);
  xnor g__187(w__883 ,w__817 ,w__793);
  xnor g__188(w__882 ,w__756 ,w__811);
  xnor g__189(w__881 ,w__820 ,w__798);
  xnor g__190(w__880 ,w__808 ,w__778);
  xnor g__191(w__896 ,w__738 ,w__802);
  xnor g__192(w__894 ,w__768 ,w__799);
  xnor g__193(w__893 ,w__772 ,w__801);
  xnor g__194(w__892 ,w__777 ,w__800);
  and g__195(w__890 ,w__829 ,w__849);
  and g__196(w__889 ,w__803 ,w__851);
  not g__197(w__877 ,w__878);
  not g__198(w__875 ,w__876);
  not g__199(w__873 ,w__874);
  and g__200(w__872 ,w__778 ,w__808);
  or g__201(w__871 ,w__756 ,w__810);
  nor g__202(w__870 ,w__755 ,w__811);
  or g__203(w__869 ,w__835 ,w__821);
  or g__204(w__868 ,w__760 ,w__834);
  or g__205(w__867 ,w__785 ,w__812);
  or g__206(w__866 ,w__769 ,w__818);
  or g__207(w__865 ,w__739 ,w__805);
  and g__208(w__864 ,w__769 ,w__818);
  or g__209(w__863 ,w__786 ,w__817);
  or g__210(w__862 ,w__759 ,w__826);
  nor g__211(w__861 ,w__787 ,w__816);
  or g__212(w__860 ,w__792 ,w__825);
  and g__213(w__879 ,w__754 ,w__833);
  and g__214(w__878 ,w__750 ,w__807);
  and g__215(w__876 ,w__780 ,w__822);
  and g__216(w__874 ,w__702 ,w__832);
  not g__217(w__858 ,w__857);
  not g__218(w__856 ,w__855);
  xnor g__219(w__8514 ,w__758 ,w__763);
  or g__220(w__854 ,w__774 ,w__809);
  and g__221(w__853 ,w__774 ,w__809);
  or g__222(w__852 ,w__778 ,w__808);
  or g__223(w__851 ,w__719 ,w__804);
  and g__224(w__850 ,w__785 ,w__812);
  or g__225(w__849 ,w__796 ,w__806);
  xnor g__226(w__848 ,w__789 ,w__544);
  xnor g__227(w__847 ,w__796 ,w__652);
  xnor g__228(w__846 ,w__651 ,w__776);
  xnor g__229(w__845 ,w__790 ,w__773);
  xnor g__230(w__844 ,w__770 ,w__715);
  xnor g__231(w__843 ,w__766 ,w__716);
  xnor g__232(w__842 ,w__769 ,w__797);
  xnor g__233(w__841 ,w__765 ,w__597);
  xnor g__234(w__859 ,w__795 ,w__761);
  xnor g__235(w__857 ,w__794 ,w__762);
  xnor g__236(w__855 ,w__779 ,w__729);
  not g__237(w__839 ,w__840);
  or g__238(w__838 ,w__585 ,w__772);
  or g__239(w__837 ,w__683 ,w__777);
  or g__240(w__836 ,w__650 ,w__776);
  nor g__241(w__835 ,w__651 ,w__775);
  and g__242(w__834 ,w__683 ,w__777);
  or g__243(w__833 ,w__743 ,w__795);
  or g__244(w__832 ,w__701 ,w__779);
  nor g__245(w__831 ,w__544 ,w__789);
  or g__246(w__830 ,w__543 ,w__788);
  or g__247(w__829 ,w__652 ,w__767);
  and g__248(w__828 ,w__716 ,w__766);
  or g__249(w__827 ,w__715 ,w__770);
  and g__250(w__826 ,w__585 ,w__772);
  and g__251(w__825 ,w__715 ,w__770);
  or g__252(w__824 ,w__716 ,w__766);
  or g__253(w__823 ,w__682 ,w__768);
  or g__254(w__822 ,w__738 ,w__781);
  and g__255(w__840 ,w__714 ,w__782);
  not g__256(w__819 ,w__820);
  not g__257(w__816 ,w__817);
  not g__258(w__813 ,w__814);
  not g__259(w__810 ,w__811);
  or g__260(w__807 ,w__751 ,w__794);
  and g__261(w__806 ,w__652 ,w__767);
  and g__262(w__805 ,w__682 ,w__768);
  and g__263(w__804 ,w__597 ,w__765);
  or g__264(w__803 ,w__597 ,w__765);
  xnor g__265(w__802 ,w__737 ,w__579);
  xnor g__266(w__801 ,w__759 ,w__585);
  xor g__267(w__800 ,w__760 ,w__683);
  xnor g__268(w__799 ,w__739 ,w__682);
  and g__269(w__821 ,w__747 ,w__764);
  xnor g__270(w__820 ,w__608 ,w__724);
  xnor g__271(w__818 ,w__757 ,w__726);
  xnor g__272(w__817 ,w__598 ,w__725);
  xnor g__273(w__815 ,w__610 ,w__723);
  xnor g__274(w__814 ,w__686 ,w__721);
  xnor g__275(w__812 ,w__616 ,w__720);
  xnor g__276(w__811 ,w__688 ,w__727);
  xnor g__277(w__809 ,w__655 ,w__722);
  xnor g__278(w__808 ,w__614 ,w__728);
  not g__279(w__788 ,w__789);
  not g__280(w__787 ,w__786);
  not g__281(w__784 ,w__783);
  or g__282(w__782 ,w__757 ,w__706);
  and g__283(w__781 ,w__579 ,w__737);
  or g__284(w__780 ,w__579 ,w__737);
  and g__285(w__798 ,w__704 ,w__742);
  and g__286(w__797 ,w__703 ,w__740);
  and g__287(w__796 ,w__672 ,w__730);
  and g__288(w__795 ,w__705 ,w__741);
  and g__289(w__794 ,w__694 ,w__744);
  and g__290(w__793 ,w__695 ,w__749);
  and g__291(w__792 ,w__690 ,w__734);
  and g__292(w__791 ,w__678 ,w__733);
  and g__293(w__790 ,w__671 ,w__732);
  and g__294(w__789 ,w__635 ,w__746);
  and g__295(w__786 ,w__699 ,w__748);
  and g__296(w__785 ,w__675 ,w__731);
  and g__297(w__783 ,w__713 ,w__752);
  not g__298(w__775 ,w__776);
  not g__299(w__774 ,w__773);
  or g__300(w__764 ,w__758 ,w__745);
  xnor g__301(w__763 ,w__612 ,w__681);
  xnor g__302(w__762 ,w__542 ,w__685);
  xnor g__303(w__761 ,w__717 ,w__607);
  xnor g__304(w__779 ,w__588 ,w__659);
  and g__305(w__778 ,w__668 ,w__753);
  xnor g__306(w__777 ,w__615 ,w__664);
  xnor g__307(w__776 ,w__623 ,w__663);
  xnor g__308(w__773 ,w__625 ,w__665);
  xnor g__309(w__772 ,w__592 ,w__667);
  xnor g__310(w__771 ,w__718 ,w__657);
  xnor g__311(w__770 ,w__617 ,w__656);
  xnor g__312(w__769 ,w__545 ,w__662);
  xnor g__313(w__768 ,w__602 ,w__658);
  xnor g__314(w__767 ,w__589 ,w__660);
  xnor g__315(w__766 ,w__599 ,w__661);
  xnor g__316(w__765 ,w__600 ,w__666);
  not g__317(w__755 ,w__756);
  or g__318(w__754 ,w__607 ,w__717);
  or g__319(w__753 ,w__595 ,w__711);
  or g__320(w__752 ,w__712 ,w__689);
  nor g__321(w__751 ,w__542 ,w__684);
  or g__322(w__750 ,w__541 ,w__685);
  or g__323(w__749 ,w__586 ,w__693);
  or g__324(w__748 ,w__687 ,w__697);
  or g__325(w__747 ,w__612 ,w__680);
  or g__326(w__746 ,w__638 ,w__718);
  nor g__327(w__745 ,w__611 ,w__681);
  or g__328(w__744 ,w__593 ,w__696);
  and g__329(w__743 ,w__607 ,w__717);
  or g__330(w__742 ,w__594 ,w__679);
  or g__331(w__741 ,w__590 ,w__698);
  or g__332(w__740 ,w__591 ,w__700);
  and g__333(w__760 ,w__644 ,w__709);
  and g__334(w__759 ,w__639 ,w__692);
  and g__335(w__758 ,w__575 ,w__708);
  and g__336(w__757 ,w__645 ,w__707);
  and g__337(w__756 ,w__646 ,w__710);
  not g__338(w__736 ,w__735);
  or g__339(w__734 ,w__624 ,w__691);
  xnor g__340(w__8513 ,w__653 ,w__626);
  or g__341(w__733 ,w__622 ,w__676);
  or g__342(w__732 ,w__570 ,w__670);
  or g__343(w__731 ,w__655 ,w__673);
  or g__344(w__730 ,w__571 ,w__669);
  xnor g__345(w__729 ,w__620 ,w__647);
  xnor g__346(w__728 ,w__622 ,w__613);
  xnor g__347(w__727 ,w__649 ,w__603);
  xnor g__348(w__726 ,w__604 ,w__648);
  xnor g__349(w__725 ,w__609 ,w__594);
  xnor g__350(w__724 ,w__601 ,w__571);
  xnor g__351(w__723 ,w__621 ,w__591);
  xnor g__352(w__722 ,w__605 ,w__606);
  xnor g__353(w__721 ,w__618 ,w__619);
  xnor g__354(w__720 ,w__624 ,w__582);
  and g__355(w__739 ,w__631 ,w__674);
  and g__356(w__738 ,w__634 ,w__677);
  xnor g__357(w__737 ,w__587 ,w__596);
  xnor g__358(w__735 ,w__569 ,w__627);
  or g__359(w__714 ,w__648 ,w__604);
  or g__360(w__713 ,w__603 ,w__649);
  and g__361(w__712 ,w__603 ,w__649);
  and g__362(w__711 ,w__562 ,w__615);
  or g__363(w__710 ,w__641 ,w__623);
  or g__364(w__709 ,w__588 ,w__642);
  or g__365(w__708 ,w__552 ,w__654);
  or g__366(w__707 ,w__592 ,w__640);
  and g__367(w__706 ,w__648 ,w__604);
  or g__368(w__705 ,w__580 ,w__602);
  or g__369(w__704 ,w__598 ,w__609);
  or g__370(w__703 ,w__610 ,w__621);
  or g__371(w__702 ,w__647 ,w__620);
  and g__372(w__701 ,w__647 ,w__620);
  and g__373(w__700 ,w__610 ,w__621);
  or g__374(w__699 ,w__619 ,w__618);
  and g__375(w__698 ,w__580 ,w__602);
  and g__376(w__697 ,w__619 ,w__618);
  and g__377(w__696 ,w__558 ,w__599);
  or g__378(w__695 ,w__583 ,w__617);
  or g__379(w__694 ,w__558 ,w__599);
  and g__380(w__693 ,w__583 ,w__617);
  or g__381(w__692 ,w__589 ,w__636);
  and g__382(w__691 ,w__582 ,w__616);
  or g__383(w__690 ,w__582 ,w__616);
  and g__384(w__719 ,w__503 ,w__630);
  and g__385(w__718 ,w__393 ,w__629);
  and g__386(w__717 ,w__402 ,w__643);
  and g__387(w__716 ,w__553 ,w__633);
  and g__388(w__715 ,w__574 ,w__637);
  not g__389(w__689 ,w__688);
  not g__390(w__687 ,w__686);
  not g__391(w__684 ,w__685);
  not g__392(w__680 ,w__681);
  and g__393(w__679 ,w__598 ,w__609);
  or g__394(w__678 ,w__613 ,w__614);
  or g__395(w__677 ,w__632 ,w__625);
  and g__396(w__676 ,w__613 ,w__614);
  or g__397(w__675 ,w__606 ,w__605);
  or g__398(w__674 ,w__545 ,w__628);
  and g__399(w__673 ,w__606 ,w__605);
  or g__400(w__672 ,w__608 ,w__601);
  or g__401(w__671 ,w__561 ,w__600);
  and g__402(w__670 ,w__561 ,w__600);
  and g__403(w__669 ,w__608 ,w__601);
  or g__404(w__668 ,w__562 ,w__615);
  xnor g__405(w__667 ,w__337 ,w__560);
  xnor g__406(w__666 ,w__570 ,w__561);
  xnor g__407(w__665 ,w__466 ,w__556);
  xnor g__408(w__664 ,w__562 ,w__595);
  xnor g__409(w__663 ,w__578 ,w__3);
  xnor g__410(w__662 ,w__559 ,w__563);
  xnor g__411(w__661 ,w__558 ,w__593);
  xnor g__412(w__660 ,w__584 ,w__581);
  xnor g__413(w__659 ,w__554 ,w__4);
  xnor g__414(w__658 ,w__590 ,w__580);
  xnor g__415(w__657 ,w__251 ,w__557);
  xnor g__416(w__656 ,w__583 ,w__586);
  xnor g__417(w__688 ,w__567 ,w__546);
  xnor g__418(w__686 ,w__467 ,w__547);
  xnor g__419(w__685 ,w__568 ,w__478);
  xor g__420(w__683 ,w__421 ,w__549);
  xnor g__421(w__682 ,w__564 ,w__470);
  xnor g__422(w__681 ,w__420 ,w__548);
  not g__423(w__654 ,w__653);
  not g__424(w__650 ,w__651);
  or g__425(w__646 ,w__3 ,w__578);
  or g__426(w__645 ,w__337 ,w__560);
  or g__427(w__644 ,w__4 ,w__554);
  or g__428(w__643 ,w__439 ,w__564);
  and g__429(w__642 ,w__4 ,w__554);
  and g__430(w__641 ,w__3 ,w__578);
  and g__431(w__640 ,w__337 ,w__560);
  or g__432(w__639 ,w__581 ,w__584);
  and g__433(w__638 ,w__251 ,w__557);
  or g__434(w__637 ,w__587 ,w__572);
  and g__435(w__636 ,w__581 ,w__584);
  or g__436(w__635 ,w__251 ,w__557);
  or g__437(w__634 ,w__465 ,w__556);
  or g__438(w__633 ,w__550 ,w__569);
  nor g__439(w__632 ,w__466 ,w__555);
  or g__440(w__631 ,w__563 ,w__559);
  or g__441(w__630 ,w__535 ,w__567);
  or g__442(w__629 ,w__427 ,w__568);
  and g__443(w__628 ,w__563 ,w__559);
  xnor g__444(w__627 ,w__253 ,w__539);
  xnor g__445(w__626 ,w__2 ,w__540);
  and g__446(w__655 ,w__395 ,w__551);
  and g__447(w__653 ,w__308 ,w__566);
  and g__448(w__652 ,w__526 ,w__577);
  or g__449(w__651 ,w__532 ,w__576);
  xnor g__450(w__649 ,w__323 ,w__498);
  xnor g__451(w__648 ,w__378 ,w__492);
  and g__452(w__647 ,w__524 ,w__573);
  not g__453(w__611 ,w__612);
  xnor g__454(w__596 ,w__275 ,w__5);
  xnor g__455(w__625 ,w__355 ,w__469);
  xnor g__456(w__624 ,w__296 ,w__473);
  xnor g__457(w__623 ,w__365 ,w__471);
  xnor g__458(w__622 ,w__360 ,w__482);
  xnor g__459(w__621 ,w__333 ,w__484);
  xnor g__460(w__620 ,w__298 ,w__483);
  xnor g__461(w__619 ,w__366 ,w__481);
  xnor g__462(w__618 ,w__361 ,w__479);
  xnor g__463(w__617 ,w__356 ,w__475);
  xnor g__464(w__616 ,w__342 ,w__500);
  xnor g__465(w__615 ,w__369 ,w__490);
  xnor g__466(w__614 ,w__282 ,w__487);
  xnor g__467(w__613 ,w__297 ,w__491);
  xnor g__468(w__612 ,w__256 ,w__495);
  xnor g__469(w__610 ,w__262 ,w__486);
  xnor g__470(w__609 ,w__285 ,w__488);
  xnor g__471(w__608 ,w__301 ,w__472);
  xnor g__472(w__607 ,w__302 ,w__493);
  xnor g__473(w__606 ,w__295 ,w__477);
  xnor g__474(w__605 ,w__423 ,w__496);
  xnor g__475(w__604 ,w__354 ,w__497);
  xnor g__476(w__603 ,w__377 ,w__480);
  xnor g__477(w__602 ,w__368 ,w__485);
  xnor g__478(w__601 ,w__364 ,w__474);
  xnor g__479(w__600 ,w__255 ,w__489);
  xnor g__480(w__599 ,w__299 ,w__476);
  xnor g__481(w__598 ,w__367 ,w__499);
  xnor g__482(w__597 ,w__1 ,w__494);
  or g__483(w__577 ,w__422 ,w__504);
  and g__484(w__576 ,w__420 ,w__501);
  or g__485(w__575 ,w__540 ,w__2);
  or g__486(w__574 ,w__275 ,w__5);
  or g__487(w__573 ,w__468 ,w__523);
  and g__488(w__572 ,w__275 ,w__5);
  and g__489(w__595 ,w__449 ,w__536);
  and g__490(w__594 ,w__388 ,w__527);
  and g__491(w__593 ,w__445 ,w__519);
  and g__492(w__592 ,w__460 ,w__525);
  and g__493(w__591 ,w__390 ,w__522);
  and g__494(w__590 ,w__399 ,w__537);
  and g__495(w__589 ,w__447 ,w__511);
  and g__496(w__588 ,w__450 ,w__531);
  and g__497(w__587 ,w__408 ,w__510);
  and g__498(w__586 ,w__428 ,w__513);
  and g__499(w__585 ,w__433 ,w__518);
  and g__500(w__584 ,w__425 ,w__512);
  and g__501(w__583 ,w__440 ,w__515);
  and g__502(w__582 ,w__456 ,w__509);
  and g__503(w__581 ,w__429 ,w__514);
  and g__504(w__580 ,w__385 ,w__505);
  and g__505(w__579 ,w__409 ,w__508);
  and g__506(w__578 ,w__400 ,w__534);
  not g__507(w__566 ,w__565);
  not g__508(w__555 ,w__556);
  or g__509(w__553 ,w__253 ,w__538);
  and g__510(w__552 ,w__540 ,w__2);
  or g__511(w__551 ,w__455 ,w__1);
  nor g__512(w__550 ,w__252 ,w__539);
  xnor g__513(w__549 ,w__344 ,w__419);
  xnor g__514(w__548 ,w__264 ,w__415);
  xnor g__515(w__547 ,w__283 ,w__416);
  xnor g__516(w__546 ,w__464 ,w__418);
  and g__517(w__571 ,w__451 ,w__530);
  and g__518(w__570 ,w__386 ,w__516);
  and g__519(w__569 ,w__413 ,w__507);
  and g__520(w__568 ,w__446 ,w__528);
  and g__521(w__567 ,w__391 ,w__502);
  xnor g__522(w__565 ,w__353 ,w__379);
  xnor g__523(w__564 ,w__370 ,w__383);
  and g__524(w__563 ,w__406 ,w__517);
  and g__525(w__562 ,w__384 ,w__520);
  and g__526(w__561 ,w__443 ,w__529);
  xnor g__527(w__560 ,w__291 ,w__382);
  and g__528(w__559 ,w__430 ,w__521);
  xnor g__529(w__558 ,w__300 ,w__381);
  xnor g__530(w__557 ,w__303 ,w__380);
  and g__531(w__556 ,w__405 ,w__533);
  and g__532(w__554 ,w__404 ,w__506);
  not g__533(w__544 ,w__543);
  not g__534(w__541 ,w__542);
  not g__535(w__538 ,w__539);
  or g__536(w__537 ,w__354 ,w__392);
  or g__537(w__536 ,w__305 ,w__448);
  nor g__538(w__535 ,w__464 ,w__417);
  or g__539(w__534 ,w__293 ,w__412);
  or g__540(w__533 ,w__294 ,w__438);
  nor g__541(w__532 ,w__264 ,w__415);
  or g__542(w__531 ,w__361 ,w__453);
  or g__543(w__530 ,w__298 ,w__442);
  or g__544(w__529 ,w__377 ,w__387);
  or g__545(w__528 ,w__299 ,w__459);
  or g__546(w__527 ,w__356 ,w__435);
  or g__547(w__526 ,w__344 ,w__419);
  or g__548(w__525 ,w__297 ,w__444);
  or g__549(w__524 ,w__283 ,w__416);
  and g__550(w__523 ,w__283 ,w__416);
  or g__551(w__522 ,w__306 ,w__434);
  or g__552(w__521 ,w__292 ,w__462);
  or g__553(w__520 ,w__367 ,w__437);
  or g__554(w__519 ,w__302 ,w__458);
  or g__555(w__518 ,w__360 ,w__441);
  or g__556(w__517 ,w__359 ,w__394);
  or g__557(w__516 ,w__307 ,w__407);
  or g__558(w__515 ,w__296 ,w__452);
  or g__559(w__514 ,w__301 ,w__389);
  or g__560(w__513 ,w__310 ,w__401);
  or g__561(w__512 ,w__364 ,w__397);
  or g__562(w__511 ,w__369 ,w__431);
  or g__563(w__510 ,w__355 ,w__436);
  or g__564(w__509 ,w__295 ,w__454);
  or g__565(w__508 ,w__457 ,w__423);
  or g__566(w__507 ,w__368 ,w__426);
  or g__567(w__506 ,w__366 ,w__411);
  or g__568(w__505 ,w__378 ,w__424);
  and g__569(w__504 ,w__344 ,w__419);
  and g__570(w__545 ,w__248 ,w__396);
  or g__571(w__543 ,w__249 ,w__410);
  or g__572(w__542 ,w__311 ,w__398);
  and g__573(w__540 ,w__316 ,w__432);
  or g__574(w__539 ,w__250 ,w__403);
  or g__575(w__503 ,w__418 ,w__463);
  or g__576(w__502 ,w__365 ,w__461);
  or g__577(w__501 ,w__263 ,w__414);
  xnor g__578(w__500 ,w__274 ,w__310);
  xnor g__579(w__499 ,w__269 ,w__279);
  xnor g__580(w__498 ,w__334 ,w__307);
  xnor g__581(w__497 ,w__326 ,w__267);
  xnor g__582(w__496 ,w__320 ,w__284);
  xnor g__583(w__495 ,w__277 ,w__293);
  xnor g__584(w__494 ,w__328 ,w__338);
  xnor g__585(w__493 ,w__276 ,w__260);
  xnor g__586(w__492 ,w__339 ,w__325);
  xnor g__587(w__491 ,w__322 ,w__336);
  xnor g__588(w__490 ,w__273 ,w__281);
  xnor g__589(w__489 ,w__329 ,w__294);
  xnor g__590(w__488 ,w__317 ,w__305);
  xnor g__591(w__487 ,w__319 ,w__306);
  xnor g__592(w__486 ,w__346 ,w__292);
  xnor g__593(w__485 ,w__261 ,w__335);
  xnor g__594(w__484 ,w__352 ,w__359);
  xnor g__595(w__483 ,w__265 ,w__332);
  xnor g__596(w__482 ,w__268 ,w__271);
  xnor g__597(w__481 ,w__278 ,w__343);
  xnor g__598(w__480 ,w__258 ,w__327);
  xnor g__599(w__479 ,w__270 ,w__259);
  xnor g__600(w__478 ,w__266 ,w__330);
  xnor g__601(w__477 ,w__321 ,w__351);
  xnor g__602(w__476 ,w__272 ,w__347);
  xnor g__603(w__475 ,w__349 ,w__257);
  xnor g__604(w__474 ,w__280 ,w__331);
  xnor g__605(w__473 ,w__324 ,w__348);
  xnor g__606(w__472 ,w__254 ,w__318);
  xnor g__607(w__471 ,w__340 ,w__287);
  xnor g__608(w__470 ,w__345 ,w__286);
  xnor g__609(w__469 ,w__350 ,w__341);
  not g__610(w__468 ,w__467);
  not g__611(w__465 ,w__466);
  not g__612(w__463 ,w__464);
  and g__613(w__462 ,w__262 ,w__346);
  and g__614(w__461 ,w__340 ,w__287);
  or g__615(w__460 ,w__322 ,w__336);
  and g__616(w__459 ,w__272 ,w__347);
  and g__617(w__458 ,w__276 ,w__260);
  and g__618(w__457 ,w__320 ,w__284);
  or g__619(w__456 ,w__321 ,w__351);
  and g__620(w__455 ,w__328 ,w__338);
  and g__621(w__454 ,w__321 ,w__351);
  and g__622(w__453 ,w__270 ,w__259);
  and g__623(w__452 ,w__324 ,w__348);
  or g__624(w__451 ,w__265 ,w__332);
  or g__625(w__450 ,w__270 ,w__259);
  or g__626(w__449 ,w__285 ,w__317);
  and g__627(w__448 ,w__285 ,w__317);
  or g__628(w__447 ,w__273 ,w__281);
  or g__629(w__446 ,w__272 ,w__347);
  or g__630(w__445 ,w__276 ,w__260);
  and g__631(w__444 ,w__322 ,w__336);
  or g__632(w__443 ,w__258 ,w__327);
  and g__633(w__442 ,w__265 ,w__332);
  and g__634(w__441 ,w__268 ,w__271);
  or g__635(w__440 ,w__324 ,w__348);
  and g__636(w__439 ,w__345 ,w__286);
  and g__637(w__438 ,w__255 ,w__329);
  and g__638(w__437 ,w__269 ,w__279);
  and g__639(w__436 ,w__350 ,w__341);
  and g__640(w__435 ,w__349 ,w__257);
  and g__641(w__434 ,w__282 ,w__319);
  or g__642(w__433 ,w__268 ,w__271);
  or g__643(w__432 ,w__353 ,w__247);
  and g__644(w__431 ,w__273 ,w__281);
  or g__645(w__430 ,w__262 ,w__346);
  or g__646(w__429 ,w__254 ,w__318);
  or g__647(w__428 ,w__274 ,w__342);
  and g__648(w__427 ,w__266 ,w__330);
  and g__649(w__426 ,w__261 ,w__335);
  or g__650(w__425 ,w__280 ,w__331);
  and g__651(w__424 ,w__339 ,w__325);
  and g__652(w__467 ,w__309 ,w__374);
  and g__653(w__466 ,w__288 ,w__358);
  and g__654(w__464 ,w__290 ,w__363);
  not g__655(w__422 ,w__421);
  not g__656(w__417 ,w__418);
  not g__657(w__414 ,w__415);
  or g__658(w__413 ,w__261 ,w__335);
  xor g__659(w__8510 ,in2[0] ,in3[0]);
  and g__660(w__412 ,w__256 ,w__277);
  and g__661(w__411 ,w__278 ,w__343);
  nor g__662(w__410 ,w__303 ,w__315);
  or g__663(w__409 ,w__320 ,w__284);
  or g__664(w__408 ,w__350 ,w__341);
  and g__665(w__407 ,w__334 ,w__323);
  or g__666(w__406 ,w__352 ,w__333);
  or g__667(w__405 ,w__255 ,w__329);
  or g__668(w__404 ,w__278 ,w__343);
  nor g__669(w__403 ,w__370 ,w__314);
  or g__670(w__402 ,w__345 ,w__286);
  and g__671(w__401 ,w__274 ,w__342);
  or g__672(w__400 ,w__256 ,w__277);
  or g__673(w__399 ,w__326 ,w__267);
  nor g__674(w__398 ,w__300 ,w__312);
  and g__675(w__397 ,w__280 ,w__331);
  or g__676(w__396 ,w__291 ,w__313);
  or g__677(w__395 ,w__328 ,w__338);
  and g__678(w__394 ,w__352 ,w__333);
  or g__679(w__393 ,w__266 ,w__330);
  and g__680(w__392 ,w__326 ,w__267);
  or g__681(w__391 ,w__340 ,w__287);
  or g__682(w__390 ,w__282 ,w__319);
  and g__683(w__389 ,w__254 ,w__318);
  or g__684(w__388 ,w__349 ,w__257);
  and g__685(w__387 ,w__258 ,w__327);
  or g__686(w__386 ,w__334 ,w__323);
  or g__687(w__385 ,w__339 ,w__325);
  or g__688(w__384 ,w__269 ,w__279);
  xnor g__689(w__383 ,in2[8] ,in3[8]);
  xnor g__690(w__382 ,in2[7] ,in3[7]);
  xnor g__691(w__381 ,in2[9] ,in3[9]);
  xnor g__692(w__380 ,in2[10] ,in3[10]);
  xnor g__693(w__379 ,in2[1] ,in3[1]);
  xnor g__694(w__423 ,in2[4] ,in3[4]);
  and g__695(w__421 ,w__372 ,w__304);
  and g__696(w__420 ,w__376 ,w__289);
  xnor g__697(w__419 ,in2[6] ,in3[6]);
  xnor g__698(w__418 ,in2[3] ,in3[3]);
  xnor g__699(w__416 ,in2[5] ,in3[5]);
  xnor g__700(w__415 ,in2[2] ,in3[2]);
  not g__701(w__376 ,w__375);
  not g__702(w__374 ,w__373);
  not g__703(w__372 ,w__371);
  not g__704(w__363 ,w__362);
  not g__705(w__358 ,w__357);
  or g__706(w__316 ,w__142 ,w__101);
  nor g__707(w__315 ,in2[10] ,in3[10]);
  nor g__708(w__314 ,in2[8] ,in3[8]);
  nor g__709(w__313 ,in2[7] ,in3[7]);
  nor g__710(w__312 ,in2[9] ,in3[9]);
  and g__711(w__311 ,in2[9] ,in3[9]);
  or g__712(w__378 ,w__70 ,w__75);
  or g__713(w__377 ,w__90 ,w__93);
  or g__714(w__375 ,w__99 ,w__145);
  or g__715(w__373 ,w__109 ,w__111);
  or g__716(w__371 ,w__32 ,w__120);
  or g__717(w__370 ,w__66 ,w__73);
  or g__718(w__369 ,w__47 ,w__38);
  or g__719(w__368 ,w__68 ,w__122);
  or g__720(w__367 ,w__133 ,w__35);
  or g__721(w__366 ,w__62 ,w__26);
  or g__722(w__365 ,w__171 ,w__124);
  or g__723(w__364 ,w__106 ,w__154);
  or g__724(w__362 ,w__118 ,w__139);
  or g__725(w__361 ,w__20 ,w__181);
  or g__726(w__360 ,w__29 ,w__59);
  or g__727(w__359 ,w__214 ,w__23);
  or g__728(w__357 ,w__80 ,w__95);
  or g__729(w__356 ,w__177 ,w__148);
  or g__730(w__355 ,w__205 ,w__37);
  or g__731(w__354 ,w__49 ,w__126);
  or g__732(w__353 ,w__35 ,w__103);
  or g__733(w__352 ,w__78 ,w__174);
  or g__734(w__351 ,w__113 ,w__140);
  or g__735(w__350 ,w__31 ,w__186);
  or g__736(w__349 ,w__29 ,w__131);
  or g__737(w__348 ,w__61 ,w__188);
  or g__738(w__347 ,w__14 ,w__168);
  or g__739(w__346 ,w__17 ,w__44);
  or g__740(w__345 ,w__86 ,w__28);
  or g__741(w__344 ,w__59 ,w__41);
  or g__742(w__343 ,w__203 ,w__184);
  or g__743(w__342 ,w__157 ,w__190);
  or g__744(w__341 ,w__43 ,w__124);
  or g__745(w__340 ,w__25 ,w__34);
  or g__746(w__339 ,w__64 ,w__174);
  or g__747(w__338 ,w__58 ,w__179);
  or g__748(w__337 ,w__8 ,w__200);
  or g__749(w__336 ,w__129 ,w__163);
  or g__750(w__335 ,w__211 ,w__83);
  or g__751(w__334 ,w__160 ,w__143);
  or g__752(w__333 ,w__115 ,w__205);
  or g__753(w__332 ,w__165 ,w__23);
  or g__754(w__331 ,w__19 ,w__22);
  or g__755(w__330 ,w__213 ,w__16);
  or g__756(w__329 ,w__56 ,w__93);
  or g__757(w__328 ,w__137 ,w__190);
  or g__758(w__327 ,w__208 ,w__146);
  or g__759(w__326 ,w__11 ,w__118);
  or g__760(w__325 ,w__88 ,w__80);
  or g__761(w__324 ,w__113 ,w__96);
  or g__762(w__323 ,w__53 ,w__181);
  or g__763(w__322 ,w__78 ,w__73);
  or g__764(w__321 ,w__120 ,w__137);
  or g__765(w__320 ,w__200 ,w__111);
  or g__766(w__319 ,w__198 ,w__41);
  or g__767(w__318 ,w__220 ,w__241);
  or g__768(w__317 ,w__217 ,w__139);
  not g__769(w__264 ,w__263);
  not g__770(w__253 ,w__252);
  nor g__771(w__250 ,w__220 ,w__211);
  nor g__772(w__249 ,w__217 ,w__214);
  or g__773(w__248 ,w__168 ,w__115);
  nor g__774(w__247 ,in2[1] ,in3[1]);
  and g__775(w__8511 ,in2[0] ,in3[0]);
  or g__776(w__310 ,w__70 ,w__149);
  and g__777(w__309 ,in2[5] ,in2[3]);
  and g__778(w__308 ,in2[1] ,in2[0]);
  or g__779(w__307 ,w__40 ,w__104);
  or g__780(w__306 ,w__68 ,w__154);
  or g__781(w__305 ,w__50 ,w__148);
  and g__782(w__304 ,in2[7] ,in2[3]);
  or g__783(w__303 ,w__13 ,w__193);
  or g__784(w__302 ,w__47 ,w__62);
  or g__785(w__301 ,w__83 ,w__151);
  or g__786(w__300 ,w__134 ,w__20);
  or g__787(w__299 ,w__50 ,w__165);
  or g__788(w__298 ,w__208 ,w__157);
  or g__789(w__297 ,w__10 ,w__99);
  or g__790(w__296 ,w__198 ,w__38);
  or g__791(w__295 ,w__166 ,w__179);
  or g__792(w__294 ,w__44 ,w__182);
  or g__793(w__293 ,w__26 ,w__149);
  or g__794(w__292 ,w__107 ,w__55);
  or g__795(w__291 ,w__196 ,w__163);
  and g__796(w__290 ,in2[3] ,in2[1]);
  and g__797(w__289 ,in3[2] ,in3[0]);
  and g__798(w__288 ,in2[4] ,in2[2]);
  or g__799(w__287 ,w__53 ,w__104);
  or g__800(w__286 ,w__133 ,w__206);
  or g__801(w__285 ,w__7 ,w__171);
  or g__802(w__284 ,w__52 ,w__191);
  or g__803(w__283 ,w__158 ,w__151);
  or g__804(w__282 ,w__88 ,w__136);
  or g__805(w__281 ,w__66 ,w__142);
  or g__806(w__280 ,w__86 ,w__184);
  or g__807(w__279 ,w__17 ,w__188);
  or g__808(w__278 ,w__201 ,w__160);
  or g__809(w__277 ,w__155 ,w__101);
  or g__810(w__276 ,w__193 ,w__203);
  or g__811(w__275 ,w__117 ,w__56);
  or g__812(w__274 ,w__128 ,w__145);
  or g__813(w__273 ,w__169 ,w__161);
  or g__814(w__272 ,w__196 ,w__64);
  or g__815(w__271 ,w__177 ,w__90);
  or g__816(w__270 ,w__8 ,w__186);
  or g__817(w__269 ,w__194 ,w__143);
  or g__818(w__268 ,w__210 ,w__152);
  or g__819(w__267 ,w__134 ,w__122);
  or g__820(w__266 ,w__14 ,w__129);
  or g__821(w__265 ,w__75 ,w__126);
  and g__822(w__263 ,in2[3] ,in2[0]);
  or g__823(w__262 ,w__11 ,w__131);
  or g__824(w__261 ,w__219 ,w__77);
  or g__825(w__260 ,w__216 ,w__32);
  or g__826(w__259 ,w__82 ,w__92);
  or g__827(w__258 ,w__136 ,w__172);
  or g__828(w__257 ,w__85 ,w__140);
  or g__829(w__256 ,w__98 ,w__96);
  or g__830(w__255 ,w__175 ,w__146);
  or g__831(w__254 ,w__109 ,w__72);
  and g__832(w__252 ,in3[9] ,in3[7]);
  or g__833(w__251 ,w__46 ,w__107);
  not g__834(w__246 ,in2[0]);
  not g__835(w__245 ,in3[0]);
  not g__836(w__244 ,in3[2]);
  not g__837(w__243 ,in3[6]);
  not g__838(w__242 ,in3[3]);
  not g__839(w__241 ,in2[3]);
  not g__840(w__240 ,in2[4]);
  not g__841(w__239 ,in2[5]);
  not g__842(w__238 ,in2[1]);
  not g__843(w__237 ,in3[1]);
  not g__844(w__236 ,in2[9]);
  not g__845(w__235 ,in2[6]);
  not g__846(w__234 ,in3[5]);
  not g__847(w__233 ,in2[2]);
  not g__848(w__232 ,in3[4]);
  not g__849(w__231 ,in3[7]);
  not g__850(w__230 ,in2[7]);
  not g__851(w__229 ,in2[8]);
  not g__852(w__228 ,in2[10]);
  not g__853(w__227 ,in3[10]);
  not g__854(w__226 ,in3[9]);
  not g__855(w__225 ,in3[8]);
  not g__856(w__222 ,w__224);
  not g__857(w__224 ,w__917);
  not g__858(w__221 ,w__223);
  not g__859(w__223 ,w__771);
  not g__860(w__220 ,w__218);
  not g__861(w__219 ,w__218);
  not g__862(w__218 ,w__229);
  not g__863(w__217 ,w__215);
  not g__864(w__216 ,w__215);
  not g__865(w__215 ,w__228);
  not g__866(w__214 ,w__212);
  not g__867(w__213 ,w__212);
  not g__868(w__212 ,w__227);
  not g__869(w__211 ,w__209);
  not g__870(w__210 ,w__209);
  not g__871(w__209 ,w__225);
  not g__872(w__208 ,w__207);
  not g__873(w__207 ,w__239);
  not g__874(w__206 ,w__204);
  not g__875(w__205 ,w__204);
  not g__876(w__204 ,w__243);
  not g__877(w__203 ,w__202);
  not g__878(w__202 ,w__230);
  not g__879(w__201 ,w__199);
  not g__880(w__200 ,w__199);
  not g__881(w__199 ,w__239);
  not g__882(w__198 ,w__197);
  not g__883(w__197 ,w__231);
  not g__884(w__196 ,w__195);
  not g__885(w__195 ,w__236);
  not g__886(w__194 ,w__192);
  not g__887(w__193 ,w__192);
  not g__888(w__192 ,w__236);
  not g__889(w__191 ,w__189);
  not g__890(w__190 ,w__189);
  not g__891(w__189 ,w__242);
  not g__892(w__188 ,w__187);
  not g__893(w__187 ,w__244);
  not g__894(w__186 ,w__185);
  not g__895(w__185 ,w__238);
  not g__896(w__184 ,w__183);
  not g__897(w__183 ,w__233);
  not g__898(w__182 ,w__180);
  not g__899(w__181 ,w__180);
  not g__900(w__180 ,w__237);
  not g__901(w__179 ,w__178);
  not g__902(w__178 ,w__245);
  not g__903(w__177 ,w__176);
  not g__904(w__176 ,w__226);
  not g__905(w__175 ,w__173);
  not g__906(w__174 ,w__173);
  not g__907(w__173 ,w__235);
  not g__908(w__172 ,w__170);
  not g__909(w__171 ,w__170);
  not g__910(w__170 ,w__233);
  not g__911(w__169 ,w__167);
  not g__912(w__168 ,w__167);
  not g__913(w__167 ,w__230);
  not g__914(w__166 ,w__164);
  not g__915(w__165 ,w__164);
  not g__916(w__164 ,w__231);
  not g__917(w__163 ,w__162);
  not g__918(w__162 ,w__240);
  not g__919(w__161 ,w__159);
  not g__920(w__160 ,w__159);
  not g__921(w__159 ,w__240);
  not g__922(w__158 ,w__156);
  not g__923(w__157 ,w__156);
  not g__924(w__156 ,w__234);
  not g__925(w__155 ,w__153);
  not g__926(w__154 ,w__153);
  not g__927(w__153 ,w__244);
  not g__928(w__152 ,w__150);
  not g__929(w__151 ,w__150);
  not g__930(w__150 ,w__232);
  not g__931(w__149 ,w__147);
  not g__932(w__148 ,w__147);
  not g__933(w__147 ,w__245);
  not g__934(w__146 ,w__144);
  not g__935(w__145 ,w__144);
  not g__936(w__144 ,w__246);
  not g__937(w__143 ,w__141);
  not g__938(w__142 ,w__141);
  not g__939(w__141 ,w__238);
  not g__940(w__140 ,w__138);
  not g__941(w__139 ,w__138);
  not g__942(w__138 ,w__246);
  not g__943(w__137 ,w__135);
  not g__944(w__136 ,w__135);
  not g__945(w__135 ,w__241);
  not g__946(w__134 ,w__132);
  not g__947(w__133 ,w__132);
  not g__948(w__132 ,w__226);
  not g__949(w__131 ,w__130);
  not g__950(w__130 ,w__241);
  not g__951(w__129 ,w__127);
  not g__952(w__128 ,w__127);
  not g__953(w__127 ,w__229);
  not g__954(w__126 ,w__125);
  not g__955(w__125 ,w__152);
  not g__956(w__124 ,w__123);
  not g__957(w__123 ,w__155);
  not g__958(w__122 ,w__121);
  not g__959(w__121 ,w__158);
  not g__960(w__120 ,w__119);
  not g__961(w__119 ,w__161);
  not g__962(w__118 ,w__116);
  not g__963(w__117 ,w__116);
  not g__964(w__116 ,w__240);
  not g__965(w__115 ,w__114);
  not g__966(w__114 ,w__166);
  not g__967(w__113 ,w__112);
  not g__968(w__112 ,w__169);
  not g__969(w__111 ,w__110);
  not g__970(w__110 ,w__172);
  not g__971(w__109 ,w__108);
  not g__972(w__108 ,w__175);
  not g__973(w__107 ,w__105);
  not g__974(w__106 ,w__105);
  not g__975(w__105 ,w__226);
  not g__976(w__104 ,w__102);
  not g__977(w__103 ,w__102);
  not g__978(w__102 ,w__245);
  not g__979(w__101 ,w__100);
  not g__980(w__100 ,w__182);
  not g__981(w__99 ,w__97);
  not g__982(w__98 ,w__97);
  not g__983(w__97 ,w__233);
  not g__984(w__96 ,w__94);
  not g__985(w__95 ,w__94);
  not g__986(w__94 ,w__238);
  not g__987(w__93 ,w__91);
  not g__988(w__92 ,w__91);
  not g__989(w__91 ,w__244);
  not g__990(w__90 ,w__89);
  not g__991(w__89 ,w__191);
  not g__992(w__88 ,w__87);
  not g__993(w__87 ,w__194);
  not g__994(w__86 ,w__84);
  not g__995(w__85 ,w__84);
  not g__996(w__84 ,w__236);
  not g__997(w__83 ,w__81);
  not g__998(w__82 ,w__81);
  not g__999(w__81 ,w__231);
  not g__1000(w__80 ,w__79);
  not g__1001(w__79 ,w__201);
  not g__1002(w__78 ,w__76);
  not g__1003(w__77 ,w__76);
  not g__1004(w__76 ,w__230);
  not g__1005(w__75 ,w__74);
  not g__1006(w__74 ,w__206);
  not g__1007(w__73 ,w__71);
  not g__1008(w__72 ,w__71);
  not g__1009(w__71 ,w__239);
  not g__1010(w__70 ,w__69);
  not g__1011(w__69 ,w__210);
  not g__1012(w__68 ,w__67);
  not g__1013(w__67 ,w__213);
  not g__1014(w__66 ,w__65);
  not g__1015(w__65 ,w__216);
  not g__1016(w__64 ,w__63);
  not g__1017(w__63 ,w__219);
  not g__1018(w__62 ,w__60);
  not g__1019(w__61 ,w__60);
  not g__1020(w__60 ,w__243);
  not g__1021(w__59 ,w__57);
  not g__1022(w__58 ,w__57);
  not g__1023(w__57 ,w__243);
  not g__1024(w__56 ,w__54);
  not g__1025(w__55 ,w__54);
  not g__1026(w__54 ,w__232);
  not g__1027(w__53 ,w__51);
  not g__1028(w__52 ,w__51);
  not g__1029(w__51 ,w__232);
  not g__1030(w__50 ,w__48);
  not g__1031(w__49 ,w__48);
  not g__1032(w__48 ,w__227);
  not g__1033(w__47 ,w__45);
  not g__1034(w__46 ,w__45);
  not g__1035(w__45 ,w__227);
  not g__1036(w__44 ,w__42);
  not g__1037(w__43 ,w__42);
  not g__1038(w__42 ,w__234);
  not g__1039(w__41 ,w__39);
  not g__1040(w__40 ,w__39);
  not g__1041(w__39 ,w__234);
  not g__1042(w__38 ,w__36);
  not g__1043(w__37 ,w__36);
  not g__1044(w__36 ,w__237);
  not g__1045(w__35 ,w__33);
  not g__1046(w__34 ,w__33);
  not g__1047(w__33 ,w__237);
  not g__1048(w__32 ,w__30);
  not g__1049(w__31 ,w__30);
  not g__1050(w__30 ,w__235);
  not g__1051(w__29 ,w__27);
  not g__1052(w__28 ,w__27);
  not g__1053(w__27 ,w__235);
  not g__1054(w__26 ,w__24);
  not g__1055(w__25 ,w__24);
  not g__1056(w__24 ,w__242);
  not g__1057(w__23 ,w__21);
  not g__1058(w__22 ,w__21);
  not g__1059(w__21 ,w__242);
  not g__1060(w__20 ,w__18);
  not g__1061(w__19 ,w__18);
  not g__1062(w__18 ,w__225);
  not g__1063(w__17 ,w__15);
  not g__1064(w__16 ,w__15);
  not g__1065(w__15 ,w__225);
  not g__1066(w__14 ,w__12);
  not g__1067(w__13 ,w__12);
  not g__1068(w__12 ,w__228);
  not g__1069(w__11 ,w__9);
  not g__1070(w__10 ,w__9);
  not g__1071(w__9 ,w__228);
  not g__1072(w__8 ,w__6);
  not g__1073(w__7 ,w__6);
  not g__1074(w__6 ,w__229);
  xor g__1075(w__8525 ,w__1050 ,w__1031);
  xor g__1076(w__8524 ,w__1048 ,w__1038);
  xor g__1077(w__8523 ,w__1046 ,w__1039);
  xor g__1078(w__8522 ,w__1044 ,w__1030);
  xor g__1079(w__8521 ,w__1042 ,w__1019);
  xor g__1080(w__8519 ,w__1023 ,w__988);
  xor g__1081(w__5 ,w__309 ,w__373);
  xnor g__1082(w__8512 ,w__308 ,w__565);
  xor g__1083(w__4 ,w__371 ,w__304);
  xor g__1084(w__3 ,w__290 ,w__362);
  xor g__1085(w__2 ,w__375 ,w__289);
  xor g__1086(w__1 ,w__288 ,w__357);
  xnor g__1087(w__8508 ,w__1737 ,w__1189);
  and g__1088(w__8509 ,w__1189 ,w__1738);
  not g__1089(w__1738 ,w__1737);
  and g__1090(w__1737 ,w__1440 ,w__1736);
  or g__1091(w__1736 ,w__1426 ,w__1735);
  and g__1092(w__1735 ,w__1536 ,w__1734);
  or g__1093(w__1734 ,w__1535 ,w__1733);
  and g__1094(w__1733 ,w__1584 ,w__1732);
  or g__1095(w__1732 ,w__1586 ,w__1731);
  and g__1096(w__1731 ,w__1641 ,w__1730);
  or g__1097(w__1730 ,w__1633 ,w__1729);
  and g__1098(w__1729 ,w__1667 ,w__1728);
  or g__1099(w__1728 ,w__1668 ,w__1727);
  and g__1100(w__1727 ,w__1675 ,w__1726);
  or g__1101(w__1726 ,w__1674 ,w__1725);
  and g__1102(w__1725 ,w__1699 ,w__1724);
  or g__1103(w__1724 ,w__1700 ,w__1723);
  and g__1104(w__1723 ,w__1706 ,w__1722);
  or g__1105(w__1722 ,w__1705 ,w__1721);
  and g__1106(w__1721 ,w__1698 ,w__1720);
  or g__1107(w__1720 ,w__1697 ,w__1719);
  and g__1108(w__1719 ,w__1696 ,w__1718);
  or g__1109(w__1718 ,w__1695 ,w__1717);
  and g__1110(w__1717 ,w__1686 ,w__1716);
  or g__1111(w__1716 ,w__1685 ,w__1715);
  and g__1112(w__1715 ,w__1672 ,w__1714);
  xnor g__1113(w__8496 ,w__1712 ,w__1679);
  or g__1114(w__1714 ,w__1666 ,w__1713);
  not g__1115(w__1713 ,w__1712);
  or g__1116(w__1712 ,w__1647 ,w__1711);
  xnor g__1117(w__8495 ,w__1710 ,w__1664);
  and g__1118(w__1711 ,w__1654 ,w__1710);
  or g__1119(w__1710 ,w__1624 ,w__1709);
  xnor g__1120(w__8494 ,w__1707 ,w__1632);
  and g__1121(w__1709 ,w__1623 ,w__1707);
  xnor g__1122(w__1708 ,w__1688 ,w__1694);
  or g__1123(w__1707 ,w__1602 ,w__1701);
  or g__1124(w__1706 ,w__1687 ,w__1693);
  nor g__1125(w__1705 ,w__1688 ,w__1694);
  xnor g__1126(w__1704 ,w__1690 ,w__1670);
  xnor g__1127(w__1703 ,w__1658 ,w__1682);
  xnor g__1128(w__1702 ,w__1660 ,w__1684);
  xnor g__1129(w__8493 ,w__1691 ,w__1610);
  and g__1130(w__1701 ,w__1601 ,w__1691);
  nor g__1131(w__1700 ,w__1690 ,w__1670);
  or g__1132(w__1699 ,w__1689 ,w__1669);
  or g__1133(w__1698 ,w__1657 ,w__1681);
  nor g__1134(w__1697 ,w__1658 ,w__1682);
  or g__1135(w__1696 ,w__1659 ,w__1683);
  nor g__1136(w__1695 ,w__1660 ,w__1684);
  not g__1137(w__1694 ,w__1693);
  xnor g__1138(w__1693 ,w__1618 ,w__1665);
  xnor g__1139(w__1692 ,w__1671 ,w__1662);
  not g__1140(w__1689 ,w__1690);
  not g__1141(w__1687 ,w__1688);
  or g__1142(w__1686 ,w__1662 ,w__1671);
  and g__1143(w__1685 ,w__1662 ,w__1671);
  or g__1144(w__1691 ,w__1571 ,w__1676);
  or g__1145(w__1690 ,w__1656 ,w__1673);
  or g__1146(w__1688 ,w__1597 ,w__1677);
  not g__1147(w__1684 ,w__1683);
  not g__1148(w__1682 ,w__1681);
  xnor g__1149(w__8492 ,w__1663 ,w__1581);
  xnor g__1150(w__1680 ,w__1648 ,w__1661);
  xnor g__1151(w__1679 ,w__1645 ,w__1652);
  xnor g__1152(w__1678 ,w__1643 ,w__1650);
  xnor g__1153(w__1683 ,w__1590 ,w__1075);
  xnor g__1154(w__1681 ,w__1653 ,w__1609);
  and g__1155(w__1677 ,w__1585 ,w__1653);
  and g__1156(w__1676 ,w__1570 ,w__1663);
  or g__1157(w__1675 ,w__1661 ,w__1648);
  and g__1158(w__1674 ,w__1661 ,w__1648);
  nor g__1159(w__1673 ,w__1618 ,w__1655);
  or g__1160(w__1672 ,w__1644 ,w__1651);
  not g__1161(w__1669 ,w__1670);
  nor g__1162(w__1668 ,w__1643 ,w__1650);
  or g__1163(w__1667 ,w__1642 ,w__1649);
  nor g__1164(w__1666 ,w__1645 ,w__1652);
  xnor g__1165(w__1665 ,w__1636 ,w__1213);
  xnor g__1166(w__1664 ,w__1616 ,w__1635);
  xnor g__1167(w__1671 ,w__1578 ,w__1631);
  xnor g__1168(w__1670 ,w__1606 ,w__1630);
  not g__1169(w__1659 ,w__1660);
  not g__1170(w__1658 ,w__1657);
  and g__1171(w__1656 ,w__1213 ,w__1636);
  nor g__1172(w__1655 ,w__1212 ,w__1636);
  or g__1173(w__1654 ,w__1616 ,w__1635);
  or g__1174(w__1663 ,w__1569 ,w__1637);
  and g__1175(w__1662 ,w__1626 ,w__1638);
  and g__1176(w__1661 ,w__1625 ,w__1640);
  or g__1177(w__1660 ,w__1621 ,w__1639);
  and g__1178(w__1657 ,w__1620 ,w__1634);
  not g__1179(w__1651 ,w__1652);
  not g__1180(w__1649 ,w__1650);
  xnor g__1181(w__8491 ,w__1628 ,w__1580);
  and g__1182(w__1647 ,w__1616 ,w__1635);
  xnor g__1183(w__1646 ,w__1617 ,w__1627);
  xnor g__1184(w__1653 ,w__1608 ,w__1221);
  xnor g__1185(w__1652 ,w__1593 ,w__1067);
  xnor g__1186(w__1650 ,w__1612 ,w__1217);
  xnor g__1187(w__1648 ,w__1561 ,w__1607);
  not g__1188(w__1645 ,w__1644);
  not g__1189(w__1643 ,w__1642);
  or g__1190(w__1641 ,w__1627 ,w__1617);
  or g__1191(w__1640 ,w__1606 ,w__1074);
  nor g__1192(w__1639 ,w__1578 ,w__1615);
  or g__1193(w__1638 ,w__1564 ,w__1622);
  and g__1194(w__1637 ,w__1568 ,w__1628);
  and g__1195(w__1644 ,w__1605 ,w__1613);
  and g__1196(w__1642 ,w__1595 ,w__1614);
  or g__1197(w__1634 ,w__1629 ,w__1619);
  xnor g__1198(w__8490 ,w__1563 ,w__1582);
  and g__1199(w__1633 ,w__1627 ,w__1617);
  xnor g__1200(w__1632 ,w__1575 ,w__1588);
  xnor g__1201(w__1631 ,w__1587 ,w__1204);
  xnor g__1202(w__1630 ,w__1591 ,w__1231);
  xnor g__1203(w__1636 ,w__1498 ,w__1583);
  xnor g__1204(w__1635 ,w__1551 ,w__1066);
  or g__1205(w__1626 ,w__1249 ,w__1593);
  or g__1206(w__1625 ,w__1262 ,w__1591);
  and g__1207(w__1624 ,w__1575 ,w__1588);
  or g__1208(w__1623 ,w__1575 ,w__1588);
  nor g__1209(w__1622 ,w__1219 ,w__1592);
  and g__1210(w__1621 ,w__1204 ,w__1587);
  or g__1211(w__1620 ,w__1554 ,w__1590);
  nor g__1212(w__1619 ,w__1555 ,w__1589);
  and g__1213(w__1629 ,w__1565 ,w__1596);
  or g__1214(w__1628 ,w__1567 ,w__1598);
  and g__1215(w__1627 ,w__1538 ,w__1599);
  nor g__1216(w__1615 ,w__1203 ,w__1587);
  or g__1217(w__1614 ,w__1561 ,w__1600);
  or g__1218(w__1613 ,w__1531 ,w__1604);
  xnor g__1219(w__1612 ,w__1579 ,w__1496);
  xnor g__1220(w__1611 ,w__1560 ,w__1553);
  xnor g__1221(w__1610 ,w__1544 ,w__1556);
  xnor g__1222(w__1609 ,w__1549 ,w__1577);
  xnor g__1223(w__1608 ,w__1562 ,w__1455);
  xnor g__1224(w__1607 ,w__1558 ,w__1234);
  and g__1225(w__1618 ,w__1513 ,w__1594);
  xnor g__1226(w__1617 ,w__1545 ,w__1224);
  or g__1227(w__1616 ,w__1574 ,w__1603);
  or g__1228(w__1605 ,w__1261 ,w__1551);
  nor g__1229(w__1604 ,w__1215 ,w__1550);
  nor g__1230(w__1603 ,w__1481 ,w__1573);
  and g__1231(w__1602 ,w__1544 ,w__1556);
  or g__1232(w__1601 ,w__1544 ,w__1556);
  nor g__1233(w__1600 ,w__1233 ,w__1558);
  or g__1234(w__1599 ,w__1073 ,w__1579);
  and g__1235(w__1598 ,w__1563 ,w__1547);
  nor g__1236(w__1597 ,w__1549 ,w__1576);
  or g__1237(w__1596 ,w__1482 ,w__1566);
  or g__1238(w__1595 ,w__1259 ,w__1557);
  or g__1239(w__1594 ,w__1072 ,w__1562);
  and g__1240(w__1606 ,w__1534 ,w__1572);
  not g__1241(w__1592 ,w__1593);
  not g__1242(w__1589 ,w__1590);
  nor g__1243(w__1586 ,w__1560 ,w__1553);
  or g__1244(w__1585 ,w__1548 ,w__1577);
  or g__1245(w__1584 ,w__1559 ,w__1552);
  xnor g__1246(w__1583 ,w__1458 ,w__1530);
  xnor g__1247(w__1582 ,w__1373 ,w__1065);
  xnor g__1248(w__1581 ,w__1477 ,w__1528);
  xnor g__1249(w__1580 ,w__1480 ,w__1526);
  xnor g__1250(w__1593 ,w__1501 ,w__1519);
  xnor g__1251(w__1591 ,w__1516 ,w__1522);
  xnor g__1252(w__1590 ,w__1517 ,w__1520);
  xnor g__1253(w__1588 ,w__1525 ,w__1521);
  xnor g__1254(w__1587 ,w__1527 ,w__1518);
  not g__1255(w__1576 ,w__1577);
  nor g__1256(w__1574 ,w__1258 ,w__1525);
  and g__1257(w__1573 ,w__1258 ,w__1525);
  or g__1258(w__1572 ,w__1530 ,w__1532);
  and g__1259(w__1571 ,w__1477 ,w__1528);
  or g__1260(w__1570 ,w__1477 ,w__1528);
  and g__1261(w__1569 ,w__1480 ,w__1526);
  or g__1262(w__1568 ,w__1480 ,w__1526);
  nor g__1263(w__1567 ,w__1373 ,w__1065);
  and g__1264(w__1566 ,w__1460 ,w__1527);
  or g__1265(w__1565 ,w__1460 ,w__1527);
  and g__1266(w__1579 ,w__1503 ,w__1539);
  and g__1267(w__1578 ,w__1505 ,w__1533);
  or g__1268(w__1577 ,w__1509 ,w__1537);
  or g__1269(w__1575 ,w__1476 ,w__1540);
  not g__1270(w__1559 ,w__1560);
  not g__1271(w__1557 ,w__1558);
  not g__1272(w__1554 ,w__1555);
  not g__1273(w__1553 ,w__1552);
  not g__1274(w__1550 ,w__1551);
  not g__1275(w__1548 ,w__1549);
  or g__1276(w__1547 ,w__1372 ,w__1529);
  xnor g__1277(w__8489 ,w__1515 ,w__1449);
  xnor g__1278(w__1546 ,w__1466 ,w__1514);
  xnor g__1279(w__1545 ,w__1500 ,w__1463);
  and g__1280(w__1564 ,w__1494 ,w__1524);
  or g__1281(w__1563 ,w__1424 ,w__1523);
  and g__1282(w__1562 ,w__1490 ,w__1542);
  and g__1283(w__1561 ,w__1511 ,w__1541);
  xnor g__1284(w__1560 ,w__1486 ,w__1226);
  xnor g__1285(w__1558 ,w__1464 ,w__1485);
  xnor g__1286(w__1556 ,w__1499 ,w__1484);
  xnor g__1287(w__1555 ,w__1454 ,w__1487);
  and g__1288(w__1552 ,w__1502 ,w__1543);
  xnor g__1289(w__1551 ,w__1456 ,w__1489);
  xnor g__1290(w__1549 ,w__1432 ,w__1488);
  or g__1291(w__1543 ,w__1500 ,w__1508);
  or g__1292(w__1542 ,w__1445 ,w__1512);
  or g__1293(w__1541 ,w__1516 ,w__1504);
  nor g__1294(w__1540 ,w__1475 ,w__1499);
  or g__1295(w__1539 ,w__1431 ,w__1495);
  or g__1296(w__1538 ,w__1257 ,w__1496);
  nor g__1297(w__1537 ,w__1507 ,w__1517);
  or g__1298(w__1536 ,w__1514 ,w__1466);
  and g__1299(w__1535 ,w__1514 ,w__1466);
  or g__1300(w__1534 ,w__1457 ,w__1498);
  or g__1301(w__1533 ,w__1510 ,w__1501);
  nor g__1302(w__1532 ,w__1458 ,w__1497);
  or g__1303(w__1544 ,w__1427 ,w__1492);
  not g__1304(w__1529 ,w__1065);
  or g__1305(w__1524 ,w__1430 ,w__1493);
  nor g__1306(w__1523 ,w__1437 ,w__1515);
  xnor g__1307(w__1522 ,w__1461 ,w__1443);
  xnor g__1308(w__1521 ,w__1481 ,w__1195);
  xnor g__1309(w__1520 ,w__1479 ,w__1210);
  xnor g__1310(w__1519 ,w__1459 ,w__1478);
  xor g__1311(w__1518 ,w__1460 ,w__1482);
  and g__1312(w__1531 ,w__1425 ,w__1491);
  and g__1313(w__1530 ,w__1470 ,w__1506);
  xnor g__1314(w__1528 ,w__1483 ,w__1064);
  xnor g__1315(w__1527 ,w__1447 ,w__1451);
  xnor g__1316(w__1526 ,w__1450 ,w__1197);
  xnor g__1317(w__1525 ,w__1467 ,w__1453);
  or g__1318(w__1513 ,w__1245 ,w__1455);
  and g__1319(w__1512 ,w__1350 ,w__1454);
  or g__1320(w__1511 ,w__1443 ,w__1461);
  and g__1321(w__1510 ,w__1478 ,w__1459);
  and g__1322(w__1509 ,w__1210 ,w__1479);
  nor g__1323(w__1508 ,w__1223 ,w__1463);
  nor g__1324(w__1507 ,w__1209 ,w__1479);
  or g__1325(w__1506 ,w__1432 ,w__1473);
  or g__1326(w__1505 ,w__1478 ,w__1459);
  and g__1327(w__1504 ,w__1443 ,w__1461);
  or g__1328(w__1503 ,w__1274 ,w__1465);
  or g__1329(w__1502 ,w__1246 ,w__1462);
  and g__1330(w__1517 ,w__1436 ,w__1472);
  and g__1331(w__1516 ,w__1339 ,w__1474);
  and g__1332(w__1514 ,w__1365 ,w__1471);
  not g__1333(w__1497 ,w__1498);
  and g__1334(w__1495 ,w__1274 ,w__1465);
  or g__1335(w__1494 ,w__1367 ,w__1456);
  and g__1336(w__1493 ,w__1367 ,w__1456);
  and g__1337(w__1492 ,w__1422 ,w__1483);
  or g__1338(w__1491 ,w__1428 ,w__1467);
  or g__1339(w__1490 ,w__1350 ,w__1454);
  xnor g__1340(w__1489 ,w__1367 ,w__1430);
  xnor g__1341(w__1488 ,w__1303 ,w__1429);
  xor g__1342(w__1487 ,w__1350 ,w__1445);
  xnor g__1343(w__1486 ,w__1446 ,w__1304);
  xnor g__1344(w__1485 ,w__1274 ,w__1431);
  xnor g__1345(w__1484 ,w__1442 ,w__1193);
  xnor g__1346(w__1501 ,w__1394 ,w__1420);
  and g__1347(w__1500 ,w__1330 ,w__1469);
  xnor g__1348(w__1499 ,w__1068 ,w__1419);
  xnor g__1349(w__1498 ,w__1444 ,w__1377);
  xnor g__1350(w__1496 ,w__1433 ,w__1381);
  nor g__1351(w__1476 ,w__1263 ,w__1442);
  and g__1352(w__1475 ,w__1263 ,w__1442);
  or g__1353(w__1474 ,w__1334 ,w__1444);
  and g__1354(w__1473 ,w__1303 ,w__1429);
  or g__1355(w__1472 ,w__1447 ,w__1441);
  or g__1356(w__1471 ,w__1069 ,w__1446);
  or g__1357(w__1470 ,w__1303 ,w__1429);
  or g__1358(w__1469 ,w__1360 ,w__1433);
  xnor g__1359(w__1468 ,w__1270 ,w__1393);
  xnor g__1360(w__1483 ,w__1351 ,w__1376);
  and g__1361(w__1482 ,w__1402 ,w__1421);
  and g__1362(w__1481 ,w__1409 ,w__1434);
  or g__1363(w__1480 ,w__1364 ,w__1435);
  xnor g__1364(w__1479 ,w__1271 ,w__1397);
  and g__1365(w__1478 ,w__1344 ,w__1423);
  or g__1366(w__1477 ,w__1413 ,w__1438);
  not g__1367(w__1465 ,w__1464);
  not g__1368(w__1462 ,w__1463);
  not g__1369(w__1457 ,w__1458);
  xnor g__1370(w__1453 ,w__1349 ,w__1392);
  xnor g__1371(w__1452 ,w__1416 ,w__1229);
  xnor g__1372(w__1451 ,w__1371 ,w__1387);
  xnor g__1373(w__1450 ,w__1071 ,w__1369);
  xnor g__1374(w__1449 ,w__1370 ,w__1417);
  xnor g__1375(w__1448 ,w__1389 ,w__1236);
  xnor g__1376(w__1467 ,w__1268 ,w__1378);
  xnor g__1377(w__1466 ,w__1396 ,w__1207);
  xnor g__1378(w__1464 ,w__1305 ,w__1383);
  xnor g__1379(w__1463 ,w__1299 ,w__1380);
  xnor g__1380(w__1461 ,w__1281 ,w__1374);
  xnor g__1381(w__1460 ,w__1276 ,w__1375);
  xnor g__1382(w__1459 ,w__1301 ,w__1386);
  xnor g__1383(w__1458 ,w__1280 ,w__1384);
  xnor g__1384(w__1456 ,w__1070 ,w__1379);
  xnor g__1385(w__1455 ,w__1300 ,w__1382);
  xnor g__1386(w__1454 ,w__1320 ,w__1385);
  and g__1387(w__1441 ,w__1371 ,w__1387);
  or g__1388(w__1440 ,w__1250 ,w__1415);
  or g__1389(w__1439 ,w__1248 ,w__1388);
  nor g__1390(w__1438 ,w__1403 ,w__1071);
  and g__1391(w__1437 ,w__1370 ,w__1418);
  or g__1392(w__1436 ,w__1371 ,w__1387);
  and g__1393(w__1435 ,w__1362 ,w__1393);
  or g__1394(w__1434 ,w__1411 ,w__1068);
  and g__1395(w__1447 ,w__1343 ,w__1405);
  and g__1396(w__1446 ,w__1359 ,w__1398);
  and g__1397(w__1445 ,w__1331 ,w__1412);
  and g__1398(w__1444 ,w__1361 ,w__1404);
  and g__1399(w__1443 ,w__1355 ,w__1410);
  and g__1400(w__1442 ,w__1337 ,w__1408);
  nor g__1401(w__1428 ,w__1349 ,w__1392);
  and g__1402(w__1427 ,w__1199 ,w__1390);
  nor g__1403(w__1426 ,w__1228 ,w__1416);
  or g__1404(w__1425 ,w__1348 ,w__1391);
  nor g__1405(w__1424 ,w__1370 ,w__1418);
  or g__1406(w__1423 ,w__1333 ,w__1070);
  or g__1407(w__1422 ,w__1199 ,w__1390);
  or g__1408(w__1421 ,w__1395 ,w__1414);
  xnor g__1409(w__1420 ,w__1312 ,w__1347);
  xnor g__1410(w__1419 ,w__1278 ,w__1368);
  and g__1411(w__1433 ,w__1354 ,w__1407);
  and g__1412(w__1432 ,w__1332 ,w__1400);
  and g__1413(w__1431 ,w__1341 ,w__1406);
  and g__1414(w__1430 ,w__1345 ,w__1399);
  and g__1415(w__1429 ,w__1357 ,w__1401);
  not g__1416(w__1418 ,w__1417);
  not g__1417(w__1416 ,w__1415);
  nor g__1418(w__1414 ,w__1311 ,w__1347);
  nor g__1419(w__1413 ,w__1247 ,w__1369);
  or g__1420(w__1412 ,w__1283 ,w__1338);
  and g__1421(w__1411 ,w__1278 ,w__1368);
  or g__1422(w__1410 ,w__1284 ,w__1353);
  or g__1423(w__1409 ,w__1278 ,w__1368);
  or g__1424(w__1407 ,w__1317 ,w__1352);
  or g__1425(w__1406 ,w__1318 ,w__1335);
  or g__1426(w__1405 ,w__1285 ,w__1342);
  or g__1427(w__1404 ,w__1291 ,w__1340);
  and g__1428(w__1403 ,w__1247 ,w__1369);
  or g__1429(w__1402 ,w__1312 ,w__1346);
  or g__1430(w__1401 ,w__1292 ,w__1358);
  or g__1431(w__1400 ,w__1320 ,w__1329);
  or g__1432(w__1399 ,w__1287 ,w__1336);
  or g__1433(w__1398 ,w__1319 ,w__1356);
  xnor g__1434(w__1397 ,w__1292 ,in4[6]);
  xnor g__1435(w__1396 ,w__1293 ,in4[10]);
  xnor g__1436(w__1417 ,w__1323 ,w__1191);
  and g__1437(w__1415 ,w__1265 ,w__1366);
  not g__1438(w__1395 ,w__1394);
  not g__1439(w__1391 ,w__1392);
  not g__1440(w__1388 ,w__1389);
  xnor g__1441(w__1386 ,w__1279 ,w__1285);
  xnor g__1442(w__1385 ,w__1266 ,w__1307);
  xnor g__1443(w__1384 ,w__1284 ,in4[7]);
  xnor g__1444(w__1383 ,w__1317 ,in4[8]);
  xnor g__1445(w__1382 ,w__1272 ,w__1291);
  xnor g__1446(w__1381 ,w__1302 ,w__1273);
  xnor g__1447(w__1380 ,w__1319 ,in4[9]);
  xnor g__1448(w__1379 ,w__1309 ,w__1310);
  xnor g__1449(w__1378 ,w__1298 ,w__1287);
  xnor g__1450(w__1377 ,w__1267 ,w__1275);
  xnor g__1451(w__1376 ,w__1277 ,w__1308);
  xnor g__1452(w__1375 ,w__1306 ,w__1283);
  xnor g__1453(w__1374 ,w__1297 ,w__1318);
  xnor g__1454(w__1394 ,w__1325 ,in4[5]);
  xnor g__1455(w__1393 ,w__1286 ,in4[2]);
  xnor g__1456(w__1392 ,w__1290 ,in4[4]);
  xnor g__1457(w__1390 ,w__1322 ,in4[3]);
  xnor g__1458(w__1389 ,w__1315 ,in4[1]);
  xnor g__1459(w__1387 ,w__1321 ,w__1295);
  not g__1460(w__1373 ,w__1372);
  or g__1461(w__1366 ,w__1293 ,w__1296);
  or g__1462(w__1365 ,w__1264 ,w__1304);
  nor g__1463(w__1364 ,w__1251 ,w__1270);
  or g__1464(w__1363 ,w__1187 ,w__1289);
  or g__1465(w__1362 ,w__1201 ,w__1269);
  or g__1466(w__1361 ,w__1272 ,w__1300);
  and g__1467(w__1360 ,w__1302 ,w__1273);
  or g__1468(w__1359 ,w__1078 ,w__1299);
  and g__1469(w__1358 ,w__1098 ,w__1271);
  or g__1470(w__1357 ,w__1102 ,w__1271);
  and g__1471(w__1356 ,w__1082 ,w__1299);
  or g__1472(w__1355 ,w__1088 ,w__1280);
  or g__1473(w__1354 ,w__1127 ,w__1305);
  and g__1474(w__1353 ,w__1092 ,w__1280);
  and g__1475(w__1352 ,w__1114 ,w__1305);
  and g__1476(w__1372 ,w__1191 ,w__1324);
  or g__1477(w__1371 ,w__1135 ,w__1325);
  or g__1478(w__1370 ,w__1145 ,w__1315);
  or g__1479(w__1369 ,w__1154 ,w__1286);
  or g__1480(w__1368 ,w__1148 ,w__1322);
  or g__1481(w__1367 ,w__1151 ,w__1290);
  not g__1482(w__1348 ,w__1349);
  not g__1483(w__1346 ,w__1347);
  or g__1484(w__1345 ,w__1268 ,w__1298);
  or g__1485(w__1344 ,w__1309 ,w__1310);
  or g__1486(w__1343 ,w__1301 ,w__1279);
  and g__1487(w__1342 ,w__1301 ,w__1279);
  or g__1488(w__1341 ,w__1297 ,w__1281);
  and g__1489(w__1340 ,w__1272 ,w__1300);
  or g__1490(w__1339 ,w__1267 ,w__1275);
  and g__1491(w__1338 ,w__1276 ,w__1306);
  or g__1492(w__1337 ,w__1277 ,w__1308);
  and g__1493(w__1336 ,w__1268 ,w__1298);
  and g__1494(w__1335 ,w__1297 ,w__1281);
  and g__1495(w__1334 ,w__1267 ,w__1275);
  and g__1496(w__1333 ,w__1309 ,w__1310);
  or g__1497(w__1332 ,w__1266 ,w__1307);
  or g__1498(w__1331 ,w__1276 ,w__1306);
  or g__1499(w__1330 ,w__1302 ,w__1273);
  and g__1500(w__1329 ,w__1266 ,w__1307);
  and g__1501(w__1351 ,w__1326 ,w__1282);
  or g__1502(w__1350 ,w__1321 ,w__1295);
  and g__1503(w__1349 ,w__1294 ,w__1314);
  and g__1504(w__1347 ,w__1316 ,w__1328);
  not g__1505(w__1328 ,w__1327);
  not g__1506(w__1324 ,w__1323);
  not g__1507(w__1314 ,w__1313);
  not g__1508(w__1312 ,w__1311);
  nor g__1509(w__1296 ,in4[10] ,w__1206);
  or g__1510(w__1327 ,w__1111 ,w__1130);
  and g__1511(w__1326 ,in4[3] ,in4[1]);
  or g__1512(w__1325 ,w__1080 ,w__1132);
  or g__1513(w__1323 ,w__1116 ,w__1162);
  or g__1514(w__1322 ,w__1137 ,w__1165);
  or g__1515(w__1321 ,w__1100 ,w__1119);
  or g__1516(w__1320 ,w__1140 ,w__1177);
  or g__1517(w__1319 ,w__1125 ,w__1090);
  or g__1518(w__1318 ,w__1108 ,w__1175);
  or g__1519(w__1317 ,w__1105 ,w__1157);
  and g__1520(w__1316 ,in4[5] ,in4[3]);
  or g__1521(w__1315 ,w__1142 ,w__1132);
  or g__1522(w__1313 ,w__1095 ,w__1130);
  and g__1523(w__1311 ,in4[8] ,in4[1]);
  or g__1524(w__1310 ,w__1085 ,w__1143);
  or g__1525(w__1309 ,w__1179 ,w__1155);
  or g__1526(w__1308 ,w__1152 ,w__1146);
  or g__1527(w__1307 ,w__1167 ,w__1122);
  or g__1528(w__1306 ,w__1113 ,w__1117);
  or g__1529(w__1305 ,w__1185 ,w__1095);
  or g__1530(w__1304 ,w__1170 ,w__1111);
  or g__1531(w__1303 ,w__1110 ,w__1120);
  or g__1532(w__1302 ,w__1140 ,w__1182);
  or g__1533(w__1301 ,w__1160 ,w__1151);
  or g__1534(w__1300 ,w__1186 ,w__1173);
  or g__1535(w__1299 ,w__1139 ,w__1167);
  or g__1536(w__1298 ,w__1137 ,w__1154);
  or g__1537(w__1297 ,w__1114 ,w__1180);
  not g__1538(w__1289 ,w__1288);
  not g__1539(w__1270 ,w__1269);
  or g__1540(w__1265 ,w__1107 ,w__1260);
  or g__1541(w__1295 ,w__1105 ,w__1162);
  and g__1542(w__1294 ,in4[4] ,in4[2]);
  or g__1543(w__1293 ,w__1104 ,w__1082);
  or g__1544(w__1292 ,w__1170 ,w__1142);
  or g__1545(w__1291 ,w__1108 ,w__1177);
  or g__1546(w__1290 ,w__1085 ,w__1165);
  or g__1547(w__1288 ,w__1163 ,w__1238);
  or g__1548(w__1287 ,w__1094 ,w__1145);
  or g__1549(w__1286 ,w__1149 ,w__1129);
  or g__1550(w__1285 ,w__1183 ,w__1155);
  or g__1551(w__1284 ,w__1171 ,w__1123);
  or g__1552(w__1283 ,w__1078 ,w__1143);
  and g__1553(w__1282 ,in4[4] ,in4[0]);
  or g__1554(w__1281 ,w__1080 ,w__1135);
  or g__1555(w__1280 ,w__1168 ,w__1157);
  or g__1556(w__1279 ,w__1102 ,w__1148);
  or g__1557(w__1278 ,w__1160 ,w__1146);
  or g__1558(w__1277 ,w__1173 ,w__1117);
  or g__1559(w__1276 ,w__1084 ,w__1149);
  or g__1560(w__1275 ,w__1077 ,w__1175);
  or g__1561(w__1274 ,w__1127 ,w__1092);
  or g__1562(w__1273 ,w__1125 ,w__1098);
  or g__1563(w__1272 ,w__1088 ,w__1158);
  or g__1564(w__1271 ,w__1090 ,w__1152);
  and g__1565(w__1269 ,in4[2] ,in4[1]);
  or g__1566(w__1268 ,w__1120 ,w__1123);
  or g__1567(w__1267 ,w__1087 ,w__1100);
  or g__1568(w__1266 ,w__1097 ,w__1134);
  not g__1569(w__1264 ,w__1226);
  not g__1570(w__1263 ,w__1193);
  not g__1571(w__1262 ,w__1231);
  not g__1572(w__1261 ,w__1215);
  not g__1573(w__1260 ,w__1207);
  not g__1574(w__1259 ,w__1234);
  not g__1575(w__1258 ,w__1195);
  not g__1576(w__1257 ,w__1217);
  not g__1577(w__1256 ,in4[0]);
  not g__1578(w__1255 ,in4[4]);
  not g__1579(w__1254 ,in4[1]);
  not g__1580(w__1253 ,in4[8]);
  not g__1581(w__1252 ,in4[9]);
  not g__1582(w__1251 ,w__1201);
  not g__1583(w__1250 ,w__1229);
  not g__1584(w__1249 ,w__1219);
  not g__1585(w__1248 ,w__1236);
  not g__1586(w__1247 ,w__1197);
  not g__1587(w__1246 ,w__1224);
  not g__1588(w__1245 ,w__1221);
  not g__1589(w__1244 ,in4[3]);
  not g__1590(w__1243 ,in4[5]);
  not g__1591(w__1242 ,in4[2]);
  not g__1592(w__1241 ,in4[7]);
  not g__1593(w__1240 ,in4[6]);
  not g__1594(w__1239 ,in4[10]);
  not g__1595(w__1236 ,w__1235);
  not g__1596(w__1235 ,w__8512);
  not g__1597(w__1234 ,w__1232);
  not g__1598(w__1233 ,w__1232);
  not g__1599(w__1232 ,w__8526);
  not g__1600(w__1231 ,w__1230);
  not g__1601(w__1230 ,w__8525);
  not g__1602(w__1229 ,w__1227);
  not g__1603(w__1228 ,w__1227);
  not g__1604(w__1227 ,w__8531);
  not g__1605(w__1226 ,w__1225);
  not g__1606(w__1225 ,w__8529);
  not g__1607(w__1224 ,w__1222);
  not g__1608(w__1223 ,w__1222);
  not g__1609(w__1222 ,w__8528);
  not g__1610(w__1221 ,w__1220);
  not g__1611(w__1220 ,w__8523);
  not g__1612(w__1219 ,w__1218);
  not g__1613(w__1218 ,w__8520);
  not g__1614(w__1217 ,w__1216);
  not g__1615(w__1216 ,w__8527);
  not g__1616(w__1215 ,w__1214);
  not g__1617(w__1214 ,w__8519);
  not g__1618(w__1213 ,w__1211);
  not g__1619(w__1212 ,w__1211);
  not g__1620(w__1211 ,w__8524);
  not g__1621(w__1210 ,w__1208);
  not g__1622(w__1209 ,w__1208);
  not g__1623(w__1208 ,w__8522);
  not g__1624(w__1207 ,w__1205);
  not g__1625(w__1206 ,w__1205);
  not g__1626(w__1205 ,w__8530);
  not g__1627(w__1204 ,w__1202);
  not g__1628(w__1203 ,w__1202);
  not g__1629(w__1202 ,w__8521);
  not g__1630(w__1201 ,w__1200);
  not g__1631(w__1200 ,w__8514);
  not g__1632(w__1199 ,w__1198);
  not g__1633(w__1198 ,w__8516);
  not g__1634(w__1197 ,w__1196);
  not g__1635(w__1196 ,w__8515);
  not g__1636(w__1195 ,w__1194);
  not g__1637(w__1194 ,w__8518);
  not g__1638(w__1193 ,w__1192);
  not g__1639(w__1192 ,w__8517);
  not g__1640(w__1191 ,w__1190);
  not g__1641(w__1190 ,w__8513);
  not g__1642(w__1189 ,w__1188);
  not g__1643(w__1188 ,w__8532);
  not g__1644(w__1238 ,w__8510);
  not g__1645(w__1187 ,w__1237);
  not g__1646(w__1237 ,w__8511);
  not g__1647(w__1186 ,w__1184);
  not g__1648(w__1185 ,w__1184);
  not g__1649(w__1184 ,w__1252);
  not g__1650(w__1183 ,w__1181);
  not g__1651(w__1182 ,w__1181);
  not g__1652(w__1181 ,w__1241);
  not g__1653(w__1180 ,w__1178);
  not g__1654(w__1179 ,w__1178);
  not g__1655(w__1178 ,w__1240);
  not g__1656(w__1177 ,w__1176);
  not g__1657(w__1176 ,w__1242);
  not g__1658(w__1175 ,w__1174);
  not g__1659(w__1174 ,w__1255);
  not g__1660(w__1173 ,w__1172);
  not g__1661(w__1172 ,w__1244);
  not g__1662(w__1171 ,w__1169);
  not g__1663(w__1170 ,w__1169);
  not g__1664(w__1169 ,w__1239);
  not g__1665(w__1168 ,w__1166);
  not g__1666(w__1167 ,w__1166);
  not g__1667(w__1166 ,w__1253);
  not g__1668(w__1165 ,w__1164);
  not g__1669(w__1164 ,w__1256);
  not g__1670(w__1163 ,w__1161);
  not g__1671(w__1162 ,w__1161);
  not g__1672(w__1161 ,w__1256);
  not g__1673(w__1160 ,w__1159);
  not g__1674(w__1159 ,w__1243);
  not g__1675(w__1158 ,w__1156);
  not g__1676(w__1157 ,w__1156);
  not g__1677(w__1156 ,w__1243);
  not g__1678(w__1155 ,w__1153);
  not g__1679(w__1154 ,w__1153);
  not g__1680(w__1153 ,w__1242);
  not g__1681(w__1152 ,w__1150);
  not g__1682(w__1151 ,w__1150);
  not g__1683(w__1150 ,w__1255);
  not g__1684(w__1149 ,w__1147);
  not g__1685(w__1148 ,w__1147);
  not g__1686(w__1147 ,w__1244);
  not g__1687(w__1146 ,w__1144);
  not g__1688(w__1145 ,w__1144);
  not g__1689(w__1144 ,w__1254);
  not g__1690(w__1143 ,w__1141);
  not g__1691(w__1142 ,w__1141);
  not g__1692(w__1141 ,w__1254);
  not g__1693(w__1140 ,w__1138);
  not g__1694(w__1139 ,w__1138);
  not g__1695(w__1138 ,w__1252);
  not g__1696(w__1137 ,w__1136);
  not g__1697(w__1136 ,w__1158);
  not g__1698(w__1135 ,w__1133);
  not g__1699(w__1134 ,w__1133);
  not g__1700(w__1133 ,w__1243);
  not g__1701(w__1132 ,w__1131);
  not g__1702(w__1131 ,w__1163);
  not g__1703(w__1130 ,w__1128);
  not g__1704(w__1129 ,w__1128);
  not g__1705(w__1128 ,w__1256);
  not g__1706(w__1127 ,w__1126);
  not g__1707(w__1126 ,w__1168);
  not g__1708(w__1125 ,w__1124);
  not g__1709(w__1124 ,w__1171);
  not g__1710(w__1123 ,w__1121);
  not g__1711(w__1122 ,w__1121);
  not g__1712(w__1121 ,w__1244);
  not g__1713(w__1120 ,w__1118);
  not g__1714(w__1119 ,w__1118);
  not g__1715(w__1118 ,w__1255);
  not g__1716(w__1117 ,w__1115);
  not g__1717(w__1116 ,w__1115);
  not g__1718(w__1115 ,w__1242);
  not g__1719(w__1114 ,w__1112);
  not g__1720(w__1113 ,w__1112);
  not g__1721(w__1112 ,w__1253);
  not g__1722(w__1111 ,w__1109);
  not g__1723(w__1110 ,w__1109);
  not g__1724(w__1109 ,w__1253);
  not g__1725(w__1108 ,w__1106);
  not g__1726(w__1107 ,w__1106);
  not g__1727(w__1106 ,w__1239);
  not g__1728(w__1105 ,w__1103);
  not g__1729(w__1104 ,w__1103);
  not g__1730(w__1103 ,w__1239);
  not g__1731(w__1102 ,w__1101);
  not g__1732(w__1101 ,w__1179);
  not g__1733(w__1100 ,w__1099);
  not g__1734(w__1099 ,w__1180);
  not g__1735(w__1098 ,w__1096);
  not g__1736(w__1097 ,w__1096);
  not g__1737(w__1096 ,w__1240);
  not g__1738(w__1095 ,w__1093);
  not g__1739(w__1094 ,w__1093);
  not g__1740(w__1093 ,w__1240);
  not g__1741(w__1092 ,w__1091);
  not g__1742(w__1091 ,w__1182);
  not g__1743(w__1090 ,w__1089);
  not g__1744(w__1089 ,w__1183);
  not g__1745(w__1088 ,w__1086);
  not g__1746(w__1087 ,w__1086);
  not g__1747(w__1086 ,w__1241);
  not g__1748(w__1085 ,w__1083);
  not g__1749(w__1084 ,w__1083);
  not g__1750(w__1083 ,w__1241);
  not g__1751(w__1082 ,w__1081);
  not g__1752(w__1081 ,w__1185);
  not g__1753(w__1080 ,w__1079);
  not g__1754(w__1079 ,w__1186);
  not g__1755(w__1078 ,w__1076);
  not g__1756(w__1077 ,w__1076);
  not g__1757(w__1076 ,w__1252);
  xor g__1758(w__8507 ,w__1735 ,w__1452);
  xor g__1759(w__8506 ,w__1733 ,w__1546);
  xor g__1760(w__8505 ,w__1731 ,w__1611);
  xor g__1761(w__8504 ,w__1729 ,w__1646);
  xor g__1762(w__8503 ,w__1727 ,w__1678);
  xor g__1763(w__8502 ,w__1725 ,w__1680);
  xor g__1764(w__8501 ,w__1723 ,w__1704);
  xor g__1765(w__8500 ,w__1721 ,w__1708);
  xor g__1766(w__8499 ,w__1719 ,w__1703);
  xor g__1767(w__8498 ,w__1717 ,w__1702);
  xor g__1768(w__8497 ,w__1715 ,w__1692);
  xor g__1769(w__1075 ,w__1555 ,w__1629);
  and g__1770(w__1074 ,w__1230 ,w__1591);
  and g__1771(w__1073 ,w__1216 ,w__1496);
  and g__1772(w__1072 ,w__1220 ,w__1455);
  xnor g__1773(w__1071 ,w__1326 ,w__1282);
  xor g__1774(w__1070 ,w__1316 ,w__1327);
  and g__1775(w__1069 ,w__1225 ,w__1304);
  xor g__1776(w__1068 ,w__1294 ,w__1313);
  xor g__1777(w__1067 ,w__1564 ,w__1218);
  xor g__1778(w__1066 ,w__1531 ,w__1214);
  xor g__1779(w__1065 ,w__1468 ,w__1200);
  xor g__1780(w__1064 ,w__1390 ,w__1198);
  xnor g__1781(w__8486 ,w__1238 ,in4[0]);
  or g__1782(w__8485 ,w__2569 ,w__2801);
  xnor g__1783(w__8484 ,w__2800 ,w__2586);
  and g__1784(w__2801 ,w__2568 ,w__2800);
  or g__1785(w__2800 ,w__2641 ,w__2799);
  xnor g__1786(w__8483 ,w__2798 ,w__2651);
  and g__1787(w__2799 ,w__2642 ,w__2798);
  or g__1788(w__2798 ,w__2692 ,w__2797);
  xnor g__1789(w__8482 ,w__2796 ,w__2704);
  and g__1790(w__2797 ,w__2699 ,w__2796);
  or g__1791(w__2796 ,w__2718 ,w__2795);
  xnor g__1792(w__8481 ,w__2794 ,w__2729);
  and g__1793(w__2795 ,w__2707 ,w__2794);
  or g__1794(w__2794 ,w__2732 ,w__2793);
  xnor g__1795(w__8480 ,w__2792 ,w__2746);
  and g__1796(w__2793 ,w__2741 ,w__2792);
  or g__1797(w__2792 ,w__2764 ,w__2791);
  xnor g__1798(w__8479 ,w__2790 ,w__2770);
  nor g__1799(w__2791 ,w__2765 ,w__2790);
  and g__1800(w__2790 ,w__2789 ,w__2766);
  or g__1801(w__2789 ,w__2758 ,w__2788);
  and g__1802(w__2788 ,w__2774 ,w__2787);
  or g__1803(w__2787 ,w__2773 ,w__2786);
  and g__1804(w__2786 ,w__2785 ,w__2775);
  or g__1805(w__2785 ,w__2772 ,w__2784);
  and g__1806(w__2784 ,w__2763 ,w__2783);
  or g__1807(w__2783 ,w__2762 ,w__2782);
  and g__1808(w__2782 ,w__2751 ,w__2781);
  or g__1809(w__2781 ,w__2752 ,w__2780);
  and g__1810(w__2780 ,w__2736 ,w__2779);
  xnor g__1811(w__8473 ,w__2778 ,w__2745);
  or g__1812(w__2779 ,w__2730 ,w__2778);
  and g__1813(w__2778 ,w__2708 ,w__2771);
  xnor g__1814(w__2777 ,w__2759 ,w__2754);
  xnor g__1815(w__2776 ,w__2760 ,w__2767);
  or g__1816(w__2775 ,w__2754 ,w__2759);
  or g__1817(w__2774 ,w__2767 ,w__2760);
  and g__1818(w__2773 ,w__2767 ,w__2760);
  and g__1819(w__2772 ,w__2754 ,w__2759);
  or g__1820(w__2771 ,w__2709 ,w__2761);
  xnor g__1821(w__2770 ,w__2756 ,w__2734);
  xnor g__1822(w__2769 ,w__2750 ,w__2755);
  xnor g__1823(w__2768 ,w__2743 ,w__2749);
  or g__1824(w__2766 ,w__2755 ,w__2750);
  and g__1825(w__2765 ,w__2756 ,w__2735);
  nor g__1826(w__2764 ,w__2756 ,w__2735);
  or g__1827(w__2763 ,w__2742 ,w__2748);
  nor g__1828(w__2762 ,w__2743 ,w__2749);
  and g__1829(w__2767 ,w__2740 ,w__2753);
  and g__1830(w__2758 ,w__2755 ,w__2750);
  xnor g__1831(w__8471 ,w__2744 ,w__2705);
  xnor g__1832(w__2757 ,w__2733 ,w__2724);
  and g__1833(w__2761 ,w__2679 ,w__2747);
  xnor g__1834(w__2760 ,w__2686 ,w__2727);
  xnor g__1835(w__2759 ,w__2723 ,w__2728);
  or g__1836(w__2753 ,w__2688 ,w__2739);
  and g__1837(w__2752 ,w__2724 ,w__2733);
  or g__1838(w__2751 ,w__2724 ,w__2733);
  and g__1839(w__2756 ,w__2694 ,w__2737);
  and g__1840(w__2755 ,w__2720 ,w__2731);
  and g__1841(w__2754 ,w__2719 ,w__2738);
  not g__1842(w__2748 ,w__2749);
  or g__1843(w__2747 ,w__2693 ,w__2744);
  xnor g__1844(w__8470 ,w__2685 ,w__2703);
  xnor g__1845(w__2746 ,w__2711 ,w__2713);
  xnor g__1846(w__2745 ,w__2682 ,w__2714);
  xnor g__1847(w__2750 ,w__2725 ,w__2706);
  xnor g__1848(w__2749 ,w__2681 ,w__2702);
  not g__1849(w__2742 ,w__2743);
  or g__1850(w__2741 ,w__2712 ,w__2710);
  or g__1851(w__2740 ,w__2654 ,w__2723);
  and g__1852(w__2739 ,w__2654 ,w__2723);
  or g__1853(w__2738 ,w__2676 ,w__2717);
  or g__1854(w__2737 ,w__2725 ,w__2691);
  or g__1855(w__2736 ,w__2682 ,w__2715);
  and g__1856(w__2744 ,w__2698 ,w__2722);
  or g__1857(w__2743 ,w__2667 ,w__2716);
  not g__1858(w__2735 ,w__2734);
  nor g__1859(w__2732 ,w__2713 ,w__2711);
  or g__1860(w__2731 ,w__2686 ,w__2721);
  and g__1861(w__2730 ,w__2682 ,w__2715);
  xnor g__1862(w__2729 ,w__2701 ,w__2655);
  xnor g__1863(w__2728 ,w__2688 ,w__2654);
  xnor g__1864(w__2727 ,w__2684 ,w__2628);
  xnor g__1865(w__2726 ,w__2683 ,w__2674);
  xnor g__1866(w__2734 ,w__2675 ,w__2677);
  xnor g__1867(w__2733 ,w__2687 ,w__2678);
  or g__1868(w__2722 ,w__2697 ,w__2685);
  and g__1869(w__2721 ,w__2628 ,w__2684);
  or g__1870(w__2720 ,w__2628 ,w__2684);
  or g__1871(w__2719 ,w__2612 ,w__2680);
  nor g__1872(w__2718 ,w__1960 ,w__2701);
  nor g__1873(w__2717 ,w__2611 ,w__2681);
  and g__1874(w__2716 ,w__2664 ,w__2687);
  and g__1875(w__2725 ,w__2665 ,w__2690);
  and g__1876(w__2724 ,w__2636 ,w__2689);
  and g__1877(w__2723 ,w__2670 ,w__2695);
  not g__1878(w__2715 ,w__2714);
  not g__1879(w__2713 ,w__2712);
  not g__1880(w__2710 ,w__2711);
  and g__1881(w__2709 ,w__2674 ,w__2683);
  or g__1882(w__2708 ,w__2674 ,w__2683);
  or g__1883(w__2707 ,w__1962 ,w__2700);
  xnor g__1884(w__2706 ,w__2662 ,w__2643);
  xnor g__1885(w__2705 ,w__2627 ,w__2661);
  xnor g__1886(w__2704 ,w__2657 ,w__2596);
  xnor g__1887(w__2703 ,w__2522 ,w__2659);
  xnor g__1888(w__2702 ,w__2676 ,w__2612);
  xnor g__1889(w__2714 ,w__2663 ,w__2649);
  xnor g__1890(w__2712 ,w__2646 ,w__2650);
  and g__1891(w__2711 ,w__2652 ,w__2696);
  not g__1892(w__2701 ,w__2700);
  or g__1893(w__2699 ,w__2595 ,w__2656);
  or g__1894(w__2698 ,w__2521 ,w__2659);
  nor g__1895(w__2697 ,w__2522 ,w__2658);
  or g__1896(w__2696 ,w__2672 ,w__2675);
  or g__1897(w__2695 ,w__2536 ,w__2669);
  or g__1898(w__2694 ,w__2643 ,w__2662);
  nor g__1899(w__2693 ,w__2626 ,w__2661);
  nor g__1900(w__2692 ,w__2596 ,w__2657);
  and g__1901(w__2691 ,w__2643 ,w__2662);
  or g__1902(w__2690 ,w__2529 ,w__2668);
  or g__1903(w__2689 ,w__2640 ,w__2663);
  or g__1904(w__2700 ,w__2637 ,w__2666);
  not g__1905(w__2680 ,w__2681);
  xnor g__1906(w__8469 ,w__2647 ,w__2620);
  or g__1907(w__2679 ,w__2627 ,w__2660);
  xnor g__1908(w__2678 ,w__2594 ,w__2645);
  xnor g__1909(w__2677 ,w__2578 ,w__2633);
  xnor g__1910(w__2688 ,w__2648 ,w__2618);
  xnor g__1911(w__2687 ,w__2525 ,w__2621);
  and g__1912(w__2686 ,w__2590 ,w__2673);
  and g__1913(w__2685 ,w__2609 ,w__2653);
  xnor g__1914(w__2684 ,w__2631 ,w__2623);
  xnor g__1915(w__2683 ,w__2634 ,w__2622);
  and g__1916(w__2682 ,w__2605 ,w__2671);
  xnor g__1917(w__2681 ,w__2630 ,w__2619);
  or g__1918(w__2673 ,w__2610 ,w__2648);
  nor g__1919(w__2672 ,w__2577 ,w__2633);
  or g__1920(w__2671 ,w__2588 ,w__2634);
  or g__1921(w__2670 ,w__2558 ,w__2629);
  nor g__1922(w__2669 ,w__2557 ,w__2630);
  and g__1923(w__2668 ,w__2553 ,w__2631);
  nor g__1924(w__2667 ,w__2593 ,w__2645);
  nor g__1925(w__2666 ,w__2635 ,w__2646);
  or g__1926(w__2665 ,w__2553 ,w__2631);
  or g__1927(w__2664 ,w__2594 ,w__2644);
  and g__1928(w__2676 ,w__2601 ,w__2639);
  and g__1929(w__2675 ,w__2604 ,w__2638);
  and g__1930(w__2674 ,w__2592 ,w__2625);
  not g__1931(w__2660 ,w__2661);
  not g__1932(w__2658 ,w__2659);
  not g__1933(w__2656 ,w__2657);
  or g__1934(w__2653 ,w__2608 ,w__2647);
  or g__1935(w__2652 ,w__2578 ,w__2632);
  xnor g__1936(w__8468 ,w__2559 ,w__2584);
  xnor g__1937(w__2651 ,w__2616 ,w__2509);
  xnor g__1938(w__2650 ,w__2473 ,w__2597);
  xnor g__1939(w__2649 ,w__2614 ,w__2552);
  xnor g__1940(w__2663 ,w__2530 ,w__2582);
  xnor g__1941(w__2662 ,w__2556 ,w__2580);
  xnor g__1942(w__2661 ,w__2547 ,w__2583);
  xnor g__1943(w__2659 ,w__2457 ,w__2579);
  and g__1944(w__2657 ,w__2562 ,w__2624);
  xnor g__1945(w__2655 ,w__2617 ,w__2581);
  xnor g__1946(w__2654 ,w__2505 ,w__2585);
  not g__1947(w__2644 ,w__2645);
  or g__1948(w__2642 ,w__1961 ,w__2615);
  nor g__1949(w__2641 ,w__1959 ,w__2616);
  nor g__1950(w__2640 ,w__2613 ,w__2552);
  or g__1951(w__2639 ,w__2531 ,w__2599);
  or g__1952(w__2638 ,w__2535 ,w__2602);
  nor g__1953(w__2637 ,w__2474 ,w__2597);
  or g__1954(w__2636 ,w__2614 ,w__2551);
  and g__1955(w__2635 ,w__2474 ,w__2597);
  and g__1956(w__2648 ,w__2575 ,w__2606);
  and g__1957(w__2647 ,w__2574 ,w__2607);
  and g__1958(w__2646 ,w__2561 ,w__2603);
  and g__1959(w__2645 ,w__2565 ,w__2598);
  and g__1960(w__2643 ,w__2576 ,w__2600);
  not g__1961(w__2633 ,w__2632);
  not g__1962(w__2629 ,w__2630);
  not g__1963(w__2626 ,w__2627);
  or g__1964(w__2625 ,w__2528 ,w__2591);
  or g__1965(w__2624 ,w__2617 ,w__2566);
  xnor g__1966(w__2623 ,w__2553 ,w__2529);
  xnor g__1967(w__2622 ,w__2550 ,w__2523);
  xnor g__1968(w__2621 ,w__2555 ,w__2531);
  xnor g__1969(w__2620 ,w__2494 ,w__2549);
  xnor g__1970(w__2619 ,w__2558 ,w__2536);
  xnor g__1971(w__2618 ,w__2546 ,w__2516);
  xnor g__1972(w__2634 ,w__2476 ,w__2540);
  xnor g__1973(w__2632 ,w__2506 ,w__2537);
  xnor g__1974(w__2631 ,w__2510 ,w__2539);
  xnor g__1975(w__2630 ,w__2515 ,w__2538);
  and g__1976(w__2628 ,w__2567 ,w__2587);
  and g__1977(w__2627 ,w__2541 ,w__2589);
  not g__1978(w__2615 ,w__2616);
  not g__1979(w__2613 ,w__2614);
  not g__1980(w__2611 ,w__2612);
  and g__1981(w__2610 ,w__2516 ,w__2546);
  or g__1982(w__2609 ,w__2494 ,w__2548);
  nor g__1983(w__2608 ,w__2493 ,w__2549);
  or g__1984(w__2607 ,w__2573 ,w__2559);
  or g__1985(w__2606 ,w__2498 ,w__2572);
  or g__1986(w__2605 ,w__2523 ,w__2550);
  or g__1987(w__2604 ,w__2507 ,w__2556);
  or g__1988(w__2603 ,w__2477 ,w__2543);
  and g__1989(w__2602 ,w__2507 ,w__2556);
  or g__1990(w__2601 ,w__2524 ,w__2555);
  or g__1991(w__2600 ,w__2497 ,w__2564);
  nor g__1992(w__2599 ,w__2525 ,w__2554);
  or g__1993(w__2598 ,w__2530 ,w__2563);
  and g__1994(w__2617 ,w__2492 ,w__2571);
  and g__1995(w__2616 ,w__2488 ,w__2545);
  and g__1996(w__2614 ,w__2518 ,w__2560);
  and g__1997(w__2612 ,w__2440 ,w__2570);
  not g__1998(w__2596 ,w__2595);
  not g__1999(w__2594 ,w__2593);
  xnor g__2000(w__8467 ,w__2496 ,w__2501);
  or g__2001(w__2592 ,w__2512 ,w__2547);
  and g__2002(w__2591 ,w__2512 ,w__2547);
  or g__2003(w__2590 ,w__2516 ,w__2546);
  or g__2004(w__2589 ,w__2457 ,w__2542);
  and g__2005(w__2588 ,w__2523 ,w__2550);
  or g__2006(w__2587 ,w__2534 ,w__2544);
  xnor g__2007(w__2586 ,w__2527 ,w__2282);
  xnor g__2008(w__2585 ,w__2534 ,w__2390);
  xnor g__2009(w__2584 ,w__2389 ,w__2514);
  xnor g__2010(w__2583 ,w__2528 ,w__2511);
  xnor g__2011(w__2582 ,w__2508 ,w__2453);
  xnor g__2012(w__2581 ,w__2504 ,w__2454);
  xnor g__2013(w__2580 ,w__2507 ,w__2535);
  xnor g__2014(w__2579 ,w__2503 ,w__2335);
  xnor g__2015(w__2597 ,w__2533 ,w__2499);
  xnor g__2016(w__2595 ,w__2532 ,w__2500);
  xnor g__2017(w__2593 ,w__2517 ,w__2467);
  not g__2018(w__2577 ,w__2578);
  or g__2019(w__2576 ,w__2323 ,w__2510);
  or g__2020(w__2575 ,w__2421 ,w__2515);
  or g__2021(w__2574 ,w__2388 ,w__2514);
  nor g__2022(w__2573 ,w__2389 ,w__2513);
  and g__2023(w__2572 ,w__2421 ,w__2515);
  or g__2024(w__2571 ,w__2481 ,w__2533);
  or g__2025(w__2570 ,w__2439 ,w__2517);
  nor g__2026(w__2569 ,w__2282 ,w__2527);
  or g__2027(w__2568 ,w__2281 ,w__2526);
  or g__2028(w__2567 ,w__2390 ,w__2505);
  and g__2029(w__2566 ,w__2454 ,w__2504);
  or g__2030(w__2565 ,w__2453 ,w__2508);
  and g__2031(w__2564 ,w__2323 ,w__2510);
  and g__2032(w__2563 ,w__2453 ,w__2508);
  or g__2033(w__2562 ,w__2454 ,w__2504);
  or g__2034(w__2561 ,w__2420 ,w__2506);
  or g__2035(w__2560 ,w__2476 ,w__2519);
  and g__2036(w__2578 ,w__2452 ,w__2520);
  not g__2037(w__2557 ,w__2558);
  not g__2038(w__2554 ,w__2555);
  not g__2039(w__2551 ,w__2552);
  not g__2040(w__2548 ,w__2549);
  or g__2041(w__2545 ,w__2489 ,w__2532);
  and g__2042(w__2544 ,w__2390 ,w__2505);
  and g__2043(w__2543 ,w__2420 ,w__2506);
  and g__2044(w__2542 ,w__2335 ,w__2503);
  or g__2045(w__2541 ,w__2335 ,w__2503);
  xnor g__2046(w__2540 ,w__2475 ,w__2317);
  xnor g__2047(w__2539 ,w__2497 ,w__2323);
  xor g__2048(w__2538 ,w__2498 ,w__2421);
  xnor g__2049(w__2537 ,w__2477 ,w__2420);
  and g__2050(w__2559 ,w__2485 ,w__2502);
  xnor g__2051(w__2558 ,w__2346 ,w__2462);
  xnor g__2052(w__2556 ,w__2495 ,w__2464);
  xnor g__2053(w__2555 ,w__2336 ,w__2463);
  xnor g__2054(w__2553 ,w__2348 ,w__2461);
  xnor g__2055(w__2552 ,w__2424 ,w__2459);
  xnor g__2056(w__2550 ,w__2354 ,w__2458);
  xnor g__2057(w__2549 ,w__2426 ,w__2465);
  xnor g__2058(w__2547 ,w__2393 ,w__2460);
  xnor g__2059(w__2546 ,w__2352 ,w__2466);
  not g__2060(w__2526 ,w__2527);
  not g__2061(w__2525 ,w__2524);
  not g__2062(w__2522 ,w__2521);
  or g__2063(w__2520 ,w__2495 ,w__2444);
  and g__2064(w__2519 ,w__2317 ,w__2475);
  or g__2065(w__2518 ,w__2317 ,w__2475);
  and g__2066(w__2536 ,w__2442 ,w__2480);
  and g__2067(w__2535 ,w__2441 ,w__2478);
  and g__2068(w__2534 ,w__2410 ,w__2468);
  and g__2069(w__2533 ,w__2443 ,w__2479);
  and g__2070(w__2532 ,w__2432 ,w__2482);
  and g__2071(w__2531 ,w__2433 ,w__2487);
  and g__2072(w__2530 ,w__2428 ,w__2472);
  and g__2073(w__2529 ,w__2416 ,w__2471);
  and g__2074(w__2528 ,w__2409 ,w__2470);
  and g__2075(w__2527 ,w__2373 ,w__2484);
  and g__2076(w__2524 ,w__2437 ,w__2486);
  and g__2077(w__2523 ,w__2413 ,w__2469);
  and g__2078(w__2521 ,w__2451 ,w__2490);
  not g__2079(w__2513 ,w__2514);
  not g__2080(w__2512 ,w__2511);
  or g__2081(w__2502 ,w__2496 ,w__2483);
  xnor g__2082(w__2501 ,w__2350 ,w__2419);
  xnor g__2083(w__2500 ,w__2280 ,w__2423);
  xnor g__2084(w__2499 ,w__2455 ,w__2345);
  xnor g__2085(w__2517 ,w__2326 ,w__2397);
  and g__2086(w__2516 ,w__2406 ,w__2491);
  xnor g__2087(w__2515 ,w__2353 ,w__2402);
  xnor g__2088(w__2514 ,w__2361 ,w__2401);
  xnor g__2089(w__2511 ,w__2363 ,w__2403);
  xnor g__2090(w__2510 ,w__2330 ,w__2405);
  xnor g__2091(w__2509 ,w__2456 ,w__2395);
  xnor g__2092(w__2508 ,w__2355 ,w__2394);
  xnor g__2093(w__2507 ,w__2283 ,w__2400);
  xnor g__2094(w__2506 ,w__2340 ,w__2396);
  xnor g__2095(w__2505 ,w__2327 ,w__2398);
  xnor g__2096(w__2504 ,w__2337 ,w__2399);
  xnor g__2097(w__2503 ,w__2338 ,w__2404);
  not g__2098(w__2493 ,w__2494);
  or g__2099(w__2492 ,w__2345 ,w__2455);
  or g__2100(w__2491 ,w__2333 ,w__2449);
  or g__2101(w__2490 ,w__2450 ,w__2427);
  nor g__2102(w__2489 ,w__2280 ,w__2422);
  or g__2103(w__2488 ,w__2279 ,w__2423);
  or g__2104(w__2487 ,w__2324 ,w__2431);
  or g__2105(w__2486 ,w__2425 ,w__2435);
  or g__2106(w__2485 ,w__2350 ,w__2418);
  or g__2107(w__2484 ,w__2376 ,w__2456);
  nor g__2108(w__2483 ,w__2349 ,w__2419);
  or g__2109(w__2482 ,w__2331 ,w__2434);
  and g__2110(w__2481 ,w__2345 ,w__2455);
  or g__2111(w__2480 ,w__2332 ,w__2417);
  or g__2112(w__2479 ,w__2328 ,w__2436);
  or g__2113(w__2478 ,w__2329 ,w__2438);
  and g__2114(w__2498 ,w__2382 ,w__2447);
  and g__2115(w__2497 ,w__2377 ,w__2430);
  and g__2116(w__2496 ,w__2313 ,w__2446);
  and g__2117(w__2495 ,w__2383 ,w__2445);
  and g__2118(w__2494 ,w__2384 ,w__2448);
  not g__2119(w__2474 ,w__2473);
  or g__2120(w__2472 ,w__2362 ,w__2429);
  xnor g__2121(w__8466 ,w__2391 ,w__2364);
  or g__2122(w__2471 ,w__2360 ,w__2414);
  or g__2123(w__2470 ,w__2308 ,w__2408);
  or g__2124(w__2469 ,w__2393 ,w__2411);
  or g__2125(w__2468 ,w__2309 ,w__2407);
  xnor g__2126(w__2467 ,w__2358 ,w__2385);
  xnor g__2127(w__2466 ,w__2360 ,w__2351);
  xnor g__2128(w__2465 ,w__2387 ,w__2341);
  xnor g__2129(w__2464 ,w__2342 ,w__2386);
  xnor g__2130(w__2463 ,w__2347 ,w__2332);
  xnor g__2131(w__2462 ,w__2339 ,w__2309);
  xnor g__2132(w__2461 ,w__2359 ,w__2329);
  xnor g__2133(w__2460 ,w__2343 ,w__2344);
  xnor g__2134(w__2459 ,w__2356 ,w__2357);
  xnor g__2135(w__2458 ,w__2362 ,w__2320);
  and g__2136(w__2477 ,w__2369 ,w__2412);
  and g__2137(w__2476 ,w__2372 ,w__2415);
  xnor g__2138(w__2475 ,w__2325 ,w__2334);
  xnor g__2139(w__2473 ,w__2307 ,w__2365);
  or g__2140(w__2452 ,w__2386 ,w__2342);
  or g__2141(w__2451 ,w__2341 ,w__2387);
  and g__2142(w__2450 ,w__2341 ,w__2387);
  and g__2143(w__2449 ,w__2300 ,w__2353);
  or g__2144(w__2448 ,w__2379 ,w__2361);
  or g__2145(w__2447 ,w__2326 ,w__2380);
  or g__2146(w__2446 ,w__2290 ,w__2392);
  or g__2147(w__2445 ,w__2330 ,w__2378);
  and g__2148(w__2444 ,w__2386 ,w__2342);
  or g__2149(w__2443 ,w__2318 ,w__2340);
  or g__2150(w__2442 ,w__2336 ,w__2347);
  or g__2151(w__2441 ,w__2348 ,w__2359);
  or g__2152(w__2440 ,w__2385 ,w__2358);
  and g__2153(w__2439 ,w__2385 ,w__2358);
  and g__2154(w__2438 ,w__2348 ,w__2359);
  or g__2155(w__2437 ,w__2357 ,w__2356);
  and g__2156(w__2436 ,w__2318 ,w__2340);
  and g__2157(w__2435 ,w__2357 ,w__2356);
  and g__2158(w__2434 ,w__2296 ,w__2337);
  or g__2159(w__2433 ,w__2321 ,w__2355);
  or g__2160(w__2432 ,w__2296 ,w__2337);
  and g__2161(w__2431 ,w__2321 ,w__2355);
  or g__2162(w__2430 ,w__2327 ,w__2374);
  and g__2163(w__2429 ,w__2320 ,w__2354);
  or g__2164(w__2428 ,w__2320 ,w__2354);
  and g__2165(w__2457 ,w__2241 ,w__2368);
  and g__2166(w__2456 ,w__2131 ,w__2367);
  and g__2167(w__2455 ,w__2140 ,w__2381);
  and g__2168(w__2454 ,w__2291 ,w__2371);
  and g__2169(w__2453 ,w__2312 ,w__2375);
  not g__2170(w__2427 ,w__2426);
  not g__2171(w__2425 ,w__2424);
  not g__2172(w__2422 ,w__2423);
  not g__2173(w__2418 ,w__2419);
  and g__2174(w__2417 ,w__2336 ,w__2347);
  or g__2175(w__2416 ,w__2351 ,w__2352);
  or g__2176(w__2415 ,w__2370 ,w__2363);
  and g__2177(w__2414 ,w__2351 ,w__2352);
  or g__2178(w__2413 ,w__2344 ,w__2343);
  or g__2179(w__2412 ,w__2283 ,w__2366);
  and g__2180(w__2411 ,w__2344 ,w__2343);
  or g__2181(w__2410 ,w__2346 ,w__2339);
  or g__2182(w__2409 ,w__2299 ,w__2338);
  and g__2183(w__2408 ,w__2299 ,w__2338);
  and g__2184(w__2407 ,w__2346 ,w__2339);
  or g__2185(w__2406 ,w__2300 ,w__2353);
  xnor g__2186(w__2405 ,w__2075 ,w__2298);
  xnor g__2187(w__2404 ,w__2308 ,w__2299);
  xnor g__2188(w__2403 ,w__2204 ,w__2294);
  xnor g__2189(w__2402 ,w__2300 ,w__2333);
  xnor g__2190(w__2401 ,w__2316 ,w__1741);
  xnor g__2191(w__2400 ,w__2297 ,w__2301);
  xnor g__2192(w__2399 ,w__2296 ,w__2331);
  xnor g__2193(w__2398 ,w__2322 ,w__2319);
  xnor g__2194(w__2397 ,w__2292 ,w__1742);
  xnor g__2195(w__2396 ,w__2328 ,w__2318);
  xnor g__2196(w__2395 ,w__1989 ,w__2295);
  xnor g__2197(w__2394 ,w__2321 ,w__2324);
  xnor g__2198(w__2426 ,w__2305 ,w__2284);
  xnor g__2199(w__2424 ,w__2205 ,w__2285);
  xnor g__2200(w__2423 ,w__2306 ,w__2216);
  xor g__2201(w__2421 ,w__2159 ,w__2287);
  xnor g__2202(w__2420 ,w__2302 ,w__2208);
  xnor g__2203(w__2419 ,w__2158 ,w__2286);
  not g__2204(w__2392 ,w__2391);
  not g__2205(w__2388 ,w__2389);
  or g__2206(w__2384 ,w__1741 ,w__2316);
  or g__2207(w__2383 ,w__2075 ,w__2298);
  or g__2208(w__2382 ,w__1742 ,w__2292);
  or g__2209(w__2381 ,w__2177 ,w__2302);
  and g__2210(w__2380 ,w__1742 ,w__2292);
  and g__2211(w__2379 ,w__1741 ,w__2316);
  and g__2212(w__2378 ,w__2075 ,w__2298);
  or g__2213(w__2377 ,w__2319 ,w__2322);
  and g__2214(w__2376 ,w__1989 ,w__2295);
  or g__2215(w__2375 ,w__2325 ,w__2310);
  and g__2216(w__2374 ,w__2319 ,w__2322);
  or g__2217(w__2373 ,w__1989 ,w__2295);
  or g__2218(w__2372 ,w__2203 ,w__2294);
  or g__2219(w__2371 ,w__2288 ,w__2307);
  nor g__2220(w__2370 ,w__2204 ,w__2293);
  or g__2221(w__2369 ,w__2301 ,w__2297);
  or g__2222(w__2368 ,w__2273 ,w__2305);
  or g__2223(w__2367 ,w__2165 ,w__2306);
  and g__2224(w__2366 ,w__2301 ,w__2297);
  xnor g__2225(w__2365 ,w__1991 ,w__2277);
  xnor g__2226(w__2364 ,w__1740 ,w__2278);
  and g__2227(w__2393 ,w__2133 ,w__2289);
  and g__2228(w__2391 ,w__2046 ,w__2304);
  and g__2229(w__2390 ,w__2264 ,w__2315);
  or g__2230(w__2389 ,w__2270 ,w__2314);
  xnor g__2231(w__2387 ,w__2061 ,w__2236);
  xnor g__2232(w__2386 ,w__2116 ,w__2230);
  and g__2233(w__2385 ,w__2262 ,w__2311);
  not g__2234(w__2349 ,w__2350);
  xnor g__2235(w__2334 ,w__2013 ,w__1743);
  xnor g__2236(w__2363 ,w__2093 ,w__2207);
  xnor g__2237(w__2362 ,w__2034 ,w__2211);
  xnor g__2238(w__2361 ,w__2103 ,w__2209);
  xnor g__2239(w__2360 ,w__2098 ,w__2220);
  xnor g__2240(w__2359 ,w__2071 ,w__2222);
  xnor g__2241(w__2358 ,w__2036 ,w__2221);
  xnor g__2242(w__2357 ,w__2104 ,w__2219);
  xnor g__2243(w__2356 ,w__2099 ,w__2217);
  xnor g__2244(w__2355 ,w__2094 ,w__2213);
  xnor g__2245(w__2354 ,w__2080 ,w__2238);
  xnor g__2246(w__2353 ,w__2107 ,w__2228);
  xnor g__2247(w__2352 ,w__2020 ,w__2225);
  xnor g__2248(w__2351 ,w__2035 ,w__2229);
  xnor g__2249(w__2350 ,w__1994 ,w__2233);
  xnor g__2250(w__2348 ,w__2000 ,w__2224);
  xnor g__2251(w__2347 ,w__2023 ,w__2226);
  xnor g__2252(w__2346 ,w__2039 ,w__2210);
  xnor g__2253(w__2345 ,w__2040 ,w__2231);
  xnor g__2254(w__2344 ,w__2033 ,w__2215);
  xnor g__2255(w__2343 ,w__2161 ,w__2234);
  xnor g__2256(w__2342 ,w__2092 ,w__2235);
  xnor g__2257(w__2341 ,w__2115 ,w__2218);
  xnor g__2258(w__2340 ,w__2106 ,w__2223);
  xnor g__2259(w__2339 ,w__2102 ,w__2212);
  xnor g__2260(w__2338 ,w__1993 ,w__2227);
  xnor g__2261(w__2337 ,w__2037 ,w__2214);
  xnor g__2262(w__2336 ,w__2105 ,w__2237);
  xnor g__2263(w__2335 ,w__1739 ,w__2232);
  or g__2264(w__2315 ,w__2160 ,w__2242);
  and g__2265(w__2314 ,w__2158 ,w__2239);
  or g__2266(w__2313 ,w__2278 ,w__1740);
  or g__2267(w__2312 ,w__2013 ,w__1743);
  or g__2268(w__2311 ,w__2206 ,w__2261);
  and g__2269(w__2310 ,w__2013 ,w__1743);
  and g__2270(w__2333 ,w__2187 ,w__2274);
  and g__2271(w__2332 ,w__2126 ,w__2265);
  and g__2272(w__2331 ,w__2183 ,w__2257);
  and g__2273(w__2330 ,w__2198 ,w__2263);
  and g__2274(w__2329 ,w__2128 ,w__2260);
  and g__2275(w__2328 ,w__2137 ,w__2275);
  and g__2276(w__2327 ,w__2185 ,w__2249);
  and g__2277(w__2326 ,w__2188 ,w__2269);
  and g__2278(w__2325 ,w__2146 ,w__2248);
  and g__2279(w__2324 ,w__2166 ,w__2251);
  and g__2280(w__2323 ,w__2171 ,w__2256);
  and g__2281(w__2322 ,w__2163 ,w__2250);
  and g__2282(w__2321 ,w__2178 ,w__2253);
  and g__2283(w__2320 ,w__2194 ,w__2247);
  and g__2284(w__2319 ,w__2167 ,w__2252);
  and g__2285(w__2318 ,w__2123 ,w__2243);
  and g__2286(w__2317 ,w__2147 ,w__2246);
  and g__2287(w__2316 ,w__2138 ,w__2272);
  not g__2288(w__2304 ,w__2303);
  not g__2289(w__2293 ,w__2294);
  or g__2290(w__2291 ,w__1991 ,w__2276);
  and g__2291(w__2290 ,w__2278 ,w__1740);
  or g__2292(w__2289 ,w__2193 ,w__1739);
  nor g__2293(w__2288 ,w__1990 ,w__2277);
  xnor g__2294(w__2287 ,w__2082 ,w__2157);
  xnor g__2295(w__2286 ,w__2002 ,w__2153);
  xnor g__2296(w__2285 ,w__2021 ,w__2154);
  xnor g__2297(w__2284 ,w__2202 ,w__2156);
  and g__2298(w__2309 ,w__2189 ,w__2268);
  and g__2299(w__2308 ,w__2124 ,w__2254);
  and g__2300(w__2307 ,w__2151 ,w__2245);
  and g__2301(w__2306 ,w__2184 ,w__2266);
  and g__2302(w__2305 ,w__2129 ,w__2240);
  xnor g__2303(w__2303 ,w__2091 ,w__2117);
  xnor g__2304(w__2302 ,w__2108 ,w__2121);
  and g__2305(w__2301 ,w__2144 ,w__2255);
  and g__2306(w__2300 ,w__2122 ,w__2258);
  and g__2307(w__2299 ,w__2181 ,w__2267);
  xnor g__2308(w__2298 ,w__2029 ,w__2120);
  and g__2309(w__2297 ,w__2168 ,w__2259);
  xnor g__2310(w__2296 ,w__2038 ,w__2119);
  xnor g__2311(w__2295 ,w__2041 ,w__2118);
  and g__2312(w__2294 ,w__2143 ,w__2271);
  and g__2313(w__2292 ,w__2142 ,w__2244);
  not g__2314(w__2282 ,w__2281);
  not g__2315(w__2279 ,w__2280);
  not g__2316(w__2276 ,w__2277);
  or g__2317(w__2275 ,w__2092 ,w__2130);
  or g__2318(w__2274 ,w__2043 ,w__2186);
  nor g__2319(w__2273 ,w__2202 ,w__2155);
  or g__2320(w__2272 ,w__2031 ,w__2150);
  or g__2321(w__2271 ,w__2032 ,w__2176);
  nor g__2322(w__2270 ,w__2002 ,w__2153);
  or g__2323(w__2269 ,w__2099 ,w__2191);
  or g__2324(w__2268 ,w__2036 ,w__2180);
  or g__2325(w__2267 ,w__2115 ,w__2125);
  or g__2326(w__2266 ,w__2037 ,w__2197);
  or g__2327(w__2265 ,w__2094 ,w__2173);
  or g__2328(w__2264 ,w__2082 ,w__2157);
  or g__2329(w__2263 ,w__2035 ,w__2182);
  or g__2330(w__2262 ,w__2021 ,w__2154);
  and g__2331(w__2261 ,w__2021 ,w__2154);
  or g__2332(w__2260 ,w__2044 ,w__2172);
  or g__2333(w__2259 ,w__2030 ,w__2200);
  or g__2334(w__2258 ,w__2105 ,w__2175);
  or g__2335(w__2257 ,w__2040 ,w__2196);
  or g__2336(w__2256 ,w__2098 ,w__2179);
  or g__2337(w__2255 ,w__2097 ,w__2132);
  or g__2338(w__2254 ,w__2045 ,w__2145);
  or g__2339(w__2253 ,w__2034 ,w__2190);
  or g__2340(w__2252 ,w__2039 ,w__2127);
  or g__2341(w__2251 ,w__2048 ,w__2139);
  or g__2342(w__2250 ,w__2102 ,w__2135);
  or g__2343(w__2249 ,w__2107 ,w__2169);
  or g__2344(w__2248 ,w__2093 ,w__2174);
  or g__2345(w__2247 ,w__2033 ,w__2192);
  or g__2346(w__2246 ,w__2195 ,w__2161);
  or g__2347(w__2245 ,w__2106 ,w__2164);
  or g__2348(w__2244 ,w__2104 ,w__2149);
  or g__2349(w__2243 ,w__2116 ,w__2162);
  and g__2350(w__2242 ,w__2082 ,w__2157);
  and g__2351(w__2283 ,w__1986 ,w__2134);
  or g__2352(w__2281 ,w__1987 ,w__2148);
  or g__2353(w__2280 ,w__2049 ,w__2136);
  and g__2354(w__2278 ,w__2054 ,w__2170);
  or g__2355(w__2277 ,w__1988 ,w__2141);
  or g__2356(w__2241 ,w__2156 ,w__2201);
  or g__2357(w__2240 ,w__2103 ,w__2199);
  or g__2358(w__2239 ,w__2001 ,w__2152);
  xnor g__2359(w__2238 ,w__2012 ,w__2048);
  xnor g__2360(w__2237 ,w__2007 ,w__2017);
  xnor g__2361(w__2236 ,w__2072 ,w__2045);
  xnor g__2362(w__2235 ,w__2064 ,w__2005);
  xnor g__2363(w__2234 ,w__2058 ,w__2022);
  xnor g__2364(w__2233 ,w__2015 ,w__2031);
  xnor g__2365(w__2232 ,w__2066 ,w__2076);
  xnor g__2366(w__2231 ,w__2014 ,w__1998);
  xnor g__2367(w__2230 ,w__2077 ,w__2063);
  xnor g__2368(w__2229 ,w__2060 ,w__2074);
  xnor g__2369(w__2228 ,w__2011 ,w__2019);
  xnor g__2370(w__2227 ,w__2067 ,w__2032);
  xnor g__2371(w__2226 ,w__2055 ,w__2043);
  xnor g__2372(w__2225 ,w__2057 ,w__2044);
  xnor g__2373(w__2224 ,w__2084 ,w__2030);
  xnor g__2374(w__2223 ,w__1999 ,w__2073);
  xnor g__2375(w__2222 ,w__2090 ,w__2097);
  xnor g__2376(w__2221 ,w__2003 ,w__2070);
  xnor g__2377(w__2220 ,w__2006 ,w__2009);
  xnor g__2378(w__2219 ,w__2016 ,w__2081);
  xnor g__2379(w__2218 ,w__1996 ,w__2065);
  xnor g__2380(w__2217 ,w__2008 ,w__1997);
  xnor g__2381(w__2216 ,w__2004 ,w__2068);
  xnor g__2382(w__2215 ,w__2059 ,w__2089);
  xnor g__2383(w__2214 ,w__2010 ,w__2085);
  xnor g__2384(w__2213 ,w__2087 ,w__1995);
  xnor g__2385(w__2212 ,w__2018 ,w__2069);
  xnor g__2386(w__2211 ,w__2062 ,w__2086);
  xnor g__2387(w__2210 ,w__1992 ,w__2056);
  xnor g__2388(w__2209 ,w__2078 ,w__2025);
  xnor g__2389(w__2208 ,w__2083 ,w__2024);
  xnor g__2390(w__2207 ,w__2088 ,w__2079);
  not g__2391(w__2206 ,w__2205);
  not g__2392(w__2203 ,w__2204);
  not g__2393(w__2201 ,w__2202);
  and g__2394(w__2200 ,w__2000 ,w__2084);
  and g__2395(w__2199 ,w__2078 ,w__2025);
  or g__2396(w__2198 ,w__2060 ,w__2074);
  and g__2397(w__2197 ,w__2010 ,w__2085);
  and g__2398(w__2196 ,w__2014 ,w__1998);
  and g__2399(w__2195 ,w__2058 ,w__2022);
  or g__2400(w__2194 ,w__2059 ,w__2089);
  and g__2401(w__2193 ,w__2066 ,w__2076);
  and g__2402(w__2192 ,w__2059 ,w__2089);
  and g__2403(w__2191 ,w__2008 ,w__1997);
  and g__2404(w__2190 ,w__2062 ,w__2086);
  or g__2405(w__2189 ,w__2003 ,w__2070);
  or g__2406(w__2188 ,w__2008 ,w__1997);
  or g__2407(w__2187 ,w__2023 ,w__2055);
  and g__2408(w__2186 ,w__2023 ,w__2055);
  or g__2409(w__2185 ,w__2011 ,w__2019);
  or g__2410(w__2184 ,w__2010 ,w__2085);
  or g__2411(w__2183 ,w__2014 ,w__1998);
  and g__2412(w__2182 ,w__2060 ,w__2074);
  or g__2413(w__2181 ,w__1996 ,w__2065);
  and g__2414(w__2180 ,w__2003 ,w__2070);
  and g__2415(w__2179 ,w__2006 ,w__2009);
  or g__2416(w__2178 ,w__2062 ,w__2086);
  and g__2417(w__2177 ,w__2083 ,w__2024);
  and g__2418(w__2176 ,w__1993 ,w__2067);
  and g__2419(w__2175 ,w__2007 ,w__2017);
  and g__2420(w__2174 ,w__2088 ,w__2079);
  and g__2421(w__2173 ,w__2087 ,w__1995);
  and g__2422(w__2172 ,w__2020 ,w__2057);
  or g__2423(w__2171 ,w__2006 ,w__2009);
  or g__2424(w__2170 ,w__2091 ,w__1985);
  and g__2425(w__2169 ,w__2011 ,w__2019);
  or g__2426(w__2168 ,w__2000 ,w__2084);
  or g__2427(w__2167 ,w__1992 ,w__2056);
  or g__2428(w__2166 ,w__2012 ,w__2080);
  and g__2429(w__2165 ,w__2004 ,w__2068);
  and g__2430(w__2164 ,w__1999 ,w__2073);
  or g__2431(w__2163 ,w__2018 ,w__2069);
  and g__2432(w__2162 ,w__2077 ,w__2063);
  and g__2433(w__2205 ,w__2047 ,w__2112);
  and g__2434(w__2204 ,w__2026 ,w__2096);
  and g__2435(w__2202 ,w__2028 ,w__2101);
  not g__2436(w__2160 ,w__2159);
  not g__2437(w__2155 ,w__2156);
  not g__2438(w__2152 ,w__2153);
  or g__2439(w__2151 ,w__1999 ,w__2073);
  xor g__2440(w__8463 ,in6[0] ,in7[0]);
  and g__2441(w__2150 ,w__1994 ,w__2015);
  and g__2442(w__2149 ,w__2016 ,w__2081);
  nor g__2443(w__2148 ,w__2041 ,w__2053);
  or g__2444(w__2147 ,w__2058 ,w__2022);
  or g__2445(w__2146 ,w__2088 ,w__2079);
  and g__2446(w__2145 ,w__2072 ,w__2061);
  or g__2447(w__2144 ,w__2090 ,w__2071);
  or g__2448(w__2143 ,w__1993 ,w__2067);
  or g__2449(w__2142 ,w__2016 ,w__2081);
  nor g__2450(w__2141 ,w__2108 ,w__2052);
  or g__2451(w__2140 ,w__2083 ,w__2024);
  and g__2452(w__2139 ,w__2012 ,w__2080);
  or g__2453(w__2138 ,w__1994 ,w__2015);
  or g__2454(w__2137 ,w__2064 ,w__2005);
  nor g__2455(w__2136 ,w__2038 ,w__2050);
  and g__2456(w__2135 ,w__2018 ,w__2069);
  or g__2457(w__2134 ,w__2029 ,w__2051);
  or g__2458(w__2133 ,w__2066 ,w__2076);
  and g__2459(w__2132 ,w__2090 ,w__2071);
  or g__2460(w__2131 ,w__2004 ,w__2068);
  and g__2461(w__2130 ,w__2064 ,w__2005);
  or g__2462(w__2129 ,w__2078 ,w__2025);
  or g__2463(w__2128 ,w__2020 ,w__2057);
  and g__2464(w__2127 ,w__1992 ,w__2056);
  or g__2465(w__2126 ,w__2087 ,w__1995);
  and g__2466(w__2125 ,w__1996 ,w__2065);
  or g__2467(w__2124 ,w__2072 ,w__2061);
  or g__2468(w__2123 ,w__2077 ,w__2063);
  or g__2469(w__2122 ,w__2007 ,w__2017);
  xnor g__2470(w__2121 ,in6[8] ,in7[8]);
  xnor g__2471(w__2120 ,in6[7] ,in7[7]);
  xnor g__2472(w__2119 ,in6[9] ,in7[9]);
  xnor g__2473(w__2118 ,in6[10] ,in7[10]);
  xnor g__2474(w__2117 ,in6[1] ,in7[1]);
  xnor g__2475(w__2161 ,in6[4] ,in7[4]);
  and g__2476(w__2159 ,w__2110 ,w__2042);
  and g__2477(w__2158 ,w__2114 ,w__2027);
  xnor g__2478(w__2157 ,in6[6] ,in7[6]);
  xnor g__2479(w__2156 ,in6[3] ,in7[3]);
  xnor g__2480(w__2154 ,in6[5] ,in7[5]);
  xnor g__2481(w__2153 ,in6[2] ,in7[2]);
  not g__2482(w__2114 ,w__2113);
  not g__2483(w__2112 ,w__2111);
  not g__2484(w__2110 ,w__2109);
  not g__2485(w__2101 ,w__2100);
  not g__2486(w__2096 ,w__2095);
  or g__2487(w__2054 ,w__1880 ,w__1839);
  nor g__2488(w__2053 ,in6[10] ,in7[10]);
  nor g__2489(w__2052 ,in6[8] ,in7[8]);
  nor g__2490(w__2051 ,in6[7] ,in7[7]);
  nor g__2491(w__2050 ,in6[9] ,in7[9]);
  and g__2492(w__2049 ,in6[9] ,in7[9]);
  or g__2493(w__2116 ,w__1808 ,w__1813);
  or g__2494(w__2115 ,w__1828 ,w__1831);
  or g__2495(w__2113 ,w__1837 ,w__1883);
  or g__2496(w__2111 ,w__1847 ,w__1849);
  or g__2497(w__2109 ,w__1770 ,w__1858);
  or g__2498(w__2108 ,w__1804 ,w__1811);
  or g__2499(w__2107 ,w__1785 ,w__1776);
  or g__2500(w__2106 ,w__1806 ,w__1860);
  or g__2501(w__2105 ,w__1871 ,w__1773);
  or g__2502(w__2104 ,w__1800 ,w__1764);
  or g__2503(w__2103 ,w__1909 ,w__1862);
  or g__2504(w__2102 ,w__1844 ,w__1892);
  or g__2505(w__2100 ,w__1856 ,w__1877);
  or g__2506(w__2099 ,w__1758 ,w__1919);
  or g__2507(w__2098 ,w__1767 ,w__1797);
  or g__2508(w__2097 ,w__1952 ,w__1761);
  or g__2509(w__2095 ,w__1818 ,w__1833);
  or g__2510(w__2094 ,w__1915 ,w__1886);
  or g__2511(w__2093 ,w__1943 ,w__1775);
  or g__2512(w__2092 ,w__1787 ,w__1864);
  or g__2513(w__2091 ,w__1773 ,w__1841);
  or g__2514(w__2090 ,w__1816 ,w__1912);
  or g__2515(w__2089 ,w__1851 ,w__1878);
  or g__2516(w__2088 ,w__1769 ,w__1924);
  or g__2517(w__2087 ,w__1767 ,w__1869);
  or g__2518(w__2086 ,w__1799 ,w__1926);
  or g__2519(w__2085 ,w__1752 ,w__1906);
  or g__2520(w__2084 ,w__1755 ,w__1782);
  or g__2521(w__2083 ,w__1824 ,w__1766);
  or g__2522(w__2082 ,w__1797 ,w__1779);
  or g__2523(w__2081 ,w__1941 ,w__1922);
  or g__2524(w__2080 ,w__1895 ,w__1928);
  or g__2525(w__2079 ,w__1781 ,w__1862);
  or g__2526(w__2078 ,w__1763 ,w__1772);
  or g__2527(w__2077 ,w__1802 ,w__1912);
  or g__2528(w__2076 ,w__1796 ,w__1917);
  or g__2529(w__2075 ,w__1746 ,w__1938);
  or g__2530(w__2074 ,w__1867 ,w__1901);
  or g__2531(w__2073 ,w__1949 ,w__1821);
  or g__2532(w__2072 ,w__1898 ,w__1881);
  or g__2533(w__2071 ,w__1853 ,w__1943);
  or g__2534(w__2070 ,w__1903 ,w__1761);
  or g__2535(w__2069 ,w__1757 ,w__1760);
  or g__2536(w__2068 ,w__1951 ,w__1754);
  or g__2537(w__2067 ,w__1794 ,w__1831);
  or g__2538(w__2066 ,w__1875 ,w__1928);
  or g__2539(w__2065 ,w__1946 ,w__1884);
  or g__2540(w__2064 ,w__1749 ,w__1856);
  or g__2541(w__2063 ,w__1826 ,w__1818);
  or g__2542(w__2062 ,w__1851 ,w__1834);
  or g__2543(w__2061 ,w__1791 ,w__1919);
  or g__2544(w__2060 ,w__1816 ,w__1811);
  or g__2545(w__2059 ,w__1858 ,w__1875);
  or g__2546(w__2058 ,w__1938 ,w__1849);
  or g__2547(w__2057 ,w__1936 ,w__1779);
  or g__2548(w__2056 ,w__1958 ,w__1979);
  or g__2549(w__2055 ,w__1955 ,w__1877);
  not g__2550(w__2002 ,w__2001);
  not g__2551(w__1991 ,w__1990);
  nor g__2552(w__1988 ,w__1958 ,w__1949);
  nor g__2553(w__1987 ,w__1955 ,w__1952);
  or g__2554(w__1986 ,w__1906 ,w__1853);
  nor g__2555(w__1985 ,in6[1] ,in7[1]);
  and g__2556(w__8464 ,in6[0] ,in7[0]);
  or g__2557(w__2048 ,w__1808 ,w__1887);
  and g__2558(w__2047 ,in6[5] ,in6[3]);
  and g__2559(w__2046 ,in6[1] ,in6[0]);
  or g__2560(w__2045 ,w__1778 ,w__1842);
  or g__2561(w__2044 ,w__1806 ,w__1892);
  or g__2562(w__2043 ,w__1788 ,w__1886);
  and g__2563(w__2042 ,in6[7] ,in6[3]);
  or g__2564(w__2041 ,w__1751 ,w__1931);
  or g__2565(w__2040 ,w__1785 ,w__1800);
  or g__2566(w__2039 ,w__1821 ,w__1889);
  or g__2567(w__2038 ,w__1872 ,w__1758);
  or g__2568(w__2037 ,w__1788 ,w__1903);
  or g__2569(w__2036 ,w__1946 ,w__1895);
  or g__2570(w__2035 ,w__1748 ,w__1837);
  or g__2571(w__2034 ,w__1936 ,w__1776);
  or g__2572(w__2033 ,w__1904 ,w__1917);
  or g__2573(w__2032 ,w__1782 ,w__1920);
  or g__2574(w__2031 ,w__1764 ,w__1887);
  or g__2575(w__2030 ,w__1845 ,w__1793);
  or g__2576(w__2029 ,w__1934 ,w__1901);
  and g__2577(w__2028 ,in6[3] ,in6[1]);
  and g__2578(w__2027 ,in7[2] ,in7[0]);
  and g__2579(w__2026 ,in6[4] ,in6[2]);
  or g__2580(w__2025 ,w__1791 ,w__1842);
  or g__2581(w__2024 ,w__1871 ,w__1944);
  or g__2582(w__2023 ,w__1745 ,w__1909);
  or g__2583(w__2022 ,w__1790 ,w__1929);
  or g__2584(w__2021 ,w__1896 ,w__1889);
  or g__2585(w__2020 ,w__1826 ,w__1874);
  or g__2586(w__2019 ,w__1804 ,w__1880);
  or g__2587(w__2018 ,w__1824 ,w__1922);
  or g__2588(w__2017 ,w__1755 ,w__1926);
  or g__2589(w__2016 ,w__1939 ,w__1898);
  or g__2590(w__2015 ,w__1893 ,w__1839);
  or g__2591(w__2014 ,w__1931 ,w__1941);
  or g__2592(w__2013 ,w__1855 ,w__1794);
  or g__2593(w__2012 ,w__1866 ,w__1883);
  or g__2594(w__2011 ,w__1907 ,w__1899);
  or g__2595(w__2010 ,w__1934 ,w__1802);
  or g__2596(w__2009 ,w__1915 ,w__1828);
  or g__2597(w__2008 ,w__1746 ,w__1924);
  or g__2598(w__2007 ,w__1932 ,w__1881);
  or g__2599(w__2006 ,w__1948 ,w__1890);
  or g__2600(w__2005 ,w__1872 ,w__1860);
  or g__2601(w__2004 ,w__1752 ,w__1867);
  or g__2602(w__2003 ,w__1813 ,w__1864);
  and g__2603(w__2001 ,in6[3] ,in6[0]);
  or g__2604(w__2000 ,w__1749 ,w__1869);
  or g__2605(w__1999 ,w__1957 ,w__1815);
  or g__2606(w__1998 ,w__1954 ,w__1770);
  or g__2607(w__1997 ,w__1820 ,w__1830);
  or g__2608(w__1996 ,w__1874 ,w__1910);
  or g__2609(w__1995 ,w__1823 ,w__1878);
  or g__2610(w__1994 ,w__1836 ,w__1834);
  or g__2611(w__1993 ,w__1913 ,w__1884);
  or g__2612(w__1992 ,w__1847 ,w__1810);
  and g__2613(w__1990 ,in7[9] ,in7[7]);
  or g__2614(w__1989 ,w__1784 ,w__1845);
  not g__2615(w__1984 ,in6[0]);
  not g__2616(w__1983 ,in7[0]);
  not g__2617(w__1982 ,in7[2]);
  not g__2618(w__1981 ,in7[6]);
  not g__2619(w__1980 ,in7[3]);
  not g__2620(w__1979 ,in6[3]);
  not g__2621(w__1978 ,in6[4]);
  not g__2622(w__1977 ,in6[5]);
  not g__2623(w__1976 ,in6[1]);
  not g__2624(w__1975 ,in7[1]);
  not g__2625(w__1974 ,in6[9]);
  not g__2626(w__1973 ,in6[6]);
  not g__2627(w__1972 ,in7[5]);
  not g__2628(w__1971 ,in6[2]);
  not g__2629(w__1970 ,in7[4]);
  not g__2630(w__1969 ,in7[7]);
  not g__2631(w__1968 ,in6[7]);
  not g__2632(w__1967 ,in6[8]);
  not g__2633(w__1966 ,in6[10]);
  not g__2634(w__1965 ,in7[10]);
  not g__2635(w__1964 ,in7[9]);
  not g__2636(w__1963 ,in7[8]);
  not g__2637(w__1960 ,w__1962);
  not g__2638(w__1962 ,w__2655);
  not g__2639(w__1959 ,w__1961);
  not g__2640(w__1961 ,w__2509);
  not g__2641(w__1958 ,w__1956);
  not g__2642(w__1957 ,w__1956);
  not g__2643(w__1956 ,w__1967);
  not g__2644(w__1955 ,w__1953);
  not g__2645(w__1954 ,w__1953);
  not g__2646(w__1953 ,w__1966);
  not g__2647(w__1952 ,w__1950);
  not g__2648(w__1951 ,w__1950);
  not g__2649(w__1950 ,w__1965);
  not g__2650(w__1949 ,w__1947);
  not g__2651(w__1948 ,w__1947);
  not g__2652(w__1947 ,w__1963);
  not g__2653(w__1946 ,w__1945);
  not g__2654(w__1945 ,w__1977);
  not g__2655(w__1944 ,w__1942);
  not g__2656(w__1943 ,w__1942);
  not g__2657(w__1942 ,w__1981);
  not g__2658(w__1941 ,w__1940);
  not g__2659(w__1940 ,w__1968);
  not g__2660(w__1939 ,w__1937);
  not g__2661(w__1938 ,w__1937);
  not g__2662(w__1937 ,w__1977);
  not g__2663(w__1936 ,w__1935);
  not g__2664(w__1935 ,w__1969);
  not g__2665(w__1934 ,w__1933);
  not g__2666(w__1933 ,w__1974);
  not g__2667(w__1932 ,w__1930);
  not g__2668(w__1931 ,w__1930);
  not g__2669(w__1930 ,w__1974);
  not g__2670(w__1929 ,w__1927);
  not g__2671(w__1928 ,w__1927);
  not g__2672(w__1927 ,w__1980);
  not g__2673(w__1926 ,w__1925);
  not g__2674(w__1925 ,w__1982);
  not g__2675(w__1924 ,w__1923);
  not g__2676(w__1923 ,w__1976);
  not g__2677(w__1922 ,w__1921);
  not g__2678(w__1921 ,w__1971);
  not g__2679(w__1920 ,w__1918);
  not g__2680(w__1919 ,w__1918);
  not g__2681(w__1918 ,w__1975);
  not g__2682(w__1917 ,w__1916);
  not g__2683(w__1916 ,w__1983);
  not g__2684(w__1915 ,w__1914);
  not g__2685(w__1914 ,w__1964);
  not g__2686(w__1913 ,w__1911);
  not g__2687(w__1912 ,w__1911);
  not g__2688(w__1911 ,w__1973);
  not g__2689(w__1910 ,w__1908);
  not g__2690(w__1909 ,w__1908);
  not g__2691(w__1908 ,w__1971);
  not g__2692(w__1907 ,w__1905);
  not g__2693(w__1906 ,w__1905);
  not g__2694(w__1905 ,w__1968);
  not g__2695(w__1904 ,w__1902);
  not g__2696(w__1903 ,w__1902);
  not g__2697(w__1902 ,w__1969);
  not g__2698(w__1901 ,w__1900);
  not g__2699(w__1900 ,w__1978);
  not g__2700(w__1899 ,w__1897);
  not g__2701(w__1898 ,w__1897);
  not g__2702(w__1897 ,w__1978);
  not g__2703(w__1896 ,w__1894);
  not g__2704(w__1895 ,w__1894);
  not g__2705(w__1894 ,w__1972);
  not g__2706(w__1893 ,w__1891);
  not g__2707(w__1892 ,w__1891);
  not g__2708(w__1891 ,w__1982);
  not g__2709(w__1890 ,w__1888);
  not g__2710(w__1889 ,w__1888);
  not g__2711(w__1888 ,w__1970);
  not g__2712(w__1887 ,w__1885);
  not g__2713(w__1886 ,w__1885);
  not g__2714(w__1885 ,w__1983);
  not g__2715(w__1884 ,w__1882);
  not g__2716(w__1883 ,w__1882);
  not g__2717(w__1882 ,w__1984);
  not g__2718(w__1881 ,w__1879);
  not g__2719(w__1880 ,w__1879);
  not g__2720(w__1879 ,w__1976);
  not g__2721(w__1878 ,w__1876);
  not g__2722(w__1877 ,w__1876);
  not g__2723(w__1876 ,w__1984);
  not g__2724(w__1875 ,w__1873);
  not g__2725(w__1874 ,w__1873);
  not g__2726(w__1873 ,w__1979);
  not g__2727(w__1872 ,w__1870);
  not g__2728(w__1871 ,w__1870);
  not g__2729(w__1870 ,w__1964);
  not g__2730(w__1869 ,w__1868);
  not g__2731(w__1868 ,w__1979);
  not g__2732(w__1867 ,w__1865);
  not g__2733(w__1866 ,w__1865);
  not g__2734(w__1865 ,w__1967);
  not g__2735(w__1864 ,w__1863);
  not g__2736(w__1863 ,w__1890);
  not g__2737(w__1862 ,w__1861);
  not g__2738(w__1861 ,w__1893);
  not g__2739(w__1860 ,w__1859);
  not g__2740(w__1859 ,w__1896);
  not g__2741(w__1858 ,w__1857);
  not g__2742(w__1857 ,w__1899);
  not g__2743(w__1856 ,w__1854);
  not g__2744(w__1855 ,w__1854);
  not g__2745(w__1854 ,w__1978);
  not g__2746(w__1853 ,w__1852);
  not g__2747(w__1852 ,w__1904);
  not g__2748(w__1851 ,w__1850);
  not g__2749(w__1850 ,w__1907);
  not g__2750(w__1849 ,w__1848);
  not g__2751(w__1848 ,w__1910);
  not g__2752(w__1847 ,w__1846);
  not g__2753(w__1846 ,w__1913);
  not g__2754(w__1845 ,w__1843);
  not g__2755(w__1844 ,w__1843);
  not g__2756(w__1843 ,w__1964);
  not g__2757(w__1842 ,w__1840);
  not g__2758(w__1841 ,w__1840);
  not g__2759(w__1840 ,w__1983);
  not g__2760(w__1839 ,w__1838);
  not g__2761(w__1838 ,w__1920);
  not g__2762(w__1837 ,w__1835);
  not g__2763(w__1836 ,w__1835);
  not g__2764(w__1835 ,w__1971);
  not g__2765(w__1834 ,w__1832);
  not g__2766(w__1833 ,w__1832);
  not g__2767(w__1832 ,w__1976);
  not g__2768(w__1831 ,w__1829);
  not g__2769(w__1830 ,w__1829);
  not g__2770(w__1829 ,w__1982);
  not g__2771(w__1828 ,w__1827);
  not g__2772(w__1827 ,w__1929);
  not g__2773(w__1826 ,w__1825);
  not g__2774(w__1825 ,w__1932);
  not g__2775(w__1824 ,w__1822);
  not g__2776(w__1823 ,w__1822);
  not g__2777(w__1822 ,w__1974);
  not g__2778(w__1821 ,w__1819);
  not g__2779(w__1820 ,w__1819);
  not g__2780(w__1819 ,w__1969);
  not g__2781(w__1818 ,w__1817);
  not g__2782(w__1817 ,w__1939);
  not g__2783(w__1816 ,w__1814);
  not g__2784(w__1815 ,w__1814);
  not g__2785(w__1814 ,w__1968);
  not g__2786(w__1813 ,w__1812);
  not g__2787(w__1812 ,w__1944);
  not g__2788(w__1811 ,w__1809);
  not g__2789(w__1810 ,w__1809);
  not g__2790(w__1809 ,w__1977);
  not g__2791(w__1808 ,w__1807);
  not g__2792(w__1807 ,w__1948);
  not g__2793(w__1806 ,w__1805);
  not g__2794(w__1805 ,w__1951);
  not g__2795(w__1804 ,w__1803);
  not g__2796(w__1803 ,w__1954);
  not g__2797(w__1802 ,w__1801);
  not g__2798(w__1801 ,w__1957);
  not g__2799(w__1800 ,w__1798);
  not g__2800(w__1799 ,w__1798);
  not g__2801(w__1798 ,w__1981);
  not g__2802(w__1797 ,w__1795);
  not g__2803(w__1796 ,w__1795);
  not g__2804(w__1795 ,w__1981);
  not g__2805(w__1794 ,w__1792);
  not g__2806(w__1793 ,w__1792);
  not g__2807(w__1792 ,w__1970);
  not g__2808(w__1791 ,w__1789);
  not g__2809(w__1790 ,w__1789);
  not g__2810(w__1789 ,w__1970);
  not g__2811(w__1788 ,w__1786);
  not g__2812(w__1787 ,w__1786);
  not g__2813(w__1786 ,w__1965);
  not g__2814(w__1785 ,w__1783);
  not g__2815(w__1784 ,w__1783);
  not g__2816(w__1783 ,w__1965);
  not g__2817(w__1782 ,w__1780);
  not g__2818(w__1781 ,w__1780);
  not g__2819(w__1780 ,w__1972);
  not g__2820(w__1779 ,w__1777);
  not g__2821(w__1778 ,w__1777);
  not g__2822(w__1777 ,w__1972);
  not g__2823(w__1776 ,w__1774);
  not g__2824(w__1775 ,w__1774);
  not g__2825(w__1774 ,w__1975);
  not g__2826(w__1773 ,w__1771);
  not g__2827(w__1772 ,w__1771);
  not g__2828(w__1771 ,w__1975);
  not g__2829(w__1770 ,w__1768);
  not g__2830(w__1769 ,w__1768);
  not g__2831(w__1768 ,w__1973);
  not g__2832(w__1767 ,w__1765);
  not g__2833(w__1766 ,w__1765);
  not g__2834(w__1765 ,w__1973);
  not g__2835(w__1764 ,w__1762);
  not g__2836(w__1763 ,w__1762);
  not g__2837(w__1762 ,w__1980);
  not g__2838(w__1761 ,w__1759);
  not g__2839(w__1760 ,w__1759);
  not g__2840(w__1759 ,w__1980);
  not g__2841(w__1758 ,w__1756);
  not g__2842(w__1757 ,w__1756);
  not g__2843(w__1756 ,w__1963);
  not g__2844(w__1755 ,w__1753);
  not g__2845(w__1754 ,w__1753);
  not g__2846(w__1753 ,w__1963);
  not g__2847(w__1752 ,w__1750);
  not g__2848(w__1751 ,w__1750);
  not g__2849(w__1750 ,w__1966);
  not g__2850(w__1749 ,w__1747);
  not g__2851(w__1748 ,w__1747);
  not g__2852(w__1747 ,w__1966);
  not g__2853(w__1746 ,w__1744);
  not g__2854(w__1745 ,w__1744);
  not g__2855(w__1744 ,w__1967);
  xor g__2856(w__8478 ,w__2788 ,w__2769);
  xor g__2857(w__8477 ,w__2786 ,w__2776);
  xor g__2858(w__8476 ,w__2784 ,w__2777);
  xor g__2859(w__8475 ,w__2782 ,w__2768);
  xor g__2860(w__8474 ,w__2780 ,w__2757);
  xor g__2861(w__8472 ,w__2761 ,w__2726);
  xor g__2862(w__1743 ,w__2047 ,w__2111);
  xnor g__2863(w__8465 ,w__2046 ,w__2303);
  xor g__2864(w__1742 ,w__2109 ,w__2042);
  xor g__2865(w__1741 ,w__2028 ,w__2100);
  xor g__2866(w__1740 ,w__2113 ,w__2027);
  xor g__2867(w__1739 ,w__2026 ,w__2095);
  xnor g__2868(w__8461 ,w__3478 ,w__2927);
  and g__2869(w__8462 ,w__2927 ,w__3479);
  not g__2870(w__3479 ,w__3478);
  and g__2871(w__3478 ,w__3180 ,w__3477);
  or g__2872(w__3477 ,w__3165 ,w__3476);
  and g__2873(w__3476 ,w__3277 ,w__3475);
  or g__2874(w__3475 ,w__3276 ,w__3474);
  and g__2875(w__3474 ,w__3325 ,w__3473);
  or g__2876(w__3473 ,w__3327 ,w__3472);
  and g__2877(w__3472 ,w__3382 ,w__3471);
  or g__2878(w__3471 ,w__3374 ,w__3470);
  and g__2879(w__3470 ,w__3408 ,w__3469);
  or g__2880(w__3469 ,w__3409 ,w__3468);
  and g__2881(w__3468 ,w__3416 ,w__3467);
  or g__2882(w__3467 ,w__3415 ,w__3466);
  and g__2883(w__3466 ,w__3440 ,w__3465);
  or g__2884(w__3465 ,w__3441 ,w__3464);
  and g__2885(w__3464 ,w__3447 ,w__3463);
  or g__2886(w__3463 ,w__3446 ,w__3462);
  and g__2887(w__3462 ,w__3439 ,w__3461);
  or g__2888(w__3461 ,w__3438 ,w__3460);
  and g__2889(w__3460 ,w__3437 ,w__3459);
  or g__2890(w__3459 ,w__3436 ,w__3458);
  and g__2891(w__3458 ,w__3427 ,w__3457);
  or g__2892(w__3457 ,w__3426 ,w__3456);
  and g__2893(w__3456 ,w__3413 ,w__3455);
  xnor g__2894(w__8449 ,w__3453 ,w__3420);
  or g__2895(w__3455 ,w__3407 ,w__3454);
  not g__2896(w__3454 ,w__3453);
  or g__2897(w__3453 ,w__3388 ,w__3452);
  xnor g__2898(w__8448 ,w__3451 ,w__3405);
  and g__2899(w__3452 ,w__3395 ,w__3451);
  or g__2900(w__3451 ,w__3365 ,w__3450);
  xnor g__2901(w__8447 ,w__3448 ,w__3373);
  and g__2902(w__3450 ,w__3364 ,w__3448);
  xnor g__2903(w__3449 ,w__3429 ,w__3435);
  or g__2904(w__3448 ,w__3343 ,w__3442);
  or g__2905(w__3447 ,w__3428 ,w__3434);
  nor g__2906(w__3446 ,w__3429 ,w__3435);
  xnor g__2907(w__3445 ,w__3431 ,w__3411);
  xnor g__2908(w__3444 ,w__3399 ,w__3423);
  xnor g__2909(w__3443 ,w__3401 ,w__3425);
  xnor g__2910(w__8446 ,w__3432 ,w__3351);
  and g__2911(w__3442 ,w__3342 ,w__3432);
  nor g__2912(w__3441 ,w__3431 ,w__3411);
  or g__2913(w__3440 ,w__3430 ,w__3410);
  or g__2914(w__3439 ,w__3398 ,w__3422);
  nor g__2915(w__3438 ,w__3399 ,w__3423);
  or g__2916(w__3437 ,w__3400 ,w__3424);
  nor g__2917(w__3436 ,w__3401 ,w__3425);
  not g__2918(w__3435 ,w__3434);
  xnor g__2919(w__3434 ,w__3359 ,w__3406);
  xnor g__2920(w__3433 ,w__3412 ,w__3403);
  not g__2921(w__3430 ,w__3431);
  not g__2922(w__3428 ,w__3429);
  or g__2923(w__3427 ,w__3403 ,w__3412);
  and g__2924(w__3426 ,w__3403 ,w__3412);
  or g__2925(w__3432 ,w__3312 ,w__3417);
  or g__2926(w__3431 ,w__3397 ,w__3414);
  or g__2927(w__3429 ,w__3338 ,w__3418);
  not g__2928(w__3425 ,w__3424);
  not g__2929(w__3423 ,w__3422);
  xnor g__2930(w__8445 ,w__3404 ,w__3322);
  xnor g__2931(w__3421 ,w__3389 ,w__3402);
  xnor g__2932(w__3420 ,w__3386 ,w__3393);
  xnor g__2933(w__3419 ,w__3384 ,w__3391);
  xnor g__2934(w__3424 ,w__3331 ,w__2813);
  xnor g__2935(w__3422 ,w__3394 ,w__3350);
  and g__2936(w__3418 ,w__3326 ,w__3394);
  and g__2937(w__3417 ,w__3311 ,w__3404);
  or g__2938(w__3416 ,w__3402 ,w__3389);
  and g__2939(w__3415 ,w__3402 ,w__3389);
  nor g__2940(w__3414 ,w__3359 ,w__3396);
  or g__2941(w__3413 ,w__3385 ,w__3392);
  not g__2942(w__3410 ,w__3411);
  nor g__2943(w__3409 ,w__3384 ,w__3391);
  or g__2944(w__3408 ,w__3383 ,w__3390);
  nor g__2945(w__3407 ,w__3386 ,w__3393);
  xnor g__2946(w__3406 ,w__3377 ,w__2951);
  xnor g__2947(w__3405 ,w__3357 ,w__3376);
  xnor g__2948(w__3412 ,w__3319 ,w__3372);
  xnor g__2949(w__3411 ,w__3347 ,w__3371);
  not g__2950(w__3400 ,w__3401);
  not g__2951(w__3399 ,w__3398);
  and g__2952(w__3397 ,w__2951 ,w__3377);
  nor g__2953(w__3396 ,w__2950 ,w__3377);
  or g__2954(w__3395 ,w__3357 ,w__3376);
  or g__2955(w__3404 ,w__3310 ,w__3378);
  and g__2956(w__3403 ,w__3367 ,w__3379);
  and g__2957(w__3402 ,w__3366 ,w__3381);
  or g__2958(w__3401 ,w__3362 ,w__3380);
  and g__2959(w__3398 ,w__3361 ,w__3375);
  not g__2960(w__3392 ,w__3393);
  not g__2961(w__3390 ,w__3391);
  xnor g__2962(w__8444 ,w__3369 ,w__3321);
  and g__2963(w__3388 ,w__3357 ,w__3376);
  xnor g__2964(w__3387 ,w__3358 ,w__3368);
  xnor g__2965(w__3394 ,w__3349 ,w__2959);
  xnor g__2966(w__3393 ,w__3334 ,w__2805);
  xnor g__2967(w__3391 ,w__3353 ,w__2955);
  xnor g__2968(w__3389 ,w__3302 ,w__3348);
  not g__2969(w__3386 ,w__3385);
  not g__2970(w__3384 ,w__3383);
  or g__2971(w__3382 ,w__3368 ,w__3358);
  or g__2972(w__3381 ,w__3347 ,w__2812);
  nor g__2973(w__3380 ,w__3319 ,w__3356);
  or g__2974(w__3379 ,w__3305 ,w__3363);
  and g__2975(w__3378 ,w__3309 ,w__3369);
  and g__2976(w__3385 ,w__3346 ,w__3354);
  and g__2977(w__3383 ,w__3336 ,w__3355);
  or g__2978(w__3375 ,w__3370 ,w__3360);
  xnor g__2979(w__8443 ,w__3304 ,w__3323);
  and g__2980(w__3374 ,w__3368 ,w__3358);
  xnor g__2981(w__3373 ,w__3316 ,w__3329);
  xnor g__2982(w__3372 ,w__3328 ,w__2942);
  xnor g__2983(w__3371 ,w__3332 ,w__2969);
  xnor g__2984(w__3377 ,w__3239 ,w__3324);
  xnor g__2985(w__3376 ,w__3292 ,w__2804);
  or g__2986(w__3367 ,w__2988 ,w__3334);
  or g__2987(w__3366 ,w__3001 ,w__3332);
  and g__2988(w__3365 ,w__3316 ,w__3329);
  or g__2989(w__3364 ,w__3316 ,w__3329);
  nor g__2990(w__3363 ,w__2957 ,w__3333);
  and g__2991(w__3362 ,w__2942 ,w__3328);
  or g__2992(w__3361 ,w__3295 ,w__3331);
  nor g__2993(w__3360 ,w__3296 ,w__3330);
  and g__2994(w__3370 ,w__3306 ,w__3337);
  or g__2995(w__3369 ,w__3308 ,w__3339);
  and g__2996(w__3368 ,w__3279 ,w__3340);
  nor g__2997(w__3356 ,w__2941 ,w__3328);
  or g__2998(w__3355 ,w__3302 ,w__3341);
  or g__2999(w__3354 ,w__3272 ,w__3345);
  xnor g__3000(w__3353 ,w__3320 ,w__3237);
  xnor g__3001(w__3352 ,w__3301 ,w__3294);
  xnor g__3002(w__3351 ,w__3285 ,w__3297);
  xnor g__3003(w__3350 ,w__3290 ,w__3318);
  xnor g__3004(w__3349 ,w__3303 ,w__3195);
  xnor g__3005(w__3348 ,w__3299 ,w__2972);
  and g__3006(w__3359 ,w__3254 ,w__3335);
  xnor g__3007(w__3358 ,w__3286 ,w__2962);
  or g__3008(w__3357 ,w__3315 ,w__3344);
  or g__3009(w__3346 ,w__3000 ,w__3292);
  nor g__3010(w__3345 ,w__2953 ,w__3291);
  nor g__3011(w__3344 ,w__3222 ,w__3314);
  and g__3012(w__3343 ,w__3285 ,w__3297);
  or g__3013(w__3342 ,w__3285 ,w__3297);
  nor g__3014(w__3341 ,w__2971 ,w__3299);
  or g__3015(w__3340 ,w__2811 ,w__3320);
  and g__3016(w__3339 ,w__3304 ,w__3288);
  nor g__3017(w__3338 ,w__3290 ,w__3317);
  or g__3018(w__3337 ,w__3223 ,w__3307);
  or g__3019(w__3336 ,w__2998 ,w__3298);
  or g__3020(w__3335 ,w__2810 ,w__3303);
  and g__3021(w__3347 ,w__3275 ,w__3313);
  not g__3022(w__3333 ,w__3334);
  not g__3023(w__3330 ,w__3331);
  nor g__3024(w__3327 ,w__3301 ,w__3294);
  or g__3025(w__3326 ,w__3289 ,w__3318);
  or g__3026(w__3325 ,w__3300 ,w__3293);
  xnor g__3027(w__3324 ,w__3198 ,w__3271);
  xnor g__3028(w__3323 ,w__3112 ,w__2803);
  xnor g__3029(w__3322 ,w__3218 ,w__3269);
  xnor g__3030(w__3321 ,w__3221 ,w__3267);
  xnor g__3031(w__3334 ,w__3242 ,w__3260);
  xnor g__3032(w__3332 ,w__3257 ,w__3263);
  xnor g__3033(w__3331 ,w__3258 ,w__3261);
  xnor g__3034(w__3329 ,w__3266 ,w__3262);
  xnor g__3035(w__3328 ,w__3268 ,w__3259);
  not g__3036(w__3317 ,w__3318);
  nor g__3037(w__3315 ,w__2997 ,w__3266);
  and g__3038(w__3314 ,w__2997 ,w__3266);
  or g__3039(w__3313 ,w__3271 ,w__3273);
  and g__3040(w__3312 ,w__3218 ,w__3269);
  or g__3041(w__3311 ,w__3218 ,w__3269);
  and g__3042(w__3310 ,w__3221 ,w__3267);
  or g__3043(w__3309 ,w__3221 ,w__3267);
  nor g__3044(w__3308 ,w__3112 ,w__2803);
  and g__3045(w__3307 ,w__3200 ,w__3268);
  or g__3046(w__3306 ,w__3200 ,w__3268);
  and g__3047(w__3320 ,w__3244 ,w__3280);
  and g__3048(w__3319 ,w__3246 ,w__3274);
  or g__3049(w__3318 ,w__3250 ,w__3278);
  or g__3050(w__3316 ,w__3217 ,w__3281);
  not g__3051(w__3300 ,w__3301);
  not g__3052(w__3298 ,w__3299);
  not g__3053(w__3295 ,w__3296);
  not g__3054(w__3294 ,w__3293);
  not g__3055(w__3291 ,w__3292);
  not g__3056(w__3289 ,w__3290);
  or g__3057(w__3288 ,w__3111 ,w__3270);
  xnor g__3058(w__8442 ,w__3256 ,w__3189);
  xnor g__3059(w__3287 ,w__3206 ,w__3255);
  xnor g__3060(w__3286 ,w__3241 ,w__3203);
  and g__3061(w__3305 ,w__3235 ,w__3265);
  or g__3062(w__3304 ,w__3163 ,w__3264);
  and g__3063(w__3303 ,w__3231 ,w__3283);
  and g__3064(w__3302 ,w__3252 ,w__3282);
  xnor g__3065(w__3301 ,w__3227 ,w__2964);
  xnor g__3066(w__3299 ,w__3204 ,w__3226);
  xnor g__3067(w__3297 ,w__3240 ,w__3225);
  xnor g__3068(w__3296 ,w__3194 ,w__3228);
  and g__3069(w__3293 ,w__3243 ,w__3284);
  xnor g__3070(w__3292 ,w__3196 ,w__3230);
  xnor g__3071(w__3290 ,w__3171 ,w__3229);
  or g__3072(w__3284 ,w__3241 ,w__3249);
  or g__3073(w__3283 ,w__3185 ,w__3253);
  or g__3074(w__3282 ,w__3257 ,w__3245);
  nor g__3075(w__3281 ,w__3216 ,w__3240);
  or g__3076(w__3280 ,w__3170 ,w__3236);
  or g__3077(w__3279 ,w__2996 ,w__3237);
  nor g__3078(w__3278 ,w__3248 ,w__3258);
  or g__3079(w__3277 ,w__3255 ,w__3206);
  and g__3080(w__3276 ,w__3255 ,w__3206);
  or g__3081(w__3275 ,w__3197 ,w__3239);
  or g__3082(w__3274 ,w__3251 ,w__3242);
  nor g__3083(w__3273 ,w__3198 ,w__3238);
  or g__3084(w__3285 ,w__3166 ,w__3233);
  not g__3085(w__3270 ,w__2803);
  or g__3086(w__3265 ,w__3169 ,w__3234);
  nor g__3087(w__3264 ,w__3177 ,w__3256);
  xor g__3088(w__8441 ,w__3106 ,w__3188);
  xnor g__3089(w__3263 ,w__3201 ,w__3183);
  xnor g__3090(w__3262 ,w__3222 ,w__2933);
  xnor g__3091(w__3261 ,w__3220 ,w__2948);
  xnor g__3092(w__3260 ,w__3199 ,w__3219);
  xor g__3093(w__3259 ,w__3200 ,w__3223);
  and g__3094(w__3272 ,w__3164 ,w__3232);
  and g__3095(w__3271 ,w__3210 ,w__3247);
  xnor g__3096(w__3269 ,w__3224 ,w__2802);
  xnor g__3097(w__3268 ,w__3187 ,w__3191);
  xnor g__3098(w__3267 ,w__3190 ,w__2935);
  xnor g__3099(w__3266 ,w__3207 ,w__3193);
  or g__3100(w__3254 ,w__2984 ,w__3195);
  and g__3101(w__3253 ,w__3089 ,w__3194);
  or g__3102(w__3252 ,w__3183 ,w__3201);
  and g__3103(w__3251 ,w__3219 ,w__3199);
  and g__3104(w__3250 ,w__2948 ,w__3220);
  nor g__3105(w__3249 ,w__2961 ,w__3203);
  nor g__3106(w__3248 ,w__2947 ,w__3220);
  or g__3107(w__3247 ,w__3171 ,w__3214);
  or g__3108(w__3246 ,w__3219 ,w__3199);
  and g__3109(w__3245 ,w__3183 ,w__3201);
  or g__3110(w__3244 ,w__3021 ,w__3205);
  or g__3111(w__3243 ,w__2985 ,w__3202);
  and g__3112(w__3258 ,w__3175 ,w__3213);
  and g__3113(w__3257 ,w__3078 ,w__3215);
  and g__3114(w__3256 ,w__3179 ,w__3211);
  and g__3115(w__3255 ,w__3103 ,w__3212);
  not g__3116(w__3238 ,w__3239);
  and g__3117(w__3236 ,w__3021 ,w__3205);
  or g__3118(w__3235 ,w__3105 ,w__3196);
  and g__3119(w__3234 ,w__3105 ,w__3196);
  and g__3120(w__3233 ,w__3161 ,w__3224);
  or g__3121(w__3232 ,w__3167 ,w__3207);
  or g__3122(w__3231 ,w__3089 ,w__3194);
  xnor g__3123(w__3230 ,w__3105 ,w__3169);
  xnor g__3124(w__3229 ,w__3042 ,w__3168);
  xor g__3125(w__3228 ,w__3089 ,w__3185);
  xnor g__3126(w__3227 ,w__3186 ,w__3043);
  xnor g__3127(w__3226 ,w__3021 ,w__3170);
  xnor g__3128(w__3225 ,w__3182 ,w__2931);
  xnor g__3129(w__3242 ,w__3133 ,w__3159);
  and g__3130(w__3241 ,w__3069 ,w__3209);
  xnor g__3131(w__3240 ,w__2806 ,w__3158);
  xnor g__3132(w__3239 ,w__3184 ,w__3116);
  xnor g__3133(w__3237 ,w__3172 ,w__3120);
  nor g__3134(w__3217 ,w__3002 ,w__3182);
  and g__3135(w__3216 ,w__3002 ,w__3182);
  or g__3136(w__3215 ,w__3073 ,w__3184);
  and g__3137(w__3214 ,w__3042 ,w__3168);
  or g__3138(w__3213 ,w__3187 ,w__3181);
  or g__3139(w__3212 ,w__2807 ,w__3186);
  or g__3140(w__3211 ,w__3106 ,w__3176);
  or g__3141(w__3210 ,w__3042 ,w__3168);
  or g__3142(w__3209 ,w__3099 ,w__3172);
  xnor g__3143(w__3208 ,w__3018 ,w__3132);
  xnor g__3144(w__3224 ,w__3090 ,w__3115);
  and g__3145(w__3223 ,w__3141 ,w__3160);
  and g__3146(w__3222 ,w__3148 ,w__3173);
  or g__3147(w__3221 ,w__3094 ,w__3174);
  xnor g__3148(w__3220 ,w__3008 ,w__3136);
  and g__3149(w__3219 ,w__3083 ,w__3162);
  or g__3150(w__3218 ,w__3152 ,w__3178);
  not g__3151(w__3205 ,w__3204);
  not g__3152(w__3202 ,w__3203);
  not g__3153(w__3197 ,w__3198);
  xnor g__3154(w__3193 ,w__3088 ,w__3131);
  xnor g__3155(w__3192 ,w__3155 ,w__2967);
  xnor g__3156(w__3191 ,w__3110 ,w__3126);
  xnor g__3157(w__3190 ,w__2808 ,w__3108);
  xnor g__3158(w__3189 ,w__3109 ,w__3156);
  xnor g__3159(w__3188 ,w__3128 ,w__2975);
  xnor g__3160(w__3207 ,w__3020 ,w__3117);
  xnor g__3161(w__3206 ,w__3135 ,w__2945);
  xnor g__3162(w__3204 ,w__3044 ,w__3122);
  xnor g__3163(w__3203 ,w__3038 ,w__3119);
  xnor g__3164(w__3201 ,w__3011 ,w__3113);
  xnor g__3165(w__3200 ,w__3013 ,w__3114);
  xnor g__3166(w__3199 ,w__3048 ,w__3125);
  xnor g__3167(w__3198 ,w__3006 ,w__3123);
  xnor g__3168(w__3196 ,w__2809 ,w__3118);
  xnor g__3169(w__3195 ,w__3039 ,w__3121);
  xnor g__3170(w__3194 ,w__3058 ,w__3124);
  and g__3171(w__3181 ,w__3110 ,w__3126);
  or g__3172(w__3180 ,w__2989 ,w__3154);
  or g__3173(w__3179 ,w__2987 ,w__3127);
  nor g__3174(w__3178 ,w__3142 ,w__2808);
  and g__3175(w__3177 ,w__3109 ,w__3157);
  nor g__3176(w__3176 ,w__2974 ,w__3128);
  or g__3177(w__3175 ,w__3110 ,w__3126);
  and g__3178(w__3174 ,w__3101 ,w__3132);
  or g__3179(w__3173 ,w__3150 ,w__2806);
  and g__3180(w__3187 ,w__3082 ,w__3144);
  and g__3181(w__3186 ,w__3098 ,w__3137);
  and g__3182(w__3185 ,w__3070 ,w__3151);
  and g__3183(w__3184 ,w__3100 ,w__3143);
  and g__3184(w__3183 ,w__3104 ,w__3149);
  and g__3185(w__3182 ,w__3076 ,w__3147);
  nor g__3186(w__3167 ,w__3088 ,w__3131);
  and g__3187(w__3166 ,w__2937 ,w__3129);
  nor g__3188(w__3165 ,w__2966 ,w__3155);
  or g__3189(w__3164 ,w__3087 ,w__3130);
  nor g__3190(w__3163 ,w__3109 ,w__3157);
  or g__3191(w__3162 ,w__3072 ,w__2809);
  or g__3192(w__3161 ,w__2937 ,w__3129);
  or g__3193(w__3160 ,w__3134 ,w__3153);
  xnor g__3194(w__3159 ,w__3051 ,w__3086);
  xnor g__3195(w__3158 ,w__3015 ,w__3107);
  and g__3196(w__3172 ,w__3093 ,w__3146);
  and g__3197(w__3171 ,w__3071 ,w__3139);
  and g__3198(w__3170 ,w__3080 ,w__3145);
  and g__3199(w__3169 ,w__3084 ,w__3138);
  and g__3200(w__3168 ,w__3096 ,w__3140);
  not g__3201(w__3157 ,w__3156);
  not g__3202(w__3155 ,w__3154);
  nor g__3203(w__3153 ,w__3050 ,w__3086);
  nor g__3204(w__3152 ,w__2986 ,w__3108);
  or g__3205(w__3151 ,w__3029 ,w__3077);
  and g__3206(w__3150 ,w__3015 ,w__3107);
  or g__3207(w__3149 ,w__3028 ,w__3092);
  or g__3208(w__3148 ,w__3015 ,w__3107);
  or g__3209(w__3146 ,w__3055 ,w__3091);
  or g__3210(w__3145 ,w__3056 ,w__3074);
  or g__3211(w__3144 ,w__3031 ,w__3081);
  or g__3212(w__3143 ,w__3024 ,w__3079);
  and g__3213(w__3142 ,w__2986 ,w__3108);
  or g__3214(w__3141 ,w__3051 ,w__3085);
  or g__3215(w__3140 ,w__3033 ,w__3097);
  or g__3216(w__3139 ,w__3058 ,w__3068);
  or g__3217(w__3138 ,w__3026 ,w__3075);
  or g__3218(w__3137 ,w__3057 ,w__3095);
  xnor g__3219(w__3136 ,w__3033 ,in5[6]);
  xnor g__3220(w__3135 ,w__3034 ,in5[10]);
  xnor g__3221(w__3156 ,w__3062 ,w__2929);
  and g__3222(w__3154 ,w__3004 ,w__3102);
  not g__3223(w__3134 ,w__3133);
  not g__3224(w__3130 ,w__3131);
  not g__3225(w__3127 ,w__3128);
  xnor g__3226(w__3125 ,w__3007 ,w__3031);
  xnor g__3227(w__3124 ,w__3012 ,w__3046);
  xnor g__3228(w__3123 ,w__3028 ,in5[7]);
  xnor g__3229(w__3122 ,w__3055 ,in5[8]);
  xnor g__3230(w__3121 ,w__3009 ,w__3024);
  xnor g__3231(w__3120 ,w__3041 ,w__3010);
  xnor g__3232(w__3119 ,w__3057 ,in5[9]);
  xnor g__3233(w__3118 ,w__3037 ,w__3049);
  xnor g__3234(w__3117 ,w__3040 ,w__3026);
  xnor g__3235(w__3116 ,w__3019 ,w__3016);
  xnor g__3236(w__3115 ,w__3014 ,w__3047);
  xnor g__3237(w__3114 ,w__3045 ,w__3029);
  xnor g__3238(w__3113 ,w__3005 ,w__3056);
  xnor g__3239(w__3133 ,w__3064 ,in5[5]);
  xnor g__3240(w__3132 ,w__3027 ,in5[2]);
  xnor g__3241(w__3131 ,w__3032 ,in5[4]);
  xnor g__3242(w__3129 ,w__3061 ,in5[3]);
  xnor g__3243(w__3128 ,w__3053 ,in5[1]);
  xnor g__3244(w__3126 ,w__3065 ,w__3022);
  not g__3245(w__3112 ,w__3111);
  or g__3246(w__3104 ,w__2826 ,w__3006);
  or g__3247(w__3103 ,w__3003 ,w__3043);
  or g__3248(w__3102 ,w__3034 ,w__3035);
  or g__3249(w__3101 ,w__2939 ,w__3017);
  or g__3250(w__3100 ,w__3009 ,w__3039);
  and g__3251(w__3099 ,w__3041 ,w__3010);
  or g__3252(w__3098 ,w__2816 ,w__3038);
  and g__3253(w__3097 ,w__2836 ,w__3008);
  or g__3254(w__3096 ,w__2840 ,w__3008);
  and g__3255(w__3095 ,w__2820 ,w__3038);
  nor g__3256(w__3094 ,w__2990 ,w__3018);
  or g__3257(w__3093 ,w__2865 ,w__3044);
  and g__3258(w__3092 ,w__2830 ,w__3006);
  and g__3259(w__3091 ,w__2852 ,w__3044);
  and g__3260(w__3111 ,w__2929 ,w__3063);
  or g__3261(w__3110 ,w__2873 ,w__3064);
  or g__3262(w__3109 ,w__2883 ,w__3053);
  or g__3263(w__3108 ,w__2892 ,w__3027);
  or g__3264(w__3107 ,w__2886 ,w__3061);
  or g__3265(w__3106 ,w__2976 ,w__3025);
  or g__3266(w__3105 ,w__2889 ,w__3032);
  not g__3267(w__3087 ,w__3088);
  not g__3268(w__3085 ,w__3086);
  and g__3269(w__8439 ,w__3025 ,w__3036);
  or g__3270(w__3084 ,w__3020 ,w__3040);
  or g__3271(w__3083 ,w__3037 ,w__3049);
  or g__3272(w__3082 ,w__3048 ,w__3007);
  and g__3273(w__3081 ,w__3048 ,w__3007);
  or g__3274(w__3080 ,w__3005 ,w__3011);
  and g__3275(w__3079 ,w__3009 ,w__3039);
  or g__3276(w__3078 ,w__3019 ,w__3016);
  and g__3277(w__3077 ,w__3013 ,w__3045);
  or g__3278(w__3076 ,w__3014 ,w__3047);
  and g__3279(w__3075 ,w__3020 ,w__3040);
  and g__3280(w__3074 ,w__3005 ,w__3011);
  and g__3281(w__3073 ,w__3019 ,w__3016);
  and g__3282(w__3072 ,w__3037 ,w__3049);
  or g__3283(w__3071 ,w__3012 ,w__3046);
  or g__3284(w__3070 ,w__3013 ,w__3045);
  or g__3285(w__3069 ,w__3041 ,w__3010);
  and g__3286(w__3068 ,w__3012 ,w__3046);
  and g__3287(w__3090 ,w__3052 ,w__3023);
  or g__3288(w__3089 ,w__3065 ,w__3022);
  and g__3289(w__3088 ,w__3030 ,w__3060);
  and g__3290(w__3086 ,w__3054 ,w__3067);
  not g__3291(w__3067 ,w__3066);
  not g__3292(w__3063 ,w__3062);
  not g__3293(w__3060 ,w__3059);
  not g__3294(w__3051 ,w__3050);
  or g__3295(w__3036 ,in5[0] ,w__2925);
  nor g__3296(w__3035 ,in5[10] ,w__2944);
  or g__3297(w__3066 ,w__2849 ,w__2868);
  or g__3298(w__3065 ,w__2838 ,w__2857);
  or g__3299(w__3064 ,w__2818 ,w__2870);
  or g__3300(w__3062 ,w__2854 ,w__2900);
  or g__3301(w__3061 ,w__2875 ,w__2903);
  or g__3302(w__3059 ,w__2833 ,w__2870);
  or g__3303(w__3058 ,w__2878 ,w__2915);
  or g__3304(w__3057 ,w__2863 ,w__2828);
  or g__3305(w__3056 ,w__2846 ,w__2913);
  or g__3306(w__3055 ,w__2843 ,w__2895);
  and g__3307(w__3054 ,in5[5] ,in5[3]);
  or g__3308(w__3053 ,w__2880 ,w__2868);
  and g__3309(w__3052 ,in5[3] ,in5[1]);
  and g__3310(w__3050 ,in5[8] ,in5[1]);
  or g__3311(w__3049 ,w__2823 ,w__2881);
  or g__3312(w__3048 ,w__2898 ,w__2890);
  or g__3313(w__3047 ,w__2858 ,w__2884);
  or g__3314(w__3046 ,w__2905 ,w__2860);
  or g__3315(w__3045 ,w__2851 ,w__2893);
  or g__3316(w__3044 ,w__2923 ,w__2917);
  or g__3317(w__3043 ,w__2908 ,w__2849);
  or g__3318(w__3042 ,w__2848 ,w__2889);
  or g__3319(w__3041 ,w__2878 ,w__2920);
  or g__3320(w__3040 ,w__2875 ,w__2855);
  or g__3321(w__3039 ,w__2924 ,w__2911);
  or g__3322(w__3038 ,w__2877 ,w__2905);
  or g__3323(w__3037 ,w__2833 ,w__2892);
  not g__3324(w__3018 ,w__3017);
  or g__3325(w__3004 ,w__2845 ,w__2999);
  or g__3326(w__3034 ,w__2843 ,w__2820);
  or g__3327(w__3033 ,w__2842 ,w__2880);
  or g__3328(w__3032 ,w__2823 ,w__2900);
  or g__3329(w__3031 ,w__2921 ,w__2915);
  and g__3330(w__3030 ,in5[4] ,in5[2]);
  or g__3331(w__3029 ,w__2816 ,w__2883);
  or g__3332(w__3028 ,w__2908 ,w__2887);
  or g__3333(w__3027 ,w__2861 ,w__2903);
  or g__3334(w__3026 ,w__2918 ,w__2881);
  or g__3335(w__3025 ,w__2901 ,w__2977);
  or g__3336(w__3024 ,w__2846 ,w__2893);
  and g__3337(w__3023 ,in5[4] ,in5[0]);
  or g__3338(w__3022 ,w__2909 ,w__2867);
  or g__3339(w__3021 ,w__2852 ,w__2822);
  or g__3340(w__3020 ,w__2913 ,w__2886);
  or g__3341(w__3019 ,w__2830 ,w__2832);
  and g__3342(w__3017 ,in5[2] ,in5[1]);
  or g__3343(w__3016 ,w__2818 ,w__2890);
  or g__3344(w__3015 ,w__2873 ,w__2884);
  or g__3345(w__3014 ,w__2911 ,w__2855);
  or g__3346(w__3013 ,w__2826 ,w__2887);
  or g__3347(w__3012 ,w__2840 ,w__2895);
  or g__3348(w__3011 ,w__2815 ,w__2898);
  or g__3349(w__3010 ,w__2863 ,w__2836);
  or g__3350(w__3009 ,w__2828 ,w__2896);
  or g__3351(w__3008 ,w__2825 ,w__2858);
  or g__3352(w__3007 ,w__2838 ,w__2861);
  or g__3353(w__3006 ,w__2906 ,w__2872);
  or g__3354(w__3005 ,w__2865 ,w__2835);
  not g__3355(w__3003 ,w__2964);
  not g__3356(w__3002 ,w__2931);
  not g__3357(w__3001 ,w__2969);
  not g__3358(w__3000 ,w__2953);
  not g__3359(w__2999 ,w__2945);
  not g__3360(w__2998 ,w__2972);
  not g__3361(w__2997 ,w__2933);
  not g__3362(w__2996 ,w__2955);
  not g__3363(w__2995 ,in5[0]);
  not g__3364(w__2994 ,in5[4]);
  not g__3365(w__2993 ,in5[1]);
  not g__3366(w__2992 ,in5[8]);
  not g__3367(w__2991 ,in5[9]);
  not g__3368(w__2990 ,w__2939);
  not g__3369(w__2989 ,w__2967);
  not g__3370(w__2988 ,w__2957);
  not g__3371(w__2987 ,w__2975);
  not g__3372(w__2986 ,w__2935);
  not g__3373(w__2985 ,w__2962);
  not g__3374(w__2984 ,w__2959);
  not g__3375(w__2983 ,in5[3]);
  not g__3376(w__2982 ,in5[5]);
  not g__3377(w__2981 ,in5[2]);
  not g__3378(w__2980 ,in5[7]);
  not g__3379(w__2979 ,in5[6]);
  not g__3380(w__2978 ,in5[10]);
  not g__3381(w__2975 ,w__2973);
  not g__3382(w__2974 ,w__2973);
  not g__3383(w__2973 ,w__8465);
  not g__3384(w__2972 ,w__2970);
  not g__3385(w__2971 ,w__2970);
  not g__3386(w__2970 ,w__8479);
  not g__3387(w__2969 ,w__2968);
  not g__3388(w__2968 ,w__8478);
  not g__3389(w__2967 ,w__2965);
  not g__3390(w__2966 ,w__2965);
  not g__3391(w__2965 ,w__8484);
  not g__3392(w__2964 ,w__2963);
  not g__3393(w__2963 ,w__8482);
  not g__3394(w__2962 ,w__2960);
  not g__3395(w__2961 ,w__2960);
  not g__3396(w__2960 ,w__8481);
  not g__3397(w__2959 ,w__2958);
  not g__3398(w__2958 ,w__8476);
  not g__3399(w__2957 ,w__2956);
  not g__3400(w__2956 ,w__8473);
  not g__3401(w__2955 ,w__2954);
  not g__3402(w__2954 ,w__8480);
  not g__3403(w__2953 ,w__2952);
  not g__3404(w__2952 ,w__8472);
  not g__3405(w__2951 ,w__2949);
  not g__3406(w__2950 ,w__2949);
  not g__3407(w__2949 ,w__8477);
  not g__3408(w__2948 ,w__2946);
  not g__3409(w__2947 ,w__2946);
  not g__3410(w__2946 ,w__8475);
  not g__3411(w__2945 ,w__2943);
  not g__3412(w__2944 ,w__2943);
  not g__3413(w__2943 ,w__8483);
  not g__3414(w__2942 ,w__2940);
  not g__3415(w__2941 ,w__2940);
  not g__3416(w__2940 ,w__8474);
  not g__3417(w__2939 ,w__2938);
  not g__3418(w__2938 ,w__8467);
  not g__3419(w__2937 ,w__2936);
  not g__3420(w__2936 ,w__8469);
  not g__3421(w__2935 ,w__2934);
  not g__3422(w__2934 ,w__8468);
  not g__3423(w__2933 ,w__2932);
  not g__3424(w__2932 ,w__8471);
  not g__3425(w__2931 ,w__2930);
  not g__3426(w__2930 ,w__8470);
  not g__3427(w__2976 ,w__8464);
  not g__3428(w__2929 ,w__2928);
  not g__3429(w__2928 ,w__8466);
  not g__3430(w__2927 ,w__2926);
  not g__3431(w__2926 ,w__8485);
  not g__3432(w__2925 ,w__2977);
  not g__3433(w__2977 ,w__8463);
  not g__3434(w__2924 ,w__2922);
  not g__3435(w__2923 ,w__2922);
  not g__3436(w__2922 ,w__2991);
  not g__3437(w__2921 ,w__2919);
  not g__3438(w__2920 ,w__2919);
  not g__3439(w__2919 ,w__2980);
  not g__3440(w__2918 ,w__2916);
  not g__3441(w__2917 ,w__2916);
  not g__3442(w__2916 ,w__2979);
  not g__3443(w__2915 ,w__2914);
  not g__3444(w__2914 ,w__2981);
  not g__3445(w__2913 ,w__2912);
  not g__3446(w__2912 ,w__2994);
  not g__3447(w__2911 ,w__2910);
  not g__3448(w__2910 ,w__2983);
  not g__3449(w__2909 ,w__2907);
  not g__3450(w__2908 ,w__2907);
  not g__3451(w__2907 ,w__2978);
  not g__3452(w__2906 ,w__2904);
  not g__3453(w__2905 ,w__2904);
  not g__3454(w__2904 ,w__2992);
  not g__3455(w__2903 ,w__2902);
  not g__3456(w__2902 ,w__2995);
  not g__3457(w__2901 ,w__2899);
  not g__3458(w__2900 ,w__2899);
  not g__3459(w__2899 ,w__2995);
  not g__3460(w__2898 ,w__2897);
  not g__3461(w__2897 ,w__2982);
  not g__3462(w__2896 ,w__2894);
  not g__3463(w__2895 ,w__2894);
  not g__3464(w__2894 ,w__2982);
  not g__3465(w__2893 ,w__2891);
  not g__3466(w__2892 ,w__2891);
  not g__3467(w__2891 ,w__2981);
  not g__3468(w__2890 ,w__2888);
  not g__3469(w__2889 ,w__2888);
  not g__3470(w__2888 ,w__2994);
  not g__3471(w__2887 ,w__2885);
  not g__3472(w__2886 ,w__2885);
  not g__3473(w__2885 ,w__2983);
  not g__3474(w__2884 ,w__2882);
  not g__3475(w__2883 ,w__2882);
  not g__3476(w__2882 ,w__2993);
  not g__3477(w__2881 ,w__2879);
  not g__3478(w__2880 ,w__2879);
  not g__3479(w__2879 ,w__2993);
  not g__3480(w__2878 ,w__2876);
  not g__3481(w__2877 ,w__2876);
  not g__3482(w__2876 ,w__2991);
  not g__3483(w__2875 ,w__2874);
  not g__3484(w__2874 ,w__2896);
  not g__3485(w__2873 ,w__2871);
  not g__3486(w__2872 ,w__2871);
  not g__3487(w__2871 ,w__2982);
  not g__3488(w__2870 ,w__2869);
  not g__3489(w__2869 ,w__2901);
  not g__3490(w__2868 ,w__2866);
  not g__3491(w__2867 ,w__2866);
  not g__3492(w__2866 ,w__2995);
  not g__3493(w__2865 ,w__2864);
  not g__3494(w__2864 ,w__2906);
  not g__3495(w__2863 ,w__2862);
  not g__3496(w__2862 ,w__2909);
  not g__3497(w__2861 ,w__2859);
  not g__3498(w__2860 ,w__2859);
  not g__3499(w__2859 ,w__2983);
  not g__3500(w__2858 ,w__2856);
  not g__3501(w__2857 ,w__2856);
  not g__3502(w__2856 ,w__2994);
  not g__3503(w__2855 ,w__2853);
  not g__3504(w__2854 ,w__2853);
  not g__3505(w__2853 ,w__2981);
  not g__3506(w__2852 ,w__2850);
  not g__3507(w__2851 ,w__2850);
  not g__3508(w__2850 ,w__2992);
  not g__3509(w__2849 ,w__2847);
  not g__3510(w__2848 ,w__2847);
  not g__3511(w__2847 ,w__2992);
  not g__3512(w__2846 ,w__2844);
  not g__3513(w__2845 ,w__2844);
  not g__3514(w__2844 ,w__2978);
  not g__3515(w__2843 ,w__2841);
  not g__3516(w__2842 ,w__2841);
  not g__3517(w__2841 ,w__2978);
  not g__3518(w__2840 ,w__2839);
  not g__3519(w__2839 ,w__2917);
  not g__3520(w__2838 ,w__2837);
  not g__3521(w__2837 ,w__2918);
  not g__3522(w__2836 ,w__2834);
  not g__3523(w__2835 ,w__2834);
  not g__3524(w__2834 ,w__2979);
  not g__3525(w__2833 ,w__2831);
  not g__3526(w__2832 ,w__2831);
  not g__3527(w__2831 ,w__2979);
  not g__3528(w__2830 ,w__2829);
  not g__3529(w__2829 ,w__2920);
  not g__3530(w__2828 ,w__2827);
  not g__3531(w__2827 ,w__2921);
  not g__3532(w__2826 ,w__2824);
  not g__3533(w__2825 ,w__2824);
  not g__3534(w__2824 ,w__2980);
  not g__3535(w__2823 ,w__2821);
  not g__3536(w__2822 ,w__2821);
  not g__3537(w__2821 ,w__2980);
  not g__3538(w__2820 ,w__2819);
  not g__3539(w__2819 ,w__2923);
  not g__3540(w__2818 ,w__2817);
  not g__3541(w__2817 ,w__2924);
  not g__3542(w__2816 ,w__2814);
  not g__3543(w__2815 ,w__2814);
  not g__3544(w__2814 ,w__2991);
  xor g__3545(w__8460 ,w__3476 ,w__3192);
  xor g__3546(w__8459 ,w__3474 ,w__3287);
  xor g__3547(w__8458 ,w__3472 ,w__3352);
  xor g__3548(w__8457 ,w__3470 ,w__3387);
  xor g__3549(w__8456 ,w__3468 ,w__3419);
  xor g__3550(w__8455 ,w__3466 ,w__3421);
  xor g__3551(w__8454 ,w__3464 ,w__3445);
  xor g__3552(w__8453 ,w__3462 ,w__3449);
  xor g__3553(w__8452 ,w__3460 ,w__3444);
  xor g__3554(w__8451 ,w__3458 ,w__3443);
  xor g__3555(w__8450 ,w__3456 ,w__3433);
  xor g__3556(w__2813 ,w__3296 ,w__3370);
  and g__3557(w__2812 ,w__2968 ,w__3332);
  and g__3558(w__2811 ,w__2954 ,w__3237);
  and g__3559(w__2810 ,w__2958 ,w__3195);
  xor g__3560(w__2809 ,w__3054 ,w__3066);
  xnor g__3561(w__2808 ,w__3052 ,w__3023);
  and g__3562(w__2807 ,w__2963 ,w__3043);
  xor g__3563(w__2806 ,w__3030 ,w__3059);
  xor g__3564(w__2805 ,w__3305 ,w__2956);
  xor g__3565(w__2804 ,w__3272 ,w__2952);
  xor g__3566(w__2803 ,w__3208 ,w__2938);
  xor g__3567(w__2802 ,w__3129 ,w__2936);
  xor g__3568(w__8440 ,w__3025 ,w__2976);
  xnor g__3569(w__8437 ,w__4153 ,w__3605);
  and g__3570(w__8438 ,w__3605 ,w__4154);
  not g__3571(w__4154 ,w__4153);
  and g__3572(w__4153 ,w__3856 ,w__4152);
  or g__3573(w__4152 ,w__3842 ,w__4151);
  and g__3574(w__4151 ,w__3952 ,w__4150);
  or g__3575(w__4150 ,w__3951 ,w__4149);
  and g__3576(w__4149 ,w__4000 ,w__4148);
  or g__3577(w__4148 ,w__4002 ,w__4147);
  and g__3578(w__4147 ,w__4057 ,w__4146);
  or g__3579(w__4146 ,w__4049 ,w__4145);
  and g__3580(w__4145 ,w__4083 ,w__4144);
  or g__3581(w__4144 ,w__4084 ,w__4143);
  and g__3582(w__4143 ,w__4091 ,w__4142);
  or g__3583(w__4142 ,w__4090 ,w__4141);
  and g__3584(w__4141 ,w__4115 ,w__4140);
  or g__3585(w__4140 ,w__4116 ,w__4139);
  and g__3586(w__4139 ,w__4122 ,w__4138);
  or g__3587(w__4138 ,w__4121 ,w__4137);
  and g__3588(w__4137 ,w__4114 ,w__4136);
  or g__3589(w__4136 ,w__4113 ,w__4135);
  and g__3590(w__4135 ,w__4112 ,w__4134);
  or g__3591(w__4134 ,w__4111 ,w__4133);
  and g__3592(w__4133 ,w__4102 ,w__4132);
  or g__3593(w__4132 ,w__4101 ,w__4131);
  and g__3594(w__4131 ,w__4088 ,w__4130);
  xnor g__3595(w__8425 ,w__4128 ,w__4095);
  or g__3596(w__4130 ,w__4082 ,w__4129);
  not g__3597(w__4129 ,w__4128);
  or g__3598(w__4128 ,w__4063 ,w__4127);
  xnor g__3599(w__8424 ,w__4126 ,w__4080);
  and g__3600(w__4127 ,w__4070 ,w__4126);
  or g__3601(w__4126 ,w__4040 ,w__4125);
  xnor g__3602(w__8423 ,w__4123 ,w__4048);
  and g__3603(w__4125 ,w__4039 ,w__4123);
  xnor g__3604(w__4124 ,w__4104 ,w__4110);
  or g__3605(w__4123 ,w__4018 ,w__4117);
  or g__3606(w__4122 ,w__4103 ,w__4109);
  nor g__3607(w__4121 ,w__4104 ,w__4110);
  xnor g__3608(w__4120 ,w__4106 ,w__4086);
  xnor g__3609(w__4119 ,w__4074 ,w__4098);
  xnor g__3610(w__4118 ,w__4076 ,w__4100);
  xnor g__3611(w__8422 ,w__4107 ,w__4026);
  and g__3612(w__4117 ,w__4017 ,w__4107);
  nor g__3613(w__4116 ,w__4106 ,w__4086);
  or g__3614(w__4115 ,w__4105 ,w__4085);
  or g__3615(w__4114 ,w__4073 ,w__4097);
  nor g__3616(w__4113 ,w__4074 ,w__4098);
  or g__3617(w__4112 ,w__4075 ,w__4099);
  nor g__3618(w__4111 ,w__4076 ,w__4100);
  not g__3619(w__4110 ,w__4109);
  xnor g__3620(w__4109 ,w__4034 ,w__4081);
  xnor g__3621(w__4108 ,w__4087 ,w__4078);
  not g__3622(w__4105 ,w__4106);
  not g__3623(w__4103 ,w__4104);
  or g__3624(w__4102 ,w__4078 ,w__4087);
  and g__3625(w__4101 ,w__4078 ,w__4087);
  or g__3626(w__4107 ,w__3987 ,w__4092);
  or g__3627(w__4106 ,w__4072 ,w__4089);
  or g__3628(w__4104 ,w__4013 ,w__4093);
  not g__3629(w__4100 ,w__4099);
  not g__3630(w__4098 ,w__4097);
  xnor g__3631(w__8421 ,w__4079 ,w__3997);
  xnor g__3632(w__4096 ,w__4064 ,w__4077);
  xnor g__3633(w__4095 ,w__4061 ,w__4068);
  xnor g__3634(w__4094 ,w__4059 ,w__4066);
  xnor g__3635(w__4099 ,w__4006 ,w__3491);
  xnor g__3636(w__4097 ,w__4069 ,w__4025);
  and g__3637(w__4093 ,w__4001 ,w__4069);
  and g__3638(w__4092 ,w__3986 ,w__4079);
  or g__3639(w__4091 ,w__4077 ,w__4064);
  and g__3640(w__4090 ,w__4077 ,w__4064);
  nor g__3641(w__4089 ,w__4034 ,w__4071);
  or g__3642(w__4088 ,w__4060 ,w__4067);
  not g__3643(w__4085 ,w__4086);
  nor g__3644(w__4084 ,w__4059 ,w__4066);
  or g__3645(w__4083 ,w__4058 ,w__4065);
  nor g__3646(w__4082 ,w__4061 ,w__4068);
  xnor g__3647(w__4081 ,w__4052 ,w__3629);
  xnor g__3648(w__4080 ,w__4032 ,w__4051);
  xnor g__3649(w__4087 ,w__3994 ,w__4047);
  xnor g__3650(w__4086 ,w__4022 ,w__4046);
  not g__3651(w__4075 ,w__4076);
  not g__3652(w__4074 ,w__4073);
  and g__3653(w__4072 ,w__3629 ,w__4052);
  nor g__3654(w__4071 ,w__3628 ,w__4052);
  or g__3655(w__4070 ,w__4032 ,w__4051);
  or g__3656(w__4079 ,w__3985 ,w__4053);
  and g__3657(w__4078 ,w__4042 ,w__4054);
  and g__3658(w__4077 ,w__4041 ,w__4056);
  or g__3659(w__4076 ,w__4037 ,w__4055);
  and g__3660(w__4073 ,w__4036 ,w__4050);
  not g__3661(w__4067 ,w__4068);
  not g__3662(w__4065 ,w__4066);
  xnor g__3663(w__8420 ,w__4044 ,w__3996);
  and g__3664(w__4063 ,w__4032 ,w__4051);
  xnor g__3665(w__4062 ,w__4033 ,w__4043);
  xnor g__3666(w__4069 ,w__4024 ,w__3637);
  xnor g__3667(w__4068 ,w__4009 ,w__3483);
  xnor g__3668(w__4066 ,w__4028 ,w__3633);
  xnor g__3669(w__4064 ,w__3977 ,w__4023);
  not g__3670(w__4061 ,w__4060);
  not g__3671(w__4059 ,w__4058);
  or g__3672(w__4057 ,w__4043 ,w__4033);
  or g__3673(w__4056 ,w__4022 ,w__3490);
  nor g__3674(w__4055 ,w__3994 ,w__4031);
  or g__3675(w__4054 ,w__3980 ,w__4038);
  and g__3676(w__4053 ,w__3984 ,w__4044);
  and g__3677(w__4060 ,w__4021 ,w__4029);
  and g__3678(w__4058 ,w__4011 ,w__4030);
  or g__3679(w__4050 ,w__4045 ,w__4035);
  xnor g__3680(w__8419 ,w__3979 ,w__3998);
  and g__3681(w__4049 ,w__4043 ,w__4033);
  xnor g__3682(w__4048 ,w__3991 ,w__4004);
  xnor g__3683(w__4047 ,w__4003 ,w__3620);
  xnor g__3684(w__4046 ,w__4007 ,w__3647);
  xnor g__3685(w__4052 ,w__3914 ,w__3999);
  xnor g__3686(w__4051 ,w__3967 ,w__3482);
  or g__3687(w__4042 ,w__3665 ,w__4009);
  or g__3688(w__4041 ,w__3678 ,w__4007);
  and g__3689(w__4040 ,w__3991 ,w__4004);
  or g__3690(w__4039 ,w__3991 ,w__4004);
  nor g__3691(w__4038 ,w__3635 ,w__4008);
  and g__3692(w__4037 ,w__3620 ,w__4003);
  or g__3693(w__4036 ,w__3970 ,w__4006);
  nor g__3694(w__4035 ,w__3971 ,w__4005);
  and g__3695(w__4045 ,w__3981 ,w__4012);
  or g__3696(w__4044 ,w__3983 ,w__4014);
  and g__3697(w__4043 ,w__3954 ,w__4015);
  nor g__3698(w__4031 ,w__3619 ,w__4003);
  or g__3699(w__4030 ,w__3977 ,w__4016);
  or g__3700(w__4029 ,w__3947 ,w__4020);
  xnor g__3701(w__4028 ,w__3995 ,w__3912);
  xnor g__3702(w__4027 ,w__3976 ,w__3969);
  xnor g__3703(w__4026 ,w__3960 ,w__3972);
  xnor g__3704(w__4025 ,w__3965 ,w__3993);
  xnor g__3705(w__4024 ,w__3978 ,w__3871);
  xnor g__3706(w__4023 ,w__3974 ,w__3650);
  and g__3707(w__4034 ,w__3929 ,w__4010);
  xnor g__3708(w__4033 ,w__3961 ,w__3640);
  or g__3709(w__4032 ,w__3990 ,w__4019);
  or g__3710(w__4021 ,w__3677 ,w__3967);
  nor g__3711(w__4020 ,w__3631 ,w__3966);
  nor g__3712(w__4019 ,w__3897 ,w__3989);
  and g__3713(w__4018 ,w__3960 ,w__3972);
  or g__3714(w__4017 ,w__3960 ,w__3972);
  nor g__3715(w__4016 ,w__3649 ,w__3974);
  or g__3716(w__4015 ,w__3489 ,w__3995);
  and g__3717(w__4014 ,w__3979 ,w__3963);
  nor g__3718(w__4013 ,w__3965 ,w__3992);
  or g__3719(w__4012 ,w__3898 ,w__3982);
  or g__3720(w__4011 ,w__3675 ,w__3973);
  or g__3721(w__4010 ,w__3488 ,w__3978);
  and g__3722(w__4022 ,w__3950 ,w__3988);
  not g__3723(w__4008 ,w__4009);
  not g__3724(w__4005 ,w__4006);
  nor g__3725(w__4002 ,w__3976 ,w__3969);
  or g__3726(w__4001 ,w__3964 ,w__3993);
  or g__3727(w__4000 ,w__3975 ,w__3968);
  xnor g__3728(w__3999 ,w__3874 ,w__3946);
  xnor g__3729(w__3998 ,w__3789 ,w__3481);
  xnor g__3730(w__3997 ,w__3893 ,w__3944);
  xnor g__3731(w__3996 ,w__3896 ,w__3942);
  xnor g__3732(w__4009 ,w__3917 ,w__3935);
  xnor g__3733(w__4007 ,w__3932 ,w__3938);
  xnor g__3734(w__4006 ,w__3933 ,w__3936);
  xnor g__3735(w__4004 ,w__3941 ,w__3937);
  xnor g__3736(w__4003 ,w__3943 ,w__3934);
  not g__3737(w__3992 ,w__3993);
  nor g__3738(w__3990 ,w__3674 ,w__3941);
  and g__3739(w__3989 ,w__3674 ,w__3941);
  or g__3740(w__3988 ,w__3946 ,w__3948);
  and g__3741(w__3987 ,w__3893 ,w__3944);
  or g__3742(w__3986 ,w__3893 ,w__3944);
  and g__3743(w__3985 ,w__3896 ,w__3942);
  or g__3744(w__3984 ,w__3896 ,w__3942);
  nor g__3745(w__3983 ,w__3789 ,w__3481);
  and g__3746(w__3982 ,w__3876 ,w__3943);
  or g__3747(w__3981 ,w__3876 ,w__3943);
  and g__3748(w__3995 ,w__3919 ,w__3955);
  and g__3749(w__3994 ,w__3921 ,w__3949);
  or g__3750(w__3993 ,w__3925 ,w__3953);
  or g__3751(w__3991 ,w__3892 ,w__3956);
  not g__3752(w__3975 ,w__3976);
  not g__3753(w__3973 ,w__3974);
  not g__3754(w__3970 ,w__3971);
  not g__3755(w__3969 ,w__3968);
  not g__3756(w__3966 ,w__3967);
  not g__3757(w__3964 ,w__3965);
  or g__3758(w__3963 ,w__3788 ,w__3945);
  xnor g__3759(w__8418 ,w__3931 ,w__3865);
  xnor g__3760(w__3962 ,w__3882 ,w__3930);
  xnor g__3761(w__3961 ,w__3916 ,w__3879);
  and g__3762(w__3980 ,w__3910 ,w__3940);
  or g__3763(w__3979 ,w__3840 ,w__3939);
  and g__3764(w__3978 ,w__3906 ,w__3958);
  and g__3765(w__3977 ,w__3927 ,w__3957);
  xnor g__3766(w__3976 ,w__3902 ,w__3642);
  xnor g__3767(w__3974 ,w__3880 ,w__3901);
  xnor g__3768(w__3972 ,w__3915 ,w__3900);
  xnor g__3769(w__3971 ,w__3870 ,w__3903);
  and g__3770(w__3968 ,w__3918 ,w__3959);
  xnor g__3771(w__3967 ,w__3872 ,w__3905);
  xnor g__3772(w__3965 ,w__3848 ,w__3904);
  or g__3773(w__3959 ,w__3916 ,w__3924);
  or g__3774(w__3958 ,w__3861 ,w__3928);
  or g__3775(w__3957 ,w__3932 ,w__3920);
  nor g__3776(w__3956 ,w__3891 ,w__3915);
  or g__3777(w__3955 ,w__3847 ,w__3911);
  or g__3778(w__3954 ,w__3673 ,w__3912);
  nor g__3779(w__3953 ,w__3923 ,w__3933);
  or g__3780(w__3952 ,w__3930 ,w__3882);
  and g__3781(w__3951 ,w__3930 ,w__3882);
  or g__3782(w__3950 ,w__3873 ,w__3914);
  or g__3783(w__3949 ,w__3926 ,w__3917);
  nor g__3784(w__3948 ,w__3874 ,w__3913);
  or g__3785(w__3960 ,w__3843 ,w__3908);
  not g__3786(w__3945 ,w__3481);
  or g__3787(w__3940 ,w__3846 ,w__3909);
  nor g__3788(w__3939 ,w__3853 ,w__3931);
  xnor g__3789(w__3938 ,w__3877 ,w__3859);
  xnor g__3790(w__3937 ,w__3897 ,w__3611);
  xnor g__3791(w__3936 ,w__3895 ,w__3626);
  xnor g__3792(w__3935 ,w__3875 ,w__3894);
  xor g__3793(w__3934 ,w__3876 ,w__3898);
  and g__3794(w__3947 ,w__3841 ,w__3907);
  and g__3795(w__3946 ,w__3886 ,w__3922);
  xnor g__3796(w__3944 ,w__3899 ,w__3480);
  xnor g__3797(w__3943 ,w__3863 ,w__3867);
  xnor g__3798(w__3942 ,w__3866 ,w__3613);
  xnor g__3799(w__3941 ,w__3883 ,w__3869);
  or g__3800(w__3929 ,w__3661 ,w__3871);
  and g__3801(w__3928 ,w__3766 ,w__3870);
  or g__3802(w__3927 ,w__3859 ,w__3877);
  and g__3803(w__3926 ,w__3894 ,w__3875);
  and g__3804(w__3925 ,w__3626 ,w__3895);
  nor g__3805(w__3924 ,w__3639 ,w__3879);
  nor g__3806(w__3923 ,w__3625 ,w__3895);
  or g__3807(w__3922 ,w__3848 ,w__3889);
  or g__3808(w__3921 ,w__3894 ,w__3875);
  and g__3809(w__3920 ,w__3859 ,w__3877);
  or g__3810(w__3919 ,w__3690 ,w__3881);
  or g__3811(w__3918 ,w__3662 ,w__3878);
  and g__3812(w__3933 ,w__3852 ,w__3888);
  and g__3813(w__3932 ,w__3755 ,w__3890);
  and g__3814(w__3930 ,w__3781 ,w__3887);
  not g__3815(w__3913 ,w__3914);
  and g__3816(w__3911 ,w__3690 ,w__3881);
  or g__3817(w__3910 ,w__3783 ,w__3872);
  and g__3818(w__3909 ,w__3783 ,w__3872);
  and g__3819(w__3908 ,w__3838 ,w__3899);
  or g__3820(w__3907 ,w__3844 ,w__3883);
  or g__3821(w__3906 ,w__3766 ,w__3870);
  xnor g__3822(w__3905 ,w__3783 ,w__3846);
  xnor g__3823(w__3904 ,w__3719 ,w__3845);
  xor g__3824(w__3903 ,w__3766 ,w__3861);
  xnor g__3825(w__3902 ,w__3862 ,w__3720);
  xnor g__3826(w__3901 ,w__3690 ,w__3847);
  xnor g__3827(w__3900 ,w__3858 ,w__3609);
  xnor g__3828(w__3917 ,w__3810 ,w__3836);
  and g__3829(w__3916 ,w__3746 ,w__3885);
  xnor g__3830(w__3915 ,w__3484 ,w__3835);
  xnor g__3831(w__3914 ,w__3860 ,w__3793);
  xnor g__3832(w__3912 ,w__3849 ,w__3797);
  nor g__3833(w__3892 ,w__3679 ,w__3858);
  and g__3834(w__3891 ,w__3679 ,w__3858);
  or g__3835(w__3890 ,w__3750 ,w__3860);
  and g__3836(w__3889 ,w__3719 ,w__3845);
  or g__3837(w__3888 ,w__3863 ,w__3857);
  or g__3838(w__3887 ,w__3485 ,w__3862);
  or g__3839(w__3886 ,w__3719 ,w__3845);
  or g__3840(w__3885 ,w__3776 ,w__3849);
  xnor g__3841(w__3884 ,w__3686 ,w__3809);
  xnor g__3842(w__3899 ,w__3767 ,w__3792);
  and g__3843(w__3898 ,w__3818 ,w__3837);
  and g__3844(w__3897 ,w__3825 ,w__3850);
  or g__3845(w__3896 ,w__3780 ,w__3851);
  xnor g__3846(w__3895 ,w__3687 ,w__3813);
  and g__3847(w__3894 ,w__3760 ,w__3839);
  or g__3848(w__3893 ,w__3829 ,w__3854);
  not g__3849(w__3881 ,w__3880);
  not g__3850(w__3878 ,w__3879);
  not g__3851(w__3873 ,w__3874);
  xnor g__3852(w__3869 ,w__3765 ,w__3808);
  xnor g__3853(w__3868 ,w__3832 ,w__3645);
  xnor g__3854(w__3867 ,w__3787 ,w__3803);
  xnor g__3855(w__3866 ,w__3487 ,w__3785);
  xnor g__3856(w__3865 ,w__3786 ,w__3833);
  xnor g__3857(w__3864 ,w__3805 ,w__3652);
  xnor g__3858(w__3883 ,w__3684 ,w__3794);
  xnor g__3859(w__3882 ,w__3812 ,w__3623);
  xnor g__3860(w__3880 ,w__3721 ,w__3799);
  xnor g__3861(w__3879 ,w__3715 ,w__3796);
  xnor g__3862(w__3877 ,w__3697 ,w__3790);
  xnor g__3863(w__3876 ,w__3692 ,w__3791);
  xnor g__3864(w__3875 ,w__3717 ,w__3802);
  xnor g__3865(w__3874 ,w__3696 ,w__3800);
  xnor g__3866(w__3872 ,w__3486 ,w__3795);
  xnor g__3867(w__3871 ,w__3716 ,w__3798);
  xnor g__3868(w__3870 ,w__3736 ,w__3801);
  and g__3869(w__3857 ,w__3787 ,w__3803);
  or g__3870(w__3856 ,w__3666 ,w__3831);
  or g__3871(w__3855 ,w__3664 ,w__3804);
  nor g__3872(w__3854 ,w__3819 ,w__3487);
  and g__3873(w__3853 ,w__3786 ,w__3834);
  or g__3874(w__3852 ,w__3787 ,w__3803);
  and g__3875(w__3851 ,w__3778 ,w__3809);
  or g__3876(w__3850 ,w__3827 ,w__3484);
  and g__3877(w__3863 ,w__3759 ,w__3821);
  and g__3878(w__3862 ,w__3775 ,w__3814);
  and g__3879(w__3861 ,w__3747 ,w__3828);
  and g__3880(w__3860 ,w__3777 ,w__3820);
  and g__3881(w__3859 ,w__3771 ,w__3826);
  and g__3882(w__3858 ,w__3753 ,w__3824);
  nor g__3883(w__3844 ,w__3765 ,w__3808);
  and g__3884(w__3843 ,w__3615 ,w__3806);
  nor g__3885(w__3842 ,w__3644 ,w__3832);
  or g__3886(w__3841 ,w__3764 ,w__3807);
  nor g__3887(w__3840 ,w__3786 ,w__3834);
  or g__3888(w__3839 ,w__3749 ,w__3486);
  or g__3889(w__3838 ,w__3615 ,w__3806);
  or g__3890(w__3837 ,w__3811 ,w__3830);
  xnor g__3891(w__3836 ,w__3728 ,w__3763);
  xnor g__3892(w__3835 ,w__3694 ,w__3784);
  and g__3893(w__3849 ,w__3770 ,w__3823);
  and g__3894(w__3848 ,w__3748 ,w__3816);
  and g__3895(w__3847 ,w__3757 ,w__3822);
  and g__3896(w__3846 ,w__3761 ,w__3815);
  and g__3897(w__3845 ,w__3773 ,w__3817);
  not g__3898(w__3834 ,w__3833);
  not g__3899(w__3832 ,w__3831);
  nor g__3900(w__3830 ,w__3727 ,w__3763);
  nor g__3901(w__3829 ,w__3663 ,w__3785);
  or g__3902(w__3828 ,w__3699 ,w__3754);
  and g__3903(w__3827 ,w__3694 ,w__3784);
  or g__3904(w__3826 ,w__3700 ,w__3769);
  or g__3905(w__3825 ,w__3694 ,w__3784);
  or g__3906(w__3823 ,w__3733 ,w__3768);
  or g__3907(w__3822 ,w__3734 ,w__3751);
  or g__3908(w__3821 ,w__3701 ,w__3758);
  or g__3909(w__3820 ,w__3707 ,w__3756);
  and g__3910(w__3819 ,w__3663 ,w__3785);
  or g__3911(w__3818 ,w__3728 ,w__3762);
  or g__3912(w__3817 ,w__3708 ,w__3774);
  or g__3913(w__3816 ,w__3736 ,w__3745);
  or g__3914(w__3815 ,w__3703 ,w__3752);
  or g__3915(w__3814 ,w__3735 ,w__3772);
  xnor g__3916(w__3813 ,w__3708 ,in1[6]);
  xnor g__3917(w__3812 ,w__3709 ,in1[10]);
  xnor g__3918(w__3833 ,w__3739 ,w__3607);
  and g__3919(w__3831 ,w__3681 ,w__3782);
  not g__3920(w__3811 ,w__3810);
  not g__3921(w__3807 ,w__3808);
  not g__3922(w__3804 ,w__3805);
  xnor g__3923(w__3802 ,w__3695 ,w__3701);
  xnor g__3924(w__3801 ,w__3682 ,w__3723);
  xnor g__3925(w__3800 ,w__3700 ,in1[7]);
  xnor g__3926(w__3799 ,w__3733 ,in1[8]);
  xnor g__3927(w__3798 ,w__3688 ,w__3707);
  xnor g__3928(w__3797 ,w__3718 ,w__3689);
  xnor g__3929(w__3796 ,w__3735 ,in1[9]);
  xnor g__3930(w__3795 ,w__3725 ,w__3726);
  xnor g__3931(w__3794 ,w__3714 ,w__3703);
  xnor g__3932(w__3793 ,w__3683 ,w__3691);
  xnor g__3933(w__3792 ,w__3693 ,w__3724);
  xnor g__3934(w__3791 ,w__3722 ,w__3699);
  xnor g__3935(w__3790 ,w__3713 ,w__3734);
  xnor g__3936(w__3810 ,w__3741 ,in1[5]);
  xnor g__3937(w__3809 ,w__3702 ,in1[2]);
  xnor g__3938(w__3808 ,w__3706 ,in1[4]);
  xnor g__3939(w__3806 ,w__3738 ,in1[3]);
  xnor g__3940(w__3805 ,w__3731 ,in1[1]);
  xnor g__3941(w__3803 ,w__3737 ,w__3711);
  not g__3942(w__3789 ,w__3788);
  or g__3943(w__3782 ,w__3709 ,w__3712);
  or g__3944(w__3781 ,w__3680 ,w__3720);
  nor g__3945(w__3780 ,w__3667 ,w__3686);
  or g__3946(w__3779 ,w__3603 ,w__3705);
  or g__3947(w__3778 ,w__3617 ,w__3685);
  or g__3948(w__3777 ,w__3688 ,w__3716);
  and g__3949(w__3776 ,w__3718 ,w__3689);
  or g__3950(w__3775 ,w__3494 ,w__3715);
  and g__3951(w__3774 ,w__3514 ,w__3687);
  or g__3952(w__3773 ,w__3518 ,w__3687);
  and g__3953(w__3772 ,w__3498 ,w__3715);
  or g__3954(w__3771 ,w__3504 ,w__3696);
  or g__3955(w__3770 ,w__3543 ,w__3721);
  and g__3956(w__3769 ,w__3508 ,w__3696);
  and g__3957(w__3768 ,w__3530 ,w__3721);
  and g__3958(w__3788 ,w__3607 ,w__3740);
  or g__3959(w__3787 ,w__3551 ,w__3741);
  or g__3960(w__3786 ,w__3561 ,w__3731);
  or g__3961(w__3785 ,w__3570 ,w__3702);
  or g__3962(w__3784 ,w__3564 ,w__3738);
  or g__3963(w__3783 ,w__3567 ,w__3706);
  not g__3964(w__3764 ,w__3765);
  not g__3965(w__3762 ,w__3763);
  or g__3966(w__3761 ,w__3684 ,w__3714);
  or g__3967(w__3760 ,w__3725 ,w__3726);
  or g__3968(w__3759 ,w__3717 ,w__3695);
  and g__3969(w__3758 ,w__3717 ,w__3695);
  or g__3970(w__3757 ,w__3713 ,w__3697);
  and g__3971(w__3756 ,w__3688 ,w__3716);
  or g__3972(w__3755 ,w__3683 ,w__3691);
  and g__3973(w__3754 ,w__3692 ,w__3722);
  or g__3974(w__3753 ,w__3693 ,w__3724);
  and g__3975(w__3752 ,w__3684 ,w__3714);
  and g__3976(w__3751 ,w__3713 ,w__3697);
  and g__3977(w__3750 ,w__3683 ,w__3691);
  and g__3978(w__3749 ,w__3725 ,w__3726);
  or g__3979(w__3748 ,w__3682 ,w__3723);
  or g__3980(w__3747 ,w__3692 ,w__3722);
  or g__3981(w__3746 ,w__3718 ,w__3689);
  and g__3982(w__3745 ,w__3682 ,w__3723);
  and g__3983(w__3767 ,w__3742 ,w__3698);
  or g__3984(w__3766 ,w__3737 ,w__3711);
  and g__3985(w__3765 ,w__3710 ,w__3730);
  and g__3986(w__3763 ,w__3732 ,w__3744);
  not g__3987(w__3744 ,w__3743);
  not g__3988(w__3740 ,w__3739);
  not g__3989(w__3730 ,w__3729);
  not g__3990(w__3728 ,w__3727);
  nor g__3991(w__3712 ,in1[10] ,w__3622);
  or g__3992(w__3743 ,w__3527 ,w__3546);
  and g__3993(w__3742 ,in1[3] ,in1[1]);
  or g__3994(w__3741 ,w__3496 ,w__3548);
  or g__3995(w__3739 ,w__3532 ,w__3578);
  or g__3996(w__3738 ,w__3553 ,w__3581);
  or g__3997(w__3737 ,w__3516 ,w__3535);
  or g__3998(w__3736 ,w__3556 ,w__3593);
  or g__3999(w__3735 ,w__3541 ,w__3506);
  or g__4000(w__3734 ,w__3524 ,w__3591);
  or g__4001(w__3733 ,w__3521 ,w__3573);
  and g__4002(w__3732 ,in1[5] ,in1[3]);
  or g__4003(w__3731 ,w__3558 ,w__3548);
  or g__4004(w__3729 ,w__3511 ,w__3546);
  and g__4005(w__3727 ,in1[8] ,in1[1]);
  or g__4006(w__3726 ,w__3501 ,w__3559);
  or g__4007(w__3725 ,w__3595 ,w__3571);
  or g__4008(w__3724 ,w__3568 ,w__3562);
  or g__4009(w__3723 ,w__3583 ,w__3538);
  or g__4010(w__3722 ,w__3529 ,w__3533);
  or g__4011(w__3721 ,w__3601 ,w__3511);
  or g__4012(w__3720 ,w__3586 ,w__3527);
  or g__4013(w__3719 ,w__3526 ,w__3536);
  or g__4014(w__3718 ,w__3556 ,w__3598);
  or g__4015(w__3717 ,w__3576 ,w__3567);
  or g__4016(w__3716 ,w__3602 ,w__3589);
  or g__4017(w__3715 ,w__3555 ,w__3583);
  or g__4018(w__3714 ,w__3553 ,w__3570);
  or g__4019(w__3713 ,w__3530 ,w__3596);
  not g__4020(w__3705 ,w__3704);
  not g__4021(w__3686 ,w__3685);
  or g__4022(w__3681 ,w__3523 ,w__3676);
  or g__4023(w__3711 ,w__3521 ,w__3578);
  and g__4024(w__3710 ,in1[4] ,in1[2]);
  or g__4025(w__3709 ,w__3520 ,w__3498);
  or g__4026(w__3708 ,w__3586 ,w__3558);
  or g__4027(w__3707 ,w__3524 ,w__3593);
  or g__4028(w__3706 ,w__3501 ,w__3581);
  or g__4029(w__3704 ,w__3579 ,w__3654);
  or g__4030(w__3703 ,w__3510 ,w__3561);
  or g__4031(w__3702 ,w__3565 ,w__3545);
  or g__4032(w__3701 ,w__3599 ,w__3571);
  or g__4033(w__3700 ,w__3587 ,w__3539);
  or g__4034(w__3699 ,w__3494 ,w__3559);
  and g__4035(w__3698 ,in1[4] ,in1[0]);
  or g__4036(w__3697 ,w__3496 ,w__3551);
  or g__4037(w__3696 ,w__3584 ,w__3573);
  or g__4038(w__3695 ,w__3518 ,w__3564);
  or g__4039(w__3694 ,w__3576 ,w__3562);
  or g__4040(w__3693 ,w__3589 ,w__3533);
  or g__4041(w__3692 ,w__3500 ,w__3565);
  or g__4042(w__3691 ,w__3493 ,w__3591);
  or g__4043(w__3690 ,w__3543 ,w__3508);
  or g__4044(w__3689 ,w__3541 ,w__3514);
  or g__4045(w__3688 ,w__3504 ,w__3574);
  or g__4046(w__3687 ,w__3506 ,w__3568);
  and g__4047(w__3685 ,in1[2] ,in1[1]);
  or g__4048(w__3684 ,w__3536 ,w__3539);
  or g__4049(w__3683 ,w__3503 ,w__3516);
  or g__4050(w__3682 ,w__3513 ,w__3550);
  not g__4051(w__3680 ,w__3642);
  not g__4052(w__3679 ,w__3609);
  not g__4053(w__3678 ,w__3647);
  not g__4054(w__3677 ,w__3631);
  not g__4055(w__3676 ,w__3623);
  not g__4056(w__3675 ,w__3650);
  not g__4057(w__3674 ,w__3611);
  not g__4058(w__3673 ,w__3633);
  not g__4059(w__3672 ,in1[0]);
  not g__4060(w__3671 ,in1[4]);
  not g__4061(w__3670 ,in1[1]);
  not g__4062(w__3669 ,in1[8]);
  not g__4063(w__3668 ,in1[9]);
  not g__4064(w__3667 ,w__3617);
  not g__4065(w__3666 ,w__3645);
  not g__4066(w__3665 ,w__3635);
  not g__4067(w__3664 ,w__3652);
  not g__4068(w__3663 ,w__3613);
  not g__4069(w__3662 ,w__3640);
  not g__4070(w__3661 ,w__3637);
  not g__4071(w__3660 ,in1[3]);
  not g__4072(w__3659 ,in1[5]);
  not g__4073(w__3658 ,in1[2]);
  not g__4074(w__3657 ,in1[7]);
  not g__4075(w__3656 ,in1[6]);
  not g__4076(w__3655 ,in1[10]);
  not g__4077(w__3652 ,w__3651);
  not g__4078(w__3651 ,w__8512);
  not g__4079(w__3650 ,w__3648);
  not g__4080(w__3649 ,w__3648);
  not g__4081(w__3648 ,w__8526);
  not g__4082(w__3647 ,w__3646);
  not g__4083(w__3646 ,w__8525);
  not g__4084(w__3645 ,w__3643);
  not g__4085(w__3644 ,w__3643);
  not g__4086(w__3643 ,w__8531);
  not g__4087(w__3642 ,w__3641);
  not g__4088(w__3641 ,w__8529);
  not g__4089(w__3640 ,w__3638);
  not g__4090(w__3639 ,w__3638);
  not g__4091(w__3638 ,w__8528);
  not g__4092(w__3637 ,w__3636);
  not g__4093(w__3636 ,w__8523);
  not g__4094(w__3635 ,w__3634);
  not g__4095(w__3634 ,w__8520);
  not g__4096(w__3633 ,w__3632);
  not g__4097(w__3632 ,w__8527);
  not g__4098(w__3631 ,w__3630);
  not g__4099(w__3630 ,w__8519);
  not g__4100(w__3629 ,w__3627);
  not g__4101(w__3628 ,w__3627);
  not g__4102(w__3627 ,w__8524);
  not g__4103(w__3626 ,w__3624);
  not g__4104(w__3625 ,w__3624);
  not g__4105(w__3624 ,w__8522);
  not g__4106(w__3623 ,w__3621);
  not g__4107(w__3622 ,w__3621);
  not g__4108(w__3621 ,w__8530);
  not g__4109(w__3620 ,w__3618);
  not g__4110(w__3619 ,w__3618);
  not g__4111(w__3618 ,w__8521);
  not g__4112(w__3617 ,w__3616);
  not g__4113(w__3616 ,w__8514);
  not g__4114(w__3615 ,w__3614);
  not g__4115(w__3614 ,w__8516);
  not g__4116(w__3613 ,w__3612);
  not g__4117(w__3612 ,w__8515);
  not g__4118(w__3611 ,w__3610);
  not g__4119(w__3610 ,w__8518);
  not g__4120(w__3609 ,w__3608);
  not g__4121(w__3608 ,w__8517);
  not g__4122(w__3607 ,w__3606);
  not g__4123(w__3606 ,w__8513);
  not g__4124(w__3605 ,w__3604);
  not g__4125(w__3604 ,w__8532);
  not g__4126(w__3654 ,w__8510);
  not g__4127(w__3603 ,w__3653);
  not g__4128(w__3653 ,w__8511);
  not g__4129(w__3602 ,w__3600);
  not g__4130(w__3601 ,w__3600);
  not g__4131(w__3600 ,w__3668);
  not g__4132(w__3599 ,w__3597);
  not g__4133(w__3598 ,w__3597);
  not g__4134(w__3597 ,w__3657);
  not g__4135(w__3596 ,w__3594);
  not g__4136(w__3595 ,w__3594);
  not g__4137(w__3594 ,w__3656);
  not g__4138(w__3593 ,w__3592);
  not g__4139(w__3592 ,w__3658);
  not g__4140(w__3591 ,w__3590);
  not g__4141(w__3590 ,w__3671);
  not g__4142(w__3589 ,w__3588);
  not g__4143(w__3588 ,w__3660);
  not g__4144(w__3587 ,w__3585);
  not g__4145(w__3586 ,w__3585);
  not g__4146(w__3585 ,w__3655);
  not g__4147(w__3584 ,w__3582);
  not g__4148(w__3583 ,w__3582);
  not g__4149(w__3582 ,w__3669);
  not g__4150(w__3581 ,w__3580);
  not g__4151(w__3580 ,w__3672);
  not g__4152(w__3579 ,w__3577);
  not g__4153(w__3578 ,w__3577);
  not g__4154(w__3577 ,w__3672);
  not g__4155(w__3576 ,w__3575);
  not g__4156(w__3575 ,w__3659);
  not g__4157(w__3574 ,w__3572);
  not g__4158(w__3573 ,w__3572);
  not g__4159(w__3572 ,w__3659);
  not g__4160(w__3571 ,w__3569);
  not g__4161(w__3570 ,w__3569);
  not g__4162(w__3569 ,w__3658);
  not g__4163(w__3568 ,w__3566);
  not g__4164(w__3567 ,w__3566);
  not g__4165(w__3566 ,w__3671);
  not g__4166(w__3565 ,w__3563);
  not g__4167(w__3564 ,w__3563);
  not g__4168(w__3563 ,w__3660);
  not g__4169(w__3562 ,w__3560);
  not g__4170(w__3561 ,w__3560);
  not g__4171(w__3560 ,w__3670);
  not g__4172(w__3559 ,w__3557);
  not g__4173(w__3558 ,w__3557);
  not g__4174(w__3557 ,w__3670);
  not g__4175(w__3556 ,w__3554);
  not g__4176(w__3555 ,w__3554);
  not g__4177(w__3554 ,w__3668);
  not g__4178(w__3553 ,w__3552);
  not g__4179(w__3552 ,w__3574);
  not g__4180(w__3551 ,w__3549);
  not g__4181(w__3550 ,w__3549);
  not g__4182(w__3549 ,w__3659);
  not g__4183(w__3548 ,w__3547);
  not g__4184(w__3547 ,w__3579);
  not g__4185(w__3546 ,w__3544);
  not g__4186(w__3545 ,w__3544);
  not g__4187(w__3544 ,w__3672);
  not g__4188(w__3543 ,w__3542);
  not g__4189(w__3542 ,w__3584);
  not g__4190(w__3541 ,w__3540);
  not g__4191(w__3540 ,w__3587);
  not g__4192(w__3539 ,w__3537);
  not g__4193(w__3538 ,w__3537);
  not g__4194(w__3537 ,w__3660);
  not g__4195(w__3536 ,w__3534);
  not g__4196(w__3535 ,w__3534);
  not g__4197(w__3534 ,w__3671);
  not g__4198(w__3533 ,w__3531);
  not g__4199(w__3532 ,w__3531);
  not g__4200(w__3531 ,w__3658);
  not g__4201(w__3530 ,w__3528);
  not g__4202(w__3529 ,w__3528);
  not g__4203(w__3528 ,w__3669);
  not g__4204(w__3527 ,w__3525);
  not g__4205(w__3526 ,w__3525);
  not g__4206(w__3525 ,w__3669);
  not g__4207(w__3524 ,w__3522);
  not g__4208(w__3523 ,w__3522);
  not g__4209(w__3522 ,w__3655);
  not g__4210(w__3521 ,w__3519);
  not g__4211(w__3520 ,w__3519);
  not g__4212(w__3519 ,w__3655);
  not g__4213(w__3518 ,w__3517);
  not g__4214(w__3517 ,w__3595);
  not g__4215(w__3516 ,w__3515);
  not g__4216(w__3515 ,w__3596);
  not g__4217(w__3514 ,w__3512);
  not g__4218(w__3513 ,w__3512);
  not g__4219(w__3512 ,w__3656);
  not g__4220(w__3511 ,w__3509);
  not g__4221(w__3510 ,w__3509);
  not g__4222(w__3509 ,w__3656);
  not g__4223(w__3508 ,w__3507);
  not g__4224(w__3507 ,w__3598);
  not g__4225(w__3506 ,w__3505);
  not g__4226(w__3505 ,w__3599);
  not g__4227(w__3504 ,w__3502);
  not g__4228(w__3503 ,w__3502);
  not g__4229(w__3502 ,w__3657);
  not g__4230(w__3501 ,w__3499);
  not g__4231(w__3500 ,w__3499);
  not g__4232(w__3499 ,w__3657);
  not g__4233(w__3498 ,w__3497);
  not g__4234(w__3497 ,w__3601);
  not g__4235(w__3496 ,w__3495);
  not g__4236(w__3495 ,w__3602);
  not g__4237(w__3494 ,w__3492);
  not g__4238(w__3493 ,w__3492);
  not g__4239(w__3492 ,w__3668);
  xor g__4240(w__8436 ,w__4151 ,w__3868);
  xor g__4241(w__8435 ,w__4149 ,w__3962);
  xor g__4242(w__8434 ,w__4147 ,w__4027);
  xor g__4243(w__8433 ,w__4145 ,w__4062);
  xor g__4244(w__8432 ,w__4143 ,w__4094);
  xor g__4245(w__8431 ,w__4141 ,w__4096);
  xor g__4246(w__8430 ,w__4139 ,w__4120);
  xor g__4247(w__8429 ,w__4137 ,w__4124);
  xor g__4248(w__8428 ,w__4135 ,w__4119);
  xor g__4249(w__8427 ,w__4133 ,w__4118);
  xor g__4250(w__8426 ,w__4131 ,w__4108);
  xor g__4251(w__3491 ,w__3971 ,w__4045);
  and g__4252(w__3490 ,w__3646 ,w__4007);
  and g__4253(w__3489 ,w__3632 ,w__3912);
  and g__4254(w__3488 ,w__3636 ,w__3871);
  xnor g__4255(w__3487 ,w__3742 ,w__3698);
  xor g__4256(w__3486 ,w__3732 ,w__3743);
  and g__4257(w__3485 ,w__3641 ,w__3720);
  xor g__4258(w__3484 ,w__3710 ,w__3729);
  xor g__4259(w__3483 ,w__3980 ,w__3634);
  xor g__4260(w__3482 ,w__3947 ,w__3630);
  xor g__4261(w__3481 ,w__3884 ,w__3616);
  xor g__4262(w__3480 ,w__3806 ,w__3614);
  xnor g__4263(w__8415 ,w__3654 ,in1[0]);
  xnor g__4264(w__8413 ,w__4831 ,w__4280);
  and g__4265(w__8414 ,w__4280 ,w__4832);
  not g__4266(w__4832 ,w__4831);
  and g__4267(w__4831 ,w__4533 ,w__4830);
  or g__4268(w__4830 ,w__4518 ,w__4829);
  and g__4269(w__4829 ,w__4630 ,w__4828);
  or g__4270(w__4828 ,w__4629 ,w__4827);
  and g__4271(w__4827 ,w__4678 ,w__4826);
  or g__4272(w__4826 ,w__4680 ,w__4825);
  and g__4273(w__4825 ,w__4735 ,w__4824);
  or g__4274(w__4824 ,w__4727 ,w__4823);
  and g__4275(w__4823 ,w__4761 ,w__4822);
  or g__4276(w__4822 ,w__4762 ,w__4821);
  and g__4277(w__4821 ,w__4769 ,w__4820);
  or g__4278(w__4820 ,w__4768 ,w__4819);
  and g__4279(w__4819 ,w__4793 ,w__4818);
  or g__4280(w__4818 ,w__4794 ,w__4817);
  and g__4281(w__4817 ,w__4800 ,w__4816);
  or g__4282(w__4816 ,w__4799 ,w__4815);
  and g__4283(w__4815 ,w__4792 ,w__4814);
  or g__4284(w__4814 ,w__4791 ,w__4813);
  and g__4285(w__4813 ,w__4790 ,w__4812);
  or g__4286(w__4812 ,w__4789 ,w__4811);
  and g__4287(w__4811 ,w__4780 ,w__4810);
  or g__4288(w__4810 ,w__4779 ,w__4809);
  and g__4289(w__4809 ,w__4766 ,w__4808);
  xnor g__4290(w__8401 ,w__4806 ,w__4773);
  or g__4291(w__4808 ,w__4760 ,w__4807);
  not g__4292(w__4807 ,w__4806);
  or g__4293(w__4806 ,w__4741 ,w__4805);
  xnor g__4294(w__8400 ,w__4804 ,w__4758);
  and g__4295(w__4805 ,w__4748 ,w__4804);
  or g__4296(w__4804 ,w__4718 ,w__4803);
  xnor g__4297(w__8399 ,w__4801 ,w__4726);
  and g__4298(w__4803 ,w__4717 ,w__4801);
  xnor g__4299(w__4802 ,w__4782 ,w__4788);
  or g__4300(w__4801 ,w__4696 ,w__4795);
  or g__4301(w__4800 ,w__4781 ,w__4787);
  nor g__4302(w__4799 ,w__4782 ,w__4788);
  xnor g__4303(w__4798 ,w__4784 ,w__4764);
  xnor g__4304(w__4797 ,w__4752 ,w__4776);
  xnor g__4305(w__4796 ,w__4754 ,w__4778);
  xnor g__4306(w__8398 ,w__4785 ,w__4704);
  and g__4307(w__4795 ,w__4695 ,w__4785);
  nor g__4308(w__4794 ,w__4784 ,w__4764);
  or g__4309(w__4793 ,w__4783 ,w__4763);
  or g__4310(w__4792 ,w__4751 ,w__4775);
  nor g__4311(w__4791 ,w__4752 ,w__4776);
  or g__4312(w__4790 ,w__4753 ,w__4777);
  nor g__4313(w__4789 ,w__4754 ,w__4778);
  not g__4314(w__4788 ,w__4787);
  xnor g__4315(w__4787 ,w__4712 ,w__4759);
  xnor g__4316(w__4786 ,w__4765 ,w__4756);
  not g__4317(w__4783 ,w__4784);
  not g__4318(w__4781 ,w__4782);
  or g__4319(w__4780 ,w__4756 ,w__4765);
  and g__4320(w__4779 ,w__4756 ,w__4765);
  or g__4321(w__4785 ,w__4665 ,w__4770);
  or g__4322(w__4784 ,w__4750 ,w__4767);
  or g__4323(w__4782 ,w__4691 ,w__4771);
  not g__4324(w__4778 ,w__4777);
  not g__4325(w__4776 ,w__4775);
  xnor g__4326(w__8397 ,w__4757 ,w__4675);
  xnor g__4327(w__4774 ,w__4742 ,w__4755);
  xnor g__4328(w__4773 ,w__4739 ,w__4746);
  xnor g__4329(w__4772 ,w__4737 ,w__4744);
  xnor g__4330(w__4777 ,w__4684 ,w__4166);
  xnor g__4331(w__4775 ,w__4747 ,w__4703);
  and g__4332(w__4771 ,w__4679 ,w__4747);
  and g__4333(w__4770 ,w__4664 ,w__4757);
  or g__4334(w__4769 ,w__4755 ,w__4742);
  and g__4335(w__4768 ,w__4755 ,w__4742);
  nor g__4336(w__4767 ,w__4712 ,w__4749);
  or g__4337(w__4766 ,w__4738 ,w__4745);
  not g__4338(w__4763 ,w__4764);
  nor g__4339(w__4762 ,w__4737 ,w__4744);
  or g__4340(w__4761 ,w__4736 ,w__4743);
  nor g__4341(w__4760 ,w__4739 ,w__4746);
  xnor g__4342(w__4759 ,w__4730 ,w__4304);
  xnor g__4343(w__4758 ,w__4710 ,w__4729);
  xnor g__4344(w__4765 ,w__4672 ,w__4725);
  xnor g__4345(w__4764 ,w__4700 ,w__4724);
  not g__4346(w__4753 ,w__4754);
  not g__4347(w__4752 ,w__4751);
  and g__4348(w__4750 ,w__4304 ,w__4730);
  nor g__4349(w__4749 ,w__4303 ,w__4730);
  or g__4350(w__4748 ,w__4710 ,w__4729);
  or g__4351(w__4757 ,w__4663 ,w__4731);
  and g__4352(w__4756 ,w__4720 ,w__4732);
  and g__4353(w__4755 ,w__4719 ,w__4734);
  or g__4354(w__4754 ,w__4715 ,w__4733);
  and g__4355(w__4751 ,w__4714 ,w__4728);
  not g__4356(w__4745 ,w__4746);
  not g__4357(w__4743 ,w__4744);
  xnor g__4358(w__8396 ,w__4722 ,w__4674);
  and g__4359(w__4741 ,w__4710 ,w__4729);
  xnor g__4360(w__4740 ,w__4711 ,w__4721);
  xnor g__4361(w__4747 ,w__4702 ,w__4312);
  xnor g__4362(w__4746 ,w__4687 ,w__4158);
  xnor g__4363(w__4744 ,w__4706 ,w__4308);
  xnor g__4364(w__4742 ,w__4655 ,w__4701);
  not g__4365(w__4739 ,w__4738);
  not g__4366(w__4737 ,w__4736);
  or g__4367(w__4735 ,w__4721 ,w__4711);
  or g__4368(w__4734 ,w__4700 ,w__4165);
  nor g__4369(w__4733 ,w__4672 ,w__4709);
  or g__4370(w__4732 ,w__4658 ,w__4716);
  and g__4371(w__4731 ,w__4662 ,w__4722);
  and g__4372(w__4738 ,w__4699 ,w__4707);
  and g__4373(w__4736 ,w__4689 ,w__4708);
  or g__4374(w__4728 ,w__4723 ,w__4713);
  xnor g__4375(w__8395 ,w__4657 ,w__4676);
  and g__4376(w__4727 ,w__4721 ,w__4711);
  xnor g__4377(w__4726 ,w__4669 ,w__4682);
  xnor g__4378(w__4725 ,w__4681 ,w__4295);
  xnor g__4379(w__4724 ,w__4685 ,w__4322);
  xnor g__4380(w__4730 ,w__4592 ,w__4677);
  xnor g__4381(w__4729 ,w__4645 ,w__4157);
  or g__4382(w__4720 ,w__4341 ,w__4687);
  or g__4383(w__4719 ,w__4354 ,w__4685);
  and g__4384(w__4718 ,w__4669 ,w__4682);
  or g__4385(w__4717 ,w__4669 ,w__4682);
  nor g__4386(w__4716 ,w__4310 ,w__4686);
  and g__4387(w__4715 ,w__4295 ,w__4681);
  or g__4388(w__4714 ,w__4648 ,w__4684);
  nor g__4389(w__4713 ,w__4649 ,w__4683);
  and g__4390(w__4723 ,w__4659 ,w__4690);
  or g__4391(w__4722 ,w__4661 ,w__4692);
  and g__4392(w__4721 ,w__4632 ,w__4693);
  nor g__4393(w__4709 ,w__4294 ,w__4681);
  or g__4394(w__4708 ,w__4655 ,w__4694);
  or g__4395(w__4707 ,w__4625 ,w__4698);
  xnor g__4396(w__4706 ,w__4673 ,w__4590);
  xnor g__4397(w__4705 ,w__4654 ,w__4647);
  xnor g__4398(w__4704 ,w__4638 ,w__4650);
  xnor g__4399(w__4703 ,w__4643 ,w__4671);
  xnor g__4400(w__4702 ,w__4656 ,w__4548);
  xnor g__4401(w__4701 ,w__4652 ,w__4325);
  and g__4402(w__4712 ,w__4607 ,w__4688);
  xnor g__4403(w__4711 ,w__4639 ,w__4315);
  or g__4404(w__4710 ,w__4668 ,w__4697);
  or g__4405(w__4699 ,w__4353 ,w__4645);
  nor g__4406(w__4698 ,w__4306 ,w__4644);
  nor g__4407(w__4697 ,w__4575 ,w__4667);
  and g__4408(w__4696 ,w__4638 ,w__4650);
  or g__4409(w__4695 ,w__4638 ,w__4650);
  nor g__4410(w__4694 ,w__4324 ,w__4652);
  or g__4411(w__4693 ,w__4164 ,w__4673);
  and g__4412(w__4692 ,w__4657 ,w__4641);
  nor g__4413(w__4691 ,w__4643 ,w__4670);
  or g__4414(w__4690 ,w__4576 ,w__4660);
  or g__4415(w__4689 ,w__4351 ,w__4651);
  or g__4416(w__4688 ,w__4163 ,w__4656);
  and g__4417(w__4700 ,w__4628 ,w__4666);
  not g__4418(w__4686 ,w__4687);
  not g__4419(w__4683 ,w__4684);
  nor g__4420(w__4680 ,w__4654 ,w__4647);
  or g__4421(w__4679 ,w__4642 ,w__4671);
  or g__4422(w__4678 ,w__4653 ,w__4646);
  xnor g__4423(w__4677 ,w__4551 ,w__4624);
  xnor g__4424(w__4676 ,w__4465 ,w__4156);
  xnor g__4425(w__4675 ,w__4571 ,w__4622);
  xnor g__4426(w__4674 ,w__4574 ,w__4620);
  xnor g__4427(w__4687 ,w__4595 ,w__4613);
  xnor g__4428(w__4685 ,w__4610 ,w__4616);
  xnor g__4429(w__4684 ,w__4611 ,w__4614);
  xnor g__4430(w__4682 ,w__4619 ,w__4615);
  xnor g__4431(w__4681 ,w__4621 ,w__4612);
  not g__4432(w__4670 ,w__4671);
  nor g__4433(w__4668 ,w__4350 ,w__4619);
  and g__4434(w__4667 ,w__4350 ,w__4619);
  or g__4435(w__4666 ,w__4624 ,w__4626);
  and g__4436(w__4665 ,w__4571 ,w__4622);
  or g__4437(w__4664 ,w__4571 ,w__4622);
  and g__4438(w__4663 ,w__4574 ,w__4620);
  or g__4439(w__4662 ,w__4574 ,w__4620);
  nor g__4440(w__4661 ,w__4465 ,w__4156);
  and g__4441(w__4660 ,w__4553 ,w__4621);
  or g__4442(w__4659 ,w__4553 ,w__4621);
  and g__4443(w__4673 ,w__4597 ,w__4633);
  and g__4444(w__4672 ,w__4599 ,w__4627);
  or g__4445(w__4671 ,w__4603 ,w__4631);
  or g__4446(w__4669 ,w__4570 ,w__4634);
  not g__4447(w__4653 ,w__4654);
  not g__4448(w__4651 ,w__4652);
  not g__4449(w__4648 ,w__4649);
  not g__4450(w__4647 ,w__4646);
  not g__4451(w__4644 ,w__4645);
  not g__4452(w__4642 ,w__4643);
  or g__4453(w__4641 ,w__4464 ,w__4623);
  xnor g__4454(w__8394 ,w__4609 ,w__4542);
  xnor g__4455(w__4640 ,w__4559 ,w__4608);
  xnor g__4456(w__4639 ,w__4594 ,w__4556);
  and g__4457(w__4658 ,w__4588 ,w__4618);
  or g__4458(w__4657 ,w__4516 ,w__4617);
  and g__4459(w__4656 ,w__4584 ,w__4636);
  and g__4460(w__4655 ,w__4605 ,w__4635);
  xnor g__4461(w__4654 ,w__4580 ,w__4317);
  xnor g__4462(w__4652 ,w__4557 ,w__4579);
  xnor g__4463(w__4650 ,w__4593 ,w__4578);
  xnor g__4464(w__4649 ,w__4547 ,w__4581);
  and g__4465(w__4646 ,w__4596 ,w__4637);
  xnor g__4466(w__4645 ,w__4549 ,w__4583);
  xnor g__4467(w__4643 ,w__4524 ,w__4582);
  or g__4468(w__4637 ,w__4594 ,w__4602);
  or g__4469(w__4636 ,w__4538 ,w__4606);
  or g__4470(w__4635 ,w__4610 ,w__4598);
  nor g__4471(w__4634 ,w__4569 ,w__4593);
  or g__4472(w__4633 ,w__4523 ,w__4589);
  or g__4473(w__4632 ,w__4349 ,w__4590);
  nor g__4474(w__4631 ,w__4601 ,w__4611);
  or g__4475(w__4630 ,w__4608 ,w__4559);
  and g__4476(w__4629 ,w__4608 ,w__4559);
  or g__4477(w__4628 ,w__4550 ,w__4592);
  or g__4478(w__4627 ,w__4604 ,w__4595);
  nor g__4479(w__4626 ,w__4551 ,w__4591);
  or g__4480(w__4638 ,w__4519 ,w__4586);
  not g__4481(w__4623 ,w__4156);
  or g__4482(w__4618 ,w__4522 ,w__4587);
  nor g__4483(w__4617 ,w__4530 ,w__4609);
  xor g__4484(w__8393 ,w__4459 ,w__4541);
  xnor g__4485(w__4616 ,w__4554 ,w__4536);
  xnor g__4486(w__4615 ,w__4575 ,w__4286);
  xnor g__4487(w__4614 ,w__4573 ,w__4301);
  xnor g__4488(w__4613 ,w__4552 ,w__4572);
  xor g__4489(w__4612 ,w__4553 ,w__4576);
  and g__4490(w__4625 ,w__4517 ,w__4585);
  and g__4491(w__4624 ,w__4563 ,w__4600);
  xnor g__4492(w__4622 ,w__4577 ,w__4155);
  xnor g__4493(w__4621 ,w__4540 ,w__4544);
  xnor g__4494(w__4620 ,w__4543 ,w__4288);
  xnor g__4495(w__4619 ,w__4560 ,w__4546);
  or g__4496(w__4607 ,w__4337 ,w__4548);
  and g__4497(w__4606 ,w__4442 ,w__4547);
  or g__4498(w__4605 ,w__4536 ,w__4554);
  and g__4499(w__4604 ,w__4572 ,w__4552);
  and g__4500(w__4603 ,w__4301 ,w__4573);
  nor g__4501(w__4602 ,w__4314 ,w__4556);
  nor g__4502(w__4601 ,w__4300 ,w__4573);
  or g__4503(w__4600 ,w__4524 ,w__4567);
  or g__4504(w__4599 ,w__4572 ,w__4552);
  and g__4505(w__4598 ,w__4536 ,w__4554);
  or g__4506(w__4597 ,w__4374 ,w__4558);
  or g__4507(w__4596 ,w__4338 ,w__4555);
  and g__4508(w__4611 ,w__4528 ,w__4566);
  and g__4509(w__4610 ,w__4431 ,w__4568);
  and g__4510(w__4609 ,w__4532 ,w__4564);
  and g__4511(w__4608 ,w__4456 ,w__4565);
  not g__4512(w__4591 ,w__4592);
  and g__4513(w__4589 ,w__4374 ,w__4558);
  or g__4514(w__4588 ,w__4458 ,w__4549);
  and g__4515(w__4587 ,w__4458 ,w__4549);
  and g__4516(w__4586 ,w__4514 ,w__4577);
  or g__4517(w__4585 ,w__4520 ,w__4560);
  or g__4518(w__4584 ,w__4442 ,w__4547);
  xnor g__4519(w__4583 ,w__4458 ,w__4522);
  xnor g__4520(w__4582 ,w__4395 ,w__4521);
  xor g__4521(w__4581 ,w__4442 ,w__4538);
  xnor g__4522(w__4580 ,w__4539 ,w__4396);
  xnor g__4523(w__4579 ,w__4374 ,w__4523);
  xnor g__4524(w__4578 ,w__4535 ,w__4284);
  xnor g__4525(w__4595 ,w__4486 ,w__4512);
  and g__4526(w__4594 ,w__4422 ,w__4562);
  xnor g__4527(w__4593 ,w__4159 ,w__4511);
  xnor g__4528(w__4592 ,w__4537 ,w__4469);
  xnor g__4529(w__4590 ,w__4525 ,w__4473);
  nor g__4530(w__4570 ,w__4355 ,w__4535);
  and g__4531(w__4569 ,w__4355 ,w__4535);
  or g__4532(w__4568 ,w__4426 ,w__4537);
  and g__4533(w__4567 ,w__4395 ,w__4521);
  or g__4534(w__4566 ,w__4540 ,w__4534);
  or g__4535(w__4565 ,w__4160 ,w__4539);
  or g__4536(w__4564 ,w__4459 ,w__4529);
  or g__4537(w__4563 ,w__4395 ,w__4521);
  or g__4538(w__4562 ,w__4452 ,w__4525);
  xnor g__4539(w__4561 ,w__4371 ,w__4485);
  xnor g__4540(w__4577 ,w__4443 ,w__4468);
  and g__4541(w__4576 ,w__4494 ,w__4513);
  and g__4542(w__4575 ,w__4501 ,w__4526);
  or g__4543(w__4574 ,w__4447 ,w__4527);
  xnor g__4544(w__4573 ,w__4361 ,w__4489);
  and g__4545(w__4572 ,w__4436 ,w__4515);
  or g__4546(w__4571 ,w__4505 ,w__4531);
  not g__4547(w__4558 ,w__4557);
  not g__4548(w__4555 ,w__4556);
  not g__4549(w__4550 ,w__4551);
  xnor g__4550(w__4546 ,w__4441 ,w__4484);
  xnor g__4551(w__4545 ,w__4508 ,w__4320);
  xnor g__4552(w__4544 ,w__4463 ,w__4479);
  xnor g__4553(w__4543 ,w__4161 ,w__4461);
  xnor g__4554(w__4542 ,w__4462 ,w__4509);
  xnor g__4555(w__4541 ,w__4481 ,w__4328);
  xnor g__4556(w__4560 ,w__4373 ,w__4470);
  xnor g__4557(w__4559 ,w__4488 ,w__4298);
  xnor g__4558(w__4557 ,w__4397 ,w__4475);
  xnor g__4559(w__4556 ,w__4391 ,w__4472);
  xnor g__4560(w__4554 ,w__4364 ,w__4466);
  xnor g__4561(w__4553 ,w__4366 ,w__4467);
  xnor g__4562(w__4552 ,w__4401 ,w__4478);
  xnor g__4563(w__4551 ,w__4359 ,w__4476);
  xnor g__4564(w__4549 ,w__4162 ,w__4471);
  xnor g__4565(w__4548 ,w__4392 ,w__4474);
  xnor g__4566(w__4547 ,w__4411 ,w__4477);
  and g__4567(w__4534 ,w__4463 ,w__4479);
  or g__4568(w__4533 ,w__4342 ,w__4507);
  or g__4569(w__4532 ,w__4340 ,w__4480);
  nor g__4570(w__4531 ,w__4495 ,w__4161);
  and g__4571(w__4530 ,w__4462 ,w__4510);
  nor g__4572(w__4529 ,w__4327 ,w__4481);
  or g__4573(w__4528 ,w__4463 ,w__4479);
  and g__4574(w__4527 ,w__4454 ,w__4485);
  or g__4575(w__4526 ,w__4503 ,w__4159);
  and g__4576(w__4540 ,w__4435 ,w__4497);
  and g__4577(w__4539 ,w__4451 ,w__4490);
  and g__4578(w__4538 ,w__4423 ,w__4504);
  and g__4579(w__4537 ,w__4453 ,w__4496);
  and g__4580(w__4536 ,w__4457 ,w__4502);
  and g__4581(w__4535 ,w__4429 ,w__4500);
  nor g__4582(w__4520 ,w__4441 ,w__4484);
  and g__4583(w__4519 ,w__4290 ,w__4482);
  nor g__4584(w__4518 ,w__4319 ,w__4508);
  or g__4585(w__4517 ,w__4440 ,w__4483);
  nor g__4586(w__4516 ,w__4462 ,w__4510);
  or g__4587(w__4515 ,w__4425 ,w__4162);
  or g__4588(w__4514 ,w__4290 ,w__4482);
  or g__4589(w__4513 ,w__4487 ,w__4506);
  xnor g__4590(w__4512 ,w__4404 ,w__4439);
  xnor g__4591(w__4511 ,w__4368 ,w__4460);
  and g__4592(w__4525 ,w__4446 ,w__4499);
  and g__4593(w__4524 ,w__4424 ,w__4492);
  and g__4594(w__4523 ,w__4433 ,w__4498);
  and g__4595(w__4522 ,w__4437 ,w__4491);
  and g__4596(w__4521 ,w__4449 ,w__4493);
  not g__4597(w__4510 ,w__4509);
  not g__4598(w__4508 ,w__4507);
  nor g__4599(w__4506 ,w__4403 ,w__4439);
  nor g__4600(w__4505 ,w__4339 ,w__4461);
  or g__4601(w__4504 ,w__4382 ,w__4430);
  and g__4602(w__4503 ,w__4368 ,w__4460);
  or g__4603(w__4502 ,w__4381 ,w__4445);
  or g__4604(w__4501 ,w__4368 ,w__4460);
  or g__4605(w__4499 ,w__4408 ,w__4444);
  or g__4606(w__4498 ,w__4409 ,w__4427);
  or g__4607(w__4497 ,w__4384 ,w__4434);
  or g__4608(w__4496 ,w__4377 ,w__4432);
  and g__4609(w__4495 ,w__4339 ,w__4461);
  or g__4610(w__4494 ,w__4404 ,w__4438);
  or g__4611(w__4493 ,w__4386 ,w__4450);
  or g__4612(w__4492 ,w__4411 ,w__4421);
  or g__4613(w__4491 ,w__4379 ,w__4428);
  or g__4614(w__4490 ,w__4410 ,w__4448);
  xnor g__4615(w__4489 ,w__4386 ,in8[6]);
  xnor g__4616(w__4488 ,w__4387 ,in8[10]);
  xnor g__4617(w__4509 ,w__4415 ,w__4282);
  and g__4618(w__4507 ,w__4357 ,w__4455);
  not g__4619(w__4487 ,w__4486);
  not g__4620(w__4483 ,w__4484);
  not g__4621(w__4480 ,w__4481);
  xnor g__4622(w__4478 ,w__4360 ,w__4384);
  xnor g__4623(w__4477 ,w__4365 ,w__4399);
  xnor g__4624(w__4476 ,w__4381 ,in8[7]);
  xnor g__4625(w__4475 ,w__4408 ,in8[8]);
  xnor g__4626(w__4474 ,w__4362 ,w__4377);
  xnor g__4627(w__4473 ,w__4394 ,w__4363);
  xnor g__4628(w__4472 ,w__4410 ,in8[9]);
  xnor g__4629(w__4471 ,w__4390 ,w__4402);
  xnor g__4630(w__4470 ,w__4393 ,w__4379);
  xnor g__4631(w__4469 ,w__4372 ,w__4369);
  xnor g__4632(w__4468 ,w__4367 ,w__4400);
  xnor g__4633(w__4467 ,w__4398 ,w__4382);
  xnor g__4634(w__4466 ,w__4358 ,w__4409);
  xnor g__4635(w__4486 ,w__4417 ,in8[5]);
  xnor g__4636(w__4485 ,w__4380 ,in8[2]);
  xnor g__4637(w__4484 ,w__4385 ,in8[4]);
  xnor g__4638(w__4482 ,w__4414 ,in8[3]);
  xnor g__4639(w__4481 ,w__4406 ,in8[1]);
  xnor g__4640(w__4479 ,w__4418 ,w__4375);
  not g__4641(w__4465 ,w__4464);
  or g__4642(w__4457 ,w__4179 ,w__4359);
  or g__4643(w__4456 ,w__4356 ,w__4396);
  or g__4644(w__4455 ,w__4387 ,w__4388);
  or g__4645(w__4454 ,w__4292 ,w__4370);
  or g__4646(w__4453 ,w__4362 ,w__4392);
  and g__4647(w__4452 ,w__4394 ,w__4363);
  or g__4648(w__4451 ,w__4169 ,w__4391);
  and g__4649(w__4450 ,w__4189 ,w__4361);
  or g__4650(w__4449 ,w__4193 ,w__4361);
  and g__4651(w__4448 ,w__4173 ,w__4391);
  nor g__4652(w__4447 ,w__4343 ,w__4371);
  or g__4653(w__4446 ,w__4218 ,w__4397);
  and g__4654(w__4445 ,w__4183 ,w__4359);
  and g__4655(w__4444 ,w__4205 ,w__4397);
  and g__4656(w__4464 ,w__4282 ,w__4416);
  or g__4657(w__4463 ,w__4226 ,w__4417);
  or g__4658(w__4462 ,w__4236 ,w__4406);
  or g__4659(w__4461 ,w__4245 ,w__4380);
  or g__4660(w__4460 ,w__4239 ,w__4414);
  or g__4661(w__4459 ,w__4329 ,w__4378);
  or g__4662(w__4458 ,w__4242 ,w__4385);
  not g__4663(w__4440 ,w__4441);
  not g__4664(w__4438 ,w__4439);
  and g__4665(w__8391 ,w__4378 ,w__4389);
  or g__4666(w__4437 ,w__4373 ,w__4393);
  or g__4667(w__4436 ,w__4390 ,w__4402);
  or g__4668(w__4435 ,w__4401 ,w__4360);
  and g__4669(w__4434 ,w__4401 ,w__4360);
  or g__4670(w__4433 ,w__4358 ,w__4364);
  and g__4671(w__4432 ,w__4362 ,w__4392);
  or g__4672(w__4431 ,w__4372 ,w__4369);
  and g__4673(w__4430 ,w__4366 ,w__4398);
  or g__4674(w__4429 ,w__4367 ,w__4400);
  and g__4675(w__4428 ,w__4373 ,w__4393);
  and g__4676(w__4427 ,w__4358 ,w__4364);
  and g__4677(w__4426 ,w__4372 ,w__4369);
  and g__4678(w__4425 ,w__4390 ,w__4402);
  or g__4679(w__4424 ,w__4365 ,w__4399);
  or g__4680(w__4423 ,w__4366 ,w__4398);
  or g__4681(w__4422 ,w__4394 ,w__4363);
  and g__4682(w__4421 ,w__4365 ,w__4399);
  and g__4683(w__4443 ,w__4405 ,w__4376);
  or g__4684(w__4442 ,w__4418 ,w__4375);
  and g__4685(w__4441 ,w__4383 ,w__4413);
  and g__4686(w__4439 ,w__4407 ,w__4420);
  not g__4687(w__4420 ,w__4419);
  not g__4688(w__4416 ,w__4415);
  not g__4689(w__4413 ,w__4412);
  not g__4690(w__4404 ,w__4403);
  or g__4691(w__4389 ,in8[0] ,w__4278);
  nor g__4692(w__4388 ,in8[10] ,w__4297);
  or g__4693(w__4419 ,w__4202 ,w__4221);
  or g__4694(w__4418 ,w__4191 ,w__4210);
  or g__4695(w__4417 ,w__4171 ,w__4223);
  or g__4696(w__4415 ,w__4207 ,w__4253);
  or g__4697(w__4414 ,w__4228 ,w__4256);
  or g__4698(w__4412 ,w__4186 ,w__4223);
  or g__4699(w__4411 ,w__4231 ,w__4268);
  or g__4700(w__4410 ,w__4216 ,w__4181);
  or g__4701(w__4409 ,w__4199 ,w__4266);
  or g__4702(w__4408 ,w__4196 ,w__4248);
  and g__4703(w__4407 ,in8[5] ,in8[3]);
  or g__4704(w__4406 ,w__4233 ,w__4221);
  and g__4705(w__4405 ,in8[3] ,in8[1]);
  and g__4706(w__4403 ,in8[8] ,in8[1]);
  or g__4707(w__4402 ,w__4176 ,w__4234);
  or g__4708(w__4401 ,w__4251 ,w__4243);
  or g__4709(w__4400 ,w__4211 ,w__4237);
  or g__4710(w__4399 ,w__4258 ,w__4213);
  or g__4711(w__4398 ,w__4204 ,w__4246);
  or g__4712(w__4397 ,w__4276 ,w__4270);
  or g__4713(w__4396 ,w__4261 ,w__4202);
  or g__4714(w__4395 ,w__4201 ,w__4242);
  or g__4715(w__4394 ,w__4231 ,w__4273);
  or g__4716(w__4393 ,w__4228 ,w__4208);
  or g__4717(w__4392 ,w__4277 ,w__4264);
  or g__4718(w__4391 ,w__4230 ,w__4258);
  or g__4719(w__4390 ,w__4186 ,w__4245);
  not g__4720(w__4371 ,w__4370);
  or g__4721(w__4357 ,w__4198 ,w__4352);
  or g__4722(w__4387 ,w__4196 ,w__4173);
  or g__4723(w__4386 ,w__4195 ,w__4233);
  or g__4724(w__4385 ,w__4176 ,w__4253);
  or g__4725(w__4384 ,w__4274 ,w__4268);
  and g__4726(w__4383 ,in8[4] ,in8[2]);
  or g__4727(w__4382 ,w__4169 ,w__4236);
  or g__4728(w__4381 ,w__4261 ,w__4240);
  or g__4729(w__4380 ,w__4214 ,w__4256);
  or g__4730(w__4379 ,w__4271 ,w__4234);
  or g__4731(w__4378 ,w__4254 ,w__4330);
  or g__4732(w__4377 ,w__4199 ,w__4246);
  and g__4733(w__4376 ,in8[4] ,in8[0]);
  or g__4734(w__4375 ,w__4262 ,w__4220);
  or g__4735(w__4374 ,w__4205 ,w__4175);
  or g__4736(w__4373 ,w__4266 ,w__4239);
  or g__4737(w__4372 ,w__4183 ,w__4185);
  and g__4738(w__4370 ,in8[2] ,in8[1]);
  or g__4739(w__4369 ,w__4171 ,w__4243);
  or g__4740(w__4368 ,w__4226 ,w__4237);
  or g__4741(w__4367 ,w__4264 ,w__4208);
  or g__4742(w__4366 ,w__4179 ,w__4240);
  or g__4743(w__4365 ,w__4193 ,w__4248);
  or g__4744(w__4364 ,w__4168 ,w__4251);
  or g__4745(w__4363 ,w__4216 ,w__4189);
  or g__4746(w__4362 ,w__4181 ,w__4249);
  or g__4747(w__4361 ,w__4178 ,w__4211);
  or g__4748(w__4360 ,w__4191 ,w__4214);
  or g__4749(w__4359 ,w__4259 ,w__4225);
  or g__4750(w__4358 ,w__4218 ,w__4188);
  not g__4751(w__4356 ,w__4317);
  not g__4752(w__4355 ,w__4284);
  not g__4753(w__4354 ,w__4322);
  not g__4754(w__4353 ,w__4306);
  not g__4755(w__4352 ,w__4298);
  not g__4756(w__4351 ,w__4325);
  not g__4757(w__4350 ,w__4286);
  not g__4758(w__4349 ,w__4308);
  not g__4759(w__4348 ,in8[0]);
  not g__4760(w__4347 ,in8[4]);
  not g__4761(w__4346 ,in8[1]);
  not g__4762(w__4345 ,in8[8]);
  not g__4763(w__4344 ,in8[9]);
  not g__4764(w__4343 ,w__4292);
  not g__4765(w__4342 ,w__4320);
  not g__4766(w__4341 ,w__4310);
  not g__4767(w__4340 ,w__4328);
  not g__4768(w__4339 ,w__4288);
  not g__4769(w__4338 ,w__4315);
  not g__4770(w__4337 ,w__4312);
  not g__4771(w__4336 ,in8[3]);
  not g__4772(w__4335 ,in8[5]);
  not g__4773(w__4334 ,in8[2]);
  not g__4774(w__4333 ,in8[7]);
  not g__4775(w__4332 ,in8[6]);
  not g__4776(w__4331 ,in8[10]);
  not g__4777(w__4328 ,w__4326);
  not g__4778(w__4327 ,w__4326);
  not g__4779(w__4326 ,w__8465);
  not g__4780(w__4325 ,w__4323);
  not g__4781(w__4324 ,w__4323);
  not g__4782(w__4323 ,w__8479);
  not g__4783(w__4322 ,w__4321);
  not g__4784(w__4321 ,w__8478);
  not g__4785(w__4320 ,w__4318);
  not g__4786(w__4319 ,w__4318);
  not g__4787(w__4318 ,w__8484);
  not g__4788(w__4317 ,w__4316);
  not g__4789(w__4316 ,w__8482);
  not g__4790(w__4315 ,w__4313);
  not g__4791(w__4314 ,w__4313);
  not g__4792(w__4313 ,w__8481);
  not g__4793(w__4312 ,w__4311);
  not g__4794(w__4311 ,w__8476);
  not g__4795(w__4310 ,w__4309);
  not g__4796(w__4309 ,w__8473);
  not g__4797(w__4308 ,w__4307);
  not g__4798(w__4307 ,w__8480);
  not g__4799(w__4306 ,w__4305);
  not g__4800(w__4305 ,w__8472);
  not g__4801(w__4304 ,w__4302);
  not g__4802(w__4303 ,w__4302);
  not g__4803(w__4302 ,w__8477);
  not g__4804(w__4301 ,w__4299);
  not g__4805(w__4300 ,w__4299);
  not g__4806(w__4299 ,w__8475);
  not g__4807(w__4298 ,w__4296);
  not g__4808(w__4297 ,w__4296);
  not g__4809(w__4296 ,w__8483);
  not g__4810(w__4295 ,w__4293);
  not g__4811(w__4294 ,w__4293);
  not g__4812(w__4293 ,w__8474);
  not g__4813(w__4292 ,w__4291);
  not g__4814(w__4291 ,w__8467);
  not g__4815(w__4290 ,w__4289);
  not g__4816(w__4289 ,w__8469);
  not g__4817(w__4288 ,w__4287);
  not g__4818(w__4287 ,w__8468);
  not g__4819(w__4286 ,w__4285);
  not g__4820(w__4285 ,w__8471);
  not g__4821(w__4284 ,w__4283);
  not g__4822(w__4283 ,w__8470);
  not g__4823(w__4329 ,w__8464);
  not g__4824(w__4282 ,w__4281);
  not g__4825(w__4281 ,w__8466);
  not g__4826(w__4280 ,w__4279);
  not g__4827(w__4279 ,w__8485);
  not g__4828(w__4278 ,w__4330);
  not g__4829(w__4330 ,w__8463);
  not g__4830(w__4277 ,w__4275);
  not g__4831(w__4276 ,w__4275);
  not g__4832(w__4275 ,w__4344);
  not g__4833(w__4274 ,w__4272);
  not g__4834(w__4273 ,w__4272);
  not g__4835(w__4272 ,w__4333);
  not g__4836(w__4271 ,w__4269);
  not g__4837(w__4270 ,w__4269);
  not g__4838(w__4269 ,w__4332);
  not g__4839(w__4268 ,w__4267);
  not g__4840(w__4267 ,w__4334);
  not g__4841(w__4266 ,w__4265);
  not g__4842(w__4265 ,w__4347);
  not g__4843(w__4264 ,w__4263);
  not g__4844(w__4263 ,w__4336);
  not g__4845(w__4262 ,w__4260);
  not g__4846(w__4261 ,w__4260);
  not g__4847(w__4260 ,w__4331);
  not g__4848(w__4259 ,w__4257);
  not g__4849(w__4258 ,w__4257);
  not g__4850(w__4257 ,w__4345);
  not g__4851(w__4256 ,w__4255);
  not g__4852(w__4255 ,w__4348);
  not g__4853(w__4254 ,w__4252);
  not g__4854(w__4253 ,w__4252);
  not g__4855(w__4252 ,w__4348);
  not g__4856(w__4251 ,w__4250);
  not g__4857(w__4250 ,w__4335);
  not g__4858(w__4249 ,w__4247);
  not g__4859(w__4248 ,w__4247);
  not g__4860(w__4247 ,w__4335);
  not g__4861(w__4246 ,w__4244);
  not g__4862(w__4245 ,w__4244);
  not g__4863(w__4244 ,w__4334);
  not g__4864(w__4243 ,w__4241);
  not g__4865(w__4242 ,w__4241);
  not g__4866(w__4241 ,w__4347);
  not g__4867(w__4240 ,w__4238);
  not g__4868(w__4239 ,w__4238);
  not g__4869(w__4238 ,w__4336);
  not g__4870(w__4237 ,w__4235);
  not g__4871(w__4236 ,w__4235);
  not g__4872(w__4235 ,w__4346);
  not g__4873(w__4234 ,w__4232);
  not g__4874(w__4233 ,w__4232);
  not g__4875(w__4232 ,w__4346);
  not g__4876(w__4231 ,w__4229);
  not g__4877(w__4230 ,w__4229);
  not g__4878(w__4229 ,w__4344);
  not g__4879(w__4228 ,w__4227);
  not g__4880(w__4227 ,w__4249);
  not g__4881(w__4226 ,w__4224);
  not g__4882(w__4225 ,w__4224);
  not g__4883(w__4224 ,w__4335);
  not g__4884(w__4223 ,w__4222);
  not g__4885(w__4222 ,w__4254);
  not g__4886(w__4221 ,w__4219);
  not g__4887(w__4220 ,w__4219);
  not g__4888(w__4219 ,w__4348);
  not g__4889(w__4218 ,w__4217);
  not g__4890(w__4217 ,w__4259);
  not g__4891(w__4216 ,w__4215);
  not g__4892(w__4215 ,w__4262);
  not g__4893(w__4214 ,w__4212);
  not g__4894(w__4213 ,w__4212);
  not g__4895(w__4212 ,w__4336);
  not g__4896(w__4211 ,w__4209);
  not g__4897(w__4210 ,w__4209);
  not g__4898(w__4209 ,w__4347);
  not g__4899(w__4208 ,w__4206);
  not g__4900(w__4207 ,w__4206);
  not g__4901(w__4206 ,w__4334);
  not g__4902(w__4205 ,w__4203);
  not g__4903(w__4204 ,w__4203);
  not g__4904(w__4203 ,w__4345);
  not g__4905(w__4202 ,w__4200);
  not g__4906(w__4201 ,w__4200);
  not g__4907(w__4200 ,w__4345);
  not g__4908(w__4199 ,w__4197);
  not g__4909(w__4198 ,w__4197);
  not g__4910(w__4197 ,w__4331);
  not g__4911(w__4196 ,w__4194);
  not g__4912(w__4195 ,w__4194);
  not g__4913(w__4194 ,w__4331);
  not g__4914(w__4193 ,w__4192);
  not g__4915(w__4192 ,w__4270);
  not g__4916(w__4191 ,w__4190);
  not g__4917(w__4190 ,w__4271);
  not g__4918(w__4189 ,w__4187);
  not g__4919(w__4188 ,w__4187);
  not g__4920(w__4187 ,w__4332);
  not g__4921(w__4186 ,w__4184);
  not g__4922(w__4185 ,w__4184);
  not g__4923(w__4184 ,w__4332);
  not g__4924(w__4183 ,w__4182);
  not g__4925(w__4182 ,w__4273);
  not g__4926(w__4181 ,w__4180);
  not g__4927(w__4180 ,w__4274);
  not g__4928(w__4179 ,w__4177);
  not g__4929(w__4178 ,w__4177);
  not g__4930(w__4177 ,w__4333);
  not g__4931(w__4176 ,w__4174);
  not g__4932(w__4175 ,w__4174);
  not g__4933(w__4174 ,w__4333);
  not g__4934(w__4173 ,w__4172);
  not g__4935(w__4172 ,w__4276);
  not g__4936(w__4171 ,w__4170);
  not g__4937(w__4170 ,w__4277);
  not g__4938(w__4169 ,w__4167);
  not g__4939(w__4168 ,w__4167);
  not g__4940(w__4167 ,w__4344);
  xor g__4941(w__8412 ,w__4829 ,w__4545);
  xor g__4942(w__8411 ,w__4827 ,w__4640);
  xor g__4943(w__8410 ,w__4825 ,w__4705);
  xor g__4944(w__8409 ,w__4823 ,w__4740);
  xor g__4945(w__8408 ,w__4821 ,w__4772);
  xor g__4946(w__8407 ,w__4819 ,w__4774);
  xor g__4947(w__8406 ,w__4817 ,w__4798);
  xor g__4948(w__8405 ,w__4815 ,w__4802);
  xor g__4949(w__8404 ,w__4813 ,w__4797);
  xor g__4950(w__8403 ,w__4811 ,w__4796);
  xor g__4951(w__8402 ,w__4809 ,w__4786);
  xor g__4952(w__4166 ,w__4649 ,w__4723);
  and g__4953(w__4165 ,w__4321 ,w__4685);
  and g__4954(w__4164 ,w__4307 ,w__4590);
  and g__4955(w__4163 ,w__4311 ,w__4548);
  xor g__4956(w__4162 ,w__4407 ,w__4419);
  xnor g__4957(w__4161 ,w__4405 ,w__4376);
  and g__4958(w__4160 ,w__4316 ,w__4396);
  xor g__4959(w__4159 ,w__4383 ,w__4412);
  xor g__4960(w__4158 ,w__4658 ,w__4309);
  xor g__4961(w__4157 ,w__4625 ,w__4305);
  xor g__4962(w__4156 ,w__4561 ,w__4291);
  xor g__4963(w__4155 ,w__4482 ,w__4289);
  xor g__4964(w__8392 ,w__4378 ,w__4329);
  or g__4965(w__8390 ,w__5663 ,w__5895);
  xnor g__4966(w__8389 ,w__5894 ,w__5680);
  and g__4967(w__5895 ,w__5662 ,w__5894);
  or g__4968(w__5894 ,w__5735 ,w__5893);
  xnor g__4969(w__8388 ,w__5892 ,w__5745);
  and g__4970(w__5893 ,w__5736 ,w__5892);
  or g__4971(w__5892 ,w__5786 ,w__5891);
  xnor g__4972(w__8387 ,w__5890 ,w__5798);
  and g__4973(w__5891 ,w__5793 ,w__5890);
  or g__4974(w__5890 ,w__5812 ,w__5889);
  xnor g__4975(w__8386 ,w__5888 ,w__5823);
  and g__4976(w__5889 ,w__5801 ,w__5888);
  or g__4977(w__5888 ,w__5826 ,w__5887);
  xnor g__4978(w__8385 ,w__5886 ,w__5840);
  and g__4979(w__5887 ,w__5835 ,w__5886);
  or g__4980(w__5886 ,w__5858 ,w__5885);
  xnor g__4981(w__8384 ,w__5884 ,w__5864);
  nor g__4982(w__5885 ,w__5859 ,w__5884);
  and g__4983(w__5884 ,w__5883 ,w__5860);
  or g__4984(w__5883 ,w__5852 ,w__5882);
  and g__4985(w__5882 ,w__5868 ,w__5881);
  or g__4986(w__5881 ,w__5867 ,w__5880);
  and g__4987(w__5880 ,w__5879 ,w__5869);
  or g__4988(w__5879 ,w__5866 ,w__5878);
  and g__4989(w__5878 ,w__5857 ,w__5877);
  or g__4990(w__5877 ,w__5856 ,w__5876);
  and g__4991(w__5876 ,w__5845 ,w__5875);
  or g__4992(w__5875 ,w__5846 ,w__5874);
  and g__4993(w__5874 ,w__5830 ,w__5873);
  xnor g__4994(w__8378 ,w__5872 ,w__5839);
  or g__4995(w__5873 ,w__5824 ,w__5872);
  and g__4996(w__5872 ,w__5802 ,w__5865);
  xnor g__4997(w__5871 ,w__5853 ,w__5848);
  xnor g__4998(w__5870 ,w__5854 ,w__5861);
  or g__4999(w__5869 ,w__5848 ,w__5853);
  or g__5000(w__5868 ,w__5861 ,w__5854);
  and g__5001(w__5867 ,w__5861 ,w__5854);
  and g__5002(w__5866 ,w__5848 ,w__5853);
  or g__5003(w__5865 ,w__5803 ,w__5855);
  xnor g__5004(w__5864 ,w__5850 ,w__5828);
  xnor g__5005(w__5863 ,w__5844 ,w__5849);
  xnor g__5006(w__5862 ,w__5837 ,w__5843);
  or g__5007(w__5860 ,w__5849 ,w__5844);
  and g__5008(w__5859 ,w__5850 ,w__5829);
  nor g__5009(w__5858 ,w__5850 ,w__5829);
  or g__5010(w__5857 ,w__5836 ,w__5842);
  nor g__5011(w__5856 ,w__5837 ,w__5843);
  and g__5012(w__5861 ,w__5834 ,w__5847);
  and g__5013(w__5852 ,w__5849 ,w__5844);
  xnor g__5014(w__8376 ,w__5838 ,w__5799);
  xnor g__5015(w__5851 ,w__5827 ,w__5818);
  and g__5016(w__5855 ,w__5773 ,w__5841);
  xnor g__5017(w__5854 ,w__5780 ,w__5821);
  xnor g__5018(w__5853 ,w__5817 ,w__5822);
  or g__5019(w__5847 ,w__5782 ,w__5833);
  and g__5020(w__5846 ,w__5818 ,w__5827);
  or g__5021(w__5845 ,w__5818 ,w__5827);
  and g__5022(w__5850 ,w__5788 ,w__5831);
  and g__5023(w__5849 ,w__5814 ,w__5825);
  and g__5024(w__5848 ,w__5813 ,w__5832);
  not g__5025(w__5842 ,w__5843);
  or g__5026(w__5841 ,w__5787 ,w__5838);
  xnor g__5027(w__8375 ,w__5779 ,w__5797);
  xnor g__5028(w__5840 ,w__5805 ,w__5807);
  xnor g__5029(w__5839 ,w__5776 ,w__5808);
  xnor g__5030(w__5844 ,w__5819 ,w__5800);
  xnor g__5031(w__5843 ,w__5775 ,w__5796);
  not g__5032(w__5836 ,w__5837);
  or g__5033(w__5835 ,w__5806 ,w__5804);
  or g__5034(w__5834 ,w__5748 ,w__5817);
  and g__5035(w__5833 ,w__5748 ,w__5817);
  or g__5036(w__5832 ,w__5770 ,w__5811);
  or g__5037(w__5831 ,w__5819 ,w__5785);
  or g__5038(w__5830 ,w__5776 ,w__5809);
  and g__5039(w__5838 ,w__5792 ,w__5816);
  or g__5040(w__5837 ,w__5761 ,w__5810);
  not g__5041(w__5829 ,w__5828);
  nor g__5042(w__5826 ,w__5807 ,w__5805);
  or g__5043(w__5825 ,w__5780 ,w__5815);
  and g__5044(w__5824 ,w__5776 ,w__5809);
  xnor g__5045(w__5823 ,w__5795 ,w__5749);
  xnor g__5046(w__5822 ,w__5782 ,w__5748);
  xnor g__5047(w__5821 ,w__5778 ,w__5722);
  xnor g__5048(w__5820 ,w__5777 ,w__5768);
  xnor g__5049(w__5828 ,w__5769 ,w__5771);
  xnor g__5050(w__5827 ,w__5781 ,w__5772);
  or g__5051(w__5816 ,w__5791 ,w__5779);
  and g__5052(w__5815 ,w__5722 ,w__5778);
  or g__5053(w__5814 ,w__5722 ,w__5778);
  or g__5054(w__5813 ,w__5706 ,w__5774);
  nor g__5055(w__5812 ,w__5054 ,w__5795);
  nor g__5056(w__5811 ,w__5705 ,w__5775);
  and g__5057(w__5810 ,w__5758 ,w__5781);
  and g__5058(w__5819 ,w__5759 ,w__5784);
  and g__5059(w__5818 ,w__5730 ,w__5783);
  and g__5060(w__5817 ,w__5764 ,w__5789);
  not g__5061(w__5809 ,w__5808);
  not g__5062(w__5807 ,w__5806);
  not g__5063(w__5804 ,w__5805);
  and g__5064(w__5803 ,w__5768 ,w__5777);
  or g__5065(w__5802 ,w__5768 ,w__5777);
  or g__5066(w__5801 ,w__5056 ,w__5794);
  xnor g__5067(w__5800 ,w__5756 ,w__5737);
  xnor g__5068(w__5799 ,w__5721 ,w__5755);
  xnor g__5069(w__5798 ,w__5751 ,w__5690);
  xnor g__5070(w__5797 ,w__5616 ,w__5753);
  xnor g__5071(w__5796 ,w__5770 ,w__5706);
  xnor g__5072(w__5808 ,w__5757 ,w__5743);
  xnor g__5073(w__5806 ,w__5740 ,w__5744);
  and g__5074(w__5805 ,w__5746 ,w__5790);
  not g__5075(w__5795 ,w__5794);
  or g__5076(w__5793 ,w__5689 ,w__5750);
  or g__5077(w__5792 ,w__5615 ,w__5753);
  nor g__5078(w__5791 ,w__5616 ,w__5752);
  or g__5079(w__5790 ,w__5766 ,w__5769);
  or g__5080(w__5789 ,w__5630 ,w__5763);
  or g__5081(w__5788 ,w__5737 ,w__5756);
  nor g__5082(w__5787 ,w__5720 ,w__5755);
  nor g__5083(w__5786 ,w__5690 ,w__5751);
  and g__5084(w__5785 ,w__5737 ,w__5756);
  or g__5085(w__5784 ,w__5623 ,w__5762);
  or g__5086(w__5783 ,w__5734 ,w__5757);
  or g__5087(w__5794 ,w__5731 ,w__5760);
  not g__5088(w__5774 ,w__5775);
  xnor g__5089(w__8374 ,w__5741 ,w__5714);
  or g__5090(w__5773 ,w__5721 ,w__5754);
  xnor g__5091(w__5772 ,w__5688 ,w__5739);
  xnor g__5092(w__5771 ,w__5672 ,w__5727);
  xnor g__5093(w__5782 ,w__5742 ,w__5712);
  xnor g__5094(w__5781 ,w__5619 ,w__5715);
  and g__5095(w__5780 ,w__5684 ,w__5767);
  and g__5096(w__5779 ,w__5703 ,w__5747);
  xnor g__5097(w__5778 ,w__5725 ,w__5717);
  xnor g__5098(w__5777 ,w__5728 ,w__5716);
  and g__5099(w__5776 ,w__5699 ,w__5765);
  xnor g__5100(w__5775 ,w__5724 ,w__5713);
  or g__5101(w__5767 ,w__5704 ,w__5742);
  nor g__5102(w__5766 ,w__5671 ,w__5727);
  or g__5103(w__5765 ,w__5682 ,w__5728);
  or g__5104(w__5764 ,w__5652 ,w__5723);
  nor g__5105(w__5763 ,w__5651 ,w__5724);
  and g__5106(w__5762 ,w__5647 ,w__5725);
  nor g__5107(w__5761 ,w__5687 ,w__5739);
  nor g__5108(w__5760 ,w__5729 ,w__5740);
  or g__5109(w__5759 ,w__5647 ,w__5725);
  or g__5110(w__5758 ,w__5688 ,w__5738);
  and g__5111(w__5770 ,w__5695 ,w__5733);
  and g__5112(w__5769 ,w__5698 ,w__5732);
  and g__5113(w__5768 ,w__5686 ,w__5719);
  not g__5114(w__5754 ,w__5755);
  not g__5115(w__5752 ,w__5753);
  not g__5116(w__5750 ,w__5751);
  or g__5117(w__5747 ,w__5702 ,w__5741);
  or g__5118(w__5746 ,w__5672 ,w__5726);
  xnor g__5119(w__8373 ,w__5653 ,w__5678);
  xnor g__5120(w__5745 ,w__5710 ,w__5603);
  xnor g__5121(w__5744 ,w__5567 ,w__5691);
  xnor g__5122(w__5743 ,w__5708 ,w__5646);
  xnor g__5123(w__5757 ,w__5624 ,w__5676);
  xnor g__5124(w__5756 ,w__5650 ,w__5674);
  xnor g__5125(w__5755 ,w__5641 ,w__5677);
  xnor g__5126(w__5753 ,w__5551 ,w__5673);
  and g__5127(w__5751 ,w__5656 ,w__5718);
  xnor g__5128(w__5749 ,w__5711 ,w__5675);
  xnor g__5129(w__5748 ,w__5599 ,w__5679);
  not g__5130(w__5738 ,w__5739);
  or g__5131(w__5736 ,w__5055 ,w__5709);
  nor g__5132(w__5735 ,w__5053 ,w__5710);
  nor g__5133(w__5734 ,w__5707 ,w__5646);
  or g__5134(w__5733 ,w__5625 ,w__5693);
  or g__5135(w__5732 ,w__5629 ,w__5696);
  nor g__5136(w__5731 ,w__5568 ,w__5691);
  or g__5137(w__5730 ,w__5708 ,w__5645);
  and g__5138(w__5729 ,w__5568 ,w__5691);
  and g__5139(w__5742 ,w__5669 ,w__5700);
  and g__5140(w__5741 ,w__5668 ,w__5701);
  and g__5141(w__5740 ,w__5655 ,w__5697);
  and g__5142(w__5739 ,w__5659 ,w__5692);
  and g__5143(w__5737 ,w__5670 ,w__5694);
  not g__5144(w__5727 ,w__5726);
  not g__5145(w__5723 ,w__5724);
  not g__5146(w__5720 ,w__5721);
  or g__5147(w__5719 ,w__5622 ,w__5685);
  or g__5148(w__5718 ,w__5711 ,w__5660);
  xnor g__5149(w__5717 ,w__5647 ,w__5623);
  xnor g__5150(w__5716 ,w__5644 ,w__5617);
  xnor g__5151(w__5715 ,w__5649 ,w__5625);
  xnor g__5152(w__5714 ,w__5588 ,w__5643);
  xnor g__5153(w__5713 ,w__5652 ,w__5630);
  xnor g__5154(w__5712 ,w__5640 ,w__5610);
  xnor g__5155(w__5728 ,w__5570 ,w__5634);
  xnor g__5156(w__5726 ,w__5600 ,w__5631);
  xnor g__5157(w__5725 ,w__5604 ,w__5633);
  xnor g__5158(w__5724 ,w__5609 ,w__5632);
  and g__5159(w__5722 ,w__5661 ,w__5681);
  and g__5160(w__5721 ,w__5635 ,w__5683);
  not g__5161(w__5709 ,w__5710);
  not g__5162(w__5707 ,w__5708);
  not g__5163(w__5705 ,w__5706);
  and g__5164(w__5704 ,w__5610 ,w__5640);
  or g__5165(w__5703 ,w__5588 ,w__5642);
  nor g__5166(w__5702 ,w__5587 ,w__5643);
  or g__5167(w__5701 ,w__5667 ,w__5653);
  or g__5168(w__5700 ,w__5592 ,w__5666);
  or g__5169(w__5699 ,w__5617 ,w__5644);
  or g__5170(w__5698 ,w__5601 ,w__5650);
  or g__5171(w__5697 ,w__5571 ,w__5637);
  and g__5172(w__5696 ,w__5601 ,w__5650);
  or g__5173(w__5695 ,w__5618 ,w__5649);
  or g__5174(w__5694 ,w__5591 ,w__5658);
  nor g__5175(w__5693 ,w__5619 ,w__5648);
  or g__5176(w__5692 ,w__5624 ,w__5657);
  and g__5177(w__5711 ,w__5586 ,w__5665);
  and g__5178(w__5710 ,w__5582 ,w__5639);
  and g__5179(w__5708 ,w__5612 ,w__5654);
  and g__5180(w__5706 ,w__5534 ,w__5664);
  not g__5181(w__5690 ,w__5689);
  not g__5182(w__5688 ,w__5687);
  xnor g__5183(w__8372 ,w__5590 ,w__5595);
  or g__5184(w__5686 ,w__5606 ,w__5641);
  and g__5185(w__5685 ,w__5606 ,w__5641);
  or g__5186(w__5684 ,w__5610 ,w__5640);
  or g__5187(w__5683 ,w__5551 ,w__5636);
  and g__5188(w__5682 ,w__5617 ,w__5644);
  or g__5189(w__5681 ,w__5628 ,w__5638);
  xnor g__5190(w__5680 ,w__5621 ,w__5376);
  xnor g__5191(w__5679 ,w__5628 ,w__5484);
  xnor g__5192(w__5678 ,w__5483 ,w__5608);
  xnor g__5193(w__5677 ,w__5622 ,w__5605);
  xnor g__5194(w__5676 ,w__5602 ,w__5547);
  xnor g__5195(w__5675 ,w__5598 ,w__5548);
  xnor g__5196(w__5674 ,w__5601 ,w__5629);
  xnor g__5197(w__5673 ,w__5597 ,w__5429);
  xnor g__5198(w__5691 ,w__5627 ,w__5593);
  xnor g__5199(w__5689 ,w__5626 ,w__5594);
  xnor g__5200(w__5687 ,w__5611 ,w__5561);
  not g__5201(w__5671 ,w__5672);
  or g__5202(w__5670 ,w__5417 ,w__5604);
  or g__5203(w__5669 ,w__5515 ,w__5609);
  or g__5204(w__5668 ,w__5482 ,w__5608);
  nor g__5205(w__5667 ,w__5483 ,w__5607);
  and g__5206(w__5666 ,w__5515 ,w__5609);
  or g__5207(w__5665 ,w__5575 ,w__5627);
  or g__5208(w__5664 ,w__5533 ,w__5611);
  nor g__5209(w__5663 ,w__5376 ,w__5621);
  or g__5210(w__5662 ,w__5375 ,w__5620);
  or g__5211(w__5661 ,w__5484 ,w__5599);
  and g__5212(w__5660 ,w__5548 ,w__5598);
  or g__5213(w__5659 ,w__5547 ,w__5602);
  and g__5214(w__5658 ,w__5417 ,w__5604);
  and g__5215(w__5657 ,w__5547 ,w__5602);
  or g__5216(w__5656 ,w__5548 ,w__5598);
  or g__5217(w__5655 ,w__5514 ,w__5600);
  or g__5218(w__5654 ,w__5570 ,w__5613);
  and g__5219(w__5672 ,w__5546 ,w__5614);
  not g__5220(w__5651 ,w__5652);
  not g__5221(w__5648 ,w__5649);
  not g__5222(w__5645 ,w__5646);
  not g__5223(w__5642 ,w__5643);
  or g__5224(w__5639 ,w__5583 ,w__5626);
  and g__5225(w__5638 ,w__5484 ,w__5599);
  and g__5226(w__5637 ,w__5514 ,w__5600);
  and g__5227(w__5636 ,w__5429 ,w__5597);
  or g__5228(w__5635 ,w__5429 ,w__5597);
  xnor g__5229(w__5634 ,w__5569 ,w__5411);
  xnor g__5230(w__5633 ,w__5591 ,w__5417);
  xor g__5231(w__5632 ,w__5592 ,w__5515);
  xnor g__5232(w__5631 ,w__5571 ,w__5514);
  and g__5233(w__5653 ,w__5579 ,w__5596);
  xnor g__5234(w__5652 ,w__5440 ,w__5556);
  xnor g__5235(w__5650 ,w__5589 ,w__5558);
  xnor g__5236(w__5649 ,w__5430 ,w__5557);
  xnor g__5237(w__5647 ,w__5442 ,w__5555);
  xnor g__5238(w__5646 ,w__5518 ,w__5553);
  xnor g__5239(w__5644 ,w__5448 ,w__5552);
  xnor g__5240(w__5643 ,w__5520 ,w__5559);
  xnor g__5241(w__5641 ,w__5487 ,w__5554);
  xnor g__5242(w__5640 ,w__5446 ,w__5560);
  not g__5243(w__5620 ,w__5621);
  not g__5244(w__5619 ,w__5618);
  not g__5245(w__5616 ,w__5615);
  or g__5246(w__5614 ,w__5589 ,w__5538);
  and g__5247(w__5613 ,w__5411 ,w__5569);
  or g__5248(w__5612 ,w__5411 ,w__5569);
  and g__5249(w__5630 ,w__5536 ,w__5574);
  and g__5250(w__5629 ,w__5535 ,w__5572);
  and g__5251(w__5628 ,w__5504 ,w__5562);
  and g__5252(w__5627 ,w__5537 ,w__5573);
  and g__5253(w__5626 ,w__5526 ,w__5576);
  and g__5254(w__5625 ,w__5527 ,w__5581);
  and g__5255(w__5624 ,w__5522 ,w__5566);
  and g__5256(w__5623 ,w__5510 ,w__5565);
  and g__5257(w__5622 ,w__5503 ,w__5564);
  and g__5258(w__5621 ,w__5467 ,w__5578);
  and g__5259(w__5618 ,w__5531 ,w__5580);
  and g__5260(w__5617 ,w__5507 ,w__5563);
  and g__5261(w__5615 ,w__5545 ,w__5584);
  not g__5262(w__5607 ,w__5608);
  not g__5263(w__5606 ,w__5605);
  or g__5264(w__5596 ,w__5590 ,w__5577);
  xnor g__5265(w__5595 ,w__5444 ,w__5513);
  xnor g__5266(w__5594 ,w__5374 ,w__5517);
  xnor g__5267(w__5593 ,w__5549 ,w__5439);
  xnor g__5268(w__5611 ,w__5420 ,w__5491);
  and g__5269(w__5610 ,w__5500 ,w__5585);
  xnor g__5270(w__5609 ,w__5447 ,w__5496);
  xnor g__5271(w__5608 ,w__5455 ,w__5495);
  xnor g__5272(w__5605 ,w__5457 ,w__5497);
  xnor g__5273(w__5604 ,w__5424 ,w__5499);
  xnor g__5274(w__5603 ,w__5550 ,w__5489);
  xnor g__5275(w__5602 ,w__5449 ,w__5488);
  xnor g__5276(w__5601 ,w__5377 ,w__5494);
  xnor g__5277(w__5600 ,w__5434 ,w__5490);
  xnor g__5278(w__5599 ,w__5421 ,w__5492);
  xnor g__5279(w__5598 ,w__5431 ,w__5493);
  xnor g__5280(w__5597 ,w__5432 ,w__5498);
  not g__5281(w__5587 ,w__5588);
  or g__5282(w__5586 ,w__5439 ,w__5549);
  or g__5283(w__5585 ,w__5427 ,w__5543);
  or g__5284(w__5584 ,w__5544 ,w__5521);
  nor g__5285(w__5583 ,w__5374 ,w__5516);
  or g__5286(w__5582 ,w__5373 ,w__5517);
  or g__5287(w__5581 ,w__5418 ,w__5525);
  or g__5288(w__5580 ,w__5519 ,w__5529);
  or g__5289(w__5579 ,w__5444 ,w__5512);
  or g__5290(w__5578 ,w__5470 ,w__5550);
  nor g__5291(w__5577 ,w__5443 ,w__5513);
  or g__5292(w__5576 ,w__5425 ,w__5528);
  and g__5293(w__5575 ,w__5439 ,w__5549);
  or g__5294(w__5574 ,w__5426 ,w__5511);
  or g__5295(w__5573 ,w__5422 ,w__5530);
  or g__5296(w__5572 ,w__5423 ,w__5532);
  and g__5297(w__5592 ,w__5476 ,w__5541);
  and g__5298(w__5591 ,w__5471 ,w__5524);
  and g__5299(w__5590 ,w__5407 ,w__5540);
  and g__5300(w__5589 ,w__5477 ,w__5539);
  and g__5301(w__5588 ,w__5478 ,w__5542);
  not g__5302(w__5568 ,w__5567);
  or g__5303(w__5566 ,w__5456 ,w__5523);
  xnor g__5304(w__8371 ,w__5485 ,w__5458);
  or g__5305(w__5565 ,w__5454 ,w__5508);
  or g__5306(w__5564 ,w__5402 ,w__5502);
  or g__5307(w__5563 ,w__5487 ,w__5505);
  or g__5308(w__5562 ,w__5403 ,w__5501);
  xnor g__5309(w__5561 ,w__5452 ,w__5479);
  xnor g__5310(w__5560 ,w__5454 ,w__5445);
  xnor g__5311(w__5559 ,w__5481 ,w__5435);
  xnor g__5312(w__5558 ,w__5436 ,w__5480);
  xnor g__5313(w__5557 ,w__5441 ,w__5426);
  xnor g__5314(w__5556 ,w__5433 ,w__5403);
  xnor g__5315(w__5555 ,w__5453 ,w__5423);
  xnor g__5316(w__5554 ,w__5437 ,w__5438);
  xnor g__5317(w__5553 ,w__5450 ,w__5451);
  xnor g__5318(w__5552 ,w__5456 ,w__5414);
  and g__5319(w__5571 ,w__5463 ,w__5506);
  and g__5320(w__5570 ,w__5466 ,w__5509);
  xnor g__5321(w__5569 ,w__5419 ,w__5428);
  xnor g__5322(w__5567 ,w__5401 ,w__5459);
  or g__5323(w__5546 ,w__5480 ,w__5436);
  or g__5324(w__5545 ,w__5435 ,w__5481);
  and g__5325(w__5544 ,w__5435 ,w__5481);
  and g__5326(w__5543 ,w__5394 ,w__5447);
  or g__5327(w__5542 ,w__5473 ,w__5455);
  or g__5328(w__5541 ,w__5420 ,w__5474);
  or g__5329(w__5540 ,w__5384 ,w__5486);
  or g__5330(w__5539 ,w__5424 ,w__5472);
  and g__5331(w__5538 ,w__5480 ,w__5436);
  or g__5332(w__5537 ,w__5412 ,w__5434);
  or g__5333(w__5536 ,w__5430 ,w__5441);
  or g__5334(w__5535 ,w__5442 ,w__5453);
  or g__5335(w__5534 ,w__5479 ,w__5452);
  and g__5336(w__5533 ,w__5479 ,w__5452);
  and g__5337(w__5532 ,w__5442 ,w__5453);
  or g__5338(w__5531 ,w__5451 ,w__5450);
  and g__5339(w__5530 ,w__5412 ,w__5434);
  and g__5340(w__5529 ,w__5451 ,w__5450);
  and g__5341(w__5528 ,w__5390 ,w__5431);
  or g__5342(w__5527 ,w__5415 ,w__5449);
  or g__5343(w__5526 ,w__5390 ,w__5431);
  and g__5344(w__5525 ,w__5415 ,w__5449);
  or g__5345(w__5524 ,w__5421 ,w__5468);
  and g__5346(w__5523 ,w__5414 ,w__5448);
  or g__5347(w__5522 ,w__5414 ,w__5448);
  and g__5348(w__5551 ,w__5335 ,w__5462);
  and g__5349(w__5550 ,w__5225 ,w__5461);
  and g__5350(w__5549 ,w__5234 ,w__5475);
  and g__5351(w__5548 ,w__5385 ,w__5465);
  and g__5352(w__5547 ,w__5406 ,w__5469);
  not g__5353(w__5521 ,w__5520);
  not g__5354(w__5519 ,w__5518);
  not g__5355(w__5516 ,w__5517);
  not g__5356(w__5512 ,w__5513);
  and g__5357(w__5511 ,w__5430 ,w__5441);
  or g__5358(w__5510 ,w__5445 ,w__5446);
  or g__5359(w__5509 ,w__5464 ,w__5457);
  and g__5360(w__5508 ,w__5445 ,w__5446);
  or g__5361(w__5507 ,w__5438 ,w__5437);
  or g__5362(w__5506 ,w__5377 ,w__5460);
  and g__5363(w__5505 ,w__5438 ,w__5437);
  or g__5364(w__5504 ,w__5440 ,w__5433);
  or g__5365(w__5503 ,w__5393 ,w__5432);
  and g__5366(w__5502 ,w__5393 ,w__5432);
  and g__5367(w__5501 ,w__5440 ,w__5433);
  or g__5368(w__5500 ,w__5394 ,w__5447);
  xnor g__5369(w__5499 ,w__5169 ,w__5392);
  xnor g__5370(w__5498 ,w__5402 ,w__5393);
  xnor g__5371(w__5497 ,w__5298 ,w__5388);
  xnor g__5372(w__5496 ,w__5394 ,w__5427);
  xnor g__5373(w__5495 ,w__5410 ,w__4835);
  xnor g__5374(w__5494 ,w__5391 ,w__5395);
  xnor g__5375(w__5493 ,w__5390 ,w__5425);
  xnor g__5376(w__5492 ,w__5416 ,w__5413);
  xnor g__5377(w__5491 ,w__5386 ,w__4836);
  xnor g__5378(w__5490 ,w__5422 ,w__5412);
  xnor g__5379(w__5489 ,w__5083 ,w__5389);
  xnor g__5380(w__5488 ,w__5415 ,w__5418);
  xnor g__5381(w__5520 ,w__5399 ,w__5378);
  xnor g__5382(w__5518 ,w__5299 ,w__5379);
  xnor g__5383(w__5517 ,w__5400 ,w__5310);
  xor g__5384(w__5515 ,w__5253 ,w__5381);
  xnor g__5385(w__5514 ,w__5396 ,w__5302);
  xnor g__5386(w__5513 ,w__5252 ,w__5380);
  not g__5387(w__5486 ,w__5485);
  not g__5388(w__5482 ,w__5483);
  or g__5389(w__5478 ,w__4835 ,w__5410);
  or g__5390(w__5477 ,w__5169 ,w__5392);
  or g__5391(w__5476 ,w__4836 ,w__5386);
  or g__5392(w__5475 ,w__5271 ,w__5396);
  and g__5393(w__5474 ,w__4836 ,w__5386);
  and g__5394(w__5473 ,w__4835 ,w__5410);
  and g__5395(w__5472 ,w__5169 ,w__5392);
  or g__5396(w__5471 ,w__5413 ,w__5416);
  and g__5397(w__5470 ,w__5083 ,w__5389);
  or g__5398(w__5469 ,w__5419 ,w__5404);
  and g__5399(w__5468 ,w__5413 ,w__5416);
  or g__5400(w__5467 ,w__5083 ,w__5389);
  or g__5401(w__5466 ,w__5297 ,w__5388);
  or g__5402(w__5465 ,w__5382 ,w__5401);
  nor g__5403(w__5464 ,w__5298 ,w__5387);
  or g__5404(w__5463 ,w__5395 ,w__5391);
  or g__5405(w__5462 ,w__5367 ,w__5399);
  or g__5406(w__5461 ,w__5259 ,w__5400);
  and g__5407(w__5460 ,w__5395 ,w__5391);
  xnor g__5408(w__5459 ,w__5085 ,w__5371);
  xnor g__5409(w__5458 ,w__4834 ,w__5372);
  and g__5410(w__5487 ,w__5227 ,w__5383);
  and g__5411(w__5485 ,w__5140 ,w__5398);
  and g__5412(w__5484 ,w__5358 ,w__5409);
  or g__5413(w__5483 ,w__5364 ,w__5408);
  xnor g__5414(w__5481 ,w__5155 ,w__5330);
  xnor g__5415(w__5480 ,w__5210 ,w__5324);
  and g__5416(w__5479 ,w__5356 ,w__5405);
  not g__5417(w__5443 ,w__5444);
  xnor g__5418(w__5428 ,w__5107 ,w__4837);
  xnor g__5419(w__5457 ,w__5187 ,w__5301);
  xnor g__5420(w__5456 ,w__5128 ,w__5305);
  xnor g__5421(w__5455 ,w__5197 ,w__5303);
  xnor g__5422(w__5454 ,w__5192 ,w__5314);
  xnor g__5423(w__5453 ,w__5165 ,w__5316);
  xnor g__5424(w__5452 ,w__5130 ,w__5315);
  xnor g__5425(w__5451 ,w__5198 ,w__5313);
  xnor g__5426(w__5450 ,w__5193 ,w__5311);
  xnor g__5427(w__5449 ,w__5188 ,w__5307);
  xnor g__5428(w__5448 ,w__5174 ,w__5332);
  xnor g__5429(w__5447 ,w__5201 ,w__5322);
  xnor g__5430(w__5446 ,w__5114 ,w__5319);
  xnor g__5431(w__5445 ,w__5129 ,w__5323);
  xnor g__5432(w__5444 ,w__5088 ,w__5327);
  xnor g__5433(w__5442 ,w__5094 ,w__5318);
  xnor g__5434(w__5441 ,w__5117 ,w__5320);
  xnor g__5435(w__5440 ,w__5133 ,w__5304);
  xnor g__5436(w__5439 ,w__5134 ,w__5325);
  xnor g__5437(w__5438 ,w__5127 ,w__5309);
  xnor g__5438(w__5437 ,w__5255 ,w__5328);
  xnor g__5439(w__5436 ,w__5186 ,w__5329);
  xnor g__5440(w__5435 ,w__5209 ,w__5312);
  xnor g__5441(w__5434 ,w__5200 ,w__5317);
  xnor g__5442(w__5433 ,w__5196 ,w__5306);
  xnor g__5443(w__5432 ,w__5087 ,w__5321);
  xnor g__5444(w__5431 ,w__5131 ,w__5308);
  xnor g__5445(w__5430 ,w__5199 ,w__5331);
  xnor g__5446(w__5429 ,w__4833 ,w__5326);
  or g__5447(w__5409 ,w__5254 ,w__5336);
  and g__5448(w__5408 ,w__5252 ,w__5333);
  or g__5449(w__5407 ,w__5372 ,w__4834);
  or g__5450(w__5406 ,w__5107 ,w__4837);
  or g__5451(w__5405 ,w__5300 ,w__5355);
  and g__5452(w__5404 ,w__5107 ,w__4837);
  and g__5453(w__5427 ,w__5281 ,w__5368);
  and g__5454(w__5426 ,w__5220 ,w__5359);
  and g__5455(w__5425 ,w__5277 ,w__5351);
  and g__5456(w__5424 ,w__5292 ,w__5357);
  and g__5457(w__5423 ,w__5222 ,w__5354);
  and g__5458(w__5422 ,w__5231 ,w__5369);
  and g__5459(w__5421 ,w__5279 ,w__5343);
  and g__5460(w__5420 ,w__5282 ,w__5363);
  and g__5461(w__5419 ,w__5240 ,w__5342);
  and g__5462(w__5418 ,w__5260 ,w__5345);
  and g__5463(w__5417 ,w__5265 ,w__5350);
  and g__5464(w__5416 ,w__5257 ,w__5344);
  and g__5465(w__5415 ,w__5272 ,w__5347);
  and g__5466(w__5414 ,w__5288 ,w__5341);
  and g__5467(w__5413 ,w__5261 ,w__5346);
  and g__5468(w__5412 ,w__5217 ,w__5337);
  and g__5469(w__5411 ,w__5241 ,w__5340);
  and g__5470(w__5410 ,w__5232 ,w__5366);
  not g__5471(w__5398 ,w__5397);
  not g__5472(w__5387 ,w__5388);
  or g__5473(w__5385 ,w__5085 ,w__5370);
  and g__5474(w__5384 ,w__5372 ,w__4834);
  or g__5475(w__5383 ,w__5287 ,w__4833);
  nor g__5476(w__5382 ,w__5084 ,w__5371);
  xnor g__5477(w__5381 ,w__5176 ,w__5251);
  xnor g__5478(w__5380 ,w__5096 ,w__5247);
  xnor g__5479(w__5379 ,w__5115 ,w__5248);
  xnor g__5480(w__5378 ,w__5296 ,w__5250);
  and g__5481(w__5403 ,w__5283 ,w__5362);
  and g__5482(w__5402 ,w__5218 ,w__5348);
  and g__5483(w__5401 ,w__5245 ,w__5339);
  and g__5484(w__5400 ,w__5278 ,w__5360);
  and g__5485(w__5399 ,w__5223 ,w__5334);
  xnor g__5486(w__5397 ,w__5185 ,w__5211);
  xnor g__5487(w__5396 ,w__5202 ,w__5215);
  and g__5488(w__5395 ,w__5238 ,w__5349);
  and g__5489(w__5394 ,w__5216 ,w__5352);
  and g__5490(w__5393 ,w__5275 ,w__5361);
  xnor g__5491(w__5392 ,w__5123 ,w__5214);
  and g__5492(w__5391 ,w__5262 ,w__5353);
  xnor g__5493(w__5390 ,w__5132 ,w__5213);
  xnor g__5494(w__5389 ,w__5135 ,w__5212);
  and g__5495(w__5388 ,w__5237 ,w__5365);
  and g__5496(w__5386 ,w__5236 ,w__5338);
  not g__5497(w__5376 ,w__5375);
  not g__5498(w__5373 ,w__5374);
  not g__5499(w__5370 ,w__5371);
  or g__5500(w__5369 ,w__5186 ,w__5224);
  or g__5501(w__5368 ,w__5137 ,w__5280);
  nor g__5502(w__5367 ,w__5296 ,w__5249);
  or g__5503(w__5366 ,w__5125 ,w__5244);
  or g__5504(w__5365 ,w__5126 ,w__5270);
  nor g__5505(w__5364 ,w__5096 ,w__5247);
  or g__5506(w__5363 ,w__5193 ,w__5285);
  or g__5507(w__5362 ,w__5130 ,w__5274);
  or g__5508(w__5361 ,w__5209 ,w__5219);
  or g__5509(w__5360 ,w__5131 ,w__5291);
  or g__5510(w__5359 ,w__5188 ,w__5267);
  or g__5511(w__5358 ,w__5176 ,w__5251);
  or g__5512(w__5357 ,w__5129 ,w__5276);
  or g__5513(w__5356 ,w__5115 ,w__5248);
  and g__5514(w__5355 ,w__5115 ,w__5248);
  or g__5515(w__5354 ,w__5138 ,w__5266);
  or g__5516(w__5353 ,w__5124 ,w__5294);
  or g__5517(w__5352 ,w__5199 ,w__5269);
  or g__5518(w__5351 ,w__5134 ,w__5290);
  or g__5519(w__5350 ,w__5192 ,w__5273);
  or g__5520(w__5349 ,w__5191 ,w__5226);
  or g__5521(w__5348 ,w__5139 ,w__5239);
  or g__5522(w__5347 ,w__5128 ,w__5284);
  or g__5523(w__5346 ,w__5133 ,w__5221);
  or g__5524(w__5345 ,w__5142 ,w__5233);
  or g__5525(w__5344 ,w__5196 ,w__5229);
  or g__5526(w__5343 ,w__5201 ,w__5263);
  or g__5527(w__5342 ,w__5187 ,w__5268);
  or g__5528(w__5341 ,w__5127 ,w__5286);
  or g__5529(w__5340 ,w__5289 ,w__5255);
  or g__5530(w__5339 ,w__5200 ,w__5258);
  or g__5531(w__5338 ,w__5198 ,w__5243);
  or g__5532(w__5337 ,w__5210 ,w__5256);
  and g__5533(w__5336 ,w__5176 ,w__5251);
  and g__5534(w__5377 ,w__5080 ,w__5228);
  or g__5535(w__5375 ,w__5081 ,w__5242);
  or g__5536(w__5374 ,w__5143 ,w__5230);
  and g__5537(w__5372 ,w__5148 ,w__5264);
  or g__5538(w__5371 ,w__5082 ,w__5235);
  or g__5539(w__5335 ,w__5250 ,w__5295);
  or g__5540(w__5334 ,w__5197 ,w__5293);
  or g__5541(w__5333 ,w__5095 ,w__5246);
  xnor g__5542(w__5332 ,w__5106 ,w__5142);
  xnor g__5543(w__5331 ,w__5101 ,w__5111);
  xnor g__5544(w__5330 ,w__5166 ,w__5139);
  xnor g__5545(w__5329 ,w__5158 ,w__5099);
  xnor g__5546(w__5328 ,w__5152 ,w__5116);
  xnor g__5547(w__5327 ,w__5109 ,w__5125);
  xnor g__5548(w__5326 ,w__5160 ,w__5170);
  xnor g__5549(w__5325 ,w__5108 ,w__5092);
  xnor g__5550(w__5324 ,w__5171 ,w__5157);
  xnor g__5551(w__5323 ,w__5154 ,w__5168);
  xnor g__5552(w__5322 ,w__5105 ,w__5113);
  xnor g__5553(w__5321 ,w__5161 ,w__5126);
  xnor g__5554(w__5320 ,w__5149 ,w__5137);
  xnor g__5555(w__5319 ,w__5151 ,w__5138);
  xnor g__5556(w__5318 ,w__5178 ,w__5124);
  xnor g__5557(w__5317 ,w__5093 ,w__5167);
  xnor g__5558(w__5316 ,w__5184 ,w__5191);
  xnor g__5559(w__5315 ,w__5097 ,w__5164);
  xnor g__5560(w__5314 ,w__5100 ,w__5103);
  xnor g__5561(w__5313 ,w__5110 ,w__5175);
  xnor g__5562(w__5312 ,w__5090 ,w__5159);
  xnor g__5563(w__5311 ,w__5102 ,w__5091);
  xnor g__5564(w__5310 ,w__5098 ,w__5162);
  xnor g__5565(w__5309 ,w__5153 ,w__5183);
  xnor g__5566(w__5308 ,w__5104 ,w__5179);
  xnor g__5567(w__5307 ,w__5181 ,w__5089);
  xnor g__5568(w__5306 ,w__5112 ,w__5163);
  xnor g__5569(w__5305 ,w__5156 ,w__5180);
  xnor g__5570(w__5304 ,w__5086 ,w__5150);
  xnor g__5571(w__5303 ,w__5172 ,w__5119);
  xnor g__5572(w__5302 ,w__5177 ,w__5118);
  xnor g__5573(w__5301 ,w__5182 ,w__5173);
  not g__5574(w__5300 ,w__5299);
  not g__5575(w__5297 ,w__5298);
  not g__5576(w__5295 ,w__5296);
  and g__5577(w__5294 ,w__5094 ,w__5178);
  and g__5578(w__5293 ,w__5172 ,w__5119);
  or g__5579(w__5292 ,w__5154 ,w__5168);
  and g__5580(w__5291 ,w__5104 ,w__5179);
  and g__5581(w__5290 ,w__5108 ,w__5092);
  and g__5582(w__5289 ,w__5152 ,w__5116);
  or g__5583(w__5288 ,w__5153 ,w__5183);
  and g__5584(w__5287 ,w__5160 ,w__5170);
  and g__5585(w__5286 ,w__5153 ,w__5183);
  and g__5586(w__5285 ,w__5102 ,w__5091);
  and g__5587(w__5284 ,w__5156 ,w__5180);
  or g__5588(w__5283 ,w__5097 ,w__5164);
  or g__5589(w__5282 ,w__5102 ,w__5091);
  or g__5590(w__5281 ,w__5117 ,w__5149);
  and g__5591(w__5280 ,w__5117 ,w__5149);
  or g__5592(w__5279 ,w__5105 ,w__5113);
  or g__5593(w__5278 ,w__5104 ,w__5179);
  or g__5594(w__5277 ,w__5108 ,w__5092);
  and g__5595(w__5276 ,w__5154 ,w__5168);
  or g__5596(w__5275 ,w__5090 ,w__5159);
  and g__5597(w__5274 ,w__5097 ,w__5164);
  and g__5598(w__5273 ,w__5100 ,w__5103);
  or g__5599(w__5272 ,w__5156 ,w__5180);
  and g__5600(w__5271 ,w__5177 ,w__5118);
  and g__5601(w__5270 ,w__5087 ,w__5161);
  and g__5602(w__5269 ,w__5101 ,w__5111);
  and g__5603(w__5268 ,w__5182 ,w__5173);
  and g__5604(w__5267 ,w__5181 ,w__5089);
  and g__5605(w__5266 ,w__5114 ,w__5151);
  or g__5606(w__5265 ,w__5100 ,w__5103);
  or g__5607(w__5264 ,w__5185 ,w__5079);
  and g__5608(w__5263 ,w__5105 ,w__5113);
  or g__5609(w__5262 ,w__5094 ,w__5178);
  or g__5610(w__5261 ,w__5086 ,w__5150);
  or g__5611(w__5260 ,w__5106 ,w__5174);
  and g__5612(w__5259 ,w__5098 ,w__5162);
  and g__5613(w__5258 ,w__5093 ,w__5167);
  or g__5614(w__5257 ,w__5112 ,w__5163);
  and g__5615(w__5256 ,w__5171 ,w__5157);
  and g__5616(w__5299 ,w__5141 ,w__5206);
  and g__5617(w__5298 ,w__5120 ,w__5190);
  and g__5618(w__5296 ,w__5122 ,w__5195);
  not g__5619(w__5254 ,w__5253);
  not g__5620(w__5249 ,w__5250);
  not g__5621(w__5246 ,w__5247);
  or g__5622(w__5245 ,w__5093 ,w__5167);
  xor g__5623(w__8368 ,in10[0] ,in11[0]);
  and g__5624(w__5244 ,w__5088 ,w__5109);
  and g__5625(w__5243 ,w__5110 ,w__5175);
  nor g__5626(w__5242 ,w__5135 ,w__5147);
  or g__5627(w__5241 ,w__5152 ,w__5116);
  or g__5628(w__5240 ,w__5182 ,w__5173);
  and g__5629(w__5239 ,w__5166 ,w__5155);
  or g__5630(w__5238 ,w__5184 ,w__5165);
  or g__5631(w__5237 ,w__5087 ,w__5161);
  or g__5632(w__5236 ,w__5110 ,w__5175);
  nor g__5633(w__5235 ,w__5202 ,w__5146);
  or g__5634(w__5234 ,w__5177 ,w__5118);
  and g__5635(w__5233 ,w__5106 ,w__5174);
  or g__5636(w__5232 ,w__5088 ,w__5109);
  or g__5637(w__5231 ,w__5158 ,w__5099);
  nor g__5638(w__5230 ,w__5132 ,w__5144);
  and g__5639(w__5229 ,w__5112 ,w__5163);
  or g__5640(w__5228 ,w__5123 ,w__5145);
  or g__5641(w__5227 ,w__5160 ,w__5170);
  and g__5642(w__5226 ,w__5184 ,w__5165);
  or g__5643(w__5225 ,w__5098 ,w__5162);
  and g__5644(w__5224 ,w__5158 ,w__5099);
  or g__5645(w__5223 ,w__5172 ,w__5119);
  or g__5646(w__5222 ,w__5114 ,w__5151);
  and g__5647(w__5221 ,w__5086 ,w__5150);
  or g__5648(w__5220 ,w__5181 ,w__5089);
  and g__5649(w__5219 ,w__5090 ,w__5159);
  or g__5650(w__5218 ,w__5166 ,w__5155);
  or g__5651(w__5217 ,w__5171 ,w__5157);
  or g__5652(w__5216 ,w__5101 ,w__5111);
  xnor g__5653(w__5215 ,in10[8] ,in11[8]);
  xnor g__5654(w__5214 ,in10[7] ,in11[7]);
  xnor g__5655(w__5213 ,in10[9] ,in11[9]);
  xnor g__5656(w__5212 ,in10[10] ,in11[10]);
  xnor g__5657(w__5211 ,in10[1] ,in11[1]);
  xnor g__5658(w__5255 ,in10[4] ,in11[4]);
  and g__5659(w__5253 ,w__5204 ,w__5136);
  and g__5660(w__5252 ,w__5208 ,w__5121);
  xnor g__5661(w__5251 ,in10[6] ,in11[6]);
  xnor g__5662(w__5250 ,in10[3] ,in11[3]);
  xnor g__5663(w__5248 ,in10[5] ,in11[5]);
  xnor g__5664(w__5247 ,in10[2] ,in11[2]);
  not g__5665(w__5208 ,w__5207);
  not g__5666(w__5206 ,w__5205);
  not g__5667(w__5204 ,w__5203);
  not g__5668(w__5195 ,w__5194);
  not g__5669(w__5190 ,w__5189);
  or g__5670(w__5148 ,w__4974 ,w__4933);
  nor g__5671(w__5147 ,in10[10] ,in11[10]);
  nor g__5672(w__5146 ,in10[8] ,in11[8]);
  nor g__5673(w__5145 ,in10[7] ,in11[7]);
  nor g__5674(w__5144 ,in10[9] ,in11[9]);
  and g__5675(w__5143 ,in10[9] ,in11[9]);
  or g__5676(w__5210 ,w__4902 ,w__4907);
  or g__5677(w__5209 ,w__4922 ,w__4925);
  or g__5678(w__5207 ,w__4931 ,w__4977);
  or g__5679(w__5205 ,w__4941 ,w__4943);
  or g__5680(w__5203 ,w__4864 ,w__4952);
  or g__5681(w__5202 ,w__4898 ,w__4905);
  or g__5682(w__5201 ,w__4879 ,w__4870);
  or g__5683(w__5200 ,w__4900 ,w__4954);
  or g__5684(w__5199 ,w__4965 ,w__4867);
  or g__5685(w__5198 ,w__4894 ,w__4858);
  or g__5686(w__5197 ,w__5003 ,w__4956);
  or g__5687(w__5196 ,w__4938 ,w__4986);
  or g__5688(w__5194 ,w__4950 ,w__4971);
  or g__5689(w__5193 ,w__4852 ,w__5013);
  or g__5690(w__5192 ,w__4861 ,w__4891);
  or g__5691(w__5191 ,w__5046 ,w__4855);
  or g__5692(w__5189 ,w__4912 ,w__4927);
  or g__5693(w__5188 ,w__5009 ,w__4980);
  or g__5694(w__5187 ,w__5037 ,w__4869);
  or g__5695(w__5186 ,w__4881 ,w__4958);
  or g__5696(w__5185 ,w__4867 ,w__4935);
  or g__5697(w__5184 ,w__4910 ,w__5006);
  or g__5698(w__5183 ,w__4945 ,w__4972);
  or g__5699(w__5182 ,w__4863 ,w__5018);
  or g__5700(w__5181 ,w__4861 ,w__4963);
  or g__5701(w__5180 ,w__4893 ,w__5020);
  or g__5702(w__5179 ,w__4846 ,w__5000);
  or g__5703(w__5178 ,w__4849 ,w__4876);
  or g__5704(w__5177 ,w__4918 ,w__4860);
  or g__5705(w__5176 ,w__4891 ,w__4873);
  or g__5706(w__5175 ,w__5035 ,w__5016);
  or g__5707(w__5174 ,w__4989 ,w__5022);
  or g__5708(w__5173 ,w__4875 ,w__4956);
  or g__5709(w__5172 ,w__4857 ,w__4866);
  or g__5710(w__5171 ,w__4896 ,w__5006);
  or g__5711(w__5170 ,w__4890 ,w__5011);
  or g__5712(w__5169 ,w__4840 ,w__5032);
  or g__5713(w__5168 ,w__4961 ,w__4995);
  or g__5714(w__5167 ,w__5043 ,w__4915);
  or g__5715(w__5166 ,w__4992 ,w__4975);
  or g__5716(w__5165 ,w__4947 ,w__5037);
  or g__5717(w__5164 ,w__4997 ,w__4855);
  or g__5718(w__5163 ,w__4851 ,w__4854);
  or g__5719(w__5162 ,w__5045 ,w__4848);
  or g__5720(w__5161 ,w__4888 ,w__4925);
  or g__5721(w__5160 ,w__4969 ,w__5022);
  or g__5722(w__5159 ,w__5040 ,w__4978);
  or g__5723(w__5158 ,w__4843 ,w__4950);
  or g__5724(w__5157 ,w__4920 ,w__4912);
  or g__5725(w__5156 ,w__4945 ,w__4928);
  or g__5726(w__5155 ,w__4885 ,w__5013);
  or g__5727(w__5154 ,w__4910 ,w__4905);
  or g__5728(w__5153 ,w__4952 ,w__4969);
  or g__5729(w__5152 ,w__5032 ,w__4943);
  or g__5730(w__5151 ,w__5030 ,w__4873);
  or g__5731(w__5150 ,w__5052 ,w__5073);
  or g__5732(w__5149 ,w__5049 ,w__4971);
  not g__5733(w__5096 ,w__5095);
  not g__5734(w__5085 ,w__5084);
  nor g__5735(w__5082 ,w__5052 ,w__5043);
  nor g__5736(w__5081 ,w__5049 ,w__5046);
  or g__5737(w__5080 ,w__5000 ,w__4947);
  nor g__5738(w__5079 ,in10[1] ,in11[1]);
  and g__5739(w__8369 ,in10[0] ,in11[0]);
  or g__5740(w__5142 ,w__4902 ,w__4981);
  and g__5741(w__5141 ,in10[5] ,in10[3]);
  and g__5742(w__5140 ,in10[1] ,in10[0]);
  or g__5743(w__5139 ,w__4872 ,w__4936);
  or g__5744(w__5138 ,w__4900 ,w__4986);
  or g__5745(w__5137 ,w__4882 ,w__4980);
  and g__5746(w__5136 ,in10[7] ,in10[3]);
  or g__5747(w__5135 ,w__4845 ,w__5025);
  or g__5748(w__5134 ,w__4879 ,w__4894);
  or g__5749(w__5133 ,w__4915 ,w__4983);
  or g__5750(w__5132 ,w__4966 ,w__4852);
  or g__5751(w__5131 ,w__4882 ,w__4997);
  or g__5752(w__5130 ,w__5040 ,w__4989);
  or g__5753(w__5129 ,w__4842 ,w__4931);
  or g__5754(w__5128 ,w__5030 ,w__4870);
  or g__5755(w__5127 ,w__4998 ,w__5011);
  or g__5756(w__5126 ,w__4876 ,w__5014);
  or g__5757(w__5125 ,w__4858 ,w__4981);
  or g__5758(w__5124 ,w__4939 ,w__4887);
  or g__5759(w__5123 ,w__5028 ,w__4995);
  and g__5760(w__5122 ,in10[3] ,in10[1]);
  and g__5761(w__5121 ,in11[2] ,in11[0]);
  and g__5762(w__5120 ,in10[4] ,in10[2]);
  or g__5763(w__5119 ,w__4885 ,w__4936);
  or g__5764(w__5118 ,w__4965 ,w__5038);
  or g__5765(w__5117 ,w__4839 ,w__5003);
  or g__5766(w__5116 ,w__4884 ,w__5023);
  or g__5767(w__5115 ,w__4990 ,w__4983);
  or g__5768(w__5114 ,w__4920 ,w__4968);
  or g__5769(w__5113 ,w__4898 ,w__4974);
  or g__5770(w__5112 ,w__4918 ,w__5016);
  or g__5771(w__5111 ,w__4849 ,w__5020);
  or g__5772(w__5110 ,w__5033 ,w__4992);
  or g__5773(w__5109 ,w__4987 ,w__4933);
  or g__5774(w__5108 ,w__5025 ,w__5035);
  or g__5775(w__5107 ,w__4949 ,w__4888);
  or g__5776(w__5106 ,w__4960 ,w__4977);
  or g__5777(w__5105 ,w__5001 ,w__4993);
  or g__5778(w__5104 ,w__5028 ,w__4896);
  or g__5779(w__5103 ,w__5009 ,w__4922);
  or g__5780(w__5102 ,w__4840 ,w__5018);
  or g__5781(w__5101 ,w__5026 ,w__4975);
  or g__5782(w__5100 ,w__5042 ,w__4984);
  or g__5783(w__5099 ,w__4966 ,w__4954);
  or g__5784(w__5098 ,w__4846 ,w__4961);
  or g__5785(w__5097 ,w__4907 ,w__4958);
  and g__5786(w__5095 ,in10[3] ,in10[0]);
  or g__5787(w__5094 ,w__4843 ,w__4963);
  or g__5788(w__5093 ,w__5051 ,w__4909);
  or g__5789(w__5092 ,w__5048 ,w__4864);
  or g__5790(w__5091 ,w__4914 ,w__4924);
  or g__5791(w__5090 ,w__4968 ,w__5004);
  or g__5792(w__5089 ,w__4917 ,w__4972);
  or g__5793(w__5088 ,w__4930 ,w__4928);
  or g__5794(w__5087 ,w__5007 ,w__4978);
  or g__5795(w__5086 ,w__4941 ,w__4904);
  and g__5796(w__5084 ,in11[9] ,in11[7]);
  or g__5797(w__5083 ,w__4878 ,w__4939);
  not g__5798(w__5078 ,in10[0]);
  not g__5799(w__5077 ,in11[0]);
  not g__5800(w__5076 ,in11[2]);
  not g__5801(w__5075 ,in11[6]);
  not g__5802(w__5074 ,in11[3]);
  not g__5803(w__5073 ,in10[3]);
  not g__5804(w__5072 ,in10[4]);
  not g__5805(w__5071 ,in10[5]);
  not g__5806(w__5070 ,in10[1]);
  not g__5807(w__5069 ,in11[1]);
  not g__5808(w__5068 ,in10[9]);
  not g__5809(w__5067 ,in10[6]);
  not g__5810(w__5066 ,in11[5]);
  not g__5811(w__5065 ,in10[2]);
  not g__5812(w__5064 ,in11[4]);
  not g__5813(w__5063 ,in11[7]);
  not g__5814(w__5062 ,in10[7]);
  not g__5815(w__5061 ,in10[8]);
  not g__5816(w__5060 ,in10[10]);
  not g__5817(w__5059 ,in11[10]);
  not g__5818(w__5058 ,in11[9]);
  not g__5819(w__5057 ,in11[8]);
  not g__5820(w__5054 ,w__5056);
  not g__5821(w__5056 ,w__5749);
  not g__5822(w__5053 ,w__5055);
  not g__5823(w__5055 ,w__5603);
  not g__5824(w__5052 ,w__5050);
  not g__5825(w__5051 ,w__5050);
  not g__5826(w__5050 ,w__5061);
  not g__5827(w__5049 ,w__5047);
  not g__5828(w__5048 ,w__5047);
  not g__5829(w__5047 ,w__5060);
  not g__5830(w__5046 ,w__5044);
  not g__5831(w__5045 ,w__5044);
  not g__5832(w__5044 ,w__5059);
  not g__5833(w__5043 ,w__5041);
  not g__5834(w__5042 ,w__5041);
  not g__5835(w__5041 ,w__5057);
  not g__5836(w__5040 ,w__5039);
  not g__5837(w__5039 ,w__5071);
  not g__5838(w__5038 ,w__5036);
  not g__5839(w__5037 ,w__5036);
  not g__5840(w__5036 ,w__5075);
  not g__5841(w__5035 ,w__5034);
  not g__5842(w__5034 ,w__5062);
  not g__5843(w__5033 ,w__5031);
  not g__5844(w__5032 ,w__5031);
  not g__5845(w__5031 ,w__5071);
  not g__5846(w__5030 ,w__5029);
  not g__5847(w__5029 ,w__5063);
  not g__5848(w__5028 ,w__5027);
  not g__5849(w__5027 ,w__5068);
  not g__5850(w__5026 ,w__5024);
  not g__5851(w__5025 ,w__5024);
  not g__5852(w__5024 ,w__5068);
  not g__5853(w__5023 ,w__5021);
  not g__5854(w__5022 ,w__5021);
  not g__5855(w__5021 ,w__5074);
  not g__5856(w__5020 ,w__5019);
  not g__5857(w__5019 ,w__5076);
  not g__5858(w__5018 ,w__5017);
  not g__5859(w__5017 ,w__5070);
  not g__5860(w__5016 ,w__5015);
  not g__5861(w__5015 ,w__5065);
  not g__5862(w__5014 ,w__5012);
  not g__5863(w__5013 ,w__5012);
  not g__5864(w__5012 ,w__5069);
  not g__5865(w__5011 ,w__5010);
  not g__5866(w__5010 ,w__5077);
  not g__5867(w__5009 ,w__5008);
  not g__5868(w__5008 ,w__5058);
  not g__5869(w__5007 ,w__5005);
  not g__5870(w__5006 ,w__5005);
  not g__5871(w__5005 ,w__5067);
  not g__5872(w__5004 ,w__5002);
  not g__5873(w__5003 ,w__5002);
  not g__5874(w__5002 ,w__5065);
  not g__5875(w__5001 ,w__4999);
  not g__5876(w__5000 ,w__4999);
  not g__5877(w__4999 ,w__5062);
  not g__5878(w__4998 ,w__4996);
  not g__5879(w__4997 ,w__4996);
  not g__5880(w__4996 ,w__5063);
  not g__5881(w__4995 ,w__4994);
  not g__5882(w__4994 ,w__5072);
  not g__5883(w__4993 ,w__4991);
  not g__5884(w__4992 ,w__4991);
  not g__5885(w__4991 ,w__5072);
  not g__5886(w__4990 ,w__4988);
  not g__5887(w__4989 ,w__4988);
  not g__5888(w__4988 ,w__5066);
  not g__5889(w__4987 ,w__4985);
  not g__5890(w__4986 ,w__4985);
  not g__5891(w__4985 ,w__5076);
  not g__5892(w__4984 ,w__4982);
  not g__5893(w__4983 ,w__4982);
  not g__5894(w__4982 ,w__5064);
  not g__5895(w__4981 ,w__4979);
  not g__5896(w__4980 ,w__4979);
  not g__5897(w__4979 ,w__5077);
  not g__5898(w__4978 ,w__4976);
  not g__5899(w__4977 ,w__4976);
  not g__5900(w__4976 ,w__5078);
  not g__5901(w__4975 ,w__4973);
  not g__5902(w__4974 ,w__4973);
  not g__5903(w__4973 ,w__5070);
  not g__5904(w__4972 ,w__4970);
  not g__5905(w__4971 ,w__4970);
  not g__5906(w__4970 ,w__5078);
  not g__5907(w__4969 ,w__4967);
  not g__5908(w__4968 ,w__4967);
  not g__5909(w__4967 ,w__5073);
  not g__5910(w__4966 ,w__4964);
  not g__5911(w__4965 ,w__4964);
  not g__5912(w__4964 ,w__5058);
  not g__5913(w__4963 ,w__4962);
  not g__5914(w__4962 ,w__5073);
  not g__5915(w__4961 ,w__4959);
  not g__5916(w__4960 ,w__4959);
  not g__5917(w__4959 ,w__5061);
  not g__5918(w__4958 ,w__4957);
  not g__5919(w__4957 ,w__4984);
  not g__5920(w__4956 ,w__4955);
  not g__5921(w__4955 ,w__4987);
  not g__5922(w__4954 ,w__4953);
  not g__5923(w__4953 ,w__4990);
  not g__5924(w__4952 ,w__4951);
  not g__5925(w__4951 ,w__4993);
  not g__5926(w__4950 ,w__4948);
  not g__5927(w__4949 ,w__4948);
  not g__5928(w__4948 ,w__5072);
  not g__5929(w__4947 ,w__4946);
  not g__5930(w__4946 ,w__4998);
  not g__5931(w__4945 ,w__4944);
  not g__5932(w__4944 ,w__5001);
  not g__5933(w__4943 ,w__4942);
  not g__5934(w__4942 ,w__5004);
  not g__5935(w__4941 ,w__4940);
  not g__5936(w__4940 ,w__5007);
  not g__5937(w__4939 ,w__4937);
  not g__5938(w__4938 ,w__4937);
  not g__5939(w__4937 ,w__5058);
  not g__5940(w__4936 ,w__4934);
  not g__5941(w__4935 ,w__4934);
  not g__5942(w__4934 ,w__5077);
  not g__5943(w__4933 ,w__4932);
  not g__5944(w__4932 ,w__5014);
  not g__5945(w__4931 ,w__4929);
  not g__5946(w__4930 ,w__4929);
  not g__5947(w__4929 ,w__5065);
  not g__5948(w__4928 ,w__4926);
  not g__5949(w__4927 ,w__4926);
  not g__5950(w__4926 ,w__5070);
  not g__5951(w__4925 ,w__4923);
  not g__5952(w__4924 ,w__4923);
  not g__5953(w__4923 ,w__5076);
  not g__5954(w__4922 ,w__4921);
  not g__5955(w__4921 ,w__5023);
  not g__5956(w__4920 ,w__4919);
  not g__5957(w__4919 ,w__5026);
  not g__5958(w__4918 ,w__4916);
  not g__5959(w__4917 ,w__4916);
  not g__5960(w__4916 ,w__5068);
  not g__5961(w__4915 ,w__4913);
  not g__5962(w__4914 ,w__4913);
  not g__5963(w__4913 ,w__5063);
  not g__5964(w__4912 ,w__4911);
  not g__5965(w__4911 ,w__5033);
  not g__5966(w__4910 ,w__4908);
  not g__5967(w__4909 ,w__4908);
  not g__5968(w__4908 ,w__5062);
  not g__5969(w__4907 ,w__4906);
  not g__5970(w__4906 ,w__5038);
  not g__5971(w__4905 ,w__4903);
  not g__5972(w__4904 ,w__4903);
  not g__5973(w__4903 ,w__5071);
  not g__5974(w__4902 ,w__4901);
  not g__5975(w__4901 ,w__5042);
  not g__5976(w__4900 ,w__4899);
  not g__5977(w__4899 ,w__5045);
  not g__5978(w__4898 ,w__4897);
  not g__5979(w__4897 ,w__5048);
  not g__5980(w__4896 ,w__4895);
  not g__5981(w__4895 ,w__5051);
  not g__5982(w__4894 ,w__4892);
  not g__5983(w__4893 ,w__4892);
  not g__5984(w__4892 ,w__5075);
  not g__5985(w__4891 ,w__4889);
  not g__5986(w__4890 ,w__4889);
  not g__5987(w__4889 ,w__5075);
  not g__5988(w__4888 ,w__4886);
  not g__5989(w__4887 ,w__4886);
  not g__5990(w__4886 ,w__5064);
  not g__5991(w__4885 ,w__4883);
  not g__5992(w__4884 ,w__4883);
  not g__5993(w__4883 ,w__5064);
  not g__5994(w__4882 ,w__4880);
  not g__5995(w__4881 ,w__4880);
  not g__5996(w__4880 ,w__5059);
  not g__5997(w__4879 ,w__4877);
  not g__5998(w__4878 ,w__4877);
  not g__5999(w__4877 ,w__5059);
  not g__6000(w__4876 ,w__4874);
  not g__6001(w__4875 ,w__4874);
  not g__6002(w__4874 ,w__5066);
  not g__6003(w__4873 ,w__4871);
  not g__6004(w__4872 ,w__4871);
  not g__6005(w__4871 ,w__5066);
  not g__6006(w__4870 ,w__4868);
  not g__6007(w__4869 ,w__4868);
  not g__6008(w__4868 ,w__5069);
  not g__6009(w__4867 ,w__4865);
  not g__6010(w__4866 ,w__4865);
  not g__6011(w__4865 ,w__5069);
  not g__6012(w__4864 ,w__4862);
  not g__6013(w__4863 ,w__4862);
  not g__6014(w__4862 ,w__5067);
  not g__6015(w__4861 ,w__4859);
  not g__6016(w__4860 ,w__4859);
  not g__6017(w__4859 ,w__5067);
  not g__6018(w__4858 ,w__4856);
  not g__6019(w__4857 ,w__4856);
  not g__6020(w__4856 ,w__5074);
  not g__6021(w__4855 ,w__4853);
  not g__6022(w__4854 ,w__4853);
  not g__6023(w__4853 ,w__5074);
  not g__6024(w__4852 ,w__4850);
  not g__6025(w__4851 ,w__4850);
  not g__6026(w__4850 ,w__5057);
  not g__6027(w__4849 ,w__4847);
  not g__6028(w__4848 ,w__4847);
  not g__6029(w__4847 ,w__5057);
  not g__6030(w__4846 ,w__4844);
  not g__6031(w__4845 ,w__4844);
  not g__6032(w__4844 ,w__5060);
  not g__6033(w__4843 ,w__4841);
  not g__6034(w__4842 ,w__4841);
  not g__6035(w__4841 ,w__5060);
  not g__6036(w__4840 ,w__4838);
  not g__6037(w__4839 ,w__4838);
  not g__6038(w__4838 ,w__5061);
  xor g__6039(w__8383 ,w__5882 ,w__5863);
  xor g__6040(w__8382 ,w__5880 ,w__5870);
  xor g__6041(w__8381 ,w__5878 ,w__5871);
  xor g__6042(w__8380 ,w__5876 ,w__5862);
  xor g__6043(w__8379 ,w__5874 ,w__5851);
  xor g__6044(w__8377 ,w__5855 ,w__5820);
  xor g__6045(w__4837 ,w__5141 ,w__5205);
  xnor g__6046(w__8370 ,w__5140 ,w__5397);
  xor g__6047(w__4836 ,w__5203 ,w__5136);
  xor g__6048(w__4835 ,w__5122 ,w__5194);
  xor g__6049(w__4834 ,w__5207 ,w__5121);
  xor g__6050(w__4833 ,w__5120 ,w__5189);
  xnor g__6051(w__8366 ,w__6572 ,w__6021);
  and g__6052(w__8367 ,w__6021 ,w__6573);
  not g__6053(w__6573 ,w__6572);
  and g__6054(w__6572 ,w__6274 ,w__6571);
  or g__6055(w__6571 ,w__6259 ,w__6570);
  and g__6056(w__6570 ,w__6371 ,w__6569);
  or g__6057(w__6569 ,w__6370 ,w__6568);
  and g__6058(w__6568 ,w__6419 ,w__6567);
  or g__6059(w__6567 ,w__6421 ,w__6566);
  and g__6060(w__6566 ,w__6476 ,w__6565);
  or g__6061(w__6565 ,w__6468 ,w__6564);
  and g__6062(w__6564 ,w__6502 ,w__6563);
  or g__6063(w__6563 ,w__6503 ,w__6562);
  and g__6064(w__6562 ,w__6510 ,w__6561);
  or g__6065(w__6561 ,w__6509 ,w__6560);
  and g__6066(w__6560 ,w__6534 ,w__6559);
  or g__6067(w__6559 ,w__6535 ,w__6558);
  and g__6068(w__6558 ,w__6541 ,w__6557);
  or g__6069(w__6557 ,w__6540 ,w__6556);
  and g__6070(w__6556 ,w__6533 ,w__6555);
  or g__6071(w__6555 ,w__6532 ,w__6554);
  and g__6072(w__6554 ,w__6531 ,w__6553);
  or g__6073(w__6553 ,w__6530 ,w__6552);
  and g__6074(w__6552 ,w__6521 ,w__6551);
  or g__6075(w__6551 ,w__6520 ,w__6550);
  and g__6076(w__6550 ,w__6507 ,w__6549);
  xnor g__6077(w__8354 ,w__6547 ,w__6514);
  or g__6078(w__6549 ,w__6501 ,w__6548);
  not g__6079(w__6548 ,w__6547);
  or g__6080(w__6547 ,w__6482 ,w__6546);
  xnor g__6081(w__8353 ,w__6545 ,w__6499);
  and g__6082(w__6546 ,w__6489 ,w__6545);
  or g__6083(w__6545 ,w__6459 ,w__6544);
  xnor g__6084(w__8352 ,w__6542 ,w__6467);
  and g__6085(w__6544 ,w__6458 ,w__6542);
  xnor g__6086(w__6543 ,w__6523 ,w__6529);
  or g__6087(w__6542 ,w__6437 ,w__6536);
  or g__6088(w__6541 ,w__6522 ,w__6528);
  nor g__6089(w__6540 ,w__6523 ,w__6529);
  xnor g__6090(w__6539 ,w__6525 ,w__6505);
  xnor g__6091(w__6538 ,w__6493 ,w__6517);
  xnor g__6092(w__6537 ,w__6495 ,w__6519);
  xnor g__6093(w__8351 ,w__6526 ,w__6445);
  and g__6094(w__6536 ,w__6436 ,w__6526);
  nor g__6095(w__6535 ,w__6525 ,w__6505);
  or g__6096(w__6534 ,w__6524 ,w__6504);
  or g__6097(w__6533 ,w__6492 ,w__6516);
  nor g__6098(w__6532 ,w__6493 ,w__6517);
  or g__6099(w__6531 ,w__6494 ,w__6518);
  nor g__6100(w__6530 ,w__6495 ,w__6519);
  not g__6101(w__6529 ,w__6528);
  xnor g__6102(w__6528 ,w__6453 ,w__6500);
  xnor g__6103(w__6527 ,w__6506 ,w__6497);
  not g__6104(w__6524 ,w__6525);
  not g__6105(w__6522 ,w__6523);
  or g__6106(w__6521 ,w__6497 ,w__6506);
  and g__6107(w__6520 ,w__6497 ,w__6506);
  or g__6108(w__6526 ,w__6406 ,w__6511);
  or g__6109(w__6525 ,w__6491 ,w__6508);
  or g__6110(w__6523 ,w__6432 ,w__6512);
  not g__6111(w__6519 ,w__6518);
  not g__6112(w__6517 ,w__6516);
  xnor g__6113(w__8350 ,w__6498 ,w__6416);
  xnor g__6114(w__6515 ,w__6483 ,w__6496);
  xnor g__6115(w__6514 ,w__6480 ,w__6487);
  xnor g__6116(w__6513 ,w__6478 ,w__6485);
  xnor g__6117(w__6518 ,w__6425 ,w__5907);
  xnor g__6118(w__6516 ,w__6488 ,w__6444);
  and g__6119(w__6512 ,w__6420 ,w__6488);
  and g__6120(w__6511 ,w__6405 ,w__6498);
  or g__6121(w__6510 ,w__6496 ,w__6483);
  and g__6122(w__6509 ,w__6496 ,w__6483);
  nor g__6123(w__6508 ,w__6453 ,w__6490);
  or g__6124(w__6507 ,w__6479 ,w__6486);
  not g__6125(w__6504 ,w__6505);
  nor g__6126(w__6503 ,w__6478 ,w__6485);
  or g__6127(w__6502 ,w__6477 ,w__6484);
  nor g__6128(w__6501 ,w__6480 ,w__6487);
  xnor g__6129(w__6500 ,w__6471 ,w__6045);
  xnor g__6130(w__6499 ,w__6451 ,w__6470);
  xnor g__6131(w__6506 ,w__6413 ,w__6466);
  xnor g__6132(w__6505 ,w__6441 ,w__6465);
  not g__6133(w__6494 ,w__6495);
  not g__6134(w__6493 ,w__6492);
  and g__6135(w__6491 ,w__6045 ,w__6471);
  nor g__6136(w__6490 ,w__6044 ,w__6471);
  or g__6137(w__6489 ,w__6451 ,w__6470);
  or g__6138(w__6498 ,w__6404 ,w__6472);
  and g__6139(w__6497 ,w__6461 ,w__6473);
  and g__6140(w__6496 ,w__6460 ,w__6475);
  or g__6141(w__6495 ,w__6456 ,w__6474);
  and g__6142(w__6492 ,w__6455 ,w__6469);
  not g__6143(w__6486 ,w__6487);
  not g__6144(w__6484 ,w__6485);
  xnor g__6145(w__8349 ,w__6463 ,w__6415);
  and g__6146(w__6482 ,w__6451 ,w__6470);
  xnor g__6147(w__6481 ,w__6452 ,w__6462);
  xnor g__6148(w__6488 ,w__6443 ,w__6053);
  xnor g__6149(w__6487 ,w__6428 ,w__5899);
  xnor g__6150(w__6485 ,w__6447 ,w__6049);
  xnor g__6151(w__6483 ,w__6396 ,w__6442);
  not g__6152(w__6480 ,w__6479);
  not g__6153(w__6478 ,w__6477);
  or g__6154(w__6476 ,w__6462 ,w__6452);
  or g__6155(w__6475 ,w__6441 ,w__5906);
  nor g__6156(w__6474 ,w__6413 ,w__6450);
  or g__6157(w__6473 ,w__6399 ,w__6457);
  and g__6158(w__6472 ,w__6403 ,w__6463);
  and g__6159(w__6479 ,w__6440 ,w__6448);
  and g__6160(w__6477 ,w__6430 ,w__6449);
  or g__6161(w__6469 ,w__6464 ,w__6454);
  xnor g__6162(w__8348 ,w__6398 ,w__6417);
  and g__6163(w__6468 ,w__6462 ,w__6452);
  xnor g__6164(w__6467 ,w__6410 ,w__6423);
  xnor g__6165(w__6466 ,w__6422 ,w__6036);
  xnor g__6166(w__6465 ,w__6426 ,w__6063);
  xnor g__6167(w__6471 ,w__6333 ,w__6418);
  xnor g__6168(w__6470 ,w__6386 ,w__5898);
  or g__6169(w__6461 ,w__6082 ,w__6428);
  or g__6170(w__6460 ,w__6095 ,w__6426);
  and g__6171(w__6459 ,w__6410 ,w__6423);
  or g__6172(w__6458 ,w__6410 ,w__6423);
  nor g__6173(w__6457 ,w__6051 ,w__6427);
  and g__6174(w__6456 ,w__6036 ,w__6422);
  or g__6175(w__6455 ,w__6389 ,w__6425);
  nor g__6176(w__6454 ,w__6390 ,w__6424);
  and g__6177(w__6464 ,w__6400 ,w__6431);
  or g__6178(w__6463 ,w__6402 ,w__6433);
  and g__6179(w__6462 ,w__6373 ,w__6434);
  nor g__6180(w__6450 ,w__6035 ,w__6422);
  or g__6181(w__6449 ,w__6396 ,w__6435);
  or g__6182(w__6448 ,w__6366 ,w__6439);
  xnor g__6183(w__6447 ,w__6414 ,w__6331);
  xnor g__6184(w__6446 ,w__6395 ,w__6388);
  xnor g__6185(w__6445 ,w__6379 ,w__6391);
  xnor g__6186(w__6444 ,w__6384 ,w__6412);
  xnor g__6187(w__6443 ,w__6397 ,w__6289);
  xnor g__6188(w__6442 ,w__6393 ,w__6066);
  and g__6189(w__6453 ,w__6348 ,w__6429);
  xnor g__6190(w__6452 ,w__6380 ,w__6056);
  or g__6191(w__6451 ,w__6409 ,w__6438);
  or g__6192(w__6440 ,w__6094 ,w__6386);
  nor g__6193(w__6439 ,w__6047 ,w__6385);
  nor g__6194(w__6438 ,w__6316 ,w__6408);
  and g__6195(w__6437 ,w__6379 ,w__6391);
  or g__6196(w__6436 ,w__6379 ,w__6391);
  nor g__6197(w__6435 ,w__6065 ,w__6393);
  or g__6198(w__6434 ,w__5905 ,w__6414);
  and g__6199(w__6433 ,w__6398 ,w__6382);
  nor g__6200(w__6432 ,w__6384 ,w__6411);
  or g__6201(w__6431 ,w__6317 ,w__6401);
  or g__6202(w__6430 ,w__6092 ,w__6392);
  or g__6203(w__6429 ,w__5904 ,w__6397);
  and g__6204(w__6441 ,w__6369 ,w__6407);
  not g__6205(w__6427 ,w__6428);
  not g__6206(w__6424 ,w__6425);
  nor g__6207(w__6421 ,w__6395 ,w__6388);
  or g__6208(w__6420 ,w__6383 ,w__6412);
  or g__6209(w__6419 ,w__6394 ,w__6387);
  xnor g__6210(w__6418 ,w__6292 ,w__6365);
  xnor g__6211(w__6417 ,w__6206 ,w__5897);
  xnor g__6212(w__6416 ,w__6312 ,w__6363);
  xnor g__6213(w__6415 ,w__6315 ,w__6361);
  xnor g__6214(w__6428 ,w__6336 ,w__6354);
  xnor g__6215(w__6426 ,w__6351 ,w__6357);
  xnor g__6216(w__6425 ,w__6352 ,w__6355);
  xnor g__6217(w__6423 ,w__6360 ,w__6356);
  xnor g__6218(w__6422 ,w__6362 ,w__6353);
  not g__6219(w__6411 ,w__6412);
  nor g__6220(w__6409 ,w__6091 ,w__6360);
  and g__6221(w__6408 ,w__6091 ,w__6360);
  or g__6222(w__6407 ,w__6365 ,w__6367);
  and g__6223(w__6406 ,w__6312 ,w__6363);
  or g__6224(w__6405 ,w__6312 ,w__6363);
  and g__6225(w__6404 ,w__6315 ,w__6361);
  or g__6226(w__6403 ,w__6315 ,w__6361);
  nor g__6227(w__6402 ,w__6206 ,w__5897);
  and g__6228(w__6401 ,w__6294 ,w__6362);
  or g__6229(w__6400 ,w__6294 ,w__6362);
  and g__6230(w__6414 ,w__6338 ,w__6374);
  and g__6231(w__6413 ,w__6340 ,w__6368);
  or g__6232(w__6412 ,w__6344 ,w__6372);
  or g__6233(w__6410 ,w__6311 ,w__6375);
  not g__6234(w__6394 ,w__6395);
  not g__6235(w__6392 ,w__6393);
  not g__6236(w__6389 ,w__6390);
  not g__6237(w__6388 ,w__6387);
  not g__6238(w__6385 ,w__6386);
  not g__6239(w__6383 ,w__6384);
  or g__6240(w__6382 ,w__6205 ,w__6364);
  xnor g__6241(w__8347 ,w__6350 ,w__6283);
  xnor g__6242(w__6381 ,w__6300 ,w__6349);
  xnor g__6243(w__6380 ,w__6335 ,w__6297);
  and g__6244(w__6399 ,w__6329 ,w__6359);
  or g__6245(w__6398 ,w__6257 ,w__6358);
  and g__6246(w__6397 ,w__6325 ,w__6377);
  and g__6247(w__6396 ,w__6346 ,w__6376);
  xnor g__6248(w__6395 ,w__6321 ,w__6058);
  xnor g__6249(w__6393 ,w__6298 ,w__6320);
  xnor g__6250(w__6391 ,w__6334 ,w__6319);
  xnor g__6251(w__6390 ,w__6288 ,w__6322);
  and g__6252(w__6387 ,w__6337 ,w__6378);
  xnor g__6253(w__6386 ,w__6290 ,w__6324);
  xnor g__6254(w__6384 ,w__6265 ,w__6323);
  or g__6255(w__6378 ,w__6335 ,w__6343);
  or g__6256(w__6377 ,w__6279 ,w__6347);
  or g__6257(w__6376 ,w__6351 ,w__6339);
  nor g__6258(w__6375 ,w__6310 ,w__6334);
  or g__6259(w__6374 ,w__6264 ,w__6330);
  or g__6260(w__6373 ,w__6090 ,w__6331);
  nor g__6261(w__6372 ,w__6342 ,w__6352);
  or g__6262(w__6371 ,w__6349 ,w__6300);
  and g__6263(w__6370 ,w__6349 ,w__6300);
  or g__6264(w__6369 ,w__6291 ,w__6333);
  or g__6265(w__6368 ,w__6345 ,w__6336);
  nor g__6266(w__6367 ,w__6292 ,w__6332);
  or g__6267(w__6379 ,w__6260 ,w__6327);
  not g__6268(w__6364 ,w__5897);
  or g__6269(w__6359 ,w__6263 ,w__6328);
  nor g__6270(w__6358 ,w__6271 ,w__6350);
  xor g__6271(w__8346 ,w__6200 ,w__6282);
  xnor g__6272(w__6357 ,w__6295 ,w__6277);
  xnor g__6273(w__6356 ,w__6316 ,w__6027);
  xnor g__6274(w__6355 ,w__6314 ,w__6042);
  xnor g__6275(w__6354 ,w__6293 ,w__6313);
  xor g__6276(w__6353 ,w__6294 ,w__6317);
  and g__6277(w__6366 ,w__6258 ,w__6326);
  and g__6278(w__6365 ,w__6304 ,w__6341);
  xnor g__6279(w__6363 ,w__6318 ,w__5896);
  xnor g__6280(w__6362 ,w__6281 ,w__6285);
  xnor g__6281(w__6361 ,w__6284 ,w__6029);
  xnor g__6282(w__6360 ,w__6301 ,w__6287);
  or g__6283(w__6348 ,w__6078 ,w__6289);
  and g__6284(w__6347 ,w__6183 ,w__6288);
  or g__6285(w__6346 ,w__6277 ,w__6295);
  and g__6286(w__6345 ,w__6313 ,w__6293);
  and g__6287(w__6344 ,w__6042 ,w__6314);
  nor g__6288(w__6343 ,w__6055 ,w__6297);
  nor g__6289(w__6342 ,w__6041 ,w__6314);
  or g__6290(w__6341 ,w__6265 ,w__6308);
  or g__6291(w__6340 ,w__6313 ,w__6293);
  and g__6292(w__6339 ,w__6277 ,w__6295);
  or g__6293(w__6338 ,w__6115 ,w__6299);
  or g__6294(w__6337 ,w__6079 ,w__6296);
  and g__6295(w__6352 ,w__6269 ,w__6307);
  and g__6296(w__6351 ,w__6172 ,w__6309);
  and g__6297(w__6350 ,w__6273 ,w__6305);
  and g__6298(w__6349 ,w__6197 ,w__6306);
  not g__6299(w__6332 ,w__6333);
  and g__6300(w__6330 ,w__6115 ,w__6299);
  or g__6301(w__6329 ,w__6199 ,w__6290);
  and g__6302(w__6328 ,w__6199 ,w__6290);
  and g__6303(w__6327 ,w__6255 ,w__6318);
  or g__6304(w__6326 ,w__6261 ,w__6301);
  or g__6305(w__6325 ,w__6183 ,w__6288);
  xnor g__6306(w__6324 ,w__6199 ,w__6263);
  xnor g__6307(w__6323 ,w__6136 ,w__6262);
  xor g__6308(w__6322 ,w__6183 ,w__6279);
  xnor g__6309(w__6321 ,w__6280 ,w__6137);
  xnor g__6310(w__6320 ,w__6115 ,w__6264);
  xnor g__6311(w__6319 ,w__6276 ,w__6025);
  xnor g__6312(w__6336 ,w__6227 ,w__6253);
  and g__6313(w__6335 ,w__6163 ,w__6303);
  xnor g__6314(w__6334 ,w__5900 ,w__6252);
  xnor g__6315(w__6333 ,w__6278 ,w__6210);
  xnor g__6316(w__6331 ,w__6266 ,w__6214);
  nor g__6317(w__6311 ,w__6096 ,w__6276);
  and g__6318(w__6310 ,w__6096 ,w__6276);
  or g__6319(w__6309 ,w__6167 ,w__6278);
  and g__6320(w__6308 ,w__6136 ,w__6262);
  or g__6321(w__6307 ,w__6281 ,w__6275);
  or g__6322(w__6306 ,w__5901 ,w__6280);
  or g__6323(w__6305 ,w__6200 ,w__6270);
  or g__6324(w__6304 ,w__6136 ,w__6262);
  or g__6325(w__6303 ,w__6193 ,w__6266);
  xnor g__6326(w__6302 ,w__6112 ,w__6226);
  xnor g__6327(w__6318 ,w__6184 ,w__6209);
  and g__6328(w__6317 ,w__6235 ,w__6254);
  and g__6329(w__6316 ,w__6242 ,w__6267);
  or g__6330(w__6315 ,w__6188 ,w__6268);
  xnor g__6331(w__6314 ,w__6102 ,w__6230);
  and g__6332(w__6313 ,w__6177 ,w__6256);
  or g__6333(w__6312 ,w__6246 ,w__6272);
  not g__6334(w__6299 ,w__6298);
  not g__6335(w__6296 ,w__6297);
  not g__6336(w__6291 ,w__6292);
  xnor g__6337(w__6287 ,w__6182 ,w__6225);
  xnor g__6338(w__6286 ,w__6249 ,w__6061);
  xnor g__6339(w__6285 ,w__6204 ,w__6220);
  xnor g__6340(w__6284 ,w__5902 ,w__6202);
  xnor g__6341(w__6283 ,w__6203 ,w__6250);
  xnor g__6342(w__6282 ,w__6222 ,w__6069);
  xnor g__6343(w__6301 ,w__6114 ,w__6211);
  xnor g__6344(w__6300 ,w__6229 ,w__6039);
  xnor g__6345(w__6298 ,w__6138 ,w__6216);
  xnor g__6346(w__6297 ,w__6132 ,w__6213);
  xnor g__6347(w__6295 ,w__6105 ,w__6207);
  xnor g__6348(w__6294 ,w__6107 ,w__6208);
  xnor g__6349(w__6293 ,w__6142 ,w__6219);
  xnor g__6350(w__6292 ,w__6100 ,w__6217);
  xnor g__6351(w__6290 ,w__5903 ,w__6212);
  xnor g__6352(w__6289 ,w__6133 ,w__6215);
  xnor g__6353(w__6288 ,w__6152 ,w__6218);
  and g__6354(w__6275 ,w__6204 ,w__6220);
  or g__6355(w__6274 ,w__6083 ,w__6248);
  or g__6356(w__6273 ,w__6081 ,w__6221);
  nor g__6357(w__6272 ,w__6236 ,w__5902);
  and g__6358(w__6271 ,w__6203 ,w__6251);
  nor g__6359(w__6270 ,w__6068 ,w__6222);
  or g__6360(w__6269 ,w__6204 ,w__6220);
  and g__6361(w__6268 ,w__6195 ,w__6226);
  or g__6362(w__6267 ,w__6244 ,w__5900);
  and g__6363(w__6281 ,w__6176 ,w__6238);
  and g__6364(w__6280 ,w__6192 ,w__6231);
  and g__6365(w__6279 ,w__6164 ,w__6245);
  and g__6366(w__6278 ,w__6194 ,w__6237);
  and g__6367(w__6277 ,w__6198 ,w__6243);
  and g__6368(w__6276 ,w__6170 ,w__6241);
  nor g__6369(w__6261 ,w__6182 ,w__6225);
  and g__6370(w__6260 ,w__6031 ,w__6223);
  nor g__6371(w__6259 ,w__6060 ,w__6249);
  or g__6372(w__6258 ,w__6181 ,w__6224);
  nor g__6373(w__6257 ,w__6203 ,w__6251);
  or g__6374(w__6256 ,w__6166 ,w__5903);
  or g__6375(w__6255 ,w__6031 ,w__6223);
  or g__6376(w__6254 ,w__6228 ,w__6247);
  xnor g__6377(w__6253 ,w__6145 ,w__6180);
  xnor g__6378(w__6252 ,w__6109 ,w__6201);
  and g__6379(w__6266 ,w__6187 ,w__6240);
  and g__6380(w__6265 ,w__6165 ,w__6233);
  and g__6381(w__6264 ,w__6174 ,w__6239);
  and g__6382(w__6263 ,w__6178 ,w__6232);
  and g__6383(w__6262 ,w__6190 ,w__6234);
  not g__6384(w__6251 ,w__6250);
  not g__6385(w__6249 ,w__6248);
  nor g__6386(w__6247 ,w__6144 ,w__6180);
  nor g__6387(w__6246 ,w__6080 ,w__6202);
  or g__6388(w__6245 ,w__6123 ,w__6171);
  and g__6389(w__6244 ,w__6109 ,w__6201);
  or g__6390(w__6243 ,w__6122 ,w__6186);
  or g__6391(w__6242 ,w__6109 ,w__6201);
  or g__6392(w__6240 ,w__6149 ,w__6185);
  or g__6393(w__6239 ,w__6150 ,w__6168);
  or g__6394(w__6238 ,w__6125 ,w__6175);
  or g__6395(w__6237 ,w__6118 ,w__6173);
  and g__6396(w__6236 ,w__6080 ,w__6202);
  or g__6397(w__6235 ,w__6145 ,w__6179);
  or g__6398(w__6234 ,w__6127 ,w__6191);
  or g__6399(w__6233 ,w__6152 ,w__6162);
  or g__6400(w__6232 ,w__6120 ,w__6169);
  or g__6401(w__6231 ,w__6151 ,w__6189);
  xnor g__6402(w__6230 ,w__6127 ,in9[6]);
  xnor g__6403(w__6229 ,w__6128 ,in9[10]);
  xnor g__6404(w__6250 ,w__6156 ,w__6023);
  and g__6405(w__6248 ,w__6098 ,w__6196);
  not g__6406(w__6228 ,w__6227);
  not g__6407(w__6224 ,w__6225);
  not g__6408(w__6221 ,w__6222);
  xnor g__6409(w__6219 ,w__6101 ,w__6125);
  xnor g__6410(w__6218 ,w__6106 ,w__6140);
  xnor g__6411(w__6217 ,w__6122 ,in9[7]);
  xnor g__6412(w__6216 ,w__6149 ,in9[8]);
  xnor g__6413(w__6215 ,w__6103 ,w__6118);
  xnor g__6414(w__6214 ,w__6135 ,w__6104);
  xnor g__6415(w__6213 ,w__6151 ,in9[9]);
  xnor g__6416(w__6212 ,w__6131 ,w__6143);
  xnor g__6417(w__6211 ,w__6134 ,w__6120);
  xnor g__6418(w__6210 ,w__6113 ,w__6110);
  xnor g__6419(w__6209 ,w__6108 ,w__6141);
  xnor g__6420(w__6208 ,w__6139 ,w__6123);
  xnor g__6421(w__6207 ,w__6099 ,w__6150);
  xnor g__6422(w__6227 ,w__6158 ,in9[5]);
  xnor g__6423(w__6226 ,w__6121 ,in9[2]);
  xnor g__6424(w__6225 ,w__6126 ,in9[4]);
  xnor g__6425(w__6223 ,w__6155 ,in9[3]);
  xnor g__6426(w__6222 ,w__6147 ,in9[1]);
  xnor g__6427(w__6220 ,w__6159 ,w__6116);
  not g__6428(w__6206 ,w__6205);
  or g__6429(w__6198 ,w__5920 ,w__6100);
  or g__6430(w__6197 ,w__6097 ,w__6137);
  or g__6431(w__6196 ,w__6128 ,w__6129);
  or g__6432(w__6195 ,w__6033 ,w__6111);
  or g__6433(w__6194 ,w__6103 ,w__6133);
  and g__6434(w__6193 ,w__6135 ,w__6104);
  or g__6435(w__6192 ,w__5910 ,w__6132);
  and g__6436(w__6191 ,w__5930 ,w__6102);
  or g__6437(w__6190 ,w__5934 ,w__6102);
  and g__6438(w__6189 ,w__5914 ,w__6132);
  nor g__6439(w__6188 ,w__6084 ,w__6112);
  or g__6440(w__6187 ,w__5959 ,w__6138);
  and g__6441(w__6186 ,w__5924 ,w__6100);
  and g__6442(w__6185 ,w__5946 ,w__6138);
  and g__6443(w__6205 ,w__6023 ,w__6157);
  or g__6444(w__6204 ,w__5967 ,w__6158);
  or g__6445(w__6203 ,w__5977 ,w__6147);
  or g__6446(w__6202 ,w__5986 ,w__6121);
  or g__6447(w__6201 ,w__5980 ,w__6155);
  or g__6448(w__6200 ,w__6070 ,w__6119);
  or g__6449(w__6199 ,w__5983 ,w__6126);
  not g__6450(w__6181 ,w__6182);
  not g__6451(w__6179 ,w__6180);
  and g__6452(w__8344 ,w__6119 ,w__6130);
  or g__6453(w__6178 ,w__6114 ,w__6134);
  or g__6454(w__6177 ,w__6131 ,w__6143);
  or g__6455(w__6176 ,w__6142 ,w__6101);
  and g__6456(w__6175 ,w__6142 ,w__6101);
  or g__6457(w__6174 ,w__6099 ,w__6105);
  and g__6458(w__6173 ,w__6103 ,w__6133);
  or g__6459(w__6172 ,w__6113 ,w__6110);
  and g__6460(w__6171 ,w__6107 ,w__6139);
  or g__6461(w__6170 ,w__6108 ,w__6141);
  and g__6462(w__6169 ,w__6114 ,w__6134);
  and g__6463(w__6168 ,w__6099 ,w__6105);
  and g__6464(w__6167 ,w__6113 ,w__6110);
  and g__6465(w__6166 ,w__6131 ,w__6143);
  or g__6466(w__6165 ,w__6106 ,w__6140);
  or g__6467(w__6164 ,w__6107 ,w__6139);
  or g__6468(w__6163 ,w__6135 ,w__6104);
  and g__6469(w__6162 ,w__6106 ,w__6140);
  and g__6470(w__6184 ,w__6146 ,w__6117);
  or g__6471(w__6183 ,w__6159 ,w__6116);
  and g__6472(w__6182 ,w__6124 ,w__6154);
  and g__6473(w__6180 ,w__6148 ,w__6161);
  not g__6474(w__6161 ,w__6160);
  not g__6475(w__6157 ,w__6156);
  not g__6476(w__6154 ,w__6153);
  not g__6477(w__6145 ,w__6144);
  or g__6478(w__6130 ,in9[0] ,w__6019);
  nor g__6479(w__6129 ,in9[10] ,w__6038);
  or g__6480(w__6160 ,w__5943 ,w__5962);
  or g__6481(w__6159 ,w__5932 ,w__5951);
  or g__6482(w__6158 ,w__5912 ,w__5964);
  or g__6483(w__6156 ,w__5948 ,w__5994);
  or g__6484(w__6155 ,w__5969 ,w__5997);
  or g__6485(w__6153 ,w__5927 ,w__5964);
  or g__6486(w__6152 ,w__5972 ,w__6009);
  or g__6487(w__6151 ,w__5957 ,w__5922);
  or g__6488(w__6150 ,w__5940 ,w__6007);
  or g__6489(w__6149 ,w__5937 ,w__5989);
  and g__6490(w__6148 ,in9[5] ,in9[3]);
  or g__6491(w__6147 ,w__5974 ,w__5962);
  and g__6492(w__6146 ,in9[3] ,in9[1]);
  and g__6493(w__6144 ,in9[8] ,in9[1]);
  or g__6494(w__6143 ,w__5917 ,w__5975);
  or g__6495(w__6142 ,w__5992 ,w__5984);
  or g__6496(w__6141 ,w__5952 ,w__5978);
  or g__6497(w__6140 ,w__5999 ,w__5954);
  or g__6498(w__6139 ,w__5945 ,w__5987);
  or g__6499(w__6138 ,w__6017 ,w__6011);
  or g__6500(w__6137 ,w__6002 ,w__5943);
  or g__6501(w__6136 ,w__5942 ,w__5983);
  or g__6502(w__6135 ,w__5972 ,w__6014);
  or g__6503(w__6134 ,w__5969 ,w__5949);
  or g__6504(w__6133 ,w__6018 ,w__6005);
  or g__6505(w__6132 ,w__5971 ,w__5999);
  or g__6506(w__6131 ,w__5927 ,w__5986);
  not g__6507(w__6112 ,w__6111);
  or g__6508(w__6098 ,w__5939 ,w__6093);
  or g__6509(w__6128 ,w__5937 ,w__5914);
  or g__6510(w__6127 ,w__5936 ,w__5974);
  or g__6511(w__6126 ,w__5917 ,w__5994);
  or g__6512(w__6125 ,w__6015 ,w__6009);
  and g__6513(w__6124 ,in9[4] ,in9[2]);
  or g__6514(w__6123 ,w__5910 ,w__5977);
  or g__6515(w__6122 ,w__6002 ,w__5981);
  or g__6516(w__6121 ,w__5955 ,w__5997);
  or g__6517(w__6120 ,w__6012 ,w__5975);
  or g__6518(w__6119 ,w__5995 ,w__6071);
  or g__6519(w__6118 ,w__5940 ,w__5987);
  and g__6520(w__6117 ,in9[4] ,in9[0]);
  or g__6521(w__6116 ,w__6003 ,w__5961);
  or g__6522(w__6115 ,w__5946 ,w__5916);
  or g__6523(w__6114 ,w__6007 ,w__5980);
  or g__6524(w__6113 ,w__5924 ,w__5926);
  and g__6525(w__6111 ,in9[2] ,in9[1]);
  or g__6526(w__6110 ,w__5912 ,w__5984);
  or g__6527(w__6109 ,w__5967 ,w__5978);
  or g__6528(w__6108 ,w__6005 ,w__5949);
  or g__6529(w__6107 ,w__5920 ,w__5981);
  or g__6530(w__6106 ,w__5934 ,w__5989);
  or g__6531(w__6105 ,w__5909 ,w__5992);
  or g__6532(w__6104 ,w__5957 ,w__5930);
  or g__6533(w__6103 ,w__5922 ,w__5990);
  or g__6534(w__6102 ,w__5919 ,w__5952);
  or g__6535(w__6101 ,w__5932 ,w__5955);
  or g__6536(w__6100 ,w__6000 ,w__5966);
  or g__6537(w__6099 ,w__5959 ,w__5929);
  not g__6538(w__6097 ,w__6058);
  not g__6539(w__6096 ,w__6025);
  not g__6540(w__6095 ,w__6063);
  not g__6541(w__6094 ,w__6047);
  not g__6542(w__6093 ,w__6039);
  not g__6543(w__6092 ,w__6066);
  not g__6544(w__6091 ,w__6027);
  not g__6545(w__6090 ,w__6049);
  not g__6546(w__6089 ,in9[0]);
  not g__6547(w__6088 ,in9[4]);
  not g__6548(w__6087 ,in9[1]);
  not g__6549(w__6086 ,in9[8]);
  not g__6550(w__6085 ,in9[9]);
  not g__6551(w__6084 ,w__6033);
  not g__6552(w__6083 ,w__6061);
  not g__6553(w__6082 ,w__6051);
  not g__6554(w__6081 ,w__6069);
  not g__6555(w__6080 ,w__6029);
  not g__6556(w__6079 ,w__6056);
  not g__6557(w__6078 ,w__6053);
  not g__6558(w__6077 ,in9[3]);
  not g__6559(w__6076 ,in9[5]);
  not g__6560(w__6075 ,in9[2]);
  not g__6561(w__6074 ,in9[7]);
  not g__6562(w__6073 ,in9[6]);
  not g__6563(w__6072 ,in9[10]);
  not g__6564(w__6069 ,w__6067);
  not g__6565(w__6068 ,w__6067);
  not g__6566(w__6067 ,w__8370);
  not g__6567(w__6066 ,w__6064);
  not g__6568(w__6065 ,w__6064);
  not g__6569(w__6064 ,w__8384);
  not g__6570(w__6063 ,w__6062);
  not g__6571(w__6062 ,w__8383);
  not g__6572(w__6061 ,w__6059);
  not g__6573(w__6060 ,w__6059);
  not g__6574(w__6059 ,w__8389);
  not g__6575(w__6058 ,w__6057);
  not g__6576(w__6057 ,w__8387);
  not g__6577(w__6056 ,w__6054);
  not g__6578(w__6055 ,w__6054);
  not g__6579(w__6054 ,w__8386);
  not g__6580(w__6053 ,w__6052);
  not g__6581(w__6052 ,w__8381);
  not g__6582(w__6051 ,w__6050);
  not g__6583(w__6050 ,w__8378);
  not g__6584(w__6049 ,w__6048);
  not g__6585(w__6048 ,w__8385);
  not g__6586(w__6047 ,w__6046);
  not g__6587(w__6046 ,w__8377);
  not g__6588(w__6045 ,w__6043);
  not g__6589(w__6044 ,w__6043);
  not g__6590(w__6043 ,w__8382);
  not g__6591(w__6042 ,w__6040);
  not g__6592(w__6041 ,w__6040);
  not g__6593(w__6040 ,w__8380);
  not g__6594(w__6039 ,w__6037);
  not g__6595(w__6038 ,w__6037);
  not g__6596(w__6037 ,w__8388);
  not g__6597(w__6036 ,w__6034);
  not g__6598(w__6035 ,w__6034);
  not g__6599(w__6034 ,w__8379);
  not g__6600(w__6033 ,w__6032);
  not g__6601(w__6032 ,w__8372);
  not g__6602(w__6031 ,w__6030);
  not g__6603(w__6030 ,w__8374);
  not g__6604(w__6029 ,w__6028);
  not g__6605(w__6028 ,w__8373);
  not g__6606(w__6027 ,w__6026);
  not g__6607(w__6026 ,w__8376);
  not g__6608(w__6025 ,w__6024);
  not g__6609(w__6024 ,w__8375);
  not g__6610(w__6070 ,w__8369);
  not g__6611(w__6023 ,w__6022);
  not g__6612(w__6022 ,w__8371);
  not g__6613(w__6021 ,w__6020);
  not g__6614(w__6020 ,w__8390);
  not g__6615(w__6019 ,w__6071);
  not g__6616(w__6071 ,w__8368);
  not g__6617(w__6018 ,w__6016);
  not g__6618(w__6017 ,w__6016);
  not g__6619(w__6016 ,w__6085);
  not g__6620(w__6015 ,w__6013);
  not g__6621(w__6014 ,w__6013);
  not g__6622(w__6013 ,w__6074);
  not g__6623(w__6012 ,w__6010);
  not g__6624(w__6011 ,w__6010);
  not g__6625(w__6010 ,w__6073);
  not g__6626(w__6009 ,w__6008);
  not g__6627(w__6008 ,w__6075);
  not g__6628(w__6007 ,w__6006);
  not g__6629(w__6006 ,w__6088);
  not g__6630(w__6005 ,w__6004);
  not g__6631(w__6004 ,w__6077);
  not g__6632(w__6003 ,w__6001);
  not g__6633(w__6002 ,w__6001);
  not g__6634(w__6001 ,w__6072);
  not g__6635(w__6000 ,w__5998);
  not g__6636(w__5999 ,w__5998);
  not g__6637(w__5998 ,w__6086);
  not g__6638(w__5997 ,w__5996);
  not g__6639(w__5996 ,w__6089);
  not g__6640(w__5995 ,w__5993);
  not g__6641(w__5994 ,w__5993);
  not g__6642(w__5993 ,w__6089);
  not g__6643(w__5992 ,w__5991);
  not g__6644(w__5991 ,w__6076);
  not g__6645(w__5990 ,w__5988);
  not g__6646(w__5989 ,w__5988);
  not g__6647(w__5988 ,w__6076);
  not g__6648(w__5987 ,w__5985);
  not g__6649(w__5986 ,w__5985);
  not g__6650(w__5985 ,w__6075);
  not g__6651(w__5984 ,w__5982);
  not g__6652(w__5983 ,w__5982);
  not g__6653(w__5982 ,w__6088);
  not g__6654(w__5981 ,w__5979);
  not g__6655(w__5980 ,w__5979);
  not g__6656(w__5979 ,w__6077);
  not g__6657(w__5978 ,w__5976);
  not g__6658(w__5977 ,w__5976);
  not g__6659(w__5976 ,w__6087);
  not g__6660(w__5975 ,w__5973);
  not g__6661(w__5974 ,w__5973);
  not g__6662(w__5973 ,w__6087);
  not g__6663(w__5972 ,w__5970);
  not g__6664(w__5971 ,w__5970);
  not g__6665(w__5970 ,w__6085);
  not g__6666(w__5969 ,w__5968);
  not g__6667(w__5968 ,w__5990);
  not g__6668(w__5967 ,w__5965);
  not g__6669(w__5966 ,w__5965);
  not g__6670(w__5965 ,w__6076);
  not g__6671(w__5964 ,w__5963);
  not g__6672(w__5963 ,w__5995);
  not g__6673(w__5962 ,w__5960);
  not g__6674(w__5961 ,w__5960);
  not g__6675(w__5960 ,w__6089);
  not g__6676(w__5959 ,w__5958);
  not g__6677(w__5958 ,w__6000);
  not g__6678(w__5957 ,w__5956);
  not g__6679(w__5956 ,w__6003);
  not g__6680(w__5955 ,w__5953);
  not g__6681(w__5954 ,w__5953);
  not g__6682(w__5953 ,w__6077);
  not g__6683(w__5952 ,w__5950);
  not g__6684(w__5951 ,w__5950);
  not g__6685(w__5950 ,w__6088);
  not g__6686(w__5949 ,w__5947);
  not g__6687(w__5948 ,w__5947);
  not g__6688(w__5947 ,w__6075);
  not g__6689(w__5946 ,w__5944);
  not g__6690(w__5945 ,w__5944);
  not g__6691(w__5944 ,w__6086);
  not g__6692(w__5943 ,w__5941);
  not g__6693(w__5942 ,w__5941);
  not g__6694(w__5941 ,w__6086);
  not g__6695(w__5940 ,w__5938);
  not g__6696(w__5939 ,w__5938);
  not g__6697(w__5938 ,w__6072);
  not g__6698(w__5937 ,w__5935);
  not g__6699(w__5936 ,w__5935);
  not g__6700(w__5935 ,w__6072);
  not g__6701(w__5934 ,w__5933);
  not g__6702(w__5933 ,w__6011);
  not g__6703(w__5932 ,w__5931);
  not g__6704(w__5931 ,w__6012);
  not g__6705(w__5930 ,w__5928);
  not g__6706(w__5929 ,w__5928);
  not g__6707(w__5928 ,w__6073);
  not g__6708(w__5927 ,w__5925);
  not g__6709(w__5926 ,w__5925);
  not g__6710(w__5925 ,w__6073);
  not g__6711(w__5924 ,w__5923);
  not g__6712(w__5923 ,w__6014);
  not g__6713(w__5922 ,w__5921);
  not g__6714(w__5921 ,w__6015);
  not g__6715(w__5920 ,w__5918);
  not g__6716(w__5919 ,w__5918);
  not g__6717(w__5918 ,w__6074);
  not g__6718(w__5917 ,w__5915);
  not g__6719(w__5916 ,w__5915);
  not g__6720(w__5915 ,w__6074);
  not g__6721(w__5914 ,w__5913);
  not g__6722(w__5913 ,w__6017);
  not g__6723(w__5912 ,w__5911);
  not g__6724(w__5911 ,w__6018);
  not g__6725(w__5910 ,w__5908);
  not g__6726(w__5909 ,w__5908);
  not g__6727(w__5908 ,w__6085);
  xor g__6728(w__8365 ,w__6570 ,w__6286);
  xor g__6729(w__8364 ,w__6568 ,w__6381);
  xor g__6730(w__8363 ,w__6566 ,w__6446);
  xor g__6731(w__8362 ,w__6564 ,w__6481);
  xor g__6732(w__8361 ,w__6562 ,w__6513);
  xor g__6733(w__8360 ,w__6560 ,w__6515);
  xor g__6734(w__8359 ,w__6558 ,w__6539);
  xor g__6735(w__8358 ,w__6556 ,w__6543);
  xor g__6736(w__8357 ,w__6554 ,w__6538);
  xor g__6737(w__8356 ,w__6552 ,w__6537);
  xor g__6738(w__8355 ,w__6550 ,w__6527);
  xor g__6739(w__5907 ,w__6390 ,w__6464);
  and g__6740(w__5906 ,w__6062 ,w__6426);
  and g__6741(w__5905 ,w__6048 ,w__6331);
  and g__6742(w__5904 ,w__6052 ,w__6289);
  xor g__6743(w__5903 ,w__6148 ,w__6160);
  xnor g__6744(w__5902 ,w__6146 ,w__6117);
  and g__6745(w__5901 ,w__6057 ,w__6137);
  xor g__6746(w__5900 ,w__6124 ,w__6153);
  xor g__6747(w__5899 ,w__6399 ,w__6050);
  xor g__6748(w__5898 ,w__6366 ,w__6046);
  xor g__6749(w__5897 ,w__6302 ,w__6032);
  xor g__6750(w__5896 ,w__6223 ,w__6030);
  xor g__6751(w__8345 ,w__6119 ,w__6070);
  xnor g__6752(w__8342 ,w__7250 ,w__6699);
  and g__6753(w__8343 ,w__6699 ,w__7251);
  not g__6754(w__7251 ,w__7250);
  and g__6755(w__7250 ,w__6952 ,w__7249);
  or g__6756(w__7249 ,w__6937 ,w__7248);
  and g__6757(w__7248 ,w__7049 ,w__7247);
  or g__6758(w__7247 ,w__7048 ,w__7246);
  and g__6759(w__7246 ,w__7097 ,w__7245);
  or g__6760(w__7245 ,w__7099 ,w__7244);
  and g__6761(w__7244 ,w__7154 ,w__7243);
  or g__6762(w__7243 ,w__7146 ,w__7242);
  and g__6763(w__7242 ,w__7180 ,w__7241);
  or g__6764(w__7241 ,w__7181 ,w__7240);
  and g__6765(w__7240 ,w__7188 ,w__7239);
  or g__6766(w__7239 ,w__7187 ,w__7238);
  and g__6767(w__7238 ,w__7212 ,w__7237);
  or g__6768(w__7237 ,w__7213 ,w__7236);
  and g__6769(w__7236 ,w__7219 ,w__7235);
  or g__6770(w__7235 ,w__7218 ,w__7234);
  and g__6771(w__7234 ,w__7211 ,w__7233);
  or g__6772(w__7233 ,w__7210 ,w__7232);
  and g__6773(w__7232 ,w__7209 ,w__7231);
  or g__6774(w__7231 ,w__7208 ,w__7230);
  and g__6775(w__7230 ,w__7199 ,w__7229);
  or g__6776(w__7229 ,w__7198 ,w__7228);
  and g__6777(w__7228 ,w__7185 ,w__7227);
  xnor g__6778(w__8330 ,w__7225 ,w__7192);
  or g__6779(w__7227 ,w__7179 ,w__7226);
  not g__6780(w__7226 ,w__7225);
  or g__6781(w__7225 ,w__7160 ,w__7224);
  xnor g__6782(w__8329 ,w__7223 ,w__7177);
  and g__6783(w__7224 ,w__7167 ,w__7223);
  or g__6784(w__7223 ,w__7137 ,w__7222);
  xnor g__6785(w__8328 ,w__7220 ,w__7145);
  and g__6786(w__7222 ,w__7136 ,w__7220);
  xnor g__6787(w__7221 ,w__7201 ,w__7207);
  or g__6788(w__7220 ,w__7115 ,w__7214);
  or g__6789(w__7219 ,w__7200 ,w__7206);
  nor g__6790(w__7218 ,w__7201 ,w__7207);
  xnor g__6791(w__7217 ,w__7203 ,w__7183);
  xnor g__6792(w__7216 ,w__7171 ,w__7195);
  xnor g__6793(w__7215 ,w__7173 ,w__7197);
  xnor g__6794(w__8327 ,w__7204 ,w__7123);
  and g__6795(w__7214 ,w__7114 ,w__7204);
  nor g__6796(w__7213 ,w__7203 ,w__7183);
  or g__6797(w__7212 ,w__7202 ,w__7182);
  or g__6798(w__7211 ,w__7170 ,w__7194);
  nor g__6799(w__7210 ,w__7171 ,w__7195);
  or g__6800(w__7209 ,w__7172 ,w__7196);
  nor g__6801(w__7208 ,w__7173 ,w__7197);
  not g__6802(w__7207 ,w__7206);
  xnor g__6803(w__7206 ,w__7131 ,w__7178);
  xnor g__6804(w__7205 ,w__7184 ,w__7175);
  not g__6805(w__7202 ,w__7203);
  not g__6806(w__7200 ,w__7201);
  or g__6807(w__7199 ,w__7175 ,w__7184);
  and g__6808(w__7198 ,w__7175 ,w__7184);
  or g__6809(w__7204 ,w__7084 ,w__7189);
  or g__6810(w__7203 ,w__7169 ,w__7186);
  or g__6811(w__7201 ,w__7110 ,w__7190);
  not g__6812(w__7197 ,w__7196);
  not g__6813(w__7195 ,w__7194);
  xnor g__6814(w__8326 ,w__7176 ,w__7094);
  xnor g__6815(w__7193 ,w__7161 ,w__7174);
  xnor g__6816(w__7192 ,w__7158 ,w__7165);
  xnor g__6817(w__7191 ,w__7156 ,w__7163);
  xnor g__6818(w__7196 ,w__7103 ,w__6585);
  xnor g__6819(w__7194 ,w__7166 ,w__7122);
  and g__6820(w__7190 ,w__7098 ,w__7166);
  and g__6821(w__7189 ,w__7083 ,w__7176);
  or g__6822(w__7188 ,w__7174 ,w__7161);
  and g__6823(w__7187 ,w__7174 ,w__7161);
  nor g__6824(w__7186 ,w__7131 ,w__7168);
  or g__6825(w__7185 ,w__7157 ,w__7164);
  not g__6826(w__7182 ,w__7183);
  nor g__6827(w__7181 ,w__7156 ,w__7163);
  or g__6828(w__7180 ,w__7155 ,w__7162);
  nor g__6829(w__7179 ,w__7158 ,w__7165);
  xnor g__6830(w__7178 ,w__7149 ,w__6723);
  xnor g__6831(w__7177 ,w__7129 ,w__7148);
  xnor g__6832(w__7184 ,w__7091 ,w__7144);
  xnor g__6833(w__7183 ,w__7119 ,w__7143);
  not g__6834(w__7172 ,w__7173);
  not g__6835(w__7171 ,w__7170);
  and g__6836(w__7169 ,w__6723 ,w__7149);
  nor g__6837(w__7168 ,w__6722 ,w__7149);
  or g__6838(w__7167 ,w__7129 ,w__7148);
  or g__6839(w__7176 ,w__7082 ,w__7150);
  and g__6840(w__7175 ,w__7139 ,w__7151);
  and g__6841(w__7174 ,w__7138 ,w__7153);
  or g__6842(w__7173 ,w__7134 ,w__7152);
  and g__6843(w__7170 ,w__7133 ,w__7147);
  not g__6844(w__7164 ,w__7165);
  not g__6845(w__7162 ,w__7163);
  xnor g__6846(w__8325 ,w__7141 ,w__7093);
  and g__6847(w__7160 ,w__7129 ,w__7148);
  xnor g__6848(w__7159 ,w__7130 ,w__7140);
  xnor g__6849(w__7166 ,w__7121 ,w__6731);
  xnor g__6850(w__7165 ,w__7106 ,w__6577);
  xnor g__6851(w__7163 ,w__7125 ,w__6727);
  xnor g__6852(w__7161 ,w__7074 ,w__7120);
  not g__6853(w__7158 ,w__7157);
  not g__6854(w__7156 ,w__7155);
  or g__6855(w__7154 ,w__7140 ,w__7130);
  or g__6856(w__7153 ,w__7119 ,w__6584);
  nor g__6857(w__7152 ,w__7091 ,w__7128);
  or g__6858(w__7151 ,w__7077 ,w__7135);
  and g__6859(w__7150 ,w__7081 ,w__7141);
  and g__6860(w__7157 ,w__7118 ,w__7126);
  and g__6861(w__7155 ,w__7108 ,w__7127);
  or g__6862(w__7147 ,w__7142 ,w__7132);
  xnor g__6863(w__8324 ,w__7076 ,w__7095);
  and g__6864(w__7146 ,w__7140 ,w__7130);
  xnor g__6865(w__7145 ,w__7088 ,w__7101);
  xnor g__6866(w__7144 ,w__7100 ,w__6714);
  xnor g__6867(w__7143 ,w__7104 ,w__6741);
  xnor g__6868(w__7149 ,w__7011 ,w__7096);
  xnor g__6869(w__7148 ,w__7064 ,w__6576);
  or g__6870(w__7139 ,w__6760 ,w__7106);
  or g__6871(w__7138 ,w__6773 ,w__7104);
  and g__6872(w__7137 ,w__7088 ,w__7101);
  or g__6873(w__7136 ,w__7088 ,w__7101);
  nor g__6874(w__7135 ,w__6729 ,w__7105);
  and g__6875(w__7134 ,w__6714 ,w__7100);
  or g__6876(w__7133 ,w__7067 ,w__7103);
  nor g__6877(w__7132 ,w__7068 ,w__7102);
  and g__6878(w__7142 ,w__7078 ,w__7109);
  or g__6879(w__7141 ,w__7080 ,w__7111);
  and g__6880(w__7140 ,w__7051 ,w__7112);
  nor g__6881(w__7128 ,w__6713 ,w__7100);
  or g__6882(w__7127 ,w__7074 ,w__7113);
  or g__6883(w__7126 ,w__7044 ,w__7117);
  xnor g__6884(w__7125 ,w__7092 ,w__7009);
  xnor g__6885(w__7124 ,w__7073 ,w__7066);
  xnor g__6886(w__7123 ,w__7057 ,w__7069);
  xnor g__6887(w__7122 ,w__7062 ,w__7090);
  xnor g__6888(w__7121 ,w__7075 ,w__6967);
  xnor g__6889(w__7120 ,w__7071 ,w__6744);
  and g__6890(w__7131 ,w__7026 ,w__7107);
  xnor g__6891(w__7130 ,w__7058 ,w__6734);
  or g__6892(w__7129 ,w__7087 ,w__7116);
  or g__6893(w__7118 ,w__6772 ,w__7064);
  nor g__6894(w__7117 ,w__6725 ,w__7063);
  nor g__6895(w__7116 ,w__6994 ,w__7086);
  and g__6896(w__7115 ,w__7057 ,w__7069);
  or g__6897(w__7114 ,w__7057 ,w__7069);
  nor g__6898(w__7113 ,w__6743 ,w__7071);
  or g__6899(w__7112 ,w__6583 ,w__7092);
  and g__6900(w__7111 ,w__7076 ,w__7060);
  nor g__6901(w__7110 ,w__7062 ,w__7089);
  or g__6902(w__7109 ,w__6995 ,w__7079);
  or g__6903(w__7108 ,w__6770 ,w__7070);
  or g__6904(w__7107 ,w__6582 ,w__7075);
  and g__6905(w__7119 ,w__7047 ,w__7085);
  not g__6906(w__7105 ,w__7106);
  not g__6907(w__7102 ,w__7103);
  nor g__6908(w__7099 ,w__7073 ,w__7066);
  or g__6909(w__7098 ,w__7061 ,w__7090);
  or g__6910(w__7097 ,w__7072 ,w__7065);
  xnor g__6911(w__7096 ,w__6970 ,w__7043);
  xnor g__6912(w__7095 ,w__6884 ,w__6575);
  xnor g__6913(w__7094 ,w__6990 ,w__7041);
  xnor g__6914(w__7093 ,w__6993 ,w__7039);
  xnor g__6915(w__7106 ,w__7014 ,w__7032);
  xnor g__6916(w__7104 ,w__7029 ,w__7035);
  xnor g__6917(w__7103 ,w__7030 ,w__7033);
  xnor g__6918(w__7101 ,w__7038 ,w__7034);
  xnor g__6919(w__7100 ,w__7040 ,w__7031);
  not g__6920(w__7089 ,w__7090);
  nor g__6921(w__7087 ,w__6769 ,w__7038);
  and g__6922(w__7086 ,w__6769 ,w__7038);
  or g__6923(w__7085 ,w__7043 ,w__7045);
  and g__6924(w__7084 ,w__6990 ,w__7041);
  or g__6925(w__7083 ,w__6990 ,w__7041);
  and g__6926(w__7082 ,w__6993 ,w__7039);
  or g__6927(w__7081 ,w__6993 ,w__7039);
  nor g__6928(w__7080 ,w__6884 ,w__6575);
  and g__6929(w__7079 ,w__6972 ,w__7040);
  or g__6930(w__7078 ,w__6972 ,w__7040);
  and g__6931(w__7092 ,w__7016 ,w__7052);
  and g__6932(w__7091 ,w__7018 ,w__7046);
  or g__6933(w__7090 ,w__7022 ,w__7050);
  or g__6934(w__7088 ,w__6989 ,w__7053);
  not g__6935(w__7072 ,w__7073);
  not g__6936(w__7070 ,w__7071);
  not g__6937(w__7067 ,w__7068);
  not g__6938(w__7066 ,w__7065);
  not g__6939(w__7063 ,w__7064);
  not g__6940(w__7061 ,w__7062);
  or g__6941(w__7060 ,w__6883 ,w__7042);
  xnor g__6942(w__8323 ,w__7028 ,w__6961);
  xnor g__6943(w__7059 ,w__6978 ,w__7027);
  xnor g__6944(w__7058 ,w__7013 ,w__6975);
  and g__6945(w__7077 ,w__7007 ,w__7037);
  or g__6946(w__7076 ,w__6935 ,w__7036);
  and g__6947(w__7075 ,w__7003 ,w__7055);
  and g__6948(w__7074 ,w__7024 ,w__7054);
  xnor g__6949(w__7073 ,w__6999 ,w__6736);
  xnor g__6950(w__7071 ,w__6976 ,w__6998);
  xnor g__6951(w__7069 ,w__7012 ,w__6997);
  xnor g__6952(w__7068 ,w__6966 ,w__7000);
  and g__6953(w__7065 ,w__7015 ,w__7056);
  xnor g__6954(w__7064 ,w__6968 ,w__7002);
  xnor g__6955(w__7062 ,w__6943 ,w__7001);
  or g__6956(w__7056 ,w__7013 ,w__7021);
  or g__6957(w__7055 ,w__6957 ,w__7025);
  or g__6958(w__7054 ,w__7029 ,w__7017);
  nor g__6959(w__7053 ,w__6988 ,w__7012);
  or g__6960(w__7052 ,w__6942 ,w__7008);
  or g__6961(w__7051 ,w__6768 ,w__7009);
  nor g__6962(w__7050 ,w__7020 ,w__7030);
  or g__6963(w__7049 ,w__7027 ,w__6978);
  and g__6964(w__7048 ,w__7027 ,w__6978);
  or g__6965(w__7047 ,w__6969 ,w__7011);
  or g__6966(w__7046 ,w__7023 ,w__7014);
  nor g__6967(w__7045 ,w__6970 ,w__7010);
  or g__6968(w__7057 ,w__6938 ,w__7005);
  not g__6969(w__7042 ,w__6575);
  or g__6970(w__7037 ,w__6941 ,w__7006);
  nor g__6971(w__7036 ,w__6949 ,w__7028);
  xor g__6972(w__8322 ,w__6878 ,w__6960);
  xnor g__6973(w__7035 ,w__6973 ,w__6955);
  xnor g__6974(w__7034 ,w__6994 ,w__6705);
  xnor g__6975(w__7033 ,w__6992 ,w__6720);
  xnor g__6976(w__7032 ,w__6971 ,w__6991);
  xor g__6977(w__7031 ,w__6972 ,w__6995);
  and g__6978(w__7044 ,w__6936 ,w__7004);
  and g__6979(w__7043 ,w__6982 ,w__7019);
  xnor g__6980(w__7041 ,w__6996 ,w__6574);
  xnor g__6981(w__7040 ,w__6959 ,w__6963);
  xnor g__6982(w__7039 ,w__6962 ,w__6707);
  xnor g__6983(w__7038 ,w__6979 ,w__6965);
  or g__6984(w__7026 ,w__6756 ,w__6967);
  and g__6985(w__7025 ,w__6861 ,w__6966);
  or g__6986(w__7024 ,w__6955 ,w__6973);
  and g__6987(w__7023 ,w__6991 ,w__6971);
  and g__6988(w__7022 ,w__6720 ,w__6992);
  nor g__6989(w__7021 ,w__6733 ,w__6975);
  nor g__6990(w__7020 ,w__6719 ,w__6992);
  or g__6991(w__7019 ,w__6943 ,w__6986);
  or g__6992(w__7018 ,w__6991 ,w__6971);
  and g__6993(w__7017 ,w__6955 ,w__6973);
  or g__6994(w__7016 ,w__6793 ,w__6977);
  or g__6995(w__7015 ,w__6757 ,w__6974);
  and g__6996(w__7030 ,w__6947 ,w__6985);
  and g__6997(w__7029 ,w__6850 ,w__6987);
  and g__6998(w__7028 ,w__6951 ,w__6983);
  and g__6999(w__7027 ,w__6875 ,w__6984);
  not g__7000(w__7010 ,w__7011);
  and g__7001(w__7008 ,w__6793 ,w__6977);
  or g__7002(w__7007 ,w__6877 ,w__6968);
  and g__7003(w__7006 ,w__6877 ,w__6968);
  and g__7004(w__7005 ,w__6933 ,w__6996);
  or g__7005(w__7004 ,w__6939 ,w__6979);
  or g__7006(w__7003 ,w__6861 ,w__6966);
  xnor g__7007(w__7002 ,w__6877 ,w__6941);
  xnor g__7008(w__7001 ,w__6814 ,w__6940);
  xor g__7009(w__7000 ,w__6861 ,w__6957);
  xnor g__7010(w__6999 ,w__6958 ,w__6815);
  xnor g__7011(w__6998 ,w__6793 ,w__6942);
  xnor g__7012(w__6997 ,w__6954 ,w__6703);
  xnor g__7013(w__7014 ,w__6905 ,w__6931);
  and g__7014(w__7013 ,w__6841 ,w__6981);
  xnor g__7015(w__7012 ,w__6578 ,w__6930);
  xnor g__7016(w__7011 ,w__6956 ,w__6888);
  xnor g__7017(w__7009 ,w__6944 ,w__6892);
  nor g__7018(w__6989 ,w__6774 ,w__6954);
  and g__7019(w__6988 ,w__6774 ,w__6954);
  or g__7020(w__6987 ,w__6845 ,w__6956);
  and g__7021(w__6986 ,w__6814 ,w__6940);
  or g__7022(w__6985 ,w__6959 ,w__6953);
  or g__7023(w__6984 ,w__6579 ,w__6958);
  or g__7024(w__6983 ,w__6878 ,w__6948);
  or g__7025(w__6982 ,w__6814 ,w__6940);
  or g__7026(w__6981 ,w__6871 ,w__6944);
  xnor g__7027(w__6980 ,w__6790 ,w__6904);
  xnor g__7028(w__6996 ,w__6862 ,w__6887);
  and g__7029(w__6995 ,w__6913 ,w__6932);
  and g__7030(w__6994 ,w__6920 ,w__6945);
  or g__7031(w__6993 ,w__6866 ,w__6946);
  xnor g__7032(w__6992 ,w__6780 ,w__6908);
  and g__7033(w__6991 ,w__6855 ,w__6934);
  or g__7034(w__6990 ,w__6924 ,w__6950);
  not g__7035(w__6977 ,w__6976);
  not g__7036(w__6974 ,w__6975);
  not g__7037(w__6969 ,w__6970);
  xnor g__7038(w__6965 ,w__6860 ,w__6903);
  xnor g__7039(w__6964 ,w__6927 ,w__6739);
  xnor g__7040(w__6963 ,w__6882 ,w__6898);
  xnor g__7041(w__6962 ,w__6580 ,w__6880);
  xnor g__7042(w__6961 ,w__6881 ,w__6928);
  xnor g__7043(w__6960 ,w__6900 ,w__6747);
  xnor g__7044(w__6979 ,w__6792 ,w__6889);
  xnor g__7045(w__6978 ,w__6907 ,w__6717);
  xnor g__7046(w__6976 ,w__6816 ,w__6894);
  xnor g__7047(w__6975 ,w__6810 ,w__6891);
  xnor g__7048(w__6973 ,w__6783 ,w__6885);
  xnor g__7049(w__6972 ,w__6785 ,w__6886);
  xnor g__7050(w__6971 ,w__6820 ,w__6897);
  xnor g__7051(w__6970 ,w__6778 ,w__6895);
  xnor g__7052(w__6968 ,w__6581 ,w__6890);
  xnor g__7053(w__6967 ,w__6811 ,w__6893);
  xnor g__7054(w__6966 ,w__6830 ,w__6896);
  and g__7055(w__6953 ,w__6882 ,w__6898);
  or g__7056(w__6952 ,w__6761 ,w__6926);
  or g__7057(w__6951 ,w__6759 ,w__6899);
  nor g__7058(w__6950 ,w__6914 ,w__6580);
  and g__7059(w__6949 ,w__6881 ,w__6929);
  nor g__7060(w__6948 ,w__6746 ,w__6900);
  or g__7061(w__6947 ,w__6882 ,w__6898);
  and g__7062(w__6946 ,w__6873 ,w__6904);
  or g__7063(w__6945 ,w__6922 ,w__6578);
  and g__7064(w__6959 ,w__6854 ,w__6916);
  and g__7065(w__6958 ,w__6870 ,w__6909);
  and g__7066(w__6957 ,w__6842 ,w__6923);
  and g__7067(w__6956 ,w__6872 ,w__6915);
  and g__7068(w__6955 ,w__6876 ,w__6921);
  and g__7069(w__6954 ,w__6848 ,w__6919);
  nor g__7070(w__6939 ,w__6860 ,w__6903);
  and g__7071(w__6938 ,w__6709 ,w__6901);
  nor g__7072(w__6937 ,w__6738 ,w__6927);
  or g__7073(w__6936 ,w__6859 ,w__6902);
  nor g__7074(w__6935 ,w__6881 ,w__6929);
  or g__7075(w__6934 ,w__6844 ,w__6581);
  or g__7076(w__6933 ,w__6709 ,w__6901);
  or g__7077(w__6932 ,w__6906 ,w__6925);
  xnor g__7078(w__6931 ,w__6823 ,w__6858);
  xnor g__7079(w__6930 ,w__6787 ,w__6879);
  and g__7080(w__6944 ,w__6865 ,w__6918);
  and g__7081(w__6943 ,w__6843 ,w__6911);
  and g__7082(w__6942 ,w__6852 ,w__6917);
  and g__7083(w__6941 ,w__6856 ,w__6910);
  and g__7084(w__6940 ,w__6868 ,w__6912);
  not g__7085(w__6929 ,w__6928);
  not g__7086(w__6927 ,w__6926);
  nor g__7087(w__6925 ,w__6822 ,w__6858);
  nor g__7088(w__6924 ,w__6758 ,w__6880);
  or g__7089(w__6923 ,w__6801 ,w__6849);
  and g__7090(w__6922 ,w__6787 ,w__6879);
  or g__7091(w__6921 ,w__6800 ,w__6864);
  or g__7092(w__6920 ,w__6787 ,w__6879);
  or g__7093(w__6918 ,w__6827 ,w__6863);
  or g__7094(w__6917 ,w__6828 ,w__6846);
  or g__7095(w__6916 ,w__6803 ,w__6853);
  or g__7096(w__6915 ,w__6796 ,w__6851);
  and g__7097(w__6914 ,w__6758 ,w__6880);
  or g__7098(w__6913 ,w__6823 ,w__6857);
  or g__7099(w__6912 ,w__6805 ,w__6869);
  or g__7100(w__6911 ,w__6830 ,w__6840);
  or g__7101(w__6910 ,w__6798 ,w__6847);
  or g__7102(w__6909 ,w__6829 ,w__6867);
  xnor g__7103(w__6908 ,w__6805 ,in12[6]);
  xnor g__7104(w__6907 ,w__6806 ,in12[10]);
  xnor g__7105(w__6928 ,w__6834 ,w__6701);
  and g__7106(w__6926 ,w__6776 ,w__6874);
  not g__7107(w__6906 ,w__6905);
  not g__7108(w__6902 ,w__6903);
  not g__7109(w__6899 ,w__6900);
  xnor g__7110(w__6897 ,w__6779 ,w__6803);
  xnor g__7111(w__6896 ,w__6784 ,w__6818);
  xnor g__7112(w__6895 ,w__6800 ,in12[7]);
  xnor g__7113(w__6894 ,w__6827 ,in12[8]);
  xnor g__7114(w__6893 ,w__6781 ,w__6796);
  xnor g__7115(w__6892 ,w__6813 ,w__6782);
  xnor g__7116(w__6891 ,w__6829 ,in12[9]);
  xnor g__7117(w__6890 ,w__6809 ,w__6821);
  xnor g__7118(w__6889 ,w__6812 ,w__6798);
  xnor g__7119(w__6888 ,w__6791 ,w__6788);
  xnor g__7120(w__6887 ,w__6786 ,w__6819);
  xnor g__7121(w__6886 ,w__6817 ,w__6801);
  xnor g__7122(w__6885 ,w__6777 ,w__6828);
  xnor g__7123(w__6905 ,w__6836 ,in12[5]);
  xnor g__7124(w__6904 ,w__6799 ,in12[2]);
  xnor g__7125(w__6903 ,w__6804 ,in12[4]);
  xnor g__7126(w__6901 ,w__6833 ,in12[3]);
  xnor g__7127(w__6900 ,w__6825 ,in12[1]);
  xnor g__7128(w__6898 ,w__6837 ,w__6794);
  not g__7129(w__6884 ,w__6883);
  or g__7130(w__6876 ,w__6598 ,w__6778);
  or g__7131(w__6875 ,w__6775 ,w__6815);
  or g__7132(w__6874 ,w__6806 ,w__6807);
  or g__7133(w__6873 ,w__6711 ,w__6789);
  or g__7134(w__6872 ,w__6781 ,w__6811);
  and g__7135(w__6871 ,w__6813 ,w__6782);
  or g__7136(w__6870 ,w__6588 ,w__6810);
  and g__7137(w__6869 ,w__6608 ,w__6780);
  or g__7138(w__6868 ,w__6612 ,w__6780);
  and g__7139(w__6867 ,w__6592 ,w__6810);
  nor g__7140(w__6866 ,w__6762 ,w__6790);
  or g__7141(w__6865 ,w__6637 ,w__6816);
  and g__7142(w__6864 ,w__6602 ,w__6778);
  and g__7143(w__6863 ,w__6624 ,w__6816);
  and g__7144(w__6883 ,w__6701 ,w__6835);
  or g__7145(w__6882 ,w__6645 ,w__6836);
  or g__7146(w__6881 ,w__6655 ,w__6825);
  or g__7147(w__6880 ,w__6664 ,w__6799);
  or g__7148(w__6879 ,w__6658 ,w__6833);
  or g__7149(w__6878 ,w__6748 ,w__6797);
  or g__7150(w__6877 ,w__6661 ,w__6804);
  not g__7151(w__6859 ,w__6860);
  not g__7152(w__6857 ,w__6858);
  and g__7153(w__8320 ,w__6797 ,w__6808);
  or g__7154(w__6856 ,w__6792 ,w__6812);
  or g__7155(w__6855 ,w__6809 ,w__6821);
  or g__7156(w__6854 ,w__6820 ,w__6779);
  and g__7157(w__6853 ,w__6820 ,w__6779);
  or g__7158(w__6852 ,w__6777 ,w__6783);
  and g__7159(w__6851 ,w__6781 ,w__6811);
  or g__7160(w__6850 ,w__6791 ,w__6788);
  and g__7161(w__6849 ,w__6785 ,w__6817);
  or g__7162(w__6848 ,w__6786 ,w__6819);
  and g__7163(w__6847 ,w__6792 ,w__6812);
  and g__7164(w__6846 ,w__6777 ,w__6783);
  and g__7165(w__6845 ,w__6791 ,w__6788);
  and g__7166(w__6844 ,w__6809 ,w__6821);
  or g__7167(w__6843 ,w__6784 ,w__6818);
  or g__7168(w__6842 ,w__6785 ,w__6817);
  or g__7169(w__6841 ,w__6813 ,w__6782);
  and g__7170(w__6840 ,w__6784 ,w__6818);
  and g__7171(w__6862 ,w__6824 ,w__6795);
  or g__7172(w__6861 ,w__6837 ,w__6794);
  and g__7173(w__6860 ,w__6802 ,w__6832);
  and g__7174(w__6858 ,w__6826 ,w__6839);
  not g__7175(w__6839 ,w__6838);
  not g__7176(w__6835 ,w__6834);
  not g__7177(w__6832 ,w__6831);
  not g__7178(w__6823 ,w__6822);
  or g__7179(w__6808 ,in12[0] ,w__6697);
  nor g__7180(w__6807 ,in12[10] ,w__6716);
  or g__7181(w__6838 ,w__6621 ,w__6640);
  or g__7182(w__6837 ,w__6610 ,w__6629);
  or g__7183(w__6836 ,w__6590 ,w__6642);
  or g__7184(w__6834 ,w__6626 ,w__6672);
  or g__7185(w__6833 ,w__6647 ,w__6675);
  or g__7186(w__6831 ,w__6605 ,w__6642);
  or g__7187(w__6830 ,w__6650 ,w__6687);
  or g__7188(w__6829 ,w__6635 ,w__6600);
  or g__7189(w__6828 ,w__6618 ,w__6685);
  or g__7190(w__6827 ,w__6615 ,w__6667);
  and g__7191(w__6826 ,in12[5] ,in12[3]);
  or g__7192(w__6825 ,w__6652 ,w__6640);
  and g__7193(w__6824 ,in12[3] ,in12[1]);
  and g__7194(w__6822 ,in12[8] ,in12[1]);
  or g__7195(w__6821 ,w__6595 ,w__6653);
  or g__7196(w__6820 ,w__6670 ,w__6662);
  or g__7197(w__6819 ,w__6630 ,w__6656);
  or g__7198(w__6818 ,w__6677 ,w__6632);
  or g__7199(w__6817 ,w__6623 ,w__6665);
  or g__7200(w__6816 ,w__6695 ,w__6689);
  or g__7201(w__6815 ,w__6680 ,w__6621);
  or g__7202(w__6814 ,w__6620 ,w__6661);
  or g__7203(w__6813 ,w__6650 ,w__6692);
  or g__7204(w__6812 ,w__6647 ,w__6627);
  or g__7205(w__6811 ,w__6696 ,w__6683);
  or g__7206(w__6810 ,w__6649 ,w__6677);
  or g__7207(w__6809 ,w__6605 ,w__6664);
  not g__7208(w__6790 ,w__6789);
  or g__7209(w__6776 ,w__6617 ,w__6771);
  or g__7210(w__6806 ,w__6615 ,w__6592);
  or g__7211(w__6805 ,w__6614 ,w__6652);
  or g__7212(w__6804 ,w__6595 ,w__6672);
  or g__7213(w__6803 ,w__6693 ,w__6687);
  and g__7214(w__6802 ,in12[4] ,in12[2]);
  or g__7215(w__6801 ,w__6588 ,w__6655);
  or g__7216(w__6800 ,w__6680 ,w__6659);
  or g__7217(w__6799 ,w__6633 ,w__6675);
  or g__7218(w__6798 ,w__6690 ,w__6653);
  or g__7219(w__6797 ,w__6673 ,w__6749);
  or g__7220(w__6796 ,w__6618 ,w__6665);
  and g__7221(w__6795 ,in12[4] ,in12[0]);
  or g__7222(w__6794 ,w__6681 ,w__6639);
  or g__7223(w__6793 ,w__6624 ,w__6594);
  or g__7224(w__6792 ,w__6685 ,w__6658);
  or g__7225(w__6791 ,w__6602 ,w__6604);
  and g__7226(w__6789 ,in12[2] ,in12[1]);
  or g__7227(w__6788 ,w__6590 ,w__6662);
  or g__7228(w__6787 ,w__6645 ,w__6656);
  or g__7229(w__6786 ,w__6683 ,w__6627);
  or g__7230(w__6785 ,w__6598 ,w__6659);
  or g__7231(w__6784 ,w__6612 ,w__6667);
  or g__7232(w__6783 ,w__6587 ,w__6670);
  or g__7233(w__6782 ,w__6635 ,w__6608);
  or g__7234(w__6781 ,w__6600 ,w__6668);
  or g__7235(w__6780 ,w__6597 ,w__6630);
  or g__7236(w__6779 ,w__6610 ,w__6633);
  or g__7237(w__6778 ,w__6678 ,w__6644);
  or g__7238(w__6777 ,w__6637 ,w__6607);
  not g__7239(w__6775 ,w__6736);
  not g__7240(w__6774 ,w__6703);
  not g__7241(w__6773 ,w__6741);
  not g__7242(w__6772 ,w__6725);
  not g__7243(w__6771 ,w__6717);
  not g__7244(w__6770 ,w__6744);
  not g__7245(w__6769 ,w__6705);
  not g__7246(w__6768 ,w__6727);
  not g__7247(w__6767 ,in12[0]);
  not g__7248(w__6766 ,in12[4]);
  not g__7249(w__6765 ,in12[1]);
  not g__7250(w__6764 ,in12[8]);
  not g__7251(w__6763 ,in12[9]);
  not g__7252(w__6762 ,w__6711);
  not g__7253(w__6761 ,w__6739);
  not g__7254(w__6760 ,w__6729);
  not g__7255(w__6759 ,w__6747);
  not g__7256(w__6758 ,w__6707);
  not g__7257(w__6757 ,w__6734);
  not g__7258(w__6756 ,w__6731);
  not g__7259(w__6755 ,in12[3]);
  not g__7260(w__6754 ,in12[5]);
  not g__7261(w__6753 ,in12[2]);
  not g__7262(w__6752 ,in12[7]);
  not g__7263(w__6751 ,in12[6]);
  not g__7264(w__6750 ,in12[10]);
  not g__7265(w__6747 ,w__6745);
  not g__7266(w__6746 ,w__6745);
  not g__7267(w__6745 ,w__8370);
  not g__7268(w__6744 ,w__6742);
  not g__7269(w__6743 ,w__6742);
  not g__7270(w__6742 ,w__8384);
  not g__7271(w__6741 ,w__6740);
  not g__7272(w__6740 ,w__8383);
  not g__7273(w__6739 ,w__6737);
  not g__7274(w__6738 ,w__6737);
  not g__7275(w__6737 ,w__8389);
  not g__7276(w__6736 ,w__6735);
  not g__7277(w__6735 ,w__8387);
  not g__7278(w__6734 ,w__6732);
  not g__7279(w__6733 ,w__6732);
  not g__7280(w__6732 ,w__8386);
  not g__7281(w__6731 ,w__6730);
  not g__7282(w__6730 ,w__8381);
  not g__7283(w__6729 ,w__6728);
  not g__7284(w__6728 ,w__8378);
  not g__7285(w__6727 ,w__6726);
  not g__7286(w__6726 ,w__8385);
  not g__7287(w__6725 ,w__6724);
  not g__7288(w__6724 ,w__8377);
  not g__7289(w__6723 ,w__6721);
  not g__7290(w__6722 ,w__6721);
  not g__7291(w__6721 ,w__8382);
  not g__7292(w__6720 ,w__6718);
  not g__7293(w__6719 ,w__6718);
  not g__7294(w__6718 ,w__8380);
  not g__7295(w__6717 ,w__6715);
  not g__7296(w__6716 ,w__6715);
  not g__7297(w__6715 ,w__8388);
  not g__7298(w__6714 ,w__6712);
  not g__7299(w__6713 ,w__6712);
  not g__7300(w__6712 ,w__8379);
  not g__7301(w__6711 ,w__6710);
  not g__7302(w__6710 ,w__8372);
  not g__7303(w__6709 ,w__6708);
  not g__7304(w__6708 ,w__8374);
  not g__7305(w__6707 ,w__6706);
  not g__7306(w__6706 ,w__8373);
  not g__7307(w__6705 ,w__6704);
  not g__7308(w__6704 ,w__8376);
  not g__7309(w__6703 ,w__6702);
  not g__7310(w__6702 ,w__8375);
  not g__7311(w__6748 ,w__8369);
  not g__7312(w__6701 ,w__6700);
  not g__7313(w__6700 ,w__8371);
  not g__7314(w__6699 ,w__6698);
  not g__7315(w__6698 ,w__8390);
  not g__7316(w__6697 ,w__6749);
  not g__7317(w__6749 ,w__8368);
  not g__7318(w__6696 ,w__6694);
  not g__7319(w__6695 ,w__6694);
  not g__7320(w__6694 ,w__6763);
  not g__7321(w__6693 ,w__6691);
  not g__7322(w__6692 ,w__6691);
  not g__7323(w__6691 ,w__6752);
  not g__7324(w__6690 ,w__6688);
  not g__7325(w__6689 ,w__6688);
  not g__7326(w__6688 ,w__6751);
  not g__7327(w__6687 ,w__6686);
  not g__7328(w__6686 ,w__6753);
  not g__7329(w__6685 ,w__6684);
  not g__7330(w__6684 ,w__6766);
  not g__7331(w__6683 ,w__6682);
  not g__7332(w__6682 ,w__6755);
  not g__7333(w__6681 ,w__6679);
  not g__7334(w__6680 ,w__6679);
  not g__7335(w__6679 ,w__6750);
  not g__7336(w__6678 ,w__6676);
  not g__7337(w__6677 ,w__6676);
  not g__7338(w__6676 ,w__6764);
  not g__7339(w__6675 ,w__6674);
  not g__7340(w__6674 ,w__6767);
  not g__7341(w__6673 ,w__6671);
  not g__7342(w__6672 ,w__6671);
  not g__7343(w__6671 ,w__6767);
  not g__7344(w__6670 ,w__6669);
  not g__7345(w__6669 ,w__6754);
  not g__7346(w__6668 ,w__6666);
  not g__7347(w__6667 ,w__6666);
  not g__7348(w__6666 ,w__6754);
  not g__7349(w__6665 ,w__6663);
  not g__7350(w__6664 ,w__6663);
  not g__7351(w__6663 ,w__6753);
  not g__7352(w__6662 ,w__6660);
  not g__7353(w__6661 ,w__6660);
  not g__7354(w__6660 ,w__6766);
  not g__7355(w__6659 ,w__6657);
  not g__7356(w__6658 ,w__6657);
  not g__7357(w__6657 ,w__6755);
  not g__7358(w__6656 ,w__6654);
  not g__7359(w__6655 ,w__6654);
  not g__7360(w__6654 ,w__6765);
  not g__7361(w__6653 ,w__6651);
  not g__7362(w__6652 ,w__6651);
  not g__7363(w__6651 ,w__6765);
  not g__7364(w__6650 ,w__6648);
  not g__7365(w__6649 ,w__6648);
  not g__7366(w__6648 ,w__6763);
  not g__7367(w__6647 ,w__6646);
  not g__7368(w__6646 ,w__6668);
  not g__7369(w__6645 ,w__6643);
  not g__7370(w__6644 ,w__6643);
  not g__7371(w__6643 ,w__6754);
  not g__7372(w__6642 ,w__6641);
  not g__7373(w__6641 ,w__6673);
  not g__7374(w__6640 ,w__6638);
  not g__7375(w__6639 ,w__6638);
  not g__7376(w__6638 ,w__6767);
  not g__7377(w__6637 ,w__6636);
  not g__7378(w__6636 ,w__6678);
  not g__7379(w__6635 ,w__6634);
  not g__7380(w__6634 ,w__6681);
  not g__7381(w__6633 ,w__6631);
  not g__7382(w__6632 ,w__6631);
  not g__7383(w__6631 ,w__6755);
  not g__7384(w__6630 ,w__6628);
  not g__7385(w__6629 ,w__6628);
  not g__7386(w__6628 ,w__6766);
  not g__7387(w__6627 ,w__6625);
  not g__7388(w__6626 ,w__6625);
  not g__7389(w__6625 ,w__6753);
  not g__7390(w__6624 ,w__6622);
  not g__7391(w__6623 ,w__6622);
  not g__7392(w__6622 ,w__6764);
  not g__7393(w__6621 ,w__6619);
  not g__7394(w__6620 ,w__6619);
  not g__7395(w__6619 ,w__6764);
  not g__7396(w__6618 ,w__6616);
  not g__7397(w__6617 ,w__6616);
  not g__7398(w__6616 ,w__6750);
  not g__7399(w__6615 ,w__6613);
  not g__7400(w__6614 ,w__6613);
  not g__7401(w__6613 ,w__6750);
  not g__7402(w__6612 ,w__6611);
  not g__7403(w__6611 ,w__6689);
  not g__7404(w__6610 ,w__6609);
  not g__7405(w__6609 ,w__6690);
  not g__7406(w__6608 ,w__6606);
  not g__7407(w__6607 ,w__6606);
  not g__7408(w__6606 ,w__6751);
  not g__7409(w__6605 ,w__6603);
  not g__7410(w__6604 ,w__6603);
  not g__7411(w__6603 ,w__6751);
  not g__7412(w__6602 ,w__6601);
  not g__7413(w__6601 ,w__6692);
  not g__7414(w__6600 ,w__6599);
  not g__7415(w__6599 ,w__6693);
  not g__7416(w__6598 ,w__6596);
  not g__7417(w__6597 ,w__6596);
  not g__7418(w__6596 ,w__6752);
  not g__7419(w__6595 ,w__6593);
  not g__7420(w__6594 ,w__6593);
  not g__7421(w__6593 ,w__6752);
  not g__7422(w__6592 ,w__6591);
  not g__7423(w__6591 ,w__6695);
  not g__7424(w__6590 ,w__6589);
  not g__7425(w__6589 ,w__6696);
  not g__7426(w__6588 ,w__6586);
  not g__7427(w__6587 ,w__6586);
  not g__7428(w__6586 ,w__6763);
  xor g__7429(w__8341 ,w__7248 ,w__6964);
  xor g__7430(w__8340 ,w__7246 ,w__7059);
  xor g__7431(w__8339 ,w__7244 ,w__7124);
  xor g__7432(w__8338 ,w__7242 ,w__7159);
  xor g__7433(w__8337 ,w__7240 ,w__7191);
  xor g__7434(w__8336 ,w__7238 ,w__7193);
  xor g__7435(w__8335 ,w__7236 ,w__7217);
  xor g__7436(w__8334 ,w__7234 ,w__7221);
  xor g__7437(w__8333 ,w__7232 ,w__7216);
  xor g__7438(w__8332 ,w__7230 ,w__7215);
  xor g__7439(w__8331 ,w__7228 ,w__7205);
  xor g__7440(w__6585 ,w__7068 ,w__7142);
  and g__7441(w__6584 ,w__6740 ,w__7104);
  and g__7442(w__6583 ,w__6726 ,w__7009);
  and g__7443(w__6582 ,w__6730 ,w__6967);
  xor g__7444(w__6581 ,w__6826 ,w__6838);
  xnor g__7445(w__6580 ,w__6824 ,w__6795);
  and g__7446(w__6579 ,w__6735 ,w__6815);
  xor g__7447(w__6578 ,w__6802 ,w__6831);
  xor g__7448(w__6577 ,w__7077 ,w__6728);
  xor g__7449(w__6576 ,w__7044 ,w__6724);
  xor g__7450(w__6575 ,w__6980 ,w__6710);
  xor g__7451(w__6574 ,w__6901 ,w__6708);
  xor g__7452(w__8321 ,w__6797 ,w__6748);
  or g__7453(out1 ,w__7359 ,w__7429);
  nor g__7454(w__7429 ,w__7346 ,w__7428);
  or g__7455(w__7428 ,w__7375 ,w__7427);
  nor g__7456(w__7427 ,w__7350 ,w__7426);
  nor g__7457(w__7426 ,w__7374 ,w__7425);
  nor g__7458(w__7425 ,w__7369 ,w__7424);
  nor g__7459(w__7424 ,w__7365 ,w__7423);
  nor g__7460(w__7423 ,w__7355 ,w__7422);
  nor g__7461(w__7422 ,w__7341 ,w__7421);
  nor g__7462(w__7421 ,w__7360 ,w__7420);
  nor g__7463(w__7420 ,w__7380 ,w__7419);
  nor g__7464(w__7419 ,w__7371 ,w__7418);
  nor g__7465(w__7418 ,w__7368 ,w__7417);
  nor g__7466(w__7417 ,w__7363 ,w__7416);
  nor g__7467(w__7416 ,w__7362 ,w__7415);
  nor g__7468(w__7415 ,w__7357 ,w__7414);
  nor g__7469(w__7414 ,w__7354 ,w__7413);
  nor g__7470(w__7413 ,w__7344 ,w__7412);
  nor g__7471(w__7412 ,w__7343 ,w__7411);
  nor g__7472(w__7411 ,w__7348 ,w__7410);
  nor g__7473(w__7410 ,w__7340 ,w__7409);
  nor g__7474(w__7409 ,w__7342 ,w__7408);
  nor g__7475(w__7408 ,w__7376 ,w__7407);
  nor g__7476(w__7407 ,w__7373 ,w__7406);
  nor g__7477(w__7406 ,w__7381 ,w__7405);
  nor g__7478(w__7405 ,w__7367 ,w__7404);
  nor g__7479(w__7404 ,w__7366 ,w__7403);
  nor g__7480(w__7403 ,w__7364 ,w__7402);
  nor g__7481(w__7402 ,w__7372 ,w__7401);
  nor g__7482(w__7401 ,w__7361 ,w__7400);
  nor g__7483(w__7400 ,w__7338 ,w__7399);
  nor g__7484(w__7399 ,w__7358 ,w__7398);
  nor g__7485(w__7398 ,w__7356 ,w__7397);
  nor g__7486(w__7397 ,w__7353 ,w__7396);
  nor g__7487(w__7396 ,w__7351 ,w__7395);
  nor g__7488(w__7395 ,w__7347 ,w__7394);
  nor g__7489(w__7394 ,w__7349 ,w__7393);
  nor g__7490(w__7393 ,w__7377 ,w__7392);
  nor g__7491(w__7392 ,w__7345 ,w__7391);
  nor g__7492(w__7391 ,w__7339 ,w__7390);
  nor g__7493(w__7390 ,w__7378 ,w__7389);
  nor g__7494(w__7389 ,w__7352 ,w__7388);
  nor g__7495(w__7388 ,w__7370 ,w__7387);
  nor g__7496(w__7387 ,w__7379 ,w__7386);
  nor g__7497(w__7386 ,w__7384 ,w__7385);
  nor g__7498(w__7385 ,w__8440 ,w__7383);
  and g__7499(w__7384 ,w__7264 ,w__7382);
  nor g__7500(w__7383 ,w__7264 ,w__7382);
  nor g__7501(w__7381 ,w__7310 ,w__7270);
  nor g__7502(w__7380 ,w__7314 ,w__7290);
  nor g__7503(w__7379 ,w__7302 ,w__7297);
  nor g__7504(w__7378 ,w__7336 ,w__7253);
  nor g__7505(w__7377 ,w__7333 ,w__7261);
  nor g__7506(w__7376 ,w__7330 ,w__7269);
  nor g__7507(w__7375 ,w__7332 ,w__7255);
  nor g__7508(w__7374 ,w__7328 ,w__7286);
  nor g__7509(w__7373 ,w__7305 ,w__7283);
  nor g__7510(w__7372 ,w__7320 ,w__7274);
  nor g__7511(w__7371 ,w__7319 ,w__7294);
  nor g__7512(w__7370 ,w__7324 ,w__7296);
  nor g__7513(w__7369 ,w__7322 ,w__7288);
  nor g__7514(w__7368 ,w__7309 ,w__7291);
  nor g__7515(w__7367 ,w__7329 ,w__7284);
  nor g__7516(w__7366 ,w__7325 ,w__7273);
  nor g__7517(w__7365 ,w__7335 ,w__7257);
  nor g__7518(w__7364 ,w__7298 ,w__7289);
  nor g__7519(w__7363 ,w__7308 ,w__7268);
  nor g__7520(w__7362 ,w__7334 ,w__7259);
  nor g__7521(w__7361 ,w__7306 ,w__7295);
  or g__7522(w__7382 ,w__7337 ,w__8486);
  nor g__7523(w__7360 ,w__7307 ,w__7292);
  nor g__7524(w__7359 ,w__7316 ,w__7265);
  nor g__7525(w__7358 ,w__7317 ,w__7272);
  and g__7526(w__7357 ,w__7259 ,w__7334);
  nor g__7527(w__7356 ,w__7299 ,w__7277);
  and g__7528(w__7355 ,w__7257 ,w__7335);
  nor g__7529(w__7354 ,w__7312 ,w__7293);
  nor g__7530(w__7353 ,w__7315 ,w__7279);
  and g__7531(w__7352 ,w__7253 ,w__7336);
  nor g__7532(w__7351 ,w__7311 ,w__7281);
  and g__7533(w__7350 ,w__7255 ,w__7332);
  and g__7534(w__7349 ,w__7261 ,w__7333);
  nor g__7535(w__7348 ,w__7326 ,w__7275);
  nor g__7536(w__7347 ,w__7313 ,w__7285);
  nor g__7537(w__7346 ,w__7321 ,w__7262);
  nor g__7538(w__7345 ,w__7323 ,w__7282);
  nor g__7539(w__7344 ,w__7304 ,w__7271);
  nor g__7540(w__7343 ,w__7327 ,w__7266);
  nor g__7541(w__7342 ,w__7303 ,w__7278);
  nor g__7542(w__7341 ,w__7331 ,w__7287);
  nor g__7543(w__7340 ,w__7300 ,w__7267);
  nor g__7544(w__7339 ,w__7301 ,w__7280);
  nor g__7545(w__7338 ,w__7318 ,w__7276);
  not g__7546(w__7337 ,w__8439);
  not g__7547(w__7336 ,w__8489);
  not g__7548(w__7335 ,w__8506);
  not g__7549(w__7334 ,w__8502);
  not g__7550(w__7333 ,w__8444);
  not g__7551(w__7332 ,w__8508);
  not g__7552(w__7297 ,w__7324);
  not g__7553(w__7324 ,w__8488);
  not g__7554(w__7296 ,w__7302);
  not g__7555(w__7302 ,w__8441);
  not g__7556(w__7295 ,w__7320);
  not g__7557(w__7320 ,w__8495);
  not g__7558(w__7294 ,w__7314);
  not g__7559(w__7314 ,w__8504);
  not g__7560(w__7293 ,w__7304);
  not g__7561(w__7304 ,w__8454);
  not g__7562(w__7292 ,w__7331);
  not g__7563(w__7331 ,w__8505);
  not g__7564(w__7291 ,w__7308);
  not g__7565(w__7308 ,w__8456);
  not g__7566(w__7290 ,w__7319);
  not g__7567(w__7319 ,w__8457);
  not g__7568(w__7289 ,w__7325);
  not g__7569(w__7325 ,w__8496);
  not g__7570(w__7288 ,w__7328);
  not g__7571(w__7328 ,w__8507);
  not g__7572(w__7287 ,w__7307);
  not g__7573(w__7307 ,w__8458);
  not g__7574(w__7286 ,w__7322);
  not g__7575(w__7322 ,w__8460);
  not g__7576(w__7285 ,w__7311);
  not g__7577(w__7311 ,w__8492);
  not g__7578(w__7284 ,w__7310);
  not g__7579(w__7310 ,w__8497);
  not g__7580(w__7283 ,w__7330);
  not g__7581(w__7330 ,w__8498);
  not g__7582(w__7282 ,w__7301);
  not g__7583(w__7301 ,w__8443);
  not g__7584(w__7281 ,w__7313);
  not g__7585(w__7313 ,w__8445);
  not g__7586(w__7280 ,w__7323);
  not g__7587(w__7323 ,w__8490);
  not g__7588(w__7279 ,w__7299);
  not g__7589(w__7299 ,w__8493);
  not g__7590(w__7278 ,w__7300);
  not g__7591(w__7300 ,w__8499);
  not g__7592(w__7277 ,w__7315);
  not g__7593(w__7315 ,w__8446);
  not g__7594(w__7276 ,w__7317);
  not g__7595(w__7317 ,w__8447);
  not g__7596(w__7275 ,w__7327);
  not g__7597(w__7327 ,w__8500);
  not g__7598(w__7274 ,w__7306);
  not g__7599(w__7306 ,w__8448);
  not g__7600(w__7273 ,w__7298);
  not g__7601(w__7298 ,w__8449);
  not g__7602(w__7272 ,w__7318);
  not g__7603(w__7318 ,w__8494);
  not g__7604(w__7271 ,w__7312);
  not g__7605(w__7312 ,w__8501);
  not g__7606(w__7270 ,w__7329);
  not g__7607(w__7329 ,w__8450);
  not g__7608(w__7269 ,w__7305);
  not g__7609(w__7305 ,w__8451);
  not g__7610(w__7268 ,w__7309);
  not g__7611(w__7309 ,w__8503);
  not g__7612(w__7267 ,w__7303);
  not g__7613(w__7303 ,w__8452);
  not g__7614(w__7266 ,w__7326);
  not g__7615(w__7326 ,w__8453);
  not g__7616(w__7265 ,w__7321);
  not g__7617(w__7321 ,w__8509);
  not g__7618(w__7264 ,w__7263);
  not g__7619(w__7263 ,w__8487);
  not g__7620(w__7262 ,w__7316);
  not g__7621(w__7316 ,w__8462);
  not g__7622(w__7261 ,w__7260);
  not g__7623(w__7260 ,w__8491);
  not g__7624(w__7259 ,w__7258);
  not g__7625(w__7258 ,w__8455);
  not g__7626(w__7257 ,w__7256);
  not g__7627(w__7256 ,w__8459);
  not g__7628(w__7255 ,w__7254);
  not g__7629(w__7254 ,w__8461);
  not g__7630(w__7253 ,w__7252);
  not g__7631(w__7252 ,w__8442);
  or g__7632(out2 ,w__7537 ,w__7607);
  nor g__7633(w__7607 ,w__7524 ,w__7606);
  or g__7634(w__7606 ,w__7553 ,w__7605);
  nor g__7635(w__7605 ,w__7528 ,w__7604);
  nor g__7636(w__7604 ,w__7552 ,w__7603);
  nor g__7637(w__7603 ,w__7547 ,w__7602);
  nor g__7638(w__7602 ,w__7543 ,w__7601);
  nor g__7639(w__7601 ,w__7533 ,w__7600);
  nor g__7640(w__7600 ,w__7519 ,w__7599);
  nor g__7641(w__7599 ,w__7538 ,w__7598);
  nor g__7642(w__7598 ,w__7558 ,w__7597);
  nor g__7643(w__7597 ,w__7549 ,w__7596);
  nor g__7644(w__7596 ,w__7546 ,w__7595);
  nor g__7645(w__7595 ,w__7541 ,w__7594);
  nor g__7646(w__7594 ,w__7540 ,w__7593);
  nor g__7647(w__7593 ,w__7535 ,w__7592);
  nor g__7648(w__7592 ,w__7532 ,w__7591);
  nor g__7649(w__7591 ,w__7522 ,w__7590);
  nor g__7650(w__7590 ,w__7521 ,w__7589);
  nor g__7651(w__7589 ,w__7526 ,w__7588);
  nor g__7652(w__7588 ,w__7518 ,w__7587);
  nor g__7653(w__7587 ,w__7520 ,w__7586);
  nor g__7654(w__7586 ,w__7554 ,w__7585);
  nor g__7655(w__7585 ,w__7551 ,w__7584);
  nor g__7656(w__7584 ,w__7559 ,w__7583);
  nor g__7657(w__7583 ,w__7545 ,w__7582);
  nor g__7658(w__7582 ,w__7544 ,w__7581);
  nor g__7659(w__7581 ,w__7542 ,w__7580);
  nor g__7660(w__7580 ,w__7550 ,w__7579);
  nor g__7661(w__7579 ,w__7539 ,w__7578);
  nor g__7662(w__7578 ,w__7516 ,w__7577);
  nor g__7663(w__7577 ,w__7536 ,w__7576);
  nor g__7664(w__7576 ,w__7534 ,w__7575);
  nor g__7665(w__7575 ,w__7531 ,w__7574);
  nor g__7666(w__7574 ,w__7529 ,w__7573);
  nor g__7667(w__7573 ,w__7525 ,w__7572);
  nor g__7668(w__7572 ,w__7527 ,w__7571);
  nor g__7669(w__7571 ,w__7555 ,w__7570);
  nor g__7670(w__7570 ,w__7523 ,w__7569);
  nor g__7671(w__7569 ,w__7517 ,w__7568);
  nor g__7672(w__7568 ,w__7556 ,w__7567);
  nor g__7673(w__7567 ,w__7530 ,w__7566);
  nor g__7674(w__7566 ,w__7548 ,w__7565);
  nor g__7675(w__7565 ,w__7557 ,w__7564);
  nor g__7676(w__7564 ,w__7562 ,w__7563);
  nor g__7677(w__7563 ,w__8392 ,w__7561);
  and g__7678(w__7562 ,w__7442 ,w__7560);
  nor g__7679(w__7561 ,w__7442 ,w__7560);
  nor g__7680(w__7559 ,w__7488 ,w__7448);
  nor g__7681(w__7558 ,w__7492 ,w__7468);
  nor g__7682(w__7557 ,w__7480 ,w__7475);
  nor g__7683(w__7556 ,w__7514 ,w__7431);
  nor g__7684(w__7555 ,w__7511 ,w__7439);
  nor g__7685(w__7554 ,w__7508 ,w__7447);
  nor g__7686(w__7553 ,w__7510 ,w__7433);
  nor g__7687(w__7552 ,w__7506 ,w__7464);
  nor g__7688(w__7551 ,w__7483 ,w__7461);
  nor g__7689(w__7550 ,w__7498 ,w__7452);
  nor g__7690(w__7549 ,w__7497 ,w__7472);
  nor g__7691(w__7548 ,w__7502 ,w__7474);
  nor g__7692(w__7547 ,w__7500 ,w__7466);
  nor g__7693(w__7546 ,w__7487 ,w__7469);
  nor g__7694(w__7545 ,w__7507 ,w__7462);
  nor g__7695(w__7544 ,w__7503 ,w__7451);
  nor g__7696(w__7543 ,w__7513 ,w__7435);
  nor g__7697(w__7542 ,w__7476 ,w__7467);
  nor g__7698(w__7541 ,w__7486 ,w__7446);
  nor g__7699(w__7540 ,w__7512 ,w__7437);
  nor g__7700(w__7539 ,w__7484 ,w__7473);
  or g__7701(w__7560 ,w__7515 ,w__8415);
  nor g__7702(w__7538 ,w__7485 ,w__7470);
  nor g__7703(w__7537 ,w__7494 ,w__7443);
  nor g__7704(w__7536 ,w__7495 ,w__7450);
  and g__7705(w__7535 ,w__7437 ,w__7512);
  nor g__7706(w__7534 ,w__7477 ,w__7455);
  and g__7707(w__7533 ,w__7435 ,w__7513);
  nor g__7708(w__7532 ,w__7490 ,w__7471);
  nor g__7709(w__7531 ,w__7493 ,w__7457);
  and g__7710(w__7530 ,w__7431 ,w__7514);
  nor g__7711(w__7529 ,w__7489 ,w__7459);
  and g__7712(w__7528 ,w__7433 ,w__7510);
  and g__7713(w__7527 ,w__7439 ,w__7511);
  nor g__7714(w__7526 ,w__7504 ,w__7453);
  nor g__7715(w__7525 ,w__7491 ,w__7463);
  nor g__7716(w__7524 ,w__7499 ,w__7440);
  nor g__7717(w__7523 ,w__7501 ,w__7460);
  nor g__7718(w__7522 ,w__7482 ,w__7449);
  nor g__7719(w__7521 ,w__7505 ,w__7444);
  nor g__7720(w__7520 ,w__7481 ,w__7456);
  nor g__7721(w__7519 ,w__7509 ,w__7465);
  nor g__7722(w__7518 ,w__7478 ,w__7445);
  nor g__7723(w__7517 ,w__7479 ,w__7458);
  nor g__7724(w__7516 ,w__7496 ,w__7454);
  not g__7725(w__7515 ,w__8391);
  not g__7726(w__7514 ,w__8418);
  not g__7727(w__7513 ,w__8435);
  not g__7728(w__7512 ,w__8431);
  not g__7729(w__7511 ,w__8396);
  not g__7730(w__7510 ,w__8437);
  not g__7731(w__7475 ,w__7502);
  not g__7732(w__7502 ,w__8417);
  not g__7733(w__7474 ,w__7480);
  not g__7734(w__7480 ,w__8393);
  not g__7735(w__7473 ,w__7498);
  not g__7736(w__7498 ,w__8424);
  not g__7737(w__7472 ,w__7492);
  not g__7738(w__7492 ,w__8433);
  not g__7739(w__7471 ,w__7482);
  not g__7740(w__7482 ,w__8406);
  not g__7741(w__7470 ,w__7509);
  not g__7742(w__7509 ,w__8434);
  not g__7743(w__7469 ,w__7486);
  not g__7744(w__7486 ,w__8408);
  not g__7745(w__7468 ,w__7497);
  not g__7746(w__7497 ,w__8409);
  not g__7747(w__7467 ,w__7503);
  not g__7748(w__7503 ,w__8425);
  not g__7749(w__7466 ,w__7506);
  not g__7750(w__7506 ,w__8436);
  not g__7751(w__7465 ,w__7485);
  not g__7752(w__7485 ,w__8410);
  not g__7753(w__7464 ,w__7500);
  not g__7754(w__7500 ,w__8412);
  not g__7755(w__7463 ,w__7489);
  not g__7756(w__7489 ,w__8421);
  not g__7757(w__7462 ,w__7488);
  not g__7758(w__7488 ,w__8426);
  not g__7759(w__7461 ,w__7508);
  not g__7760(w__7508 ,w__8427);
  not g__7761(w__7460 ,w__7479);
  not g__7762(w__7479 ,w__8395);
  not g__7763(w__7459 ,w__7491);
  not g__7764(w__7491 ,w__8397);
  not g__7765(w__7458 ,w__7501);
  not g__7766(w__7501 ,w__8419);
  not g__7767(w__7457 ,w__7477);
  not g__7768(w__7477 ,w__8422);
  not g__7769(w__7456 ,w__7478);
  not g__7770(w__7478 ,w__8428);
  not g__7771(w__7455 ,w__7493);
  not g__7772(w__7493 ,w__8398);
  not g__7773(w__7454 ,w__7495);
  not g__7774(w__7495 ,w__8399);
  not g__7775(w__7453 ,w__7505);
  not g__7776(w__7505 ,w__8429);
  not g__7777(w__7452 ,w__7484);
  not g__7778(w__7484 ,w__8400);
  not g__7779(w__7451 ,w__7476);
  not g__7780(w__7476 ,w__8401);
  not g__7781(w__7450 ,w__7496);
  not g__7782(w__7496 ,w__8423);
  not g__7783(w__7449 ,w__7490);
  not g__7784(w__7490 ,w__8430);
  not g__7785(w__7448 ,w__7507);
  not g__7786(w__7507 ,w__8402);
  not g__7787(w__7447 ,w__7483);
  not g__7788(w__7483 ,w__8403);
  not g__7789(w__7446 ,w__7487);
  not g__7790(w__7487 ,w__8432);
  not g__7791(w__7445 ,w__7481);
  not g__7792(w__7481 ,w__8404);
  not g__7793(w__7444 ,w__7504);
  not g__7794(w__7504 ,w__8405);
  not g__7795(w__7443 ,w__7499);
  not g__7796(w__7499 ,w__8438);
  not g__7797(w__7442 ,w__7441);
  not g__7798(w__7441 ,w__8416);
  not g__7799(w__7440 ,w__7494);
  not g__7800(w__7494 ,w__8414);
  not g__7801(w__7439 ,w__7438);
  not g__7802(w__7438 ,w__8420);
  not g__7803(w__7437 ,w__7436);
  not g__7804(w__7436 ,w__8407);
  not g__7805(w__7435 ,w__7434);
  not g__7806(w__7434 ,w__8411);
  not g__7807(w__7433 ,w__7432);
  not g__7808(w__7432 ,w__8413);
  not g__7809(w__7431 ,w__7430);
  not g__7810(w__7430 ,w__8394);
  or g__7811(out3 ,w__7715 ,w__7785);
  nor g__7812(w__7785 ,w__7702 ,w__7784);
  or g__7813(w__7784 ,w__7731 ,w__7783);
  nor g__7814(w__7783 ,w__7706 ,w__7782);
  nor g__7815(w__7782 ,w__7730 ,w__7781);
  nor g__7816(w__7781 ,w__7725 ,w__7780);
  nor g__7817(w__7780 ,w__7721 ,w__7779);
  nor g__7818(w__7779 ,w__7711 ,w__7778);
  nor g__7819(w__7778 ,w__7697 ,w__7777);
  nor g__7820(w__7777 ,w__7716 ,w__7776);
  nor g__7821(w__7776 ,w__7736 ,w__7775);
  nor g__7822(w__7775 ,w__7727 ,w__7774);
  nor g__7823(w__7774 ,w__7724 ,w__7773);
  nor g__7824(w__7773 ,w__7719 ,w__7772);
  nor g__7825(w__7772 ,w__7718 ,w__7771);
  nor g__7826(w__7771 ,w__7713 ,w__7770);
  nor g__7827(w__7770 ,w__7710 ,w__7769);
  nor g__7828(w__7769 ,w__7700 ,w__7768);
  nor g__7829(w__7768 ,w__7699 ,w__7767);
  nor g__7830(w__7767 ,w__7704 ,w__7766);
  nor g__7831(w__7766 ,w__7696 ,w__7765);
  nor g__7832(w__7765 ,w__7698 ,w__7764);
  nor g__7833(w__7764 ,w__7732 ,w__7763);
  nor g__7834(w__7763 ,w__7729 ,w__7762);
  nor g__7835(w__7762 ,w__7737 ,w__7761);
  nor g__7836(w__7761 ,w__7723 ,w__7760);
  nor g__7837(w__7760 ,w__7722 ,w__7759);
  nor g__7838(w__7759 ,w__7720 ,w__7758);
  nor g__7839(w__7758 ,w__7728 ,w__7757);
  nor g__7840(w__7757 ,w__7717 ,w__7756);
  nor g__7841(w__7756 ,w__7694 ,w__7755);
  nor g__7842(w__7755 ,w__7714 ,w__7754);
  nor g__7843(w__7754 ,w__7712 ,w__7753);
  nor g__7844(w__7753 ,w__7709 ,w__7752);
  nor g__7845(w__7752 ,w__7707 ,w__7751);
  nor g__7846(w__7751 ,w__7703 ,w__7750);
  nor g__7847(w__7750 ,w__7705 ,w__7749);
  nor g__7848(w__7749 ,w__7733 ,w__7748);
  nor g__7849(w__7748 ,w__7701 ,w__7747);
  nor g__7850(w__7747 ,w__7695 ,w__7746);
  nor g__7851(w__7746 ,w__7734 ,w__7745);
  nor g__7852(w__7745 ,w__7708 ,w__7744);
  nor g__7853(w__7744 ,w__7726 ,w__7743);
  nor g__7854(w__7743 ,w__7735 ,w__7742);
  nor g__7855(w__7742 ,w__7740 ,w__7741);
  nor g__7856(w__7741 ,w__8392 ,w__7739);
  and g__7857(w__7740 ,w__7620 ,w__7738);
  nor g__7858(w__7739 ,w__7620 ,w__7738);
  nor g__7859(w__7737 ,w__7666 ,w__7626);
  nor g__7860(w__7736 ,w__7670 ,w__7646);
  nor g__7861(w__7735 ,w__7658 ,w__7653);
  nor g__7862(w__7734 ,w__7692 ,w__7609);
  nor g__7863(w__7733 ,w__7689 ,w__7617);
  nor g__7864(w__7732 ,w__7686 ,w__7625);
  nor g__7865(w__7731 ,w__7688 ,w__7611);
  nor g__7866(w__7730 ,w__7684 ,w__7642);
  nor g__7867(w__7729 ,w__7661 ,w__7639);
  nor g__7868(w__7728 ,w__7676 ,w__7630);
  nor g__7869(w__7727 ,w__7675 ,w__7650);
  nor g__7870(w__7726 ,w__7680 ,w__7652);
  nor g__7871(w__7725 ,w__7678 ,w__7644);
  nor g__7872(w__7724 ,w__7665 ,w__7647);
  nor g__7873(w__7723 ,w__7685 ,w__7640);
  nor g__7874(w__7722 ,w__7681 ,w__7629);
  nor g__7875(w__7721 ,w__7691 ,w__7613);
  nor g__7876(w__7720 ,w__7654 ,w__7645);
  nor g__7877(w__7719 ,w__7664 ,w__7624);
  nor g__7878(w__7718 ,w__7690 ,w__7615);
  nor g__7879(w__7717 ,w__7662 ,w__7651);
  or g__7880(w__7738 ,w__7693 ,w__8344);
  nor g__7881(w__7716 ,w__7663 ,w__7648);
  nor g__7882(w__7715 ,w__7672 ,w__7621);
  nor g__7883(w__7714 ,w__7673 ,w__7628);
  and g__7884(w__7713 ,w__7615 ,w__7690);
  nor g__7885(w__7712 ,w__7655 ,w__7633);
  and g__7886(w__7711 ,w__7613 ,w__7691);
  nor g__7887(w__7710 ,w__7668 ,w__7649);
  nor g__7888(w__7709 ,w__7671 ,w__7635);
  and g__7889(w__7708 ,w__7609 ,w__7692);
  nor g__7890(w__7707 ,w__7667 ,w__7637);
  and g__7891(w__7706 ,w__7611 ,w__7688);
  and g__7892(w__7705 ,w__7617 ,w__7689);
  nor g__7893(w__7704 ,w__7682 ,w__7631);
  nor g__7894(w__7703 ,w__7669 ,w__7641);
  nor g__7895(w__7702 ,w__7677 ,w__7618);
  nor g__7896(w__7701 ,w__7679 ,w__7638);
  nor g__7897(w__7700 ,w__7660 ,w__7627);
  nor g__7898(w__7699 ,w__7683 ,w__7622);
  nor g__7899(w__7698 ,w__7659 ,w__7634);
  nor g__7900(w__7697 ,w__7687 ,w__7643);
  nor g__7901(w__7696 ,w__7656 ,w__7623);
  nor g__7902(w__7695 ,w__7657 ,w__7636);
  nor g__7903(w__7694 ,w__7674 ,w__7632);
  not g__7904(w__7693 ,w__8391);
  not g__7905(w__7692 ,w__8347);
  not g__7906(w__7691 ,w__8364);
  not g__7907(w__7690 ,w__8360);
  not g__7908(w__7689 ,w__8396);
  not g__7909(w__7688 ,w__8366);
  not g__7910(w__7653 ,w__7680);
  not g__7911(w__7680 ,w__8346);
  not g__7912(w__7652 ,w__7658);
  not g__7913(w__7658 ,w__8393);
  not g__7914(w__7651 ,w__7676);
  not g__7915(w__7676 ,w__8353);
  not g__7916(w__7650 ,w__7670);
  not g__7917(w__7670 ,w__8362);
  not g__7918(w__7649 ,w__7660);
  not g__7919(w__7660 ,w__8406);
  not g__7920(w__7648 ,w__7687);
  not g__7921(w__7687 ,w__8363);
  not g__7922(w__7647 ,w__7664);
  not g__7923(w__7664 ,w__8408);
  not g__7924(w__7646 ,w__7675);
  not g__7925(w__7675 ,w__8409);
  not g__7926(w__7645 ,w__7681);
  not g__7927(w__7681 ,w__8354);
  not g__7928(w__7644 ,w__7684);
  not g__7929(w__7684 ,w__8365);
  not g__7930(w__7643 ,w__7663);
  not g__7931(w__7663 ,w__8410);
  not g__7932(w__7642 ,w__7678);
  not g__7933(w__7678 ,w__8412);
  not g__7934(w__7641 ,w__7667);
  not g__7935(w__7667 ,w__8350);
  not g__7936(w__7640 ,w__7666);
  not g__7937(w__7666 ,w__8355);
  not g__7938(w__7639 ,w__7686);
  not g__7939(w__7686 ,w__8356);
  not g__7940(w__7638 ,w__7657);
  not g__7941(w__7657 ,w__8395);
  not g__7942(w__7637 ,w__7669);
  not g__7943(w__7669 ,w__8397);
  not g__7944(w__7636 ,w__7679);
  not g__7945(w__7679 ,w__8348);
  not g__7946(w__7635 ,w__7655);
  not g__7947(w__7655 ,w__8351);
  not g__7948(w__7634 ,w__7656);
  not g__7949(w__7656 ,w__8357);
  not g__7950(w__7633 ,w__7671);
  not g__7951(w__7671 ,w__8398);
  not g__7952(w__7632 ,w__7673);
  not g__7953(w__7673 ,w__8399);
  not g__7954(w__7631 ,w__7683);
  not g__7955(w__7683 ,w__8358);
  not g__7956(w__7630 ,w__7662);
  not g__7957(w__7662 ,w__8400);
  not g__7958(w__7629 ,w__7654);
  not g__7959(w__7654 ,w__8401);
  not g__7960(w__7628 ,w__7674);
  not g__7961(w__7674 ,w__8352);
  not g__7962(w__7627 ,w__7668);
  not g__7963(w__7668 ,w__8359);
  not g__7964(w__7626 ,w__7685);
  not g__7965(w__7685 ,w__8402);
  not g__7966(w__7625 ,w__7661);
  not g__7967(w__7661 ,w__8403);
  not g__7968(w__7624 ,w__7665);
  not g__7969(w__7665 ,w__8361);
  not g__7970(w__7623 ,w__7659);
  not g__7971(w__7659 ,w__8404);
  not g__7972(w__7622 ,w__7682);
  not g__7973(w__7682 ,w__8405);
  not g__7974(w__7621 ,w__7677);
  not g__7975(w__7677 ,w__8367);
  not g__7976(w__7620 ,w__7619);
  not g__7977(w__7619 ,w__8345);
  not g__7978(w__7618 ,w__7672);
  not g__7979(w__7672 ,w__8414);
  not g__7980(w__7617 ,w__7616);
  not g__7981(w__7616 ,w__8349);
  not g__7982(w__7615 ,w__7614);
  not g__7983(w__7614 ,w__8407);
  not g__7984(w__7613 ,w__7612);
  not g__7985(w__7612 ,w__8411);
  not g__7986(w__7611 ,w__7610);
  not g__7987(w__7610 ,w__8413);
  not g__7988(w__7609 ,w__7608);
  not g__7989(w__7608 ,w__8394);
  or g__7990(out4 ,w__7893 ,w__7963);
  nor g__7991(w__7963 ,w__7880 ,w__7962);
  or g__7992(w__7962 ,w__7909 ,w__7961);
  nor g__7993(w__7961 ,w__7884 ,w__7960);
  nor g__7994(w__7960 ,w__7908 ,w__7959);
  nor g__7995(w__7959 ,w__7903 ,w__7958);
  nor g__7996(w__7958 ,w__7899 ,w__7957);
  nor g__7997(w__7957 ,w__7889 ,w__7956);
  nor g__7998(w__7956 ,w__7875 ,w__7955);
  nor g__7999(w__7955 ,w__7894 ,w__7954);
  nor g__8000(w__7954 ,w__7914 ,w__7953);
  nor g__8001(w__7953 ,w__7905 ,w__7952);
  nor g__8002(w__7952 ,w__7902 ,w__7951);
  nor g__8003(w__7951 ,w__7897 ,w__7950);
  nor g__8004(w__7950 ,w__7896 ,w__7949);
  nor g__8005(w__7949 ,w__7891 ,w__7948);
  nor g__8006(w__7948 ,w__7888 ,w__7947);
  nor g__8007(w__7947 ,w__7878 ,w__7946);
  nor g__8008(w__7946 ,w__7877 ,w__7945);
  nor g__8009(w__7945 ,w__7882 ,w__7944);
  nor g__8010(w__7944 ,w__7874 ,w__7943);
  nor g__8011(w__7943 ,w__7876 ,w__7942);
  nor g__8012(w__7942 ,w__7910 ,w__7941);
  nor g__8013(w__7941 ,w__7907 ,w__7940);
  nor g__8014(w__7940 ,w__7915 ,w__7939);
  nor g__8015(w__7939 ,w__7901 ,w__7938);
  nor g__8016(w__7938 ,w__7900 ,w__7937);
  nor g__8017(w__7937 ,w__7898 ,w__7936);
  nor g__8018(w__7936 ,w__7906 ,w__7935);
  nor g__8019(w__7935 ,w__7895 ,w__7934);
  nor g__8020(w__7934 ,w__7872 ,w__7933);
  nor g__8021(w__7933 ,w__7892 ,w__7932);
  nor g__8022(w__7932 ,w__7890 ,w__7931);
  nor g__8023(w__7931 ,w__7887 ,w__7930);
  nor g__8024(w__7930 ,w__7885 ,w__7929);
  nor g__8025(w__7929 ,w__7881 ,w__7928);
  nor g__8026(w__7928 ,w__7883 ,w__7927);
  nor g__8027(w__7927 ,w__7911 ,w__7926);
  nor g__8028(w__7926 ,w__7879 ,w__7925);
  nor g__8029(w__7925 ,w__7873 ,w__7924);
  nor g__8030(w__7924 ,w__7912 ,w__7923);
  nor g__8031(w__7923 ,w__7886 ,w__7922);
  nor g__8032(w__7922 ,w__7904 ,w__7921);
  nor g__8033(w__7921 ,w__7913 ,w__7920);
  nor g__8034(w__7920 ,w__7918 ,w__7919);
  nor g__8035(w__7919 ,w__8321 ,w__7917);
  and g__8036(w__7918 ,w__7798 ,w__7916);
  nor g__8037(w__7917 ,w__7798 ,w__7916);
  nor g__8038(w__7915 ,w__7844 ,w__7804);
  nor g__8039(w__7914 ,w__7848 ,w__7824);
  nor g__8040(w__7913 ,w__7836 ,w__7831);
  nor g__8041(w__7912 ,w__7870 ,w__7787);
  nor g__8042(w__7911 ,w__7867 ,w__7795);
  nor g__8043(w__7910 ,w__7864 ,w__7803);
  nor g__8044(w__7909 ,w__7866 ,w__7789);
  nor g__8045(w__7908 ,w__7862 ,w__7820);
  nor g__8046(w__7907 ,w__7839 ,w__7817);
  nor g__8047(w__7906 ,w__7854 ,w__7808);
  nor g__8048(w__7905 ,w__7853 ,w__7828);
  nor g__8049(w__7904 ,w__7858 ,w__7830);
  nor g__8050(w__7903 ,w__7856 ,w__7822);
  nor g__8051(w__7902 ,w__7843 ,w__7825);
  nor g__8052(w__7901 ,w__7863 ,w__7818);
  nor g__8053(w__7900 ,w__7859 ,w__7807);
  nor g__8054(w__7899 ,w__7869 ,w__7791);
  nor g__8055(w__7898 ,w__7832 ,w__7823);
  nor g__8056(w__7897 ,w__7842 ,w__7802);
  nor g__8057(w__7896 ,w__7868 ,w__7793);
  nor g__8058(w__7895 ,w__7840 ,w__7829);
  or g__8059(w__7916 ,w__7871 ,w__8486);
  nor g__8060(w__7894 ,w__7841 ,w__7826);
  nor g__8061(w__7893 ,w__7850 ,w__7799);
  nor g__8062(w__7892 ,w__7851 ,w__7806);
  and g__8063(w__7891 ,w__7793 ,w__7868);
  nor g__8064(w__7890 ,w__7833 ,w__7811);
  and g__8065(w__7889 ,w__7791 ,w__7869);
  nor g__8066(w__7888 ,w__7846 ,w__7827);
  nor g__8067(w__7887 ,w__7849 ,w__7813);
  and g__8068(w__7886 ,w__7787 ,w__7870);
  nor g__8069(w__7885 ,w__7845 ,w__7815);
  and g__8070(w__7884 ,w__7789 ,w__7866);
  and g__8071(w__7883 ,w__7795 ,w__7867);
  nor g__8072(w__7882 ,w__7860 ,w__7809);
  nor g__8073(w__7881 ,w__7847 ,w__7819);
  nor g__8074(w__7880 ,w__7855 ,w__7796);
  nor g__8075(w__7879 ,w__7857 ,w__7816);
  nor g__8076(w__7878 ,w__7838 ,w__7805);
  nor g__8077(w__7877 ,w__7861 ,w__7800);
  nor g__8078(w__7876 ,w__7837 ,w__7812);
  nor g__8079(w__7875 ,w__7865 ,w__7821);
  nor g__8080(w__7874 ,w__7834 ,w__7801);
  nor g__8081(w__7873 ,w__7835 ,w__7814);
  nor g__8082(w__7872 ,w__7852 ,w__7810);
  not g__8083(w__7871 ,w__8320);
  not g__8084(w__7870 ,w__8489);
  not g__8085(w__7869 ,w__8506);
  not g__8086(w__7868 ,w__8502);
  not g__8087(w__7867 ,w__8325);
  not g__8088(w__7866 ,w__8508);
  not g__8089(w__7831 ,w__7858);
  not g__8090(w__7858 ,w__8488);
  not g__8091(w__7830 ,w__7836);
  not g__8092(w__7836 ,w__8322);
  not g__8093(w__7829 ,w__7854);
  not g__8094(w__7854 ,w__8495);
  not g__8095(w__7828 ,w__7848);
  not g__8096(w__7848 ,w__8504);
  not g__8097(w__7827 ,w__7838);
  not g__8098(w__7838 ,w__8335);
  not g__8099(w__7826 ,w__7865);
  not g__8100(w__7865 ,w__8505);
  not g__8101(w__7825 ,w__7842);
  not g__8102(w__7842 ,w__8337);
  not g__8103(w__7824 ,w__7853);
  not g__8104(w__7853 ,w__8338);
  not g__8105(w__7823 ,w__7859);
  not g__8106(w__7859 ,w__8496);
  not g__8107(w__7822 ,w__7862);
  not g__8108(w__7862 ,w__8507);
  not g__8109(w__7821 ,w__7841);
  not g__8110(w__7841 ,w__8339);
  not g__8111(w__7820 ,w__7856);
  not g__8112(w__7856 ,w__8341);
  not g__8113(w__7819 ,w__7845);
  not g__8114(w__7845 ,w__8492);
  not g__8115(w__7818 ,w__7844);
  not g__8116(w__7844 ,w__8497);
  not g__8117(w__7817 ,w__7864);
  not g__8118(w__7864 ,w__8498);
  not g__8119(w__7816 ,w__7835);
  not g__8120(w__7835 ,w__8324);
  not g__8121(w__7815 ,w__7847);
  not g__8122(w__7847 ,w__8326);
  not g__8123(w__7814 ,w__7857);
  not g__8124(w__7857 ,w__8490);
  not g__8125(w__7813 ,w__7833);
  not g__8126(w__7833 ,w__8493);
  not g__8127(w__7812 ,w__7834);
  not g__8128(w__7834 ,w__8499);
  not g__8129(w__7811 ,w__7849);
  not g__8130(w__7849 ,w__8327);
  not g__8131(w__7810 ,w__7851);
  not g__8132(w__7851 ,w__8328);
  not g__8133(w__7809 ,w__7861);
  not g__8134(w__7861 ,w__8500);
  not g__8135(w__7808 ,w__7840);
  not g__8136(w__7840 ,w__8329);
  not g__8137(w__7807 ,w__7832);
  not g__8138(w__7832 ,w__8330);
  not g__8139(w__7806 ,w__7852);
  not g__8140(w__7852 ,w__8494);
  not g__8141(w__7805 ,w__7846);
  not g__8142(w__7846 ,w__8501);
  not g__8143(w__7804 ,w__7863);
  not g__8144(w__7863 ,w__8331);
  not g__8145(w__7803 ,w__7839);
  not g__8146(w__7839 ,w__8332);
  not g__8147(w__7802 ,w__7843);
  not g__8148(w__7843 ,w__8503);
  not g__8149(w__7801 ,w__7837);
  not g__8150(w__7837 ,w__8333);
  not g__8151(w__7800 ,w__7860);
  not g__8152(w__7860 ,w__8334);
  not g__8153(w__7799 ,w__7855);
  not g__8154(w__7855 ,w__8509);
  not g__8155(w__7798 ,w__7797);
  not g__8156(w__7797 ,w__8487);
  not g__8157(w__7796 ,w__7850);
  not g__8158(w__7850 ,w__8343);
  not g__8159(w__7795 ,w__7794);
  not g__8160(w__7794 ,w__8491);
  not g__8161(w__7793 ,w__7792);
  not g__8162(w__7792 ,w__8336);
  not g__8163(w__7791 ,w__7790);
  not g__8164(w__7790 ,w__8340);
  not g__8165(w__7789 ,w__7788);
  not g__8166(w__7788 ,w__8342);
  not g__8167(w__7787 ,w__7786);
  not g__8168(w__7786 ,w__8323);
  or g__8169(out5 ,w__8071 ,w__8141);
  nor g__8170(w__8141 ,w__8058 ,w__8140);
  or g__8171(w__8140 ,w__8087 ,w__8139);
  nor g__8172(w__8139 ,w__8062 ,w__8138);
  nor g__8173(w__8138 ,w__8086 ,w__8137);
  nor g__8174(w__8137 ,w__8081 ,w__8136);
  nor g__8175(w__8136 ,w__8077 ,w__8135);
  nor g__8176(w__8135 ,w__8067 ,w__8134);
  nor g__8177(w__8134 ,w__8053 ,w__8133);
  nor g__8178(w__8133 ,w__8072 ,w__8132);
  nor g__8179(w__8132 ,w__8092 ,w__8131);
  nor g__8180(w__8131 ,w__8083 ,w__8130);
  nor g__8181(w__8130 ,w__8080 ,w__8129);
  nor g__8182(w__8129 ,w__8075 ,w__8128);
  nor g__8183(w__8128 ,w__8074 ,w__8127);
  nor g__8184(w__8127 ,w__8069 ,w__8126);
  nor g__8185(w__8126 ,w__8066 ,w__8125);
  nor g__8186(w__8125 ,w__8056 ,w__8124);
  nor g__8187(w__8124 ,w__8055 ,w__8123);
  nor g__8188(w__8123 ,w__8060 ,w__8122);
  nor g__8189(w__8122 ,w__8052 ,w__8121);
  nor g__8190(w__8121 ,w__8054 ,w__8120);
  nor g__8191(w__8120 ,w__8088 ,w__8119);
  nor g__8192(w__8119 ,w__8085 ,w__8118);
  nor g__8193(w__8118 ,w__8093 ,w__8117);
  nor g__8194(w__8117 ,w__8079 ,w__8116);
  nor g__8195(w__8116 ,w__8078 ,w__8115);
  nor g__8196(w__8115 ,w__8076 ,w__8114);
  nor g__8197(w__8114 ,w__8084 ,w__8113);
  nor g__8198(w__8113 ,w__8073 ,w__8112);
  nor g__8199(w__8112 ,w__8050 ,w__8111);
  nor g__8200(w__8111 ,w__8070 ,w__8110);
  nor g__8201(w__8110 ,w__8068 ,w__8109);
  nor g__8202(w__8109 ,w__8065 ,w__8108);
  nor g__8203(w__8108 ,w__8063 ,w__8107);
  nor g__8204(w__8107 ,w__8059 ,w__8106);
  nor g__8205(w__8106 ,w__8061 ,w__8105);
  nor g__8206(w__8105 ,w__8089 ,w__8104);
  nor g__8207(w__8104 ,w__8057 ,w__8103);
  nor g__8208(w__8103 ,w__8051 ,w__8102);
  nor g__8209(w__8102 ,w__8090 ,w__8101);
  nor g__8210(w__8101 ,w__8064 ,w__8100);
  nor g__8211(w__8100 ,w__8082 ,w__8099);
  nor g__8212(w__8099 ,w__8091 ,w__8098);
  nor g__8213(w__8098 ,w__8096 ,w__8097);
  nor g__8214(w__8097 ,w__8440 ,w__8095);
  and g__8215(w__8096 ,w__7976 ,w__8094);
  nor g__8216(w__8095 ,w__7976 ,w__8094);
  nor g__8217(w__8093 ,w__8022 ,w__7982);
  nor g__8218(w__8092 ,w__8026 ,w__8002);
  nor g__8219(w__8091 ,w__8014 ,w__8009);
  nor g__8220(w__8090 ,w__8048 ,w__7965);
  nor g__8221(w__8089 ,w__8045 ,w__7973);
  nor g__8222(w__8088 ,w__8042 ,w__7981);
  nor g__8223(w__8087 ,w__8044 ,w__7967);
  nor g__8224(w__8086 ,w__8040 ,w__7998);
  nor g__8225(w__8085 ,w__8017 ,w__7995);
  nor g__8226(w__8084 ,w__8032 ,w__7986);
  nor g__8227(w__8083 ,w__8031 ,w__8006);
  nor g__8228(w__8082 ,w__8036 ,w__8008);
  nor g__8229(w__8081 ,w__8034 ,w__8000);
  nor g__8230(w__8080 ,w__8021 ,w__8003);
  nor g__8231(w__8079 ,w__8041 ,w__7996);
  nor g__8232(w__8078 ,w__8037 ,w__7985);
  nor g__8233(w__8077 ,w__8047 ,w__7969);
  nor g__8234(w__8076 ,w__8010 ,w__8001);
  nor g__8235(w__8075 ,w__8020 ,w__7980);
  nor g__8236(w__8074 ,w__8046 ,w__7971);
  nor g__8237(w__8073 ,w__8018 ,w__8007);
  or g__8238(w__8094 ,w__8049 ,w__8320);
  nor g__8239(w__8072 ,w__8019 ,w__8004);
  nor g__8240(w__8071 ,w__8028 ,w__7977);
  nor g__8241(w__8070 ,w__8029 ,w__7984);
  and g__8242(w__8069 ,w__7971 ,w__8046);
  nor g__8243(w__8068 ,w__8011 ,w__7989);
  and g__8244(w__8067 ,w__7969 ,w__8047);
  nor g__8245(w__8066 ,w__8024 ,w__8005);
  nor g__8246(w__8065 ,w__8027 ,w__7991);
  and g__8247(w__8064 ,w__7965 ,w__8048);
  nor g__8248(w__8063 ,w__8023 ,w__7993);
  and g__8249(w__8062 ,w__7967 ,w__8044);
  and g__8250(w__8061 ,w__7973 ,w__8045);
  nor g__8251(w__8060 ,w__8038 ,w__7987);
  nor g__8252(w__8059 ,w__8025 ,w__7997);
  nor g__8253(w__8058 ,w__8033 ,w__7974);
  nor g__8254(w__8057 ,w__8035 ,w__7994);
  nor g__8255(w__8056 ,w__8016 ,w__7983);
  nor g__8256(w__8055 ,w__8039 ,w__7978);
  nor g__8257(w__8054 ,w__8015 ,w__7990);
  nor g__8258(w__8053 ,w__8043 ,w__7999);
  nor g__8259(w__8052 ,w__8012 ,w__7979);
  nor g__8260(w__8051 ,w__8013 ,w__7992);
  nor g__8261(w__8050 ,w__8030 ,w__7988);
  not g__8262(w__8049 ,w__8439);
  not g__8263(w__8048 ,w__8323);
  not g__8264(w__8047 ,w__8340);
  not g__8265(w__8046 ,w__8336);
  not g__8266(w__8045 ,w__8444);
  not g__8267(w__8044 ,w__8342);
  not g__8268(w__8009 ,w__8036);
  not g__8269(w__8036 ,w__8322);
  not g__8270(w__8008 ,w__8014);
  not g__8271(w__8014 ,w__8441);
  not g__8272(w__8007 ,w__8032);
  not g__8273(w__8032 ,w__8329);
  not g__8274(w__8006 ,w__8026);
  not g__8275(w__8026 ,w__8338);
  not g__8276(w__8005 ,w__8016);
  not g__8277(w__8016 ,w__8454);
  not g__8278(w__8004 ,w__8043);
  not g__8279(w__8043 ,w__8339);
  not g__8280(w__8003 ,w__8020);
  not g__8281(w__8020 ,w__8456);
  not g__8282(w__8002 ,w__8031);
  not g__8283(w__8031 ,w__8457);
  not g__8284(w__8001 ,w__8037);
  not g__8285(w__8037 ,w__8330);
  not g__8286(w__8000 ,w__8040);
  not g__8287(w__8040 ,w__8341);
  not g__8288(w__7999 ,w__8019);
  not g__8289(w__8019 ,w__8458);
  not g__8290(w__7998 ,w__8034);
  not g__8291(w__8034 ,w__8460);
  not g__8292(w__7997 ,w__8023);
  not g__8293(w__8023 ,w__8326);
  not g__8294(w__7996 ,w__8022);
  not g__8295(w__8022 ,w__8331);
  not g__8296(w__7995 ,w__8042);
  not g__8297(w__8042 ,w__8332);
  not g__8298(w__7994 ,w__8013);
  not g__8299(w__8013 ,w__8443);
  not g__8300(w__7993 ,w__8025);
  not g__8301(w__8025 ,w__8445);
  not g__8302(w__7992 ,w__8035);
  not g__8303(w__8035 ,w__8324);
  not g__8304(w__7991 ,w__8011);
  not g__8305(w__8011 ,w__8327);
  not g__8306(w__7990 ,w__8012);
  not g__8307(w__8012 ,w__8333);
  not g__8308(w__7989 ,w__8027);
  not g__8309(w__8027 ,w__8446);
  not g__8310(w__7988 ,w__8029);
  not g__8311(w__8029 ,w__8447);
  not g__8312(w__7987 ,w__8039);
  not g__8313(w__8039 ,w__8334);
  not g__8314(w__7986 ,w__8018);
  not g__8315(w__8018 ,w__8448);
  not g__8316(w__7985 ,w__8010);
  not g__8317(w__8010 ,w__8449);
  not g__8318(w__7984 ,w__8030);
  not g__8319(w__8030 ,w__8328);
  not g__8320(w__7983 ,w__8024);
  not g__8321(w__8024 ,w__8335);
  not g__8322(w__7982 ,w__8041);
  not g__8323(w__8041 ,w__8450);
  not g__8324(w__7981 ,w__8017);
  not g__8325(w__8017 ,w__8451);
  not g__8326(w__7980 ,w__8021);
  not g__8327(w__8021 ,w__8337);
  not g__8328(w__7979 ,w__8015);
  not g__8329(w__8015 ,w__8452);
  not g__8330(w__7978 ,w__8038);
  not g__8331(w__8038 ,w__8453);
  not g__8332(w__7977 ,w__8033);
  not g__8333(w__8033 ,w__8343);
  not g__8334(w__7976 ,w__7975);
  not g__8335(w__7975 ,w__8321);
  not g__8336(w__7974 ,w__8028);
  not g__8337(w__8028 ,w__8462);
  not g__8338(w__7973 ,w__7972);
  not g__8339(w__7972 ,w__8325);
  not g__8340(w__7971 ,w__7970);
  not g__8341(w__7970 ,w__8455);
  not g__8342(w__7969 ,w__7968);
  not g__8343(w__7968 ,w__8459);
  not g__8344(w__7967 ,w__7966);
  not g__8345(w__7966 ,w__8461);
  not g__8346(w__7965 ,w__7964);
  not g__8347(w__7964 ,w__8442);
  or g__8348(out6 ,w__8249 ,w__8319);
  nor g__8349(w__8319 ,w__8236 ,w__8318);
  or g__8350(w__8318 ,w__8265 ,w__8317);
  nor g__8351(w__8317 ,w__8240 ,w__8316);
  nor g__8352(w__8316 ,w__8264 ,w__8315);
  nor g__8353(w__8315 ,w__8259 ,w__8314);
  nor g__8354(w__8314 ,w__8255 ,w__8313);
  nor g__8355(w__8313 ,w__8245 ,w__8312);
  nor g__8356(w__8312 ,w__8231 ,w__8311);
  nor g__8357(w__8311 ,w__8250 ,w__8310);
  nor g__8358(w__8310 ,w__8270 ,w__8309);
  nor g__8359(w__8309 ,w__8261 ,w__8308);
  nor g__8360(w__8308 ,w__8258 ,w__8307);
  nor g__8361(w__8307 ,w__8253 ,w__8306);
  nor g__8362(w__8306 ,w__8252 ,w__8305);
  nor g__8363(w__8305 ,w__8247 ,w__8304);
  nor g__8364(w__8304 ,w__8244 ,w__8303);
  nor g__8365(w__8303 ,w__8234 ,w__8302);
  nor g__8366(w__8302 ,w__8233 ,w__8301);
  nor g__8367(w__8301 ,w__8238 ,w__8300);
  nor g__8368(w__8300 ,w__8230 ,w__8299);
  nor g__8369(w__8299 ,w__8232 ,w__8298);
  nor g__8370(w__8298 ,w__8266 ,w__8297);
  nor g__8371(w__8297 ,w__8263 ,w__8296);
  nor g__8372(w__8296 ,w__8271 ,w__8295);
  nor g__8373(w__8295 ,w__8257 ,w__8294);
  nor g__8374(w__8294 ,w__8256 ,w__8293);
  nor g__8375(w__8293 ,w__8254 ,w__8292);
  nor g__8376(w__8292 ,w__8262 ,w__8291);
  nor g__8377(w__8291 ,w__8251 ,w__8290);
  nor g__8378(w__8290 ,w__8228 ,w__8289);
  nor g__8379(w__8289 ,w__8248 ,w__8288);
  nor g__8380(w__8288 ,w__8246 ,w__8287);
  nor g__8381(w__8287 ,w__8243 ,w__8286);
  nor g__8382(w__8286 ,w__8241 ,w__8285);
  nor g__8383(w__8285 ,w__8237 ,w__8284);
  nor g__8384(w__8284 ,w__8239 ,w__8283);
  nor g__8385(w__8283 ,w__8267 ,w__8282);
  nor g__8386(w__8282 ,w__8235 ,w__8281);
  nor g__8387(w__8281 ,w__8229 ,w__8280);
  nor g__8388(w__8280 ,w__8268 ,w__8279);
  nor g__8389(w__8279 ,w__8242 ,w__8278);
  nor g__8390(w__8278 ,w__8260 ,w__8277);
  nor g__8391(w__8277 ,w__8269 ,w__8276);
  nor g__8392(w__8276 ,w__8274 ,w__8275);
  nor g__8393(w__8275 ,w__8345 ,w__8273);
  and g__8394(w__8274 ,w__8154 ,w__8272);
  nor g__8395(w__8273 ,w__8154 ,w__8272);
  nor g__8396(w__8271 ,w__8200 ,w__8160);
  nor g__8397(w__8270 ,w__8204 ,w__8180);
  nor g__8398(w__8269 ,w__8192 ,w__8187);
  nor g__8399(w__8268 ,w__8226 ,w__8143);
  nor g__8400(w__8267 ,w__8223 ,w__8151);
  nor g__8401(w__8266 ,w__8220 ,w__8159);
  nor g__8402(w__8265 ,w__8222 ,w__8145);
  nor g__8403(w__8264 ,w__8218 ,w__8176);
  nor g__8404(w__8263 ,w__8195 ,w__8173);
  nor g__8405(w__8262 ,w__8210 ,w__8164);
  nor g__8406(w__8261 ,w__8209 ,w__8184);
  nor g__8407(w__8260 ,w__8214 ,w__8186);
  nor g__8408(w__8259 ,w__8212 ,w__8178);
  nor g__8409(w__8258 ,w__8199 ,w__8181);
  nor g__8410(w__8257 ,w__8219 ,w__8174);
  nor g__8411(w__8256 ,w__8215 ,w__8163);
  nor g__8412(w__8255 ,w__8225 ,w__8147);
  nor g__8413(w__8254 ,w__8188 ,w__8179);
  nor g__8414(w__8253 ,w__8198 ,w__8158);
  nor g__8415(w__8252 ,w__8224 ,w__8149);
  nor g__8416(w__8251 ,w__8196 ,w__8185);
  or g__8417(w__8272 ,w__8227 ,w__8415);
  nor g__8418(w__8250 ,w__8197 ,w__8182);
  nor g__8419(w__8249 ,w__8206 ,w__8155);
  nor g__8420(w__8248 ,w__8207 ,w__8162);
  and g__8421(w__8247 ,w__8149 ,w__8224);
  nor g__8422(w__8246 ,w__8189 ,w__8167);
  and g__8423(w__8245 ,w__8147 ,w__8225);
  nor g__8424(w__8244 ,w__8202 ,w__8183);
  nor g__8425(w__8243 ,w__8205 ,w__8169);
  and g__8426(w__8242 ,w__8143 ,w__8226);
  nor g__8427(w__8241 ,w__8201 ,w__8171);
  and g__8428(w__8240 ,w__8145 ,w__8222);
  and g__8429(w__8239 ,w__8151 ,w__8223);
  nor g__8430(w__8238 ,w__8216 ,w__8165);
  nor g__8431(w__8237 ,w__8203 ,w__8175);
  nor g__8432(w__8236 ,w__8211 ,w__8152);
  nor g__8433(w__8235 ,w__8213 ,w__8172);
  nor g__8434(w__8234 ,w__8194 ,w__8161);
  nor g__8435(w__8233 ,w__8217 ,w__8156);
  nor g__8436(w__8232 ,w__8193 ,w__8168);
  nor g__8437(w__8231 ,w__8221 ,w__8177);
  nor g__8438(w__8230 ,w__8190 ,w__8157);
  nor g__8439(w__8229 ,w__8191 ,w__8170);
  nor g__8440(w__8228 ,w__8208 ,w__8166);
  not g__8441(w__8227 ,w__8344);
  not g__8442(w__8226 ,w__8418);
  not g__8443(w__8225 ,w__8435);
  not g__8444(w__8224 ,w__8431);
  not g__8445(w__8223 ,w__8349);
  not g__8446(w__8222 ,w__8437);
  not g__8447(w__8187 ,w__8214);
  not g__8448(w__8214 ,w__8417);
  not g__8449(w__8186 ,w__8192);
  not g__8450(w__8192 ,w__8346);
  not g__8451(w__8185 ,w__8210);
  not g__8452(w__8210 ,w__8424);
  not g__8453(w__8184 ,w__8204);
  not g__8454(w__8204 ,w__8433);
  not g__8455(w__8183 ,w__8194);
  not g__8456(w__8194 ,w__8359);
  not g__8457(w__8182 ,w__8221);
  not g__8458(w__8221 ,w__8434);
  not g__8459(w__8181 ,w__8198);
  not g__8460(w__8198 ,w__8361);
  not g__8461(w__8180 ,w__8209);
  not g__8462(w__8209 ,w__8362);
  not g__8463(w__8179 ,w__8215);
  not g__8464(w__8215 ,w__8425);
  not g__8465(w__8178 ,w__8218);
  not g__8466(w__8218 ,w__8436);
  not g__8467(w__8177 ,w__8197);
  not g__8468(w__8197 ,w__8363);
  not g__8469(w__8176 ,w__8212);
  not g__8470(w__8212 ,w__8365);
  not g__8471(w__8175 ,w__8201);
  not g__8472(w__8201 ,w__8421);
  not g__8473(w__8174 ,w__8200);
  not g__8474(w__8200 ,w__8426);
  not g__8475(w__8173 ,w__8220);
  not g__8476(w__8220 ,w__8427);
  not g__8477(w__8172 ,w__8191);
  not g__8478(w__8191 ,w__8348);
  not g__8479(w__8171 ,w__8203);
  not g__8480(w__8203 ,w__8350);
  not g__8481(w__8170 ,w__8213);
  not g__8482(w__8213 ,w__8419);
  not g__8483(w__8169 ,w__8189);
  not g__8484(w__8189 ,w__8422);
  not g__8485(w__8168 ,w__8190);
  not g__8486(w__8190 ,w__8428);
  not g__8487(w__8167 ,w__8205);
  not g__8488(w__8205 ,w__8351);
  not g__8489(w__8166 ,w__8207);
  not g__8490(w__8207 ,w__8352);
  not g__8491(w__8165 ,w__8217);
  not g__8492(w__8217 ,w__8429);
  not g__8493(w__8164 ,w__8196);
  not g__8494(w__8196 ,w__8353);
  not g__8495(w__8163 ,w__8188);
  not g__8496(w__8188 ,w__8354);
  not g__8497(w__8162 ,w__8208);
  not g__8498(w__8208 ,w__8423);
  not g__8499(w__8161 ,w__8202);
  not g__8500(w__8202 ,w__8430);
  not g__8501(w__8160 ,w__8219);
  not g__8502(w__8219 ,w__8355);
  not g__8503(w__8159 ,w__8195);
  not g__8504(w__8195 ,w__8356);
  not g__8505(w__8158 ,w__8199);
  not g__8506(w__8199 ,w__8432);
  not g__8507(w__8157 ,w__8193);
  not g__8508(w__8193 ,w__8357);
  not g__8509(w__8156 ,w__8216);
  not g__8510(w__8216 ,w__8358);
  not g__8511(w__8155 ,w__8211);
  not g__8512(w__8211 ,w__8438);
  not g__8513(w__8154 ,w__8153);
  not g__8514(w__8153 ,w__8416);
  not g__8515(w__8152 ,w__8206);
  not g__8516(w__8206 ,w__8367);
  not g__8517(w__8151 ,w__8150);
  not g__8518(w__8150 ,w__8420);
  not g__8519(w__8149 ,w__8148);
  not g__8520(w__8148 ,w__8360);
  not g__8521(w__8147 ,w__8146);
  not g__8522(w__8146 ,w__8364);
  not g__8523(w__8145 ,w__8144);
  not g__8524(w__8144 ,w__8366);
  not g__8525(w__8143 ,w__8142);
  not g__8526(w__8142 ,w__8347);
  not g__8527(w__1408 ,w__1351);
  not g__8528(w__3147 ,w__3090);
  not g__8529(w__3824 ,w__3767);
  not g__8530(w__4500 ,w__4443);
  not g__8531(w__6241 ,w__6184);
  not g__8532(w__6919 ,w__6862);
  buf g__8533(w__8487 ,w__1363);
  buf g__8534(w__8416 ,w__3779);
  not g__8535(w__8488 ,w__1448);
  not g__8536(w__8417 ,w__3864);
  buf g__8537(w__1515 ,w__1439);
  buf g__8538(w__3931 ,w__3855);
endmodule
