// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.

module WT_USP_KS_8x8_noX(
        input logic [7:0] IN1,
        input logic [7:0] IN2,
        output logic [15:0] result);
    
    
// Creating Partial Products 

    wire logic [7:0] pp0;
    wire logic [7:0] pp1;
    wire logic [7:0] pp2;
    wire logic [7:0] pp3;
    wire logic [7:0] pp4;
    wire logic [7:0] pp5;
    wire logic [7:0] pp6;
    wire logic [7:0] pp7;
    assign pp0 = {8{IN1[0]}} & IN2;
    assign pp1 = {8{IN1[1]}} & IN2;
    assign pp2 = {8{IN1[2]}} & IN2;
    assign pp3 = {8{IN1[3]}} & IN2;
    assign pp4 = {8{IN1[4]}} & IN2;
    assign pp5 = {8{IN1[5]}} & IN2;
    assign pp6 = {8{IN1[6]}} & IN2;
    assign pp7 = {8{IN1[7]}} & IN2;
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp0[0] pp0[1] pp0[2] pp0[3] pp0[4] pp0[5] pp0[6] pp0[7]   --     --     --     --     --     --     --   
     //   --   pp1[0] pp1[1] pp1[2] pp1[3] pp1[4] pp1[5] pp1[6] pp1[7]   --     --     --     --     --     --   
     //   --     --   pp2[0] pp2[1] pp2[2] pp2[3] pp2[4] pp2[5] pp2[6] pp2[7]   --     --     --     --     --   
     //   --     --     --   pp3[0] pp3[1] pp3[2] pp3[3] pp3[4] pp3[5] pp3[6] pp3[7]   --     --     --     --   
     //   --     --     --     --   pp4[0] pp4[1] pp4[2] pp4[3] pp4[4] pp4[5] pp4[6] pp4[7]   --     --     --   
     //   --     --     --     --     --   pp5[0] pp5[1] pp5[2] pp5[3] pp5[4] pp5[5] pp5[6] pp5[7]   --     --   
     //   --     --     --     --     --     --   pp6[0] pp6[1] pp6[2] pp6[3] pp6[4] pp6[5] pp6[6] pp6[7]   --   
     //   --     --     --     --     --     --     --   pp7[0] pp7[1] pp7[2] pp7[3] pp7[4] pp7[5] pp7[6] pp7[7] 
    
// Creating Summation Tree 

    
    // Wallace Summation Stage 1
    logic s0 ,c0;
    ha ha0 (pp0[1], pp1[0], s0, c0);
    logic s1 ,c1; 
    fa fa1 (pp0[2], pp1[1], pp2[0], s1, c1);
    logic s2 ,c2; 
    fa fa2 (pp0[3], pp1[2], pp2[1], s2, c2);
    logic s3 ,c3; 
    fa fa3 (pp0[4], pp1[3], pp2[2], s3, c3);
    logic s4 ,c4;
    ha ha4 (pp3[1], pp4[0], s4, c4);
    logic s5 ,c5; 
    fa fa5 (pp0[5], pp1[4], pp2[3], s5, c5);
    logic s6 ,c6; 
    fa fa6 (pp3[2], pp4[1], pp5[0], s6, c6);
    logic s7 ,c7; 
    fa fa7 (pp0[6], pp1[5], pp2[4], s7, c7);
    logic s8 ,c8; 
    fa fa8 (pp3[3], pp4[2], pp5[1], s8, c8);
    logic s9 ,c9; 
    fa fa9 (pp0[7], pp1[6], pp2[5], s9, c9);
    logic s10 ,c10; 
    fa fa10 (pp3[4], pp4[3], pp5[2], s10, c10);
    logic s11 ,c11;
    ha ha11 (pp6[1], pp7[0], s11, c11);
    logic s12 ,c12; 
    fa fa12 (pp1[7], pp2[6], pp3[5], s12, c12);
    logic s13 ,c13; 
    fa fa13 (pp4[4], pp5[3], pp6[2], s13, c13);
    logic s14 ,c14; 
    fa fa14 (pp2[7], pp3[6], pp4[5], s14, c14);
    logic s15 ,c15; 
    fa fa15 (pp5[4], pp6[3], pp7[2], s15, c15);
    logic s16 ,c16; 
    fa fa16 (pp3[7], pp4[6], pp5[5], s16, c16);
    logic s17 ,c17;
    ha ha17 (pp6[4], pp7[3], s17, c17);
    logic s18 ,c18; 
    fa fa18 (pp4[7], pp5[6], pp6[5], s18, c18);
    logic s19 ,c19; 
    fa fa19 (pp5[7], pp6[6], pp7[5], s19, c19);
    logic s20 ,c20;
    ha ha20 (pp6[7], pp7[6], s20, c20);
    
    // Wallace Summation Stage 2
    logic s21 ,c21;
    ha ha21 (c0, s1, s21, c21);
    logic s22 ,c22; 
    fa fa22 (pp3[0], c1, s2, s22, c22);
    logic s23 ,c23; 
    fa fa23 (c2, s3, s4, s23, c23);
    logic s24 ,c24; 
    fa fa24 (c3, c4, s5, s24, c24);
    logic s25 ,c25; 
    fa fa25 (pp6[0], c5, c6, s25, c25);
    logic s26 ,c26;
    ha ha26 (s7, s8, s26, c26);
    logic s27 ,c27; 
    fa fa27 (c7, c8, s9, s27, c27);
    logic s28 ,c28;
    ha ha28 (s10, s11, s28, c28);
    logic s29 ,c29; 
    fa fa29 (pp7[1], c9, c10, s29, c29);
    logic s30 ,c30; 
    fa fa30 (c11, s12, s13, s30, c30);
    logic s31 ,c31; 
    fa fa31 (c12, c13, s14, s31, c31);
    logic s32 ,c32; 
    fa fa32 (c14, c15, s16, s32, c32);
    logic s33 ,c33; 
    fa fa33 (pp7[4], c16, c17, s33, c33);
    logic s34 ,c34;
    ha ha34 (c18, s19, s34, c34);
    logic s35 ,c35;
    ha ha35 (c19, s20, s35, c35);
    logic s36 ,c36;
    ha ha36 (pp7[7], c20, s36, c36);
    
    // Wallace Summation Stage 3
    logic s37 ,c37;
    ha ha37 (c21, s22, s37, c37);
    logic s38 ,c38;
    ha ha38 (c22, s23, s38, c38);
    logic s39 ,c39; 
    fa fa39 (s6, c23, s24, s39, c39);
    logic s40 ,c40; 
    fa fa40 (c24, s25, s26, s40, c40);
    logic s41 ,c41; 
    fa fa41 (c25, c26, s27, s41, c41);
    logic s42 ,c42; 
    fa fa42 (c27, c28, s29, s42, c42);
    logic s43 ,c43; 
    fa fa43 (s15, c29, c30, s43, c43);
    logic s44 ,c44; 
    fa fa44 (s17, c31, s32, s44, c44);
    logic s45 ,c45; 
    fa fa45 (s18, c32, s33, s45, c45);
    logic s46 ,c46;
    ha ha46 (c33, s34, s46, c46);
    logic s47 ,c47;
    ha ha47 (c34, s35, s47, c47);
    logic s48 ,c48;
    ha ha48 (c35, s36, s48, c48);
    
    // Wallace Summation Stage 4
    logic s49 ,c49;
    ha ha49 (c37, s38, s49, c49);
    logic s50 ,c50;
    ha ha50 (c38, s39, s50, c50);
    logic s51 ,c51;
    ha ha51 (c39, s40, s51, c51);
    logic s52 ,c52; 
    fa fa52 (s28, c40, s41, s52, c52);
    logic s53 ,c53; 
    fa fa53 (s30, c41, s42, s53, c53);
    logic s54 ,c54; 
    fa fa54 (s31, c42, s43, s54, c54);
    logic s55 ,c55;
    ha ha55 (c43, s44, s55, c55);
    logic s56 ,c56;
    ha ha56 (c44, s45, s56, c56);
    logic s57 ,c57;
    ha ha57 (c45, s46, s57, c57);
    logic s58 ,c58;
    ha ha58 (c46, s47, s58, c58);
    logic s59 ,c59;
    ha ha59 (c47, s48, s59, c59);
    logic s60 ,c60;
    ha ha60 (c36, c48, s60, c60);
    
    assign result[0] = pp0[0];
    assign result[1] = s0;
    assign result[2] = s21;
    assign result[3] = s37;
    assign result[4] = s49;
    logic [11:0] adder_result;
    KS_11 final_adder ({c59, c58, c57, c56, c55, c54, c53, c52, c51, c50, c49 }, {s60, s59, s58, s57, s56, s55, s54, s53, s52, s51, s50 }, adder_result );
    assign result[15:5] = adder_result[10:0];
endmodule



module KS_11 ( 
        input logic [10:0] IN1,
        input logic [10:0] IN2,
        output logic [11:0] OUT);
    
    wire logic [10:0] p_0;
    wire logic [10:0] g_0;
    assign g_0 = IN1 & IN2;
    assign p_0 = IN1 ^ IN2;
    
// Kogge-Stone Adder 

    
    // KS stage 1
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_2;
    wire logic g_1_2;
    assign p_1_2 = p_0[2] & p_0[1];
    assign g_1_2 = (p_0[2] & g_0[1]) | g_0[2];
    wire logic p_1_3;
    wire logic g_1_3;
    assign p_1_3 = p_0[3] & p_0[2];
    assign g_1_3 = (p_0[3] & g_0[2]) | g_0[3];
    wire logic p_1_4;
    wire logic g_1_4;
    assign p_1_4 = p_0[4] & p_0[3];
    assign g_1_4 = (p_0[4] & g_0[3]) | g_0[4];
    wire logic p_1_5;
    wire logic g_1_5;
    assign p_1_5 = p_0[5] & p_0[4];
    assign g_1_5 = (p_0[5] & g_0[4]) | g_0[5];
    wire logic p_1_6;
    wire logic g_1_6;
    assign p_1_6 = p_0[6] & p_0[5];
    assign g_1_6 = (p_0[6] & g_0[5]) | g_0[6];
    wire logic p_1_7;
    wire logic g_1_7;
    assign p_1_7 = p_0[7] & p_0[6];
    assign g_1_7 = (p_0[7] & g_0[6]) | g_0[7];
    wire logic p_1_8;
    wire logic g_1_8;
    assign p_1_8 = p_0[8] & p_0[7];
    assign g_1_8 = (p_0[8] & g_0[7]) | g_0[8];
    wire logic p_1_9;
    wire logic g_1_9;
    assign p_1_9 = p_0[9] & p_0[8];
    assign g_1_9 = (p_0[9] & g_0[8]) | g_0[9];
    wire logic p_1_10;
    wire logic g_1_10;
    assign p_1_10 = p_0[10] & p_0[9];
    assign g_1_10 = (p_0[10] & g_0[9]) | g_0[10];
    
    // KS stage 2
    wire logic p_2_2;
    wire logic g_2_2;
    assign p_2_2 = p_1_2 & p_0[0];
    assign g_2_2 = (p_1_2 & g_0[0]) | g_1_2;
    wire logic p_2_3;
    wire logic g_2_3;
    assign p_2_3 = p_1_3 & p_1_1;
    assign g_2_3 = (p_1_3 & g_1_1) | g_1_3;
    wire logic p_2_4;
    wire logic g_2_4;
    assign p_2_4 = p_1_4 & p_1_2;
    assign g_2_4 = (p_1_4 & g_1_2) | g_1_4;
    wire logic p_2_5;
    wire logic g_2_5;
    assign p_2_5 = p_1_5 & p_1_3;
    assign g_2_5 = (p_1_5 & g_1_3) | g_1_5;
    wire logic p_2_6;
    wire logic g_2_6;
    assign p_2_6 = p_1_6 & p_1_4;
    assign g_2_6 = (p_1_6 & g_1_4) | g_1_6;
    wire logic p_2_7;
    wire logic g_2_7;
    assign p_2_7 = p_1_7 & p_1_5;
    assign g_2_7 = (p_1_7 & g_1_5) | g_1_7;
    wire logic p_2_8;
    wire logic g_2_8;
    assign p_2_8 = p_1_8 & p_1_6;
    assign g_2_8 = (p_1_8 & g_1_6) | g_1_8;
    wire logic p_2_9;
    wire logic g_2_9;
    assign p_2_9 = p_1_9 & p_1_7;
    assign g_2_9 = (p_1_9 & g_1_7) | g_1_9;
    wire logic p_2_10;
    wire logic g_2_10;
    assign p_2_10 = p_1_10 & p_1_8;
    assign g_2_10 = (p_1_10 & g_1_8) | g_1_10;
    
    // KS stage 3
    wire logic p_3_4;
    wire logic g_3_4;
    assign p_3_4 = p_2_4 & p_0[0];
    assign g_3_4 = (p_2_4 & g_0[0]) | g_2_4;
    wire logic p_3_5;
    wire logic g_3_5;
    assign p_3_5 = p_2_5 & p_1_1;
    assign g_3_5 = (p_2_5 & g_1_1) | g_2_5;
    wire logic p_3_6;
    wire logic g_3_6;
    assign p_3_6 = p_2_6 & p_2_2;
    assign g_3_6 = (p_2_6 & g_2_2) | g_2_6;
    wire logic p_3_7;
    wire logic g_3_7;
    assign p_3_7 = p_2_7 & p_2_3;
    assign g_3_7 = (p_2_7 & g_2_3) | g_2_7;
    wire logic p_3_8;
    wire logic g_3_8;
    assign p_3_8 = p_2_8 & p_2_4;
    assign g_3_8 = (p_2_8 & g_2_4) | g_2_8;
    wire logic p_3_9;
    wire logic g_3_9;
    assign p_3_9 = p_2_9 & p_2_5;
    assign g_3_9 = (p_2_9 & g_2_5) | g_2_9;
    wire logic p_3_10;
    wire logic g_3_10;
    assign p_3_10 = p_2_10 & p_2_6;
    assign g_3_10 = (p_2_10 & g_2_6) | g_2_10;
    
    // KS stage 4
    wire logic p_4_8;
    wire logic g_4_8;
    assign p_4_8 = p_3_8 & p_0[0];
    assign g_4_8 = (p_3_8 & g_0[0]) | g_3_8;
    wire logic p_4_9;
    wire logic g_4_9;
    assign p_4_9 = p_3_9 & p_1_1;
    assign g_4_9 = (p_3_9 & g_1_1) | g_3_9;
    wire logic p_4_10;
    wire logic g_4_10;
    assign p_4_10 = p_3_10 & p_2_2;
    assign g_4_10 = (p_3_10 & g_2_2) | g_3_10;
    
    // KS postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = p_0[3] ^ g_2_2;
    assign OUT[4] = p_0[4] ^ g_2_3;
    assign OUT[5] = p_0[5] ^ g_3_4;
    assign OUT[6] = p_0[6] ^ g_3_5;
    assign OUT[7] = p_0[7] ^ g_3_6;
    assign OUT[8] = p_0[8] ^ g_3_7;
    assign OUT[9] = p_0[9] ^ g_4_8;
    assign OUT[10] = p_0[10] ^ g_4_9;
    assign OUT[11] = g_4_10;
endmodule

module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule

module Four2Two 
        #(parameter WIDTH=1) (
        input logic [WIDTH-1:0] in1,
        input logic [WIDTH-1:0] in2,
        input logic [WIDTH-1:0] in3,
        input logic [WIDTH-1:0] in4,
        input logic cin,
        output logic [WIDTH-1:0] sum,
        output logic [WIDTH-1:0] carry,
        output logic cout);
    
    wire logic [WIDTH:0] temp1;
    assign temp1 = {((in1 ^ in2)&in3 | in1 & ~(in1^in2)),cin};
    assign sum = ((in1 ^ in2) ^ in3 ^ in4) ^ temp1[WIDTH-1:0];
    assign carry = ((in1 ^ in2) ^ in3 ^ in4) & temp1[WIDTH-1:0] | in4 & ~((in1 ^ in2) ^ in3 ^ in4);
    assign cout = temp1[WIDTH];
endmodule




