module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, out1);
  input [6:0] in1, in2, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31;
  input in3, in4;
  output [12:0] out1;
  wire [6:0] in1, in2, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31;
  wire in3, in4;
  wire [12:0] out1;
  wire csa_tree_sub001036_groupi_n_0, csa_tree_sub001036_groupi_n_1, csa_tree_sub001036_groupi_n_2, csa_tree_sub001036_groupi_n_3, csa_tree_sub001036_groupi_n_4, csa_tree_sub001036_groupi_n_5, csa_tree_sub001036_groupi_n_8, csa_tree_sub001036_groupi_n_9;
  wire csa_tree_sub001036_groupi_n_10, csa_tree_sub001036_groupi_n_11, csa_tree_sub001036_groupi_n_12, csa_tree_sub001036_groupi_n_13, csa_tree_sub001036_groupi_n_14, csa_tree_sub001036_groupi_n_15, csa_tree_sub001036_groupi_n_16, csa_tree_sub001036_groupi_n_17;
  wire csa_tree_sub001036_groupi_n_18, csa_tree_sub001036_groupi_n_19, csa_tree_sub001036_groupi_n_20, csa_tree_sub001036_groupi_n_21, csa_tree_sub001036_groupi_n_22, csa_tree_sub001036_groupi_n_23, csa_tree_sub001036_groupi_n_24, csa_tree_sub001036_groupi_n_25;
  wire csa_tree_sub001036_groupi_n_26, csa_tree_sub001036_groupi_n_27, csa_tree_sub001036_groupi_n_28, csa_tree_sub001036_groupi_n_29, csa_tree_sub001036_groupi_n_30, csa_tree_sub001036_groupi_n_31, csa_tree_sub001036_groupi_n_32, csa_tree_sub001036_groupi_n_33;
  wire csa_tree_sub001036_groupi_n_34, csa_tree_sub001036_groupi_n_35, csa_tree_sub001036_groupi_n_36, csa_tree_sub001036_groupi_n_37, csa_tree_sub001036_groupi_n_38, csa_tree_sub001036_groupi_n_39, csa_tree_sub001036_groupi_n_40, csa_tree_sub001036_groupi_n_41;
  wire csa_tree_sub001036_groupi_n_42, csa_tree_sub001036_groupi_n_43, csa_tree_sub001036_groupi_n_44, csa_tree_sub001036_groupi_n_45, csa_tree_sub001036_groupi_n_46, csa_tree_sub001036_groupi_n_47, csa_tree_sub001036_groupi_n_48, csa_tree_sub001036_groupi_n_49;
  wire csa_tree_sub001036_groupi_n_50, csa_tree_sub001036_groupi_n_51, csa_tree_sub001036_groupi_n_52, csa_tree_sub001036_groupi_n_53, csa_tree_sub001036_groupi_n_54, csa_tree_sub001036_groupi_n_55, csa_tree_sub001036_groupi_n_56, csa_tree_sub001036_groupi_n_57;
  wire csa_tree_sub001036_groupi_n_58, csa_tree_sub001036_groupi_n_59, csa_tree_sub001036_groupi_n_60, csa_tree_sub001036_groupi_n_61, csa_tree_sub001036_groupi_n_62, csa_tree_sub001036_groupi_n_63, csa_tree_sub001036_groupi_n_64, csa_tree_sub001036_groupi_n_65;
  wire csa_tree_sub001036_groupi_n_66, csa_tree_sub001036_groupi_n_67, csa_tree_sub001036_groupi_n_68, csa_tree_sub001036_groupi_n_69, csa_tree_sub001036_groupi_n_70, csa_tree_sub001036_groupi_n_71, csa_tree_sub001036_groupi_n_72, csa_tree_sub001036_groupi_n_73;
  wire csa_tree_sub001036_groupi_n_74, csa_tree_sub001036_groupi_n_75, csa_tree_sub001036_groupi_n_76, csa_tree_sub001036_groupi_n_77, csa_tree_sub001036_groupi_n_78, csa_tree_sub001036_groupi_n_79, csa_tree_sub001036_groupi_n_80, csa_tree_sub001036_groupi_n_81;
  wire csa_tree_sub001036_groupi_n_82, csa_tree_sub001036_groupi_n_83, csa_tree_sub001036_groupi_n_84, csa_tree_sub001036_groupi_n_85, csa_tree_sub001036_groupi_n_86, csa_tree_sub001036_groupi_n_87, csa_tree_sub001036_groupi_n_88, csa_tree_sub001036_groupi_n_89;
  wire csa_tree_sub001036_groupi_n_90, csa_tree_sub001036_groupi_n_91, csa_tree_sub001036_groupi_n_92, csa_tree_sub001036_groupi_n_93, csa_tree_sub001036_groupi_n_94, csa_tree_sub001036_groupi_n_95, csa_tree_sub001036_groupi_n_96, csa_tree_sub001036_groupi_n_97;
  wire csa_tree_sub001036_groupi_n_98, csa_tree_sub001036_groupi_n_99, csa_tree_sub001036_groupi_n_100, csa_tree_sub001036_groupi_n_101, csa_tree_sub001036_groupi_n_102, csa_tree_sub001036_groupi_n_103, csa_tree_sub001036_groupi_n_104, csa_tree_sub001036_groupi_n_105;
  wire csa_tree_sub001036_groupi_n_106, csa_tree_sub001036_groupi_n_107, csa_tree_sub001036_groupi_n_108, csa_tree_sub001036_groupi_n_109, csa_tree_sub001036_groupi_n_110, csa_tree_sub001036_groupi_n_111, csa_tree_sub001036_groupi_n_112, csa_tree_sub001036_groupi_n_113;
  wire csa_tree_sub001036_groupi_n_114, csa_tree_sub001036_groupi_n_115, csa_tree_sub001036_groupi_n_116, csa_tree_sub001036_groupi_n_117, csa_tree_sub001036_groupi_n_118, csa_tree_sub001036_groupi_n_119, csa_tree_sub001036_groupi_n_120, csa_tree_sub001036_groupi_n_121;
  wire csa_tree_sub001036_groupi_n_122, csa_tree_sub001036_groupi_n_123, csa_tree_sub001036_groupi_n_124, csa_tree_sub001036_groupi_n_125, csa_tree_sub001036_groupi_n_126, csa_tree_sub001036_groupi_n_127, csa_tree_sub001036_groupi_n_128, csa_tree_sub001036_groupi_n_129;
  wire csa_tree_sub001036_groupi_n_130, csa_tree_sub001036_groupi_n_131, csa_tree_sub001036_groupi_n_132, csa_tree_sub001036_groupi_n_133, csa_tree_sub001036_groupi_n_134, csa_tree_sub001036_groupi_n_135, csa_tree_sub001036_groupi_n_136, csa_tree_sub001036_groupi_n_137;
  wire csa_tree_sub001036_groupi_n_138, csa_tree_sub001036_groupi_n_139, csa_tree_sub001036_groupi_n_140, csa_tree_sub001036_groupi_n_141, csa_tree_sub001036_groupi_n_142, csa_tree_sub001036_groupi_n_143, csa_tree_sub001036_groupi_n_144, csa_tree_sub001036_groupi_n_145;
  wire csa_tree_sub001036_groupi_n_146, csa_tree_sub001036_groupi_n_147, csa_tree_sub001036_groupi_n_148, csa_tree_sub001036_groupi_n_149, csa_tree_sub001036_groupi_n_150, csa_tree_sub001036_groupi_n_151, csa_tree_sub001036_groupi_n_152, csa_tree_sub001036_groupi_n_153;
  wire csa_tree_sub001036_groupi_n_154, csa_tree_sub001036_groupi_n_155, csa_tree_sub001036_groupi_n_156, csa_tree_sub001036_groupi_n_157, csa_tree_sub001036_groupi_n_158, csa_tree_sub001036_groupi_n_159, csa_tree_sub001036_groupi_n_160, csa_tree_sub001036_groupi_n_161;
  wire csa_tree_sub001036_groupi_n_162, csa_tree_sub001036_groupi_n_163, csa_tree_sub001036_groupi_n_164, csa_tree_sub001036_groupi_n_165, csa_tree_sub001036_groupi_n_166, csa_tree_sub001036_groupi_n_167, csa_tree_sub001036_groupi_n_168, csa_tree_sub001036_groupi_n_169;
  wire csa_tree_sub001036_groupi_n_170, csa_tree_sub001036_groupi_n_171, csa_tree_sub001036_groupi_n_172, csa_tree_sub001036_groupi_n_173, csa_tree_sub001036_groupi_n_174, csa_tree_sub001036_groupi_n_175, csa_tree_sub001036_groupi_n_176, csa_tree_sub001036_groupi_n_177;
  wire csa_tree_sub001036_groupi_n_178, csa_tree_sub001036_groupi_n_179, csa_tree_sub001036_groupi_n_180, csa_tree_sub001036_groupi_n_181, csa_tree_sub001036_groupi_n_182, csa_tree_sub001036_groupi_n_183, csa_tree_sub001036_groupi_n_184, csa_tree_sub001036_groupi_n_185;
  wire csa_tree_sub001036_groupi_n_186, csa_tree_sub001036_groupi_n_187, csa_tree_sub001036_groupi_n_188, csa_tree_sub001036_groupi_n_189, csa_tree_sub001036_groupi_n_190, csa_tree_sub001036_groupi_n_191, csa_tree_sub001036_groupi_n_192, csa_tree_sub001036_groupi_n_193;
  wire csa_tree_sub001036_groupi_n_194, csa_tree_sub001036_groupi_n_195, csa_tree_sub001036_groupi_n_196, csa_tree_sub001036_groupi_n_197, csa_tree_sub001036_groupi_n_198, csa_tree_sub001036_groupi_n_199, csa_tree_sub001036_groupi_n_200, csa_tree_sub001036_groupi_n_201;
  wire csa_tree_sub001036_groupi_n_202, csa_tree_sub001036_groupi_n_203, csa_tree_sub001036_groupi_n_204, csa_tree_sub001036_groupi_n_205, csa_tree_sub001036_groupi_n_206, csa_tree_sub001036_groupi_n_207, csa_tree_sub001036_groupi_n_208, csa_tree_sub001036_groupi_n_209;
  wire csa_tree_sub001036_groupi_n_210, csa_tree_sub001036_groupi_n_211, csa_tree_sub001036_groupi_n_212, csa_tree_sub001036_groupi_n_213, csa_tree_sub001036_groupi_n_214, csa_tree_sub001036_groupi_n_215, csa_tree_sub001036_groupi_n_216, csa_tree_sub001036_groupi_n_217;
  wire csa_tree_sub001036_groupi_n_218, csa_tree_sub001036_groupi_n_219, csa_tree_sub001036_groupi_n_220, csa_tree_sub001036_groupi_n_221, csa_tree_sub001036_groupi_n_222, csa_tree_sub001036_groupi_n_223, csa_tree_sub001036_groupi_n_224, csa_tree_sub001036_groupi_n_225;
  wire csa_tree_sub001036_groupi_n_226, csa_tree_sub001036_groupi_n_227, csa_tree_sub001036_groupi_n_228, csa_tree_sub001036_groupi_n_229, csa_tree_sub001036_groupi_n_230, csa_tree_sub001036_groupi_n_231, csa_tree_sub001036_groupi_n_232, csa_tree_sub001036_groupi_n_233;
  wire csa_tree_sub001036_groupi_n_234, csa_tree_sub001036_groupi_n_235, csa_tree_sub001036_groupi_n_236, csa_tree_sub001036_groupi_n_237, csa_tree_sub001036_groupi_n_238, csa_tree_sub001036_groupi_n_239, csa_tree_sub001036_groupi_n_240, csa_tree_sub001036_groupi_n_241;
  wire csa_tree_sub001036_groupi_n_242, csa_tree_sub001036_groupi_n_243, csa_tree_sub001036_groupi_n_244, csa_tree_sub001036_groupi_n_245, csa_tree_sub001036_groupi_n_246, csa_tree_sub001036_groupi_n_247, csa_tree_sub001036_groupi_n_248, csa_tree_sub001036_groupi_n_249;
  wire csa_tree_sub001036_groupi_n_250, csa_tree_sub001036_groupi_n_251, csa_tree_sub001036_groupi_n_252, csa_tree_sub001036_groupi_n_253, csa_tree_sub001036_groupi_n_254, csa_tree_sub001036_groupi_n_255, csa_tree_sub001036_groupi_n_256, csa_tree_sub001036_groupi_n_257;
  wire csa_tree_sub001036_groupi_n_258, csa_tree_sub001036_groupi_n_259, csa_tree_sub001036_groupi_n_260, csa_tree_sub001036_groupi_n_261, csa_tree_sub001036_groupi_n_262, csa_tree_sub001036_groupi_n_263, csa_tree_sub001036_groupi_n_264, csa_tree_sub001036_groupi_n_265;
  wire csa_tree_sub001036_groupi_n_266, csa_tree_sub001036_groupi_n_267, csa_tree_sub001036_groupi_n_268, csa_tree_sub001036_groupi_n_269, csa_tree_sub001036_groupi_n_270, csa_tree_sub001036_groupi_n_271, csa_tree_sub001036_groupi_n_272, csa_tree_sub001036_groupi_n_273;
  wire csa_tree_sub001036_groupi_n_274, csa_tree_sub001036_groupi_n_275, csa_tree_sub001036_groupi_n_276, csa_tree_sub001036_groupi_n_277, csa_tree_sub001036_groupi_n_278, csa_tree_sub001036_groupi_n_279, csa_tree_sub001036_groupi_n_280, csa_tree_sub001036_groupi_n_281;
  wire csa_tree_sub001036_groupi_n_282, csa_tree_sub001036_groupi_n_283, csa_tree_sub001036_groupi_n_284, csa_tree_sub001036_groupi_n_285, csa_tree_sub001036_groupi_n_286, csa_tree_sub001036_groupi_n_287, csa_tree_sub001036_groupi_n_288, csa_tree_sub001036_groupi_n_289;
  wire csa_tree_sub001036_groupi_n_290, csa_tree_sub001036_groupi_n_291, csa_tree_sub001036_groupi_n_292, csa_tree_sub001036_groupi_n_293, csa_tree_sub001036_groupi_n_294, csa_tree_sub001036_groupi_n_295, csa_tree_sub001036_groupi_n_296, csa_tree_sub001036_groupi_n_297;
  wire csa_tree_sub001036_groupi_n_298, csa_tree_sub001036_groupi_n_299, csa_tree_sub001036_groupi_n_300, csa_tree_sub001036_groupi_n_301, csa_tree_sub001036_groupi_n_302, csa_tree_sub001036_groupi_n_303, csa_tree_sub001036_groupi_n_304, csa_tree_sub001036_groupi_n_305;
  wire csa_tree_sub001036_groupi_n_306, csa_tree_sub001036_groupi_n_307, csa_tree_sub001036_groupi_n_308, csa_tree_sub001036_groupi_n_309, csa_tree_sub001036_groupi_n_310, csa_tree_sub001036_groupi_n_311, csa_tree_sub001036_groupi_n_312, csa_tree_sub001036_groupi_n_313;
  wire csa_tree_sub001036_groupi_n_314, csa_tree_sub001036_groupi_n_315, csa_tree_sub001036_groupi_n_316, csa_tree_sub001036_groupi_n_317, csa_tree_sub001036_groupi_n_318, csa_tree_sub001036_groupi_n_319, csa_tree_sub001036_groupi_n_320, csa_tree_sub001036_groupi_n_321;
  wire csa_tree_sub001036_groupi_n_322, csa_tree_sub001036_groupi_n_323, csa_tree_sub001036_groupi_n_324, csa_tree_sub001036_groupi_n_325, csa_tree_sub001036_groupi_n_326, csa_tree_sub001036_groupi_n_327, csa_tree_sub001036_groupi_n_328, csa_tree_sub001036_groupi_n_329;
  wire csa_tree_sub001036_groupi_n_330, csa_tree_sub001036_groupi_n_331, csa_tree_sub001036_groupi_n_332, csa_tree_sub001036_groupi_n_333, csa_tree_sub001036_groupi_n_334, csa_tree_sub001036_groupi_n_335, csa_tree_sub001036_groupi_n_336, csa_tree_sub001036_groupi_n_337;
  wire csa_tree_sub001036_groupi_n_338, csa_tree_sub001036_groupi_n_339, csa_tree_sub001036_groupi_n_340, csa_tree_sub001036_groupi_n_341, csa_tree_sub001036_groupi_n_342, csa_tree_sub001036_groupi_n_343, csa_tree_sub001036_groupi_n_344, csa_tree_sub001036_groupi_n_345;
  wire csa_tree_sub001036_groupi_n_346, csa_tree_sub001036_groupi_n_347, csa_tree_sub001036_groupi_n_348, csa_tree_sub001036_groupi_n_349, csa_tree_sub001036_groupi_n_350, csa_tree_sub001036_groupi_n_351, csa_tree_sub001036_groupi_n_352, csa_tree_sub001036_groupi_n_353;
  wire csa_tree_sub001036_groupi_n_354, csa_tree_sub001036_groupi_n_355, csa_tree_sub001036_groupi_n_356, csa_tree_sub001036_groupi_n_357, csa_tree_sub001036_groupi_n_358, csa_tree_sub001036_groupi_n_359, csa_tree_sub001036_groupi_n_360, csa_tree_sub001036_groupi_n_361;
  wire csa_tree_sub001036_groupi_n_362, csa_tree_sub001036_groupi_n_363, csa_tree_sub001036_groupi_n_364, csa_tree_sub001036_groupi_n_365, csa_tree_sub001036_groupi_n_366, csa_tree_sub001036_groupi_n_367, csa_tree_sub001036_groupi_n_368, csa_tree_sub001036_groupi_n_369;
  wire csa_tree_sub001036_groupi_n_370, csa_tree_sub001036_groupi_n_371, csa_tree_sub001036_groupi_n_372, csa_tree_sub001036_groupi_n_373, csa_tree_sub001036_groupi_n_374, csa_tree_sub001036_groupi_n_375, csa_tree_sub001036_groupi_n_376, csa_tree_sub001036_groupi_n_377;
  wire csa_tree_sub001036_groupi_n_378, csa_tree_sub001036_groupi_n_379, csa_tree_sub001036_groupi_n_380, csa_tree_sub001036_groupi_n_381, csa_tree_sub001036_groupi_n_382, csa_tree_sub001036_groupi_n_383, csa_tree_sub001036_groupi_n_384, csa_tree_sub001036_groupi_n_385;
  wire csa_tree_sub001036_groupi_n_386, csa_tree_sub001036_groupi_n_387, csa_tree_sub001036_groupi_n_388, csa_tree_sub001036_groupi_n_389, csa_tree_sub001036_groupi_n_390, csa_tree_sub001036_groupi_n_391, csa_tree_sub001036_groupi_n_392, csa_tree_sub001036_groupi_n_393;
  wire csa_tree_sub001036_groupi_n_394, csa_tree_sub001036_groupi_n_395, csa_tree_sub001036_groupi_n_396, csa_tree_sub001036_groupi_n_397, csa_tree_sub001036_groupi_n_398, csa_tree_sub001036_groupi_n_399, csa_tree_sub001036_groupi_n_400, csa_tree_sub001036_groupi_n_401;
  wire csa_tree_sub001036_groupi_n_402, csa_tree_sub001036_groupi_n_403, csa_tree_sub001036_groupi_n_404, csa_tree_sub001036_groupi_n_405, csa_tree_sub001036_groupi_n_406, csa_tree_sub001036_groupi_n_407, csa_tree_sub001036_groupi_n_408, csa_tree_sub001036_groupi_n_409;
  wire csa_tree_sub001036_groupi_n_410, csa_tree_sub001036_groupi_n_411, csa_tree_sub001036_groupi_n_412, csa_tree_sub001036_groupi_n_413, csa_tree_sub001036_groupi_n_414, csa_tree_sub001036_groupi_n_415, csa_tree_sub001036_groupi_n_416, csa_tree_sub001036_groupi_n_417;
  wire csa_tree_sub001036_groupi_n_418, csa_tree_sub001036_groupi_n_419, csa_tree_sub001036_groupi_n_420, csa_tree_sub001036_groupi_n_421, csa_tree_sub001036_groupi_n_422, csa_tree_sub001036_groupi_n_423, csa_tree_sub001036_groupi_n_424, csa_tree_sub001036_groupi_n_425;
  wire csa_tree_sub001036_groupi_n_426, csa_tree_sub001036_groupi_n_427, csa_tree_sub001036_groupi_n_428, csa_tree_sub001036_groupi_n_429, csa_tree_sub001036_groupi_n_430, csa_tree_sub001036_groupi_n_431, csa_tree_sub001036_groupi_n_432, csa_tree_sub001036_groupi_n_433;
  wire csa_tree_sub001036_groupi_n_434, csa_tree_sub001036_groupi_n_435, csa_tree_sub001036_groupi_n_436, csa_tree_sub001036_groupi_n_437, csa_tree_sub001036_groupi_n_438, csa_tree_sub001036_groupi_n_439, csa_tree_sub001036_groupi_n_440, csa_tree_sub001036_groupi_n_441;
  wire csa_tree_sub001036_groupi_n_442, csa_tree_sub001036_groupi_n_443, csa_tree_sub001036_groupi_n_444, csa_tree_sub001036_groupi_n_445, csa_tree_sub001036_groupi_n_446, csa_tree_sub001036_groupi_n_447, csa_tree_sub001036_groupi_n_448, csa_tree_sub001036_groupi_n_449;
  wire csa_tree_sub001036_groupi_n_450, csa_tree_sub001036_groupi_n_451, csa_tree_sub001036_groupi_n_452, csa_tree_sub001036_groupi_n_453, csa_tree_sub001036_groupi_n_454, csa_tree_sub001036_groupi_n_455, csa_tree_sub001036_groupi_n_456, csa_tree_sub001036_groupi_n_457;
  wire csa_tree_sub001036_groupi_n_458, csa_tree_sub001036_groupi_n_459, csa_tree_sub001036_groupi_n_460, csa_tree_sub001036_groupi_n_461, csa_tree_sub001036_groupi_n_462, csa_tree_sub001036_groupi_n_463, csa_tree_sub001036_groupi_n_464, csa_tree_sub001036_groupi_n_465;
  wire csa_tree_sub001036_groupi_n_466, csa_tree_sub001036_groupi_n_467, csa_tree_sub001036_groupi_n_468, csa_tree_sub001036_groupi_n_469, csa_tree_sub001036_groupi_n_470, csa_tree_sub001036_groupi_n_471, csa_tree_sub001036_groupi_n_472, csa_tree_sub001036_groupi_n_473;
  wire csa_tree_sub001036_groupi_n_474, csa_tree_sub001036_groupi_n_475, csa_tree_sub001036_groupi_n_476, csa_tree_sub001036_groupi_n_477, csa_tree_sub001036_groupi_n_478, csa_tree_sub001036_groupi_n_479, csa_tree_sub001036_groupi_n_480, csa_tree_sub001036_groupi_n_481;
  wire csa_tree_sub001036_groupi_n_482, csa_tree_sub001036_groupi_n_483, csa_tree_sub001036_groupi_n_484, csa_tree_sub001036_groupi_n_485, csa_tree_sub001036_groupi_n_486, csa_tree_sub001036_groupi_n_487, csa_tree_sub001036_groupi_n_488, csa_tree_sub001036_groupi_n_489;
  wire csa_tree_sub001036_groupi_n_490, csa_tree_sub001036_groupi_n_491, csa_tree_sub001036_groupi_n_492, csa_tree_sub001036_groupi_n_493, csa_tree_sub001036_groupi_n_494, csa_tree_sub001036_groupi_n_495, csa_tree_sub001036_groupi_n_496, csa_tree_sub001036_groupi_n_497;
  wire csa_tree_sub001036_groupi_n_498, csa_tree_sub001036_groupi_n_499, csa_tree_sub001036_groupi_n_500, csa_tree_sub001036_groupi_n_501, csa_tree_sub001036_groupi_n_502, csa_tree_sub001036_groupi_n_503, csa_tree_sub001036_groupi_n_504, csa_tree_sub001036_groupi_n_505;
  wire csa_tree_sub001036_groupi_n_506, csa_tree_sub001036_groupi_n_507, csa_tree_sub001036_groupi_n_508, csa_tree_sub001036_groupi_n_509, csa_tree_sub001036_groupi_n_510, csa_tree_sub001036_groupi_n_511, csa_tree_sub001036_groupi_n_512, csa_tree_sub001036_groupi_n_513;
  wire csa_tree_sub001036_groupi_n_514, csa_tree_sub001036_groupi_n_515, csa_tree_sub001036_groupi_n_516, csa_tree_sub001036_groupi_n_517, csa_tree_sub001036_groupi_n_518, csa_tree_sub001036_groupi_n_519, csa_tree_sub001036_groupi_n_520, csa_tree_sub001036_groupi_n_521;
  wire csa_tree_sub001036_groupi_n_522, csa_tree_sub001036_groupi_n_523, csa_tree_sub001036_groupi_n_524, csa_tree_sub001036_groupi_n_525, csa_tree_sub001036_groupi_n_526, csa_tree_sub001036_groupi_n_527, csa_tree_sub001036_groupi_n_528, csa_tree_sub001036_groupi_n_529;
  wire csa_tree_sub001036_groupi_n_530, csa_tree_sub001036_groupi_n_531, csa_tree_sub001036_groupi_n_532, csa_tree_sub001036_groupi_n_533, csa_tree_sub001036_groupi_n_534, csa_tree_sub001036_groupi_n_535, csa_tree_sub001036_groupi_n_536, csa_tree_sub001036_groupi_n_537;
  wire csa_tree_sub001036_groupi_n_538, csa_tree_sub001036_groupi_n_539, csa_tree_sub001036_groupi_n_540, csa_tree_sub001036_groupi_n_541, csa_tree_sub001036_groupi_n_542, csa_tree_sub001036_groupi_n_543, csa_tree_sub001036_groupi_n_544, csa_tree_sub001036_groupi_n_545;
  wire csa_tree_sub001036_groupi_n_546, csa_tree_sub001036_groupi_n_547, csa_tree_sub001036_groupi_n_548, csa_tree_sub001036_groupi_n_549, csa_tree_sub001036_groupi_n_550, csa_tree_sub001036_groupi_n_551, csa_tree_sub001036_groupi_n_552, csa_tree_sub001036_groupi_n_553;
  wire csa_tree_sub001036_groupi_n_554, csa_tree_sub001036_groupi_n_555, csa_tree_sub001036_groupi_n_556, csa_tree_sub001036_groupi_n_557, csa_tree_sub001036_groupi_n_558, csa_tree_sub001036_groupi_n_559, csa_tree_sub001036_groupi_n_560, csa_tree_sub001036_groupi_n_561;
  wire csa_tree_sub001036_groupi_n_562, csa_tree_sub001036_groupi_n_563, csa_tree_sub001036_groupi_n_564, csa_tree_sub001036_groupi_n_565, csa_tree_sub001036_groupi_n_566, csa_tree_sub001036_groupi_n_567, csa_tree_sub001036_groupi_n_568, csa_tree_sub001036_groupi_n_569;
  wire csa_tree_sub001036_groupi_n_570, csa_tree_sub001036_groupi_n_571, csa_tree_sub001036_groupi_n_572, csa_tree_sub001036_groupi_n_573, csa_tree_sub001036_groupi_n_574, csa_tree_sub001036_groupi_n_575, csa_tree_sub001036_groupi_n_576, csa_tree_sub001036_groupi_n_577;
  wire csa_tree_sub001036_groupi_n_578, csa_tree_sub001036_groupi_n_579, csa_tree_sub001036_groupi_n_580, csa_tree_sub001036_groupi_n_581, csa_tree_sub001036_groupi_n_582, csa_tree_sub001036_groupi_n_583, csa_tree_sub001036_groupi_n_584, csa_tree_sub001036_groupi_n_585;
  wire csa_tree_sub001036_groupi_n_586, csa_tree_sub001036_groupi_n_587, csa_tree_sub001036_groupi_n_588, csa_tree_sub001036_groupi_n_589, csa_tree_sub001036_groupi_n_590, csa_tree_sub001036_groupi_n_591, csa_tree_sub001036_groupi_n_592, csa_tree_sub001036_groupi_n_593;
  wire csa_tree_sub001036_groupi_n_594, csa_tree_sub001036_groupi_n_595, csa_tree_sub001036_groupi_n_596, csa_tree_sub001036_groupi_n_597, csa_tree_sub001036_groupi_n_598, csa_tree_sub001036_groupi_n_599, csa_tree_sub001036_groupi_n_600, csa_tree_sub001036_groupi_n_601;
  wire csa_tree_sub001036_groupi_n_602, csa_tree_sub001036_groupi_n_603, csa_tree_sub001036_groupi_n_604, csa_tree_sub001036_groupi_n_605, csa_tree_sub001036_groupi_n_606, csa_tree_sub001036_groupi_n_607, csa_tree_sub001036_groupi_n_608, csa_tree_sub001036_groupi_n_609;
  wire csa_tree_sub001036_groupi_n_610, csa_tree_sub001036_groupi_n_611, csa_tree_sub001036_groupi_n_612, csa_tree_sub001036_groupi_n_613, csa_tree_sub001036_groupi_n_614, csa_tree_sub001036_groupi_n_615, csa_tree_sub001036_groupi_n_616, csa_tree_sub001036_groupi_n_617;
  wire csa_tree_sub001036_groupi_n_618, csa_tree_sub001036_groupi_n_619, csa_tree_sub001036_groupi_n_620, csa_tree_sub001036_groupi_n_621, csa_tree_sub001036_groupi_n_622, csa_tree_sub001036_groupi_n_623, csa_tree_sub001036_groupi_n_624, csa_tree_sub001036_groupi_n_625;
  wire csa_tree_sub001036_groupi_n_626, csa_tree_sub001036_groupi_n_627, csa_tree_sub001036_groupi_n_628, csa_tree_sub001036_groupi_n_629, csa_tree_sub001036_groupi_n_630, csa_tree_sub001036_groupi_n_631, csa_tree_sub001036_groupi_n_632, csa_tree_sub001036_groupi_n_633;
  wire csa_tree_sub001036_groupi_n_634, csa_tree_sub001036_groupi_n_635, csa_tree_sub001036_groupi_n_636, csa_tree_sub001036_groupi_n_637, csa_tree_sub001036_groupi_n_638, csa_tree_sub001036_groupi_n_639, csa_tree_sub001036_groupi_n_640, csa_tree_sub001036_groupi_n_641;
  wire csa_tree_sub001036_groupi_n_642, csa_tree_sub001036_groupi_n_643, csa_tree_sub001036_groupi_n_644, csa_tree_sub001036_groupi_n_645, csa_tree_sub001036_groupi_n_646, csa_tree_sub001036_groupi_n_647, csa_tree_sub001036_groupi_n_648, csa_tree_sub001036_groupi_n_649;
  wire csa_tree_sub001036_groupi_n_650, csa_tree_sub001036_groupi_n_651, csa_tree_sub001036_groupi_n_652, csa_tree_sub001036_groupi_n_653, csa_tree_sub001036_groupi_n_654, csa_tree_sub001036_groupi_n_655, csa_tree_sub001036_groupi_n_656, csa_tree_sub001036_groupi_n_657;
  wire csa_tree_sub001036_groupi_n_658, csa_tree_sub001036_groupi_n_659, csa_tree_sub001036_groupi_n_660, csa_tree_sub001036_groupi_n_661, csa_tree_sub001036_groupi_n_662, csa_tree_sub001036_groupi_n_663, csa_tree_sub001036_groupi_n_664, csa_tree_sub001036_groupi_n_665;
  wire csa_tree_sub001036_groupi_n_666, csa_tree_sub001036_groupi_n_667, csa_tree_sub001036_groupi_n_668, csa_tree_sub001036_groupi_n_669, csa_tree_sub001036_groupi_n_670, csa_tree_sub001036_groupi_n_671, csa_tree_sub001036_groupi_n_672, csa_tree_sub001036_groupi_n_673;
  wire csa_tree_sub001036_groupi_n_674, csa_tree_sub001036_groupi_n_675, csa_tree_sub001036_groupi_n_676, csa_tree_sub001036_groupi_n_677, csa_tree_sub001036_groupi_n_678, csa_tree_sub001036_groupi_n_679, csa_tree_sub001036_groupi_n_680, csa_tree_sub001036_groupi_n_681;
  wire csa_tree_sub001036_groupi_n_682, csa_tree_sub001036_groupi_n_683, csa_tree_sub001036_groupi_n_684, csa_tree_sub001036_groupi_n_685, csa_tree_sub001036_groupi_n_686, csa_tree_sub001036_groupi_n_687, csa_tree_sub001036_groupi_n_688, csa_tree_sub001036_groupi_n_689;
  wire csa_tree_sub001036_groupi_n_690, csa_tree_sub001036_groupi_n_691, csa_tree_sub001036_groupi_n_692, csa_tree_sub001036_groupi_n_693, csa_tree_sub001036_groupi_n_694, csa_tree_sub001036_groupi_n_695, csa_tree_sub001036_groupi_n_696, csa_tree_sub001036_groupi_n_697;
  wire csa_tree_sub001036_groupi_n_698, csa_tree_sub001036_groupi_n_699, csa_tree_sub001036_groupi_n_700, csa_tree_sub001036_groupi_n_701, csa_tree_sub001036_groupi_n_702, csa_tree_sub001036_groupi_n_703, csa_tree_sub001036_groupi_n_704, csa_tree_sub001036_groupi_n_705;
  wire csa_tree_sub001036_groupi_n_706, csa_tree_sub001036_groupi_n_707, csa_tree_sub001036_groupi_n_708, csa_tree_sub001036_groupi_n_709, csa_tree_sub001036_groupi_n_710, csa_tree_sub001036_groupi_n_711, csa_tree_sub001036_groupi_n_712, csa_tree_sub001036_groupi_n_713;
  wire csa_tree_sub001036_groupi_n_714, csa_tree_sub001036_groupi_n_715, csa_tree_sub001036_groupi_n_716, csa_tree_sub001036_groupi_n_717, csa_tree_sub001036_groupi_n_718, csa_tree_sub001036_groupi_n_719, csa_tree_sub001036_groupi_n_720, csa_tree_sub001036_groupi_n_721;
  wire csa_tree_sub001036_groupi_n_722, csa_tree_sub001036_groupi_n_723, csa_tree_sub001036_groupi_n_724, csa_tree_sub001036_groupi_n_725, csa_tree_sub001036_groupi_n_726, csa_tree_sub001036_groupi_n_727, csa_tree_sub001036_groupi_n_728, csa_tree_sub001036_groupi_n_729;
  wire csa_tree_sub001036_groupi_n_730, csa_tree_sub001036_groupi_n_731, csa_tree_sub001036_groupi_n_732, csa_tree_sub001036_groupi_n_733, csa_tree_sub001036_groupi_n_734, csa_tree_sub001036_groupi_n_735, csa_tree_sub001036_groupi_n_736, csa_tree_sub001036_groupi_n_737;
  wire csa_tree_sub001036_groupi_n_738, csa_tree_sub001036_groupi_n_739, csa_tree_sub001036_groupi_n_740, csa_tree_sub001036_groupi_n_741, csa_tree_sub001036_groupi_n_742, csa_tree_sub001036_groupi_n_743, csa_tree_sub001036_groupi_n_744, csa_tree_sub001036_groupi_n_745;
  wire csa_tree_sub001036_groupi_n_746, csa_tree_sub001036_groupi_n_747, csa_tree_sub001036_groupi_n_748, csa_tree_sub001036_groupi_n_749, csa_tree_sub001036_groupi_n_750, csa_tree_sub001036_groupi_n_751, csa_tree_sub001036_groupi_n_752, csa_tree_sub001036_groupi_n_753;
  wire csa_tree_sub001036_groupi_n_754, csa_tree_sub001036_groupi_n_755, csa_tree_sub001036_groupi_n_756, csa_tree_sub001036_groupi_n_757, csa_tree_sub001036_groupi_n_758, csa_tree_sub001036_groupi_n_759, csa_tree_sub001036_groupi_n_760, csa_tree_sub001036_groupi_n_761;
  wire csa_tree_sub001036_groupi_n_762, csa_tree_sub001036_groupi_n_763, csa_tree_sub001036_groupi_n_764, csa_tree_sub001036_groupi_n_765, csa_tree_sub001036_groupi_n_766, csa_tree_sub001036_groupi_n_767, csa_tree_sub001036_groupi_n_768, csa_tree_sub001036_groupi_n_769;
  wire csa_tree_sub001036_groupi_n_770, csa_tree_sub001036_groupi_n_771, csa_tree_sub001036_groupi_n_772, csa_tree_sub001036_groupi_n_773, csa_tree_sub001036_groupi_n_774, csa_tree_sub001036_groupi_n_775, csa_tree_sub001036_groupi_n_776, csa_tree_sub001036_groupi_n_777;
  wire csa_tree_sub001036_groupi_n_778, csa_tree_sub001036_groupi_n_779, csa_tree_sub001036_groupi_n_780, csa_tree_sub001036_groupi_n_781, csa_tree_sub001036_groupi_n_782, csa_tree_sub001036_groupi_n_783, csa_tree_sub001036_groupi_n_784, csa_tree_sub001036_groupi_n_785;
  wire csa_tree_sub001036_groupi_n_786, csa_tree_sub001036_groupi_n_787, csa_tree_sub001036_groupi_n_789, csa_tree_sub001036_groupi_n_790, csa_tree_sub001036_groupi_n_791, csa_tree_sub001036_groupi_n_792, csa_tree_sub001036_groupi_n_793, csa_tree_sub001036_groupi_n_794;
  wire csa_tree_sub001036_groupi_n_795, csa_tree_sub001036_groupi_n_796, csa_tree_sub001036_groupi_n_797, csa_tree_sub001036_groupi_n_798, csa_tree_sub001036_groupi_n_799, csa_tree_sub001036_groupi_n_800, csa_tree_sub001036_groupi_n_801, csa_tree_sub001036_groupi_n_802;
  wire csa_tree_sub001036_groupi_n_803, csa_tree_sub001036_groupi_n_804, csa_tree_sub001036_groupi_n_805, csa_tree_sub001036_groupi_n_806, csa_tree_sub001036_groupi_n_807, csa_tree_sub001036_groupi_n_808, csa_tree_sub001036_groupi_n_809, csa_tree_sub001036_groupi_n_810;
  wire csa_tree_sub001036_groupi_n_811, csa_tree_sub001036_groupi_n_812, csa_tree_sub001036_groupi_n_813, csa_tree_sub001036_groupi_n_814, csa_tree_sub001036_groupi_n_815, csa_tree_sub001036_groupi_n_816, csa_tree_sub001036_groupi_n_817, csa_tree_sub001036_groupi_n_818;
  wire csa_tree_sub001036_groupi_n_819, csa_tree_sub001036_groupi_n_820, csa_tree_sub001036_groupi_n_821, csa_tree_sub001036_groupi_n_822, csa_tree_sub001036_groupi_n_823, csa_tree_sub001036_groupi_n_824, csa_tree_sub001036_groupi_n_825, csa_tree_sub001036_groupi_n_826;
  wire csa_tree_sub001036_groupi_n_827, csa_tree_sub001036_groupi_n_828, csa_tree_sub001036_groupi_n_829, csa_tree_sub001036_groupi_n_830, csa_tree_sub001036_groupi_n_831, csa_tree_sub001036_groupi_n_832, csa_tree_sub001036_groupi_n_833, csa_tree_sub001036_groupi_n_834;
  wire csa_tree_sub001036_groupi_n_835, csa_tree_sub001036_groupi_n_836, csa_tree_sub001036_groupi_n_837, csa_tree_sub001036_groupi_n_838, csa_tree_sub001036_groupi_n_839, csa_tree_sub001036_groupi_n_840, csa_tree_sub001036_groupi_n_841, csa_tree_sub001036_groupi_n_842;
  wire csa_tree_sub001036_groupi_n_843, csa_tree_sub001036_groupi_n_844, csa_tree_sub001036_groupi_n_845, csa_tree_sub001036_groupi_n_846, csa_tree_sub001036_groupi_n_847, csa_tree_sub001036_groupi_n_848, csa_tree_sub001036_groupi_n_849, csa_tree_sub001036_groupi_n_850;
  wire csa_tree_sub001036_groupi_n_851, csa_tree_sub001036_groupi_n_852, csa_tree_sub001036_groupi_n_853, csa_tree_sub001036_groupi_n_854, csa_tree_sub001036_groupi_n_855, csa_tree_sub001036_groupi_n_856, csa_tree_sub001036_groupi_n_857, csa_tree_sub001036_groupi_n_858;
  wire csa_tree_sub001036_groupi_n_859, csa_tree_sub001036_groupi_n_860, csa_tree_sub001036_groupi_n_861, csa_tree_sub001036_groupi_n_862, csa_tree_sub001036_groupi_n_863, csa_tree_sub001036_groupi_n_864, csa_tree_sub001036_groupi_n_865, csa_tree_sub001036_groupi_n_866;
  wire csa_tree_sub001036_groupi_n_867, csa_tree_sub001036_groupi_n_868, csa_tree_sub001036_groupi_n_869, csa_tree_sub001036_groupi_n_870, csa_tree_sub001036_groupi_n_871, csa_tree_sub001036_groupi_n_872, csa_tree_sub001036_groupi_n_873, csa_tree_sub001036_groupi_n_874;
  wire csa_tree_sub001036_groupi_n_875, csa_tree_sub001036_groupi_n_876, csa_tree_sub001036_groupi_n_877, csa_tree_sub001036_groupi_n_878, csa_tree_sub001036_groupi_n_879, csa_tree_sub001036_groupi_n_880, csa_tree_sub001036_groupi_n_881, csa_tree_sub001036_groupi_n_882;
  wire csa_tree_sub001036_groupi_n_883, csa_tree_sub001036_groupi_n_884, csa_tree_sub001036_groupi_n_885, csa_tree_sub001036_groupi_n_886, csa_tree_sub001036_groupi_n_887, csa_tree_sub001036_groupi_n_888, csa_tree_sub001036_groupi_n_889, csa_tree_sub001036_groupi_n_890;
  wire csa_tree_sub001036_groupi_n_891, csa_tree_sub001036_groupi_n_892, csa_tree_sub001036_groupi_n_893, csa_tree_sub001036_groupi_n_894, csa_tree_sub001036_groupi_n_895, csa_tree_sub001036_groupi_n_896, csa_tree_sub001036_groupi_n_897, csa_tree_sub001036_groupi_n_898;
  wire csa_tree_sub001036_groupi_n_899, csa_tree_sub001036_groupi_n_900, csa_tree_sub001036_groupi_n_901, csa_tree_sub001036_groupi_n_902, csa_tree_sub001036_groupi_n_903, csa_tree_sub001036_groupi_n_904, csa_tree_sub001036_groupi_n_905, csa_tree_sub001036_groupi_n_906;
  wire csa_tree_sub001036_groupi_n_907, csa_tree_sub001036_groupi_n_908, csa_tree_sub001036_groupi_n_909, csa_tree_sub001036_groupi_n_910, csa_tree_sub001036_groupi_n_911, csa_tree_sub001036_groupi_n_912, csa_tree_sub001036_groupi_n_913, csa_tree_sub001036_groupi_n_914;
  wire csa_tree_sub001036_groupi_n_915, csa_tree_sub001036_groupi_n_916, csa_tree_sub001036_groupi_n_917, csa_tree_sub001036_groupi_n_918, csa_tree_sub001036_groupi_n_919, csa_tree_sub001036_groupi_n_920, csa_tree_sub001036_groupi_n_921, csa_tree_sub001036_groupi_n_922;
  wire csa_tree_sub001036_groupi_n_923, csa_tree_sub001036_groupi_n_924, csa_tree_sub001036_groupi_n_925, csa_tree_sub001036_groupi_n_926, csa_tree_sub001036_groupi_n_927, csa_tree_sub001036_groupi_n_928, csa_tree_sub001036_groupi_n_929, csa_tree_sub001036_groupi_n_930;
  wire csa_tree_sub001036_groupi_n_931, csa_tree_sub001036_groupi_n_932, csa_tree_sub001036_groupi_n_933, csa_tree_sub001036_groupi_n_934, csa_tree_sub001036_groupi_n_935, csa_tree_sub001036_groupi_n_936, csa_tree_sub001036_groupi_n_937, csa_tree_sub001036_groupi_n_938;
  wire csa_tree_sub001036_groupi_n_939, csa_tree_sub001036_groupi_n_940, csa_tree_sub001036_groupi_n_941, csa_tree_sub001036_groupi_n_942, csa_tree_sub001036_groupi_n_943, csa_tree_sub001036_groupi_n_944, csa_tree_sub001036_groupi_n_945, csa_tree_sub001036_groupi_n_946;
  wire csa_tree_sub001036_groupi_n_947, csa_tree_sub001036_groupi_n_948, csa_tree_sub001036_groupi_n_949, csa_tree_sub001036_groupi_n_950, csa_tree_sub001036_groupi_n_951, csa_tree_sub001036_groupi_n_952, csa_tree_sub001036_groupi_n_953, csa_tree_sub001036_groupi_n_954;
  wire csa_tree_sub001036_groupi_n_955, csa_tree_sub001036_groupi_n_956, csa_tree_sub001036_groupi_n_957, csa_tree_sub001036_groupi_n_958, csa_tree_sub001036_groupi_n_959, csa_tree_sub001036_groupi_n_960, csa_tree_sub001036_groupi_n_961, csa_tree_sub001036_groupi_n_962;
  wire csa_tree_sub001036_groupi_n_963, csa_tree_sub001036_groupi_n_964, csa_tree_sub001036_groupi_n_965, csa_tree_sub001036_groupi_n_966, csa_tree_sub001036_groupi_n_967, csa_tree_sub001036_groupi_n_968, csa_tree_sub001036_groupi_n_969, csa_tree_sub001036_groupi_n_970;
  wire csa_tree_sub001036_groupi_n_971, csa_tree_sub001036_groupi_n_972, csa_tree_sub001036_groupi_n_973, csa_tree_sub001036_groupi_n_974, csa_tree_sub001036_groupi_n_975, csa_tree_sub001036_groupi_n_976, csa_tree_sub001036_groupi_n_977, csa_tree_sub001036_groupi_n_978;
  wire csa_tree_sub001036_groupi_n_979, csa_tree_sub001036_groupi_n_980, csa_tree_sub001036_groupi_n_981, csa_tree_sub001036_groupi_n_982, csa_tree_sub001036_groupi_n_983, csa_tree_sub001036_groupi_n_984, csa_tree_sub001036_groupi_n_985, csa_tree_sub001036_groupi_n_986;
  wire csa_tree_sub001036_groupi_n_987, csa_tree_sub001036_groupi_n_988, csa_tree_sub001036_groupi_n_989, csa_tree_sub001036_groupi_n_990, csa_tree_sub001036_groupi_n_991, csa_tree_sub001036_groupi_n_992, csa_tree_sub001036_groupi_n_993, csa_tree_sub001036_groupi_n_994;
  wire csa_tree_sub001036_groupi_n_995, csa_tree_sub001036_groupi_n_996, csa_tree_sub001036_groupi_n_997, csa_tree_sub001036_groupi_n_998, csa_tree_sub001036_groupi_n_999, csa_tree_sub001036_groupi_n_1000, csa_tree_sub001036_groupi_n_1001, csa_tree_sub001036_groupi_n_1002;
  wire csa_tree_sub001036_groupi_n_1003, csa_tree_sub001036_groupi_n_1004, csa_tree_sub001036_groupi_n_1005, csa_tree_sub001036_groupi_n_1006, csa_tree_sub001036_groupi_n_1007, csa_tree_sub001036_groupi_n_1008, csa_tree_sub001036_groupi_n_1009, csa_tree_sub001036_groupi_n_1010;
  wire csa_tree_sub001036_groupi_n_1011, csa_tree_sub001036_groupi_n_1012, csa_tree_sub001036_groupi_n_1013, csa_tree_sub001036_groupi_n_1014, csa_tree_sub001036_groupi_n_1015, csa_tree_sub001036_groupi_n_1016, csa_tree_sub001036_groupi_n_1017, csa_tree_sub001036_groupi_n_1018;
  wire csa_tree_sub001036_groupi_n_1019, csa_tree_sub001036_groupi_n_1020, csa_tree_sub001036_groupi_n_1021, csa_tree_sub001036_groupi_n_1022, csa_tree_sub001036_groupi_n_1023, csa_tree_sub001036_groupi_n_1024, csa_tree_sub001036_groupi_n_1025, csa_tree_sub001036_groupi_n_1026;
  wire csa_tree_sub001036_groupi_n_1027, csa_tree_sub001036_groupi_n_1028, csa_tree_sub001036_groupi_n_1029, csa_tree_sub001036_groupi_n_1030, csa_tree_sub001036_groupi_n_1031, csa_tree_sub001036_groupi_n_1032, csa_tree_sub001036_groupi_n_1033, csa_tree_sub001036_groupi_n_1034;
  wire csa_tree_sub001036_groupi_n_1035, csa_tree_sub001036_groupi_n_1036, csa_tree_sub001036_groupi_n_1037, csa_tree_sub001036_groupi_n_1038, csa_tree_sub001036_groupi_n_1039, csa_tree_sub001036_groupi_n_1040, csa_tree_sub001036_groupi_n_1041, csa_tree_sub001036_groupi_n_1042;
  wire csa_tree_sub001036_groupi_n_1043, csa_tree_sub001036_groupi_n_1044, csa_tree_sub001036_groupi_n_1045, csa_tree_sub001036_groupi_n_1046, csa_tree_sub001036_groupi_n_1047, csa_tree_sub001036_groupi_n_1048, csa_tree_sub001036_groupi_n_1049, csa_tree_sub001036_groupi_n_1050;
  wire csa_tree_sub001036_groupi_n_1051, csa_tree_sub001036_groupi_n_1052, csa_tree_sub001036_groupi_n_1053, csa_tree_sub001036_groupi_n_1054, csa_tree_sub001036_groupi_n_1055, csa_tree_sub001036_groupi_n_1056, csa_tree_sub001036_groupi_n_1057, csa_tree_sub001036_groupi_n_1058;
  wire csa_tree_sub001036_groupi_n_1059, csa_tree_sub001036_groupi_n_1060, csa_tree_sub001036_groupi_n_1061, csa_tree_sub001036_groupi_n_1062, csa_tree_sub001036_groupi_n_1063, csa_tree_sub001036_groupi_n_1064, csa_tree_sub001036_groupi_n_1065, csa_tree_sub001036_groupi_n_1066;
  wire csa_tree_sub001036_groupi_n_1067, csa_tree_sub001036_groupi_n_1068, csa_tree_sub001036_groupi_n_1069, csa_tree_sub001036_groupi_n_1070, csa_tree_sub001036_groupi_n_1071, csa_tree_sub001036_groupi_n_1072, csa_tree_sub001036_groupi_n_1073, csa_tree_sub001036_groupi_n_1074;
  wire csa_tree_sub001036_groupi_n_1075, csa_tree_sub001036_groupi_n_1076, csa_tree_sub001036_groupi_n_1077, csa_tree_sub001036_groupi_n_1078, csa_tree_sub001036_groupi_n_1079, csa_tree_sub001036_groupi_n_1080, csa_tree_sub001036_groupi_n_1081, csa_tree_sub001036_groupi_n_1082;
  wire csa_tree_sub001036_groupi_n_1083, csa_tree_sub001036_groupi_n_1084, csa_tree_sub001036_groupi_n_1085, csa_tree_sub001036_groupi_n_1086, csa_tree_sub001036_groupi_n_1087, csa_tree_sub001036_groupi_n_1088, csa_tree_sub001036_groupi_n_1089, csa_tree_sub001036_groupi_n_1090;
  wire csa_tree_sub001036_groupi_n_1091, csa_tree_sub001036_groupi_n_1092, csa_tree_sub001036_groupi_n_1093, csa_tree_sub001036_groupi_n_1094, csa_tree_sub001036_groupi_n_1095, csa_tree_sub001036_groupi_n_1096, csa_tree_sub001036_groupi_n_1097, csa_tree_sub001036_groupi_n_1098;
  wire csa_tree_sub001036_groupi_n_1099, csa_tree_sub001036_groupi_n_1100, csa_tree_sub001036_groupi_n_1101, csa_tree_sub001036_groupi_n_1102, csa_tree_sub001036_groupi_n_1103, csa_tree_sub001036_groupi_n_1104, csa_tree_sub001036_groupi_n_1105, csa_tree_sub001036_groupi_n_1106;
  wire csa_tree_sub001036_groupi_n_1107, csa_tree_sub001036_groupi_n_1108, csa_tree_sub001036_groupi_n_1109, csa_tree_sub001036_groupi_n_1110, csa_tree_sub001036_groupi_n_1111, csa_tree_sub001036_groupi_n_1112, csa_tree_sub001036_groupi_n_1113, csa_tree_sub001036_groupi_n_1114;
  wire csa_tree_sub001036_groupi_n_1115, csa_tree_sub001036_groupi_n_1116, csa_tree_sub001036_groupi_n_1117, csa_tree_sub001036_groupi_n_1118, csa_tree_sub001036_groupi_n_1119, csa_tree_sub001036_groupi_n_1120, csa_tree_sub001036_groupi_n_1121, csa_tree_sub001036_groupi_n_1122;
  wire csa_tree_sub001036_groupi_n_1123, csa_tree_sub001036_groupi_n_1124, csa_tree_sub001036_groupi_n_1125, csa_tree_sub001036_groupi_n_1126, csa_tree_sub001036_groupi_n_1127, csa_tree_sub001036_groupi_n_1128, csa_tree_sub001036_groupi_n_1129, csa_tree_sub001036_groupi_n_1130;
  wire csa_tree_sub001036_groupi_n_1131, csa_tree_sub001036_groupi_n_1132, csa_tree_sub001036_groupi_n_1133, csa_tree_sub001036_groupi_n_1134, csa_tree_sub001036_groupi_n_1135, csa_tree_sub001036_groupi_n_1136, csa_tree_sub001036_groupi_n_1137, csa_tree_sub001036_groupi_n_1138;
  wire csa_tree_sub001036_groupi_n_1139, csa_tree_sub001036_groupi_n_1140, csa_tree_sub001036_groupi_n_1141, csa_tree_sub001036_groupi_n_1142, csa_tree_sub001036_groupi_n_1144, csa_tree_sub001036_groupi_n_1145, csa_tree_sub001036_groupi_n_1146, csa_tree_sub001036_groupi_n_1147;
  wire csa_tree_sub001036_groupi_n_1148, csa_tree_sub001036_groupi_n_1149, csa_tree_sub001036_groupi_n_1150, csa_tree_sub001036_groupi_n_1151, csa_tree_sub001036_groupi_n_1152, csa_tree_sub001036_groupi_n_1153, csa_tree_sub001036_groupi_n_1154, csa_tree_sub001036_groupi_n_1155;
  wire csa_tree_sub001036_groupi_n_1156, csa_tree_sub001036_groupi_n_1157, csa_tree_sub001036_groupi_n_1158, csa_tree_sub001036_groupi_n_1159, csa_tree_sub001036_groupi_n_1160, csa_tree_sub001036_groupi_n_1161, csa_tree_sub001036_groupi_n_1162, csa_tree_sub001036_groupi_n_1163;
  wire csa_tree_sub001036_groupi_n_1164, csa_tree_sub001036_groupi_n_1165, csa_tree_sub001036_groupi_n_1166, csa_tree_sub001036_groupi_n_1167, csa_tree_sub001036_groupi_n_1168, csa_tree_sub001036_groupi_n_1169, csa_tree_sub001036_groupi_n_1170, csa_tree_sub001036_groupi_n_1171;
  wire csa_tree_sub001036_groupi_n_1172, csa_tree_sub001036_groupi_n_1173, csa_tree_sub001036_groupi_n_1174, csa_tree_sub001036_groupi_n_1175, csa_tree_sub001036_groupi_n_1176, csa_tree_sub001036_groupi_n_1177, csa_tree_sub001036_groupi_n_1178, csa_tree_sub001036_groupi_n_1179;
  wire csa_tree_sub001036_groupi_n_1180, csa_tree_sub001036_groupi_n_1181, csa_tree_sub001036_groupi_n_1182, csa_tree_sub001036_groupi_n_1183, csa_tree_sub001036_groupi_n_1184, csa_tree_sub001036_groupi_n_1185, csa_tree_sub001036_groupi_n_1186, csa_tree_sub001036_groupi_n_1187;
  wire csa_tree_sub001036_groupi_n_1188, csa_tree_sub001036_groupi_n_1189, csa_tree_sub001036_groupi_n_1190, csa_tree_sub001036_groupi_n_1191, csa_tree_sub001036_groupi_n_1192, csa_tree_sub001036_groupi_n_1193, csa_tree_sub001036_groupi_n_1194, csa_tree_sub001036_groupi_n_1195;
  wire csa_tree_sub001036_groupi_n_1196, csa_tree_sub001036_groupi_n_1197, csa_tree_sub001036_groupi_n_1198, csa_tree_sub001036_groupi_n_1199, csa_tree_sub001036_groupi_n_1200, csa_tree_sub001036_groupi_n_1201, csa_tree_sub001036_groupi_n_1202, csa_tree_sub001036_groupi_n_1203;
  wire csa_tree_sub001036_groupi_n_1204, csa_tree_sub001036_groupi_n_1205, csa_tree_sub001036_groupi_n_1206, csa_tree_sub001036_groupi_n_1207, csa_tree_sub001036_groupi_n_1208, csa_tree_sub001036_groupi_n_1209, csa_tree_sub001036_groupi_n_1210, csa_tree_sub001036_groupi_n_1211;
  wire csa_tree_sub001036_groupi_n_1212, csa_tree_sub001036_groupi_n_1213, csa_tree_sub001036_groupi_n_1214, csa_tree_sub001036_groupi_n_1215, csa_tree_sub001036_groupi_n_1216, csa_tree_sub001036_groupi_n_1217, csa_tree_sub001036_groupi_n_1218, csa_tree_sub001036_groupi_n_1219;
  wire csa_tree_sub001036_groupi_n_1220, csa_tree_sub001036_groupi_n_1221, csa_tree_sub001036_groupi_n_1222, csa_tree_sub001036_groupi_n_1223, csa_tree_sub001036_groupi_n_1224, csa_tree_sub001036_groupi_n_1225, csa_tree_sub001036_groupi_n_1226, csa_tree_sub001036_groupi_n_1227;
  wire csa_tree_sub001036_groupi_n_1228, csa_tree_sub001036_groupi_n_1229, csa_tree_sub001036_groupi_n_1230, csa_tree_sub001036_groupi_n_1231, csa_tree_sub001036_groupi_n_1232, csa_tree_sub001036_groupi_n_1233, csa_tree_sub001036_groupi_n_1234, csa_tree_sub001036_groupi_n_1235;
  wire csa_tree_sub001036_groupi_n_1236, csa_tree_sub001036_groupi_n_1237, csa_tree_sub001036_groupi_n_1238, csa_tree_sub001036_groupi_n_1239, csa_tree_sub001036_groupi_n_1240, csa_tree_sub001036_groupi_n_1241, csa_tree_sub001036_groupi_n_1242, csa_tree_sub001036_groupi_n_1243;
  wire csa_tree_sub001036_groupi_n_1244, csa_tree_sub001036_groupi_n_1245, csa_tree_sub001036_groupi_n_1246, csa_tree_sub001036_groupi_n_1247, csa_tree_sub001036_groupi_n_1248, csa_tree_sub001036_groupi_n_1249, csa_tree_sub001036_groupi_n_1250, csa_tree_sub001036_groupi_n_1251;
  wire csa_tree_sub001036_groupi_n_1252, csa_tree_sub001036_groupi_n_1253, csa_tree_sub001036_groupi_n_1254, csa_tree_sub001036_groupi_n_1255, csa_tree_sub001036_groupi_n_1256, csa_tree_sub001036_groupi_n_1257, csa_tree_sub001036_groupi_n_1258, csa_tree_sub001036_groupi_n_1259;
  wire csa_tree_sub001036_groupi_n_1260, csa_tree_sub001036_groupi_n_1261, csa_tree_sub001036_groupi_n_1262, csa_tree_sub001036_groupi_n_1263, csa_tree_sub001036_groupi_n_1264, csa_tree_sub001036_groupi_n_1265, csa_tree_sub001036_groupi_n_1266, csa_tree_sub001036_groupi_n_1267;
  wire csa_tree_sub001036_groupi_n_1268, csa_tree_sub001036_groupi_n_1269, csa_tree_sub001036_groupi_n_1270, csa_tree_sub001036_groupi_n_1271, csa_tree_sub001036_groupi_n_1272, csa_tree_sub001036_groupi_n_1273, csa_tree_sub001036_groupi_n_1274, csa_tree_sub001036_groupi_n_1275;
  wire csa_tree_sub001036_groupi_n_1276, csa_tree_sub001036_groupi_n_1277, csa_tree_sub001036_groupi_n_1278, csa_tree_sub001036_groupi_n_1279, csa_tree_sub001036_groupi_n_1280, csa_tree_sub001036_groupi_n_1281, csa_tree_sub001036_groupi_n_1282, csa_tree_sub001036_groupi_n_1283;
  wire csa_tree_sub001036_groupi_n_1284, csa_tree_sub001036_groupi_n_1285, csa_tree_sub001036_groupi_n_1286, csa_tree_sub001036_groupi_n_1287, csa_tree_sub001036_groupi_n_1288, csa_tree_sub001036_groupi_n_1289, csa_tree_sub001036_groupi_n_1290, csa_tree_sub001036_groupi_n_1291;
  wire csa_tree_sub001036_groupi_n_1292, csa_tree_sub001036_groupi_n_1293, csa_tree_sub001036_groupi_n_1294, csa_tree_sub001036_groupi_n_1295, csa_tree_sub001036_groupi_n_1296, csa_tree_sub001036_groupi_n_1297, csa_tree_sub001036_groupi_n_1298, csa_tree_sub001036_groupi_n_1299;
  wire csa_tree_sub001036_groupi_n_1300, csa_tree_sub001036_groupi_n_1301, csa_tree_sub001036_groupi_n_1302, csa_tree_sub001036_groupi_n_1303, csa_tree_sub001036_groupi_n_1304, csa_tree_sub001036_groupi_n_1305, csa_tree_sub001036_groupi_n_1306, csa_tree_sub001036_groupi_n_1307;
  wire csa_tree_sub001036_groupi_n_1308, csa_tree_sub001036_groupi_n_1309, csa_tree_sub001036_groupi_n_1310, csa_tree_sub001036_groupi_n_1311, csa_tree_sub001036_groupi_n_1312, csa_tree_sub001036_groupi_n_1313, csa_tree_sub001036_groupi_n_1314, csa_tree_sub001036_groupi_n_1315;
  wire csa_tree_sub001036_groupi_n_1316, csa_tree_sub001036_groupi_n_1317, csa_tree_sub001036_groupi_n_1318, csa_tree_sub001036_groupi_n_1319, csa_tree_sub001036_groupi_n_1320, csa_tree_sub001036_groupi_n_1321, csa_tree_sub001036_groupi_n_1322, csa_tree_sub001036_groupi_n_1323;
  wire csa_tree_sub001036_groupi_n_1324, csa_tree_sub001036_groupi_n_1325, csa_tree_sub001036_groupi_n_1326, csa_tree_sub001036_groupi_n_1327, csa_tree_sub001036_groupi_n_1328, csa_tree_sub001036_groupi_n_1329, csa_tree_sub001036_groupi_n_1330, csa_tree_sub001036_groupi_n_1331;
  wire csa_tree_sub001036_groupi_n_1332, csa_tree_sub001036_groupi_n_1333, csa_tree_sub001036_groupi_n_1334, csa_tree_sub001036_groupi_n_1335, csa_tree_sub001036_groupi_n_1336, csa_tree_sub001036_groupi_n_1337, csa_tree_sub001036_groupi_n_1338, csa_tree_sub001036_groupi_n_1339;
  wire csa_tree_sub001036_groupi_n_1340, csa_tree_sub001036_groupi_n_1341, csa_tree_sub001036_groupi_n_1342, csa_tree_sub001036_groupi_n_1344, csa_tree_sub001036_groupi_n_1345, csa_tree_sub001036_groupi_n_1346, csa_tree_sub001036_groupi_n_1347, csa_tree_sub001036_groupi_n_1348;
  wire csa_tree_sub001036_groupi_n_1349, csa_tree_sub001036_groupi_n_1350, csa_tree_sub001036_groupi_n_1351, csa_tree_sub001036_groupi_n_1352, csa_tree_sub001036_groupi_n_1353, csa_tree_sub001036_groupi_n_1354, csa_tree_sub001036_groupi_n_1355, csa_tree_sub001036_groupi_n_1356;
  wire csa_tree_sub001036_groupi_n_1357, csa_tree_sub001036_groupi_n_1358, csa_tree_sub001036_groupi_n_1359, csa_tree_sub001036_groupi_n_1360, csa_tree_sub001036_groupi_n_1361, csa_tree_sub001036_groupi_n_1362, csa_tree_sub001036_groupi_n_1363, csa_tree_sub001036_groupi_n_1364;
  wire csa_tree_sub001036_groupi_n_1365, csa_tree_sub001036_groupi_n_1366, csa_tree_sub001036_groupi_n_1367, csa_tree_sub001036_groupi_n_1368, csa_tree_sub001036_groupi_n_1369, csa_tree_sub001036_groupi_n_1370, csa_tree_sub001036_groupi_n_1371, csa_tree_sub001036_groupi_n_1372;
  wire csa_tree_sub001036_groupi_n_1373, csa_tree_sub001036_groupi_n_1374, csa_tree_sub001036_groupi_n_1375, csa_tree_sub001036_groupi_n_1376, csa_tree_sub001036_groupi_n_1377, csa_tree_sub001036_groupi_n_1378, csa_tree_sub001036_groupi_n_1379, csa_tree_sub001036_groupi_n_1380;
  wire csa_tree_sub001036_groupi_n_1381, csa_tree_sub001036_groupi_n_1382, csa_tree_sub001036_groupi_n_1383, csa_tree_sub001036_groupi_n_1384, csa_tree_sub001036_groupi_n_1385, csa_tree_sub001036_groupi_n_1386, csa_tree_sub001036_groupi_n_1387, csa_tree_sub001036_groupi_n_1388;
  wire csa_tree_sub001036_groupi_n_1389, csa_tree_sub001036_groupi_n_1390, csa_tree_sub001036_groupi_n_1391, csa_tree_sub001036_groupi_n_1392, csa_tree_sub001036_groupi_n_1393, csa_tree_sub001036_groupi_n_1394, csa_tree_sub001036_groupi_n_1395, csa_tree_sub001036_groupi_n_1396;
  wire csa_tree_sub001036_groupi_n_1397, csa_tree_sub001036_groupi_n_1398, csa_tree_sub001036_groupi_n_1399, csa_tree_sub001036_groupi_n_1400, csa_tree_sub001036_groupi_n_1401, csa_tree_sub001036_groupi_n_1403, csa_tree_sub001036_groupi_n_1404, csa_tree_sub001036_groupi_n_1405;
  wire csa_tree_sub001036_groupi_n_1406, csa_tree_sub001036_groupi_n_1407, csa_tree_sub001036_groupi_n_1408, csa_tree_sub001036_groupi_n_1409, csa_tree_sub001036_groupi_n_1410, csa_tree_sub001036_groupi_n_1411, csa_tree_sub001036_groupi_n_1412, csa_tree_sub001036_groupi_n_1413;
  wire csa_tree_sub001036_groupi_n_1414, csa_tree_sub001036_groupi_n_1415, csa_tree_sub001036_groupi_n_1416, csa_tree_sub001036_groupi_n_1417, csa_tree_sub001036_groupi_n_1418, csa_tree_sub001036_groupi_n_1419, csa_tree_sub001036_groupi_n_1420, csa_tree_sub001036_groupi_n_1421;
  wire csa_tree_sub001036_groupi_n_1422, csa_tree_sub001036_groupi_n_1423, csa_tree_sub001036_groupi_n_1424, csa_tree_sub001036_groupi_n_1425, csa_tree_sub001036_groupi_n_1426, csa_tree_sub001036_groupi_n_1427, csa_tree_sub001036_groupi_n_1428, csa_tree_sub001036_groupi_n_1429;
  wire csa_tree_sub001036_groupi_n_1430, csa_tree_sub001036_groupi_n_1431, csa_tree_sub001036_groupi_n_1432, csa_tree_sub001036_groupi_n_1434, csa_tree_sub001036_groupi_n_1435, csa_tree_sub001036_groupi_n_1436, csa_tree_sub001036_groupi_n_1437, csa_tree_sub001036_groupi_n_1438;
  wire csa_tree_sub001036_groupi_n_1439, csa_tree_sub001036_groupi_n_1440, csa_tree_sub001036_groupi_n_1441, csa_tree_sub001036_groupi_n_1442, csa_tree_sub001036_groupi_n_1443, csa_tree_sub001036_groupi_n_1444, csa_tree_sub001036_groupi_n_1445, csa_tree_sub001036_groupi_n_1446;
  wire csa_tree_sub001036_groupi_n_1448, csa_tree_sub001036_groupi_n_1449, csa_tree_sub001036_groupi_n_1450, csa_tree_sub001036_groupi_n_1451, csa_tree_sub001036_groupi_n_1452, csa_tree_sub001036_groupi_n_1453, csa_tree_sub001036_groupi_n_1454, csa_tree_sub001036_groupi_n_1455;
  wire csa_tree_sub001036_groupi_n_1456, csa_tree_sub001036_groupi_n_1457, csa_tree_sub001036_groupi_n_1458, csa_tree_sub001036_groupi_n_1459, csa_tree_sub001036_groupi_n_1461, csa_tree_sub001036_groupi_n_1462, csa_tree_sub001036_groupi_n_1463, csa_tree_sub001036_groupi_n_1464;
  wire csa_tree_sub001036_groupi_n_1466, csa_tree_sub001036_groupi_n_1467, csa_tree_sub001036_groupi_n_1468, csa_tree_sub001036_groupi_n_1470, csa_tree_sub001036_groupi_n_1471, csa_tree_sub001036_groupi_n_1472, csa_tree_sub001036_groupi_n_1473, csa_tree_sub001036_groupi_n_1474;
  wire csa_tree_sub001036_groupi_n_1475, csa_tree_sub001036_groupi_n_1477, n_0, n_1, n_2, n_3, n_4, n_5;
  wire n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13;
  wire n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21;
  wire n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93;
  wire n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  or g514__2398(n_118 ,n_66 ,n_94);
  or g515__5107(n_138 ,n_77 ,n_101);
  or g516__6260(n_135 ,n_81 ,n_108);
  or g517__4319(n_114 ,n_80 ,n_107);
  or g518__8428(n_129 ,n_82 ,n_109);
  or g519__5526(n_128 ,n_79 ,n_106);
  or g520__6783(n_120 ,n_75 ,n_103);
  or g521__3680(n_127 ,n_76 ,n_105);
  or g522__1617(n_126 ,n_74 ,n_104);
  or g523__2802(n_137 ,n_68 ,n_96);
  or g524__1705(n_119 ,n_71 ,n_100);
  or g525__5122(n_125 ,n_72 ,n_102);
  or g526__8246(n_124 ,n_70 ,n_99);
  or g527__7098(n_141 ,n_73 ,n_111);
  or g528__6131(n_130 ,n_57 ,n_85);
  or g529__1881(n_140 ,n_83 ,n_98);
  or g530__5115(n_139 ,n_78 ,n_90);
  or g531__7482(n_122 ,n_65 ,n_95);
  or g532__4733(n_121 ,n_63 ,n_93);
  or g533__6161(n_136 ,n_60 ,n_112);
  or g534__9315(n_117 ,n_62 ,n_92);
  or g535__9945(n_134 ,n_61 ,n_91);
  or g536__2883(n_116 ,n_58 ,n_87);
  or g537__2346(n_133 ,n_59 ,n_89);
  or g538__1666(n_132 ,n_84 ,n_88);
  or g539__7410(n_115 ,n_67 ,n_110);
  or g540__6417(n_131 ,n_64 ,n_86);
  or g541__5477(n_123 ,n_69 ,n_97);
  and g542__2398(n_112 ,in6[1] ,n_39);
  and g543__5107(n_111 ,in6[6] ,n_28);
  and g544__6260(n_110 ,in21[1] ,n_43);
  and g545__4319(n_109 ,in5[1] ,n_39);
  and g546__8428(n_108 ,in6[0] ,n_24);
  and g547__5526(n_107 ,in21[0] ,n_45);
  and g548__6783(n_106 ,in5[0] ,n_46);
  and g549__3680(n_105 ,in22[6] ,n_46);
  and g550__1617(n_104 ,in22[5] ,n_45);
  and g551__2802(n_103 ,in21[6] ,n_33);
  and g552__1705(n_102 ,in22[4] ,n_31);
  and g553__5122(n_101 ,in6[3] ,n_34);
  and g554__8246(n_100 ,in21[5] ,n_28);
  and g555__7098(n_99 ,in22[3] ,n_31);
  and g556__6131(n_98 ,in6[5] ,n_43);
  and g557__1881(n_97 ,in22[2] ,n_40);
  and g558__5115(n_96 ,in6[2] ,n_42);
  and g559__7482(n_95 ,in22[1] ,n_30);
  and g560__4733(n_94 ,in21[4] ,n_27);
  and g561__6161(n_93 ,in22[0] ,n_27);
  and g562__9315(n_92 ,in21[3] ,n_34);
  and g563__9945(n_91 ,in5[6] ,n_33);
  and g564__2883(n_90 ,in6[4] ,n_25);
  and g565__2346(n_89 ,in5[5] ,n_42);
  and g566__1666(n_88 ,in5[4] ,n_40);
  and g567__7410(n_87 ,in21[2] ,n_30);
  and g568__6417(n_86 ,in5[3] ,n_25);
  and g569__5477(n_85 ,in5[2] ,n_24);
  and g570__2398(n_84 ,in1[4] ,n_18);
  and g571__5107(n_83 ,in2[5] ,n_7);
  and g572__6260(n_82 ,in1[1] ,n_21);
  and g573__4319(n_81 ,in2[0] ,n_19);
  and g574__8428(n_80 ,n_4 ,in19[0]);
  and g575__5526(n_79 ,in1[0] ,n_1);
  and g576__6783(n_78 ,in2[4] ,n_11);
  and g577__3680(n_77 ,in2[3] ,n_11);
  and g578__1617(n_76 ,n_4 ,in20[6]);
  and g579__2802(n_75 ,n_21 ,in19[6]);
  and g580__1705(n_74 ,n_5 ,in20[5]);
  and g581__5122(n_73 ,in2[6] ,n_2);
  and g582__8246(n_72 ,n_8 ,in20[4]);
  and g583__7098(n_71 ,n_1 ,in19[5]);
  and g584__6131(n_70 ,n_2 ,in20[3]);
  and g585__1881(n_69 ,n_22 ,in20[2]);
  and g586__5115(n_68 ,in2[2] ,n_10);
  and g587__7482(n_67 ,n_5 ,in19[1]);
  and g588__4733(n_66 ,n_10 ,in19[4]);
  and g589__6161(n_65 ,n_7 ,in20[1]);
  and g590__9315(n_64 ,in1[3] ,n_13);
  and g591__9945(n_63 ,n_8 ,in20[0]);
  and g592__2883(n_62 ,n_22 ,in19[3]);
  and g593__2346(n_61 ,in1[6] ,n_18);
  and g594__1666(n_60 ,in2[1] ,n_14);
  and g595__7410(n_59 ,in1[5] ,n_19);
  and g596__6417(n_58 ,n_47 ,in19[2]);
  and g597__5477(n_57 ,in1[2] ,n_14);
  not g598(n_56 ,n_16);
  not g600(n_55 ,n_54);
  not g601(n_53 ,n_51);
  not g602(n_52 ,n_51);
  not g603(n_51 ,n_16);
  not g607(n_50 ,n_54);
  not g608(n_54 ,in3);
  not drc_bufs630(n_47 ,n_49);
  not drc_bufs632(n_49 ,n_55);
  not drc_bufs638(n_46 ,n_44);
  not drc_bufs639(n_45 ,n_44);
  not drc_bufs640(n_44 ,n_49);
  not drc_bufs642(n_43 ,n_41);
  not drc_bufs643(n_42 ,n_41);
  not drc_bufs644(n_41 ,n_48);
  not drc_bufs646(n_40 ,n_38);
  not drc_bufs647(n_39 ,n_38);
  not drc_bufs648(n_38 ,n_48);
  not drc_bufs650(n_37 ,n_36);
  not drc_bufs652(n_36 ,n_56);
  not drc_bufs655(n_35 ,n_36);
  not drc_bufs660(n_34 ,n_32);
  not drc_bufs661(n_33 ,n_32);
  not drc_bufs662(n_32 ,n_52);
  not drc_bufs664(n_31 ,n_29);
  not drc_bufs665(n_30 ,n_29);
  not drc_bufs666(n_29 ,n_53);
  not drc_bufs668(n_28 ,n_26);
  not drc_bufs669(n_27 ,n_26);
  not drc_bufs670(n_26 ,n_52);
  not drc_bufs672(n_25 ,n_23);
  not drc_bufs673(n_24 ,n_23);
  not drc_bufs674(n_23 ,n_53);
  not drc_bufs676(n_22 ,n_20);
  not drc_bufs677(n_21 ,n_20);
  not drc_bufs678(n_20 ,n_50);
  not drc_bufs680(n_19 ,n_17);
  not drc_bufs681(n_18 ,n_17);
  not drc_bufs682(n_17 ,n_50);
  not drc_bufs684(n_16 ,n_15);
  not drc_bufs685(n_48 ,n_15);
  not drc_bufs686(n_15 ,n_54);
  not drc_bufs688(n_14 ,n_12);
  not drc_bufs689(n_13 ,n_12);
  not drc_bufs690(n_12 ,n_55);
  not drc_bufs692(n_11 ,n_9);
  not drc_bufs693(n_10 ,n_9);
  not drc_bufs694(n_9 ,n_37);
  not drc_bufs696(n_8 ,n_6);
  not drc_bufs697(n_7 ,n_6);
  not drc_bufs698(n_6 ,n_35);
  not drc_bufs700(n_5 ,n_3);
  not drc_bufs701(n_4 ,n_3);
  not drc_bufs702(n_3 ,n_35);
  not drc_bufs704(n_2 ,n_0);
  not drc_bufs705(n_1 ,n_0);
  not drc_bufs706(n_0 ,n_37);
  xnor csa_tree_sub001036_groupi_g4522__2398(out1[12] ,csa_tree_sub001036_groupi_n_1362 ,csa_tree_sub001036_groupi_n_1477);
  nor csa_tree_sub001036_groupi_g4523__5107(csa_tree_sub001036_groupi_n_1477 ,csa_tree_sub001036_groupi_n_1475 ,csa_tree_sub001036_groupi_n_1431);
  xnor csa_tree_sub001036_groupi_g4524__6260(out1[11] ,csa_tree_sub001036_groupi_n_1474 ,csa_tree_sub001036_groupi_n_1435);
  nor csa_tree_sub001036_groupi_g4525__4319(csa_tree_sub001036_groupi_n_1475 ,csa_tree_sub001036_groupi_n_1474 ,csa_tree_sub001036_groupi_n_1430);
  and csa_tree_sub001036_groupi_g4526__8428(csa_tree_sub001036_groupi_n_1474 ,csa_tree_sub001036_groupi_n_1473 ,csa_tree_sub001036_groupi_n_1448);
  or csa_tree_sub001036_groupi_g4528__5526(csa_tree_sub001036_groupi_n_1473 ,csa_tree_sub001036_groupi_n_1472 ,csa_tree_sub001036_groupi_n_1449);
  and csa_tree_sub001036_groupi_g4530__6783(csa_tree_sub001036_groupi_n_1472 ,csa_tree_sub001036_groupi_n_1471 ,csa_tree_sub001036_groupi_n_1457);
  or csa_tree_sub001036_groupi_g4532__3680(csa_tree_sub001036_groupi_n_1471 ,csa_tree_sub001036_groupi_n_1470 ,csa_tree_sub001036_groupi_n_1455);
  and csa_tree_sub001036_groupi_g4534__1617(csa_tree_sub001036_groupi_n_1470 ,csa_tree_sub001036_groupi_n_1468 ,csa_tree_sub001036_groupi_n_1456);
  xnor csa_tree_sub001036_groupi_g4535__2802(out1[8] ,csa_tree_sub001036_groupi_n_1466 ,csa_tree_sub001036_groupi_n_1462);
  or csa_tree_sub001036_groupi_g4536__1705(csa_tree_sub001036_groupi_n_1468 ,csa_tree_sub001036_groupi_n_1459 ,csa_tree_sub001036_groupi_n_1467);
  not csa_tree_sub001036_groupi_g4537(csa_tree_sub001036_groupi_n_1467 ,csa_tree_sub001036_groupi_n_1466);
  or csa_tree_sub001036_groupi_g4538__5122(csa_tree_sub001036_groupi_n_1466 ,csa_tree_sub001036_groupi_n_1452 ,csa_tree_sub001036_groupi_n_1464);
  xnor csa_tree_sub001036_groupi_g4539__8246(out1[7] ,csa_tree_sub001036_groupi_n_1463 ,csa_tree_sub001036_groupi_n_1454);
  and csa_tree_sub001036_groupi_g4540__7098(csa_tree_sub001036_groupi_n_1464 ,csa_tree_sub001036_groupi_n_1451 ,csa_tree_sub001036_groupi_n_1463);
  or csa_tree_sub001036_groupi_g4541__6131(csa_tree_sub001036_groupi_n_1463 ,csa_tree_sub001036_groupi_n_1427 ,csa_tree_sub001036_groupi_n_1458);
  xnor csa_tree_sub001036_groupi_g4542__1881(csa_tree_sub001036_groupi_n_1462 ,csa_tree_sub001036_groupi_n_1440 ,csa_tree_sub001036_groupi_n_1446);
  xnor csa_tree_sub001036_groupi_g4543__5115(csa_tree_sub001036_groupi_n_1461 ,csa_tree_sub001036_groupi_n_1437 ,csa_tree_sub001036_groupi_n_1444);
  xnor csa_tree_sub001036_groupi_g4544__7482(out1[6] ,csa_tree_sub001036_groupi_n_1450 ,csa_tree_sub001036_groupi_n_1434);
  nor csa_tree_sub001036_groupi_g4545__4733(csa_tree_sub001036_groupi_n_1459 ,csa_tree_sub001036_groupi_n_1440 ,csa_tree_sub001036_groupi_n_1446);
  nor csa_tree_sub001036_groupi_g4546__6161(csa_tree_sub001036_groupi_n_1458 ,csa_tree_sub001036_groupi_n_1450 ,csa_tree_sub001036_groupi_n_1423);
  or csa_tree_sub001036_groupi_g4547__9315(csa_tree_sub001036_groupi_n_1457 ,csa_tree_sub001036_groupi_n_1436 ,csa_tree_sub001036_groupi_n_1443);
  or csa_tree_sub001036_groupi_g4548__9945(csa_tree_sub001036_groupi_n_1456 ,csa_tree_sub001036_groupi_n_1439 ,csa_tree_sub001036_groupi_n_1445);
  nor csa_tree_sub001036_groupi_g4549__2883(csa_tree_sub001036_groupi_n_1455 ,csa_tree_sub001036_groupi_n_1437 ,csa_tree_sub001036_groupi_n_1444);
  xnor csa_tree_sub001036_groupi_g4550__2346(csa_tree_sub001036_groupi_n_1454 ,csa_tree_sub001036_groupi_n_1432 ,csa_tree_sub001036_groupi_n_1417);
  xnor csa_tree_sub001036_groupi_g4551__1666(csa_tree_sub001036_groupi_n_1453 ,csa_tree_sub001036_groupi_n_1408 ,csa_tree_sub001036_groupi_n_1442);
  and csa_tree_sub001036_groupi_g4552__7410(csa_tree_sub001036_groupi_n_1452 ,csa_tree_sub001036_groupi_n_1432 ,csa_tree_sub001036_groupi_n_1417);
  or csa_tree_sub001036_groupi_g4553__6417(csa_tree_sub001036_groupi_n_1451 ,csa_tree_sub001036_groupi_n_1432 ,csa_tree_sub001036_groupi_n_1417);
  and csa_tree_sub001036_groupi_g4554__5477(csa_tree_sub001036_groupi_n_1450 ,csa_tree_sub001036_groupi_n_1438 ,csa_tree_sub001036_groupi_n_1403);
  nor csa_tree_sub001036_groupi_g4555__2398(csa_tree_sub001036_groupi_n_1449 ,csa_tree_sub001036_groupi_n_1408 ,csa_tree_sub001036_groupi_n_1442);
  or csa_tree_sub001036_groupi_g4556__5107(csa_tree_sub001036_groupi_n_1448 ,csa_tree_sub001036_groupi_n_1407 ,csa_tree_sub001036_groupi_n_1441);
  xnor csa_tree_sub001036_groupi_g4557__6260(out1[5] ,csa_tree_sub001036_groupi_n_1425 ,csa_tree_sub001036_groupi_n_1422);
  not csa_tree_sub001036_groupi_g4558(csa_tree_sub001036_groupi_n_1446 ,csa_tree_sub001036_groupi_n_1445);
  xnor csa_tree_sub001036_groupi_g4559__4319(csa_tree_sub001036_groupi_n_1445 ,csa_tree_sub001036_groupi_n_1388 ,csa_tree_sub001036_groupi_n_1421);
  not csa_tree_sub001036_groupi_g4560(csa_tree_sub001036_groupi_n_1444 ,csa_tree_sub001036_groupi_n_1443);
  xnor csa_tree_sub001036_groupi_g4561__8428(csa_tree_sub001036_groupi_n_1443 ,csa_tree_sub001036_groupi_n_1383 ,csa_tree_sub001036_groupi_n_1420);
  not csa_tree_sub001036_groupi_g4562(csa_tree_sub001036_groupi_n_1442 ,csa_tree_sub001036_groupi_n_1441);
  and csa_tree_sub001036_groupi_g4563__5526(csa_tree_sub001036_groupi_n_1441 ,csa_tree_sub001036_groupi_n_1410 ,csa_tree_sub001036_groupi_n_1429);
  not csa_tree_sub001036_groupi_g4564(csa_tree_sub001036_groupi_n_1440 ,csa_tree_sub001036_groupi_n_1439);
  and csa_tree_sub001036_groupi_g4565__6783(csa_tree_sub001036_groupi_n_1439 ,csa_tree_sub001036_groupi_n_1428 ,csa_tree_sub001036_groupi_n_1414);
  or csa_tree_sub001036_groupi_g4566__3680(csa_tree_sub001036_groupi_n_1438 ,csa_tree_sub001036_groupi_n_1426 ,csa_tree_sub001036_groupi_n_1406);
  not csa_tree_sub001036_groupi_g4567(csa_tree_sub001036_groupi_n_1437 ,csa_tree_sub001036_groupi_n_1436);
  and csa_tree_sub001036_groupi_g4568__1617(csa_tree_sub001036_groupi_n_1436 ,csa_tree_sub001036_groupi_n_1424 ,csa_tree_sub001036_groupi_n_1404);
  xnor csa_tree_sub001036_groupi_g4569__2802(csa_tree_sub001036_groupi_n_1435 ,csa_tree_sub001036_groupi_n_1320 ,csa_tree_sub001036_groupi_n_1416);
  xnor csa_tree_sub001036_groupi_g4570__1705(csa_tree_sub001036_groupi_n_1434 ,csa_tree_sub001036_groupi_n_1409 ,csa_tree_sub001036_groupi_n_1418);
  xnor csa_tree_sub001036_groupi_g4571__5122(out1[4] ,csa_tree_sub001036_groupi_n_1386 ,csa_tree_sub001036_groupi_n_1400);
  xnor csa_tree_sub001036_groupi_g4572__8246(csa_tree_sub001036_groupi_n_1432 ,csa_tree_sub001036_groupi_n_4 ,csa_tree_sub001036_groupi_n_1401);
  and csa_tree_sub001036_groupi_g4573__7098(csa_tree_sub001036_groupi_n_1431 ,csa_tree_sub001036_groupi_n_1319 ,csa_tree_sub001036_groupi_n_1416);
  and csa_tree_sub001036_groupi_g4574__6131(csa_tree_sub001036_groupi_n_1430 ,csa_tree_sub001036_groupi_n_1320 ,csa_tree_sub001036_groupi_n_1415);
  or csa_tree_sub001036_groupi_g4575__1881(csa_tree_sub001036_groupi_n_1429 ,csa_tree_sub001036_groupi_n_1413 ,csa_tree_sub001036_groupi_n_1383);
  or csa_tree_sub001036_groupi_g4576__5115(csa_tree_sub001036_groupi_n_1428 ,csa_tree_sub001036_groupi_n_1389 ,csa_tree_sub001036_groupi_n_1411);
  nor csa_tree_sub001036_groupi_g4577__7482(csa_tree_sub001036_groupi_n_1427 ,csa_tree_sub001036_groupi_n_1409 ,csa_tree_sub001036_groupi_n_1419);
  not csa_tree_sub001036_groupi_g4578(csa_tree_sub001036_groupi_n_1426 ,csa_tree_sub001036_groupi_n_1425);
  or csa_tree_sub001036_groupi_g4579__4733(csa_tree_sub001036_groupi_n_1424 ,csa_tree_sub001036_groupi_n_1388 ,csa_tree_sub001036_groupi_n_1405);
  and csa_tree_sub001036_groupi_g4580__6161(csa_tree_sub001036_groupi_n_1423 ,csa_tree_sub001036_groupi_n_1409 ,csa_tree_sub001036_groupi_n_1419);
  xnor csa_tree_sub001036_groupi_g4581__9315(csa_tree_sub001036_groupi_n_1422 ,csa_tree_sub001036_groupi_n_1393 ,csa_tree_sub001036_groupi_n_1381);
  xnor csa_tree_sub001036_groupi_g4582__9945(csa_tree_sub001036_groupi_n_1421 ,csa_tree_sub001036_groupi_n_1394 ,csa_tree_sub001036_groupi_n_1367);
  xnor csa_tree_sub001036_groupi_g4583__2883(csa_tree_sub001036_groupi_n_1420 ,csa_tree_sub001036_groupi_n_1358 ,csa_tree_sub001036_groupi_n_1391);
  or csa_tree_sub001036_groupi_g4584__2346(csa_tree_sub001036_groupi_n_1425 ,csa_tree_sub001036_groupi_n_1396 ,csa_tree_sub001036_groupi_n_1412);
  not csa_tree_sub001036_groupi_g4585(csa_tree_sub001036_groupi_n_1419 ,csa_tree_sub001036_groupi_n_1418);
  not csa_tree_sub001036_groupi_g4586(csa_tree_sub001036_groupi_n_1415 ,csa_tree_sub001036_groupi_n_1416);
  or csa_tree_sub001036_groupi_g4587__1666(csa_tree_sub001036_groupi_n_1414 ,csa_tree_sub001036_groupi_n_4 ,csa_tree_sub001036_groupi_n_1365);
  nor csa_tree_sub001036_groupi_g4588__7410(csa_tree_sub001036_groupi_n_1413 ,csa_tree_sub001036_groupi_n_1358 ,csa_tree_sub001036_groupi_n_1391);
  and csa_tree_sub001036_groupi_g4589__6417(csa_tree_sub001036_groupi_n_1412 ,csa_tree_sub001036_groupi_n_1395 ,csa_tree_sub001036_groupi_n_1386);
  and csa_tree_sub001036_groupi_g4590__5477(csa_tree_sub001036_groupi_n_1411 ,csa_tree_sub001036_groupi_n_4 ,csa_tree_sub001036_groupi_n_1365);
  or csa_tree_sub001036_groupi_g4591__2398(csa_tree_sub001036_groupi_n_1410 ,csa_tree_sub001036_groupi_n_1357 ,csa_tree_sub001036_groupi_n_1390);
  or csa_tree_sub001036_groupi_g4592__5107(csa_tree_sub001036_groupi_n_1418 ,csa_tree_sub001036_groupi_n_1385 ,csa_tree_sub001036_groupi_n_1397);
  or csa_tree_sub001036_groupi_g4593__6260(csa_tree_sub001036_groupi_n_1417 ,csa_tree_sub001036_groupi_n_1398 ,csa_tree_sub001036_groupi_n_1376);
  or csa_tree_sub001036_groupi_g4594__4319(csa_tree_sub001036_groupi_n_1416 ,csa_tree_sub001036_groupi_n_1351 ,csa_tree_sub001036_groupi_n_1399);
  not csa_tree_sub001036_groupi_g4595(csa_tree_sub001036_groupi_n_1408 ,csa_tree_sub001036_groupi_n_1407);
  nor csa_tree_sub001036_groupi_g4596__8428(csa_tree_sub001036_groupi_n_1406 ,csa_tree_sub001036_groupi_n_1393 ,csa_tree_sub001036_groupi_n_1381);
  nor csa_tree_sub001036_groupi_g4597__5526(csa_tree_sub001036_groupi_n_1405 ,csa_tree_sub001036_groupi_n_1394 ,csa_tree_sub001036_groupi_n_1367);
  or csa_tree_sub001036_groupi_g4598__6783(csa_tree_sub001036_groupi_n_1404 ,csa_tree_sub001036_groupi_n_5 ,csa_tree_sub001036_groupi_n_1366);
  or csa_tree_sub001036_groupi_g4599__3680(csa_tree_sub001036_groupi_n_1403 ,csa_tree_sub001036_groupi_n_1392 ,csa_tree_sub001036_groupi_n_1380);
  xnor csa_tree_sub001036_groupi_g4600__1617(out1[3] ,csa_tree_sub001036_groupi_n_1308 ,csa_tree_sub001036_groupi_n_1378);
  xor csa_tree_sub001036_groupi_g4601__2802(csa_tree_sub001036_groupi_n_1401 ,csa_tree_sub001036_groupi_n_1365 ,csa_tree_sub001036_groupi_n_1389);
  xnor csa_tree_sub001036_groupi_g4602__1705(csa_tree_sub001036_groupi_n_1400 ,csa_tree_sub001036_groupi_n_1336 ,csa_tree_sub001036_groupi_n_1379);
  xnor csa_tree_sub001036_groupi_g4603__5122(csa_tree_sub001036_groupi_n_1409 ,csa_tree_sub001036_groupi_n_1382 ,csa_tree_sub001036_groupi_n_1377);
  xnor csa_tree_sub001036_groupi_g4604__8246(csa_tree_sub001036_groupi_n_1407 ,csa_tree_sub001036_groupi_n_1387 ,csa_tree_sub001036_groupi_n_1364);
  and csa_tree_sub001036_groupi_g4605__7098(csa_tree_sub001036_groupi_n_1399 ,csa_tree_sub001036_groupi_n_1350 ,csa_tree_sub001036_groupi_n_1387);
  nor csa_tree_sub001036_groupi_g4606__6131(csa_tree_sub001036_groupi_n_1398 ,csa_tree_sub001036_groupi_n_1373 ,csa_tree_sub001036_groupi_n_1382);
  nor csa_tree_sub001036_groupi_g4607__1881(csa_tree_sub001036_groupi_n_1397 ,csa_tree_sub001036_groupi_n_1337 ,csa_tree_sub001036_groupi_n_1384);
  and csa_tree_sub001036_groupi_g4608__5115(csa_tree_sub001036_groupi_n_1396 ,csa_tree_sub001036_groupi_n_1336 ,csa_tree_sub001036_groupi_n_1379);
  or csa_tree_sub001036_groupi_g4609__7482(csa_tree_sub001036_groupi_n_1395 ,csa_tree_sub001036_groupi_n_1336 ,csa_tree_sub001036_groupi_n_1379);
  not csa_tree_sub001036_groupi_g4611(csa_tree_sub001036_groupi_n_1394 ,csa_tree_sub001036_groupi_n_5);
  not csa_tree_sub001036_groupi_g4613(csa_tree_sub001036_groupi_n_1393 ,csa_tree_sub001036_groupi_n_1392);
  xnor csa_tree_sub001036_groupi_g4614__4733(csa_tree_sub001036_groupi_n_1392 ,csa_tree_sub001036_groupi_n_1368 ,csa_tree_sub001036_groupi_n_1359);
  not csa_tree_sub001036_groupi_g4615(csa_tree_sub001036_groupi_n_1391 ,csa_tree_sub001036_groupi_n_1390);
  xnor csa_tree_sub001036_groupi_g4616__6161(csa_tree_sub001036_groupi_n_1390 ,csa_tree_sub001036_groupi_n_1311 ,csa_tree_sub001036_groupi_n_1360);
  nor csa_tree_sub001036_groupi_g4617__9315(csa_tree_sub001036_groupi_n_1385 ,csa_tree_sub001036_groupi_n_1325 ,csa_tree_sub001036_groupi_n_1368);
  and csa_tree_sub001036_groupi_g4618__9945(csa_tree_sub001036_groupi_n_1384 ,csa_tree_sub001036_groupi_n_1325 ,csa_tree_sub001036_groupi_n_1368);
  and csa_tree_sub001036_groupi_g4619__2883(csa_tree_sub001036_groupi_n_1389 ,csa_tree_sub001036_groupi_n_1356 ,csa_tree_sub001036_groupi_n_1374);
  and csa_tree_sub001036_groupi_g4620__2346(csa_tree_sub001036_groupi_n_1388 ,csa_tree_sub001036_groupi_n_1353 ,csa_tree_sub001036_groupi_n_1372);
  or csa_tree_sub001036_groupi_g4621__1666(csa_tree_sub001036_groupi_n_1387 ,csa_tree_sub001036_groupi_n_1354 ,csa_tree_sub001036_groupi_n_1375);
  or csa_tree_sub001036_groupi_g4622__7410(csa_tree_sub001036_groupi_n_1386 ,csa_tree_sub001036_groupi_n_1331 ,csa_tree_sub001036_groupi_n_1371);
  not csa_tree_sub001036_groupi_g4623(csa_tree_sub001036_groupi_n_1381 ,csa_tree_sub001036_groupi_n_1380);
  xnor csa_tree_sub001036_groupi_g4624__6417(csa_tree_sub001036_groupi_n_1378 ,csa_tree_sub001036_groupi_n_1247 ,csa_tree_sub001036_groupi_n_1347);
  xnor csa_tree_sub001036_groupi_g4625__5477(csa_tree_sub001036_groupi_n_1377 ,csa_tree_sub001036_groupi_n_1344 ,csa_tree_sub001036_groupi_n_1345);
  and csa_tree_sub001036_groupi_g4626__2398(csa_tree_sub001036_groupi_n_1383 ,csa_tree_sub001036_groupi_n_1341 ,csa_tree_sub001036_groupi_n_1369);
  xnor csa_tree_sub001036_groupi_g4627__5107(csa_tree_sub001036_groupi_n_1382 ,csa_tree_sub001036_groupi_n_1327 ,csa_tree_sub001036_groupi_n_1339);
  and csa_tree_sub001036_groupi_g4628__6260(csa_tree_sub001036_groupi_n_1380 ,csa_tree_sub001036_groupi_n_1316 ,csa_tree_sub001036_groupi_n_1370);
  xnor csa_tree_sub001036_groupi_g4629__4319(csa_tree_sub001036_groupi_n_1379 ,csa_tree_sub001036_groupi_n_1348 ,csa_tree_sub001036_groupi_n_1340);
  and csa_tree_sub001036_groupi_g4630__8428(csa_tree_sub001036_groupi_n_1376 ,csa_tree_sub001036_groupi_n_1344 ,csa_tree_sub001036_groupi_n_1345);
  and csa_tree_sub001036_groupi_g4631__5526(csa_tree_sub001036_groupi_n_1375 ,csa_tree_sub001036_groupi_n_1311 ,csa_tree_sub001036_groupi_n_1352);
  or csa_tree_sub001036_groupi_g4632__6783(csa_tree_sub001036_groupi_n_1374 ,csa_tree_sub001036_groupi_n_1297 ,csa_tree_sub001036_groupi_n_1349);
  nor csa_tree_sub001036_groupi_g4633__3680(csa_tree_sub001036_groupi_n_1373 ,csa_tree_sub001036_groupi_n_1344 ,csa_tree_sub001036_groupi_n_1345);
  or csa_tree_sub001036_groupi_g4634__1617(csa_tree_sub001036_groupi_n_1372 ,csa_tree_sub001036_groupi_n_1338 ,csa_tree_sub001036_groupi_n_1355);
  and csa_tree_sub001036_groupi_g4635__2802(csa_tree_sub001036_groupi_n_1371 ,csa_tree_sub001036_groupi_n_1332 ,csa_tree_sub001036_groupi_n_1347);
  or csa_tree_sub001036_groupi_g4636__1705(csa_tree_sub001036_groupi_n_1370 ,csa_tree_sub001036_groupi_n_1315 ,csa_tree_sub001036_groupi_n_1348);
  or csa_tree_sub001036_groupi_g4637__5122(csa_tree_sub001036_groupi_n_1369 ,csa_tree_sub001036_groupi_n_1342 ,csa_tree_sub001036_groupi_n_1346);
  not csa_tree_sub001036_groupi_g4638(csa_tree_sub001036_groupi_n_1367 ,csa_tree_sub001036_groupi_n_1366);
  xnor csa_tree_sub001036_groupi_g4639__8246(csa_tree_sub001036_groupi_n_1364 ,csa_tree_sub001036_groupi_n_1296 ,csa_tree_sub001036_groupi_n_1335);
  xnor csa_tree_sub001036_groupi_g4640__7098(csa_tree_sub001036_groupi_n_1363 ,csa_tree_sub001036_groupi_n_1310 ,csa_tree_sub001036_groupi_n_1324);
  xnor csa_tree_sub001036_groupi_g4641__6131(csa_tree_sub001036_groupi_n_1362 ,csa_tree_sub001036_groupi_n_1328 ,csa_tree_sub001036_groupi_n_505);
  xnor csa_tree_sub001036_groupi_g4642__1881(csa_tree_sub001036_groupi_n_1361 ,csa_tree_sub001036_groupi_n_1306 ,csa_tree_sub001036_groupi_n_1318);
  xnor csa_tree_sub001036_groupi_g4643__5115(csa_tree_sub001036_groupi_n_1360 ,csa_tree_sub001036_groupi_n_1222 ,csa_tree_sub001036_groupi_n_1322);
  xnor csa_tree_sub001036_groupi_g4644__7482(csa_tree_sub001036_groupi_n_1359 ,csa_tree_sub001036_groupi_n_1325 ,csa_tree_sub001036_groupi_n_1337);
  xnor csa_tree_sub001036_groupi_g4645__4733(csa_tree_sub001036_groupi_n_1368 ,csa_tree_sub001036_groupi_n_1269 ,csa_tree_sub001036_groupi_n_1314);
  xnor csa_tree_sub001036_groupi_g4646__6161(csa_tree_sub001036_groupi_n_1366 ,csa_tree_sub001036_groupi_n_1261 ,csa_tree_sub001036_groupi_n_1313);
  xnor csa_tree_sub001036_groupi_g4647__9315(csa_tree_sub001036_groupi_n_1365 ,csa_tree_sub001036_groupi_n_1282 ,csa_tree_sub001036_groupi_n_1312);
  not csa_tree_sub001036_groupi_g4648(csa_tree_sub001036_groupi_n_1357 ,csa_tree_sub001036_groupi_n_1358);
  or csa_tree_sub001036_groupi_g4649__9945(csa_tree_sub001036_groupi_n_1356 ,csa_tree_sub001036_groupi_n_1266 ,csa_tree_sub001036_groupi_n_1326);
  nor csa_tree_sub001036_groupi_g4650__2883(csa_tree_sub001036_groupi_n_1355 ,csa_tree_sub001036_groupi_n_1310 ,csa_tree_sub001036_groupi_n_1323);
  nor csa_tree_sub001036_groupi_g4651__2346(csa_tree_sub001036_groupi_n_1354 ,csa_tree_sub001036_groupi_n_1221 ,csa_tree_sub001036_groupi_n_1322);
  or csa_tree_sub001036_groupi_g4652__1666(csa_tree_sub001036_groupi_n_1353 ,csa_tree_sub001036_groupi_n_1309 ,csa_tree_sub001036_groupi_n_1324);
  or csa_tree_sub001036_groupi_g4653__7410(csa_tree_sub001036_groupi_n_1352 ,csa_tree_sub001036_groupi_n_1222 ,csa_tree_sub001036_groupi_n_1321);
  nor csa_tree_sub001036_groupi_g4654__6417(csa_tree_sub001036_groupi_n_1351 ,csa_tree_sub001036_groupi_n_1296 ,csa_tree_sub001036_groupi_n_1334);
  or csa_tree_sub001036_groupi_g4655__5477(csa_tree_sub001036_groupi_n_1350 ,csa_tree_sub001036_groupi_n_1295 ,csa_tree_sub001036_groupi_n_1335);
  nor csa_tree_sub001036_groupi_g4656__2398(csa_tree_sub001036_groupi_n_1349 ,csa_tree_sub001036_groupi_n_1267 ,csa_tree_sub001036_groupi_n_1327);
  or csa_tree_sub001036_groupi_g4657__5107(csa_tree_sub001036_groupi_n_1358 ,csa_tree_sub001036_groupi_n_1300 ,csa_tree_sub001036_groupi_n_1333);
  xnor csa_tree_sub001036_groupi_g4659__6260(out1[2] ,csa_tree_sub001036_groupi_n_1128 ,csa_tree_sub001036_groupi_n_3);
  nor csa_tree_sub001036_groupi_g4660__4319(csa_tree_sub001036_groupi_n_1342 ,csa_tree_sub001036_groupi_n_1305 ,csa_tree_sub001036_groupi_n_1318);
  or csa_tree_sub001036_groupi_g4661__8428(csa_tree_sub001036_groupi_n_1341 ,csa_tree_sub001036_groupi_n_1306 ,csa_tree_sub001036_groupi_n_1317);
  xnor csa_tree_sub001036_groupi_g4662__5526(csa_tree_sub001036_groupi_n_1340 ,csa_tree_sub001036_groupi_n_1265 ,csa_tree_sub001036_groupi_n_1294);
  xnor csa_tree_sub001036_groupi_g4663__6783(csa_tree_sub001036_groupi_n_1339 ,csa_tree_sub001036_groupi_n_1267 ,csa_tree_sub001036_groupi_n_1297);
  xnor csa_tree_sub001036_groupi_g4664__3680(csa_tree_sub001036_groupi_n_1348 ,csa_tree_sub001036_groupi_n_1245 ,csa_tree_sub001036_groupi_n_1287);
  xnor csa_tree_sub001036_groupi_g4665__1617(csa_tree_sub001036_groupi_n_1347 ,csa_tree_sub001036_groupi_n_1270 ,csa_tree_sub001036_groupi_n_1288);
  and csa_tree_sub001036_groupi_g4666__2802(csa_tree_sub001036_groupi_n_1346 ,csa_tree_sub001036_groupi_n_1303 ,csa_tree_sub001036_groupi_n_1330);
  xnor csa_tree_sub001036_groupi_g4667__1705(csa_tree_sub001036_groupi_n_1345 ,csa_tree_sub001036_groupi_n_1253 ,csa_tree_sub001036_groupi_n_1286);
  or csa_tree_sub001036_groupi_g4668__5122(csa_tree_sub001036_groupi_n_1344 ,csa_tree_sub001036_groupi_n_1290 ,csa_tree_sub001036_groupi_n_1329);
  not csa_tree_sub001036_groupi_g4670(csa_tree_sub001036_groupi_n_1334 ,csa_tree_sub001036_groupi_n_1335);
  nor csa_tree_sub001036_groupi_g4671__8246(csa_tree_sub001036_groupi_n_1333 ,csa_tree_sub001036_groupi_n_1284 ,csa_tree_sub001036_groupi_n_1304);
  or csa_tree_sub001036_groupi_g4672__7098(csa_tree_sub001036_groupi_n_1332 ,csa_tree_sub001036_groupi_n_1246 ,csa_tree_sub001036_groupi_n_1307);
  nor csa_tree_sub001036_groupi_g4673__6131(csa_tree_sub001036_groupi_n_1331 ,csa_tree_sub001036_groupi_n_1247 ,csa_tree_sub001036_groupi_n_1308);
  or csa_tree_sub001036_groupi_g4674__1881(csa_tree_sub001036_groupi_n_1330 ,csa_tree_sub001036_groupi_n_1283 ,csa_tree_sub001036_groupi_n_1289);
  nor csa_tree_sub001036_groupi_g4675__5115(csa_tree_sub001036_groupi_n_1329 ,csa_tree_sub001036_groupi_n_1252 ,csa_tree_sub001036_groupi_n_1291);
  or csa_tree_sub001036_groupi_g4676__7482(csa_tree_sub001036_groupi_n_1328 ,csa_tree_sub001036_groupi_n_1197 ,csa_tree_sub001036_groupi_n_1299);
  and csa_tree_sub001036_groupi_g4677__4733(csa_tree_sub001036_groupi_n_1338 ,csa_tree_sub001036_groupi_n_1273 ,csa_tree_sub001036_groupi_n_1301);
  and csa_tree_sub001036_groupi_g4678__6161(csa_tree_sub001036_groupi_n_1337 ,csa_tree_sub001036_groupi_n_1277 ,csa_tree_sub001036_groupi_n_1302);
  or csa_tree_sub001036_groupi_g4679__9315(csa_tree_sub001036_groupi_n_1336 ,csa_tree_sub001036_groupi_n_1275 ,csa_tree_sub001036_groupi_n_1292);
  or csa_tree_sub001036_groupi_g4680__9945(csa_tree_sub001036_groupi_n_1335 ,csa_tree_sub001036_groupi_n_1260 ,csa_tree_sub001036_groupi_n_1298);
  not csa_tree_sub001036_groupi_g4681(csa_tree_sub001036_groupi_n_1327 ,csa_tree_sub001036_groupi_n_1326);
  not csa_tree_sub001036_groupi_g4682(csa_tree_sub001036_groupi_n_1324 ,csa_tree_sub001036_groupi_n_1323);
  not csa_tree_sub001036_groupi_g4683(csa_tree_sub001036_groupi_n_1322 ,csa_tree_sub001036_groupi_n_1321);
  not csa_tree_sub001036_groupi_g4684(csa_tree_sub001036_groupi_n_1319 ,csa_tree_sub001036_groupi_n_1320);
  not csa_tree_sub001036_groupi_g4685(csa_tree_sub001036_groupi_n_1318 ,csa_tree_sub001036_groupi_n_1317);
  or csa_tree_sub001036_groupi_g4686__2883(csa_tree_sub001036_groupi_n_1316 ,csa_tree_sub001036_groupi_n_1265 ,csa_tree_sub001036_groupi_n_1293);
  nor csa_tree_sub001036_groupi_g4687__2346(csa_tree_sub001036_groupi_n_1315 ,csa_tree_sub001036_groupi_n_1264 ,csa_tree_sub001036_groupi_n_1294);
  xnor csa_tree_sub001036_groupi_g4688__1666(csa_tree_sub001036_groupi_n_1314 ,csa_tree_sub001036_groupi_n_1252 ,csa_tree_sub001036_groupi_n_1268);
  xor csa_tree_sub001036_groupi_g4689__7410(csa_tree_sub001036_groupi_n_1313 ,csa_tree_sub001036_groupi_n_1225 ,csa_tree_sub001036_groupi_n_1284);
  xnor csa_tree_sub001036_groupi_g4690__6417(csa_tree_sub001036_groupi_n_1312 ,csa_tree_sub001036_groupi_n_1227 ,csa_tree_sub001036_groupi_n_1262);
  xnor csa_tree_sub001036_groupi_g4691__5477(csa_tree_sub001036_groupi_n_1326 ,csa_tree_sub001036_groupi_n_1213 ,csa_tree_sub001036_groupi_n_1254);
  xnor csa_tree_sub001036_groupi_g4692__2398(csa_tree_sub001036_groupi_n_1325 ,csa_tree_sub001036_groupi_n_1233 ,csa_tree_sub001036_groupi_n_1258);
  xnor csa_tree_sub001036_groupi_g4693__5107(csa_tree_sub001036_groupi_n_1323 ,csa_tree_sub001036_groupi_n_1251 ,csa_tree_sub001036_groupi_n_1257);
  xnor csa_tree_sub001036_groupi_g4694__6260(csa_tree_sub001036_groupi_n_1321 ,csa_tree_sub001036_groupi_n_1230 ,csa_tree_sub001036_groupi_n_1256);
  xnor csa_tree_sub001036_groupi_g4695__4319(csa_tree_sub001036_groupi_n_1320 ,csa_tree_sub001036_groupi_n_1285 ,csa_tree_sub001036_groupi_n_1216);
  xnor csa_tree_sub001036_groupi_g4696__8428(csa_tree_sub001036_groupi_n_1317 ,csa_tree_sub001036_groupi_n_1250 ,csa_tree_sub001036_groupi_n_1255);
  not csa_tree_sub001036_groupi_g4697(csa_tree_sub001036_groupi_n_1309 ,csa_tree_sub001036_groupi_n_1310);
  not csa_tree_sub001036_groupi_g4698(csa_tree_sub001036_groupi_n_1307 ,csa_tree_sub001036_groupi_n_1308);
  not csa_tree_sub001036_groupi_g4699(csa_tree_sub001036_groupi_n_1306 ,csa_tree_sub001036_groupi_n_1305);
  and csa_tree_sub001036_groupi_g4700__5526(csa_tree_sub001036_groupi_n_1304 ,csa_tree_sub001036_groupi_n_1226 ,csa_tree_sub001036_groupi_n_1261);
  or csa_tree_sub001036_groupi_g4701__6783(csa_tree_sub001036_groupi_n_1303 ,csa_tree_sub001036_groupi_n_1227 ,csa_tree_sub001036_groupi_n_1263);
  or csa_tree_sub001036_groupi_g4702__3680(csa_tree_sub001036_groupi_n_1302 ,csa_tree_sub001036_groupi_n_1214 ,csa_tree_sub001036_groupi_n_1276);
  or csa_tree_sub001036_groupi_g4703__1617(csa_tree_sub001036_groupi_n_1301 ,csa_tree_sub001036_groupi_n_1253 ,csa_tree_sub001036_groupi_n_1278);
  nor csa_tree_sub001036_groupi_g4704__2802(csa_tree_sub001036_groupi_n_1300 ,csa_tree_sub001036_groupi_n_1226 ,csa_tree_sub001036_groupi_n_1261);
  and csa_tree_sub001036_groupi_g4705__1705(csa_tree_sub001036_groupi_n_1299 ,csa_tree_sub001036_groupi_n_1187 ,csa_tree_sub001036_groupi_n_1285);
  and csa_tree_sub001036_groupi_g4706__5122(csa_tree_sub001036_groupi_n_1298 ,csa_tree_sub001036_groupi_n_1196 ,csa_tree_sub001036_groupi_n_1281);
  or csa_tree_sub001036_groupi_g4707__8246(csa_tree_sub001036_groupi_n_1311 ,csa_tree_sub001036_groupi_n_1219 ,csa_tree_sub001036_groupi_n_1271);
  or csa_tree_sub001036_groupi_g4708__7098(csa_tree_sub001036_groupi_n_1310 ,csa_tree_sub001036_groupi_n_1240 ,csa_tree_sub001036_groupi_n_1280);
  and csa_tree_sub001036_groupi_g4709__6131(csa_tree_sub001036_groupi_n_1308 ,csa_tree_sub001036_groupi_n_1142 ,csa_tree_sub001036_groupi_n_1272);
  or csa_tree_sub001036_groupi_g4710__1881(csa_tree_sub001036_groupi_n_1305 ,csa_tree_sub001036_groupi_n_1243 ,csa_tree_sub001036_groupi_n_1279);
  not csa_tree_sub001036_groupi_g4711(csa_tree_sub001036_groupi_n_1296 ,csa_tree_sub001036_groupi_n_1295);
  not csa_tree_sub001036_groupi_g4712(csa_tree_sub001036_groupi_n_1294 ,csa_tree_sub001036_groupi_n_1293);
  nor csa_tree_sub001036_groupi_g4713__5115(csa_tree_sub001036_groupi_n_1292 ,csa_tree_sub001036_groupi_n_1274 ,csa_tree_sub001036_groupi_n_1270);
  nor csa_tree_sub001036_groupi_g4714__7482(csa_tree_sub001036_groupi_n_1291 ,csa_tree_sub001036_groupi_n_1269 ,csa_tree_sub001036_groupi_n_1268);
  and csa_tree_sub001036_groupi_g4715__4733(csa_tree_sub001036_groupi_n_1290 ,csa_tree_sub001036_groupi_n_1269 ,csa_tree_sub001036_groupi_n_1268);
  and csa_tree_sub001036_groupi_g4716__6161(csa_tree_sub001036_groupi_n_1289 ,csa_tree_sub001036_groupi_n_1227 ,csa_tree_sub001036_groupi_n_1263);
  xnor csa_tree_sub001036_groupi_g4717__9315(csa_tree_sub001036_groupi_n_1288 ,csa_tree_sub001036_groupi_n_1153 ,csa_tree_sub001036_groupi_n_1223);
  xnor csa_tree_sub001036_groupi_g4718__9945(csa_tree_sub001036_groupi_n_1287 ,csa_tree_sub001036_groupi_n_1214 ,csa_tree_sub001036_groupi_n_1232);
  xnor csa_tree_sub001036_groupi_g4720__2883(csa_tree_sub001036_groupi_n_1286 ,csa_tree_sub001036_groupi_n_1249 ,csa_tree_sub001036_groupi_n_1229);
  and csa_tree_sub001036_groupi_g4721__2346(csa_tree_sub001036_groupi_n_1297 ,csa_tree_sub001036_groupi_n_1242 ,csa_tree_sub001036_groupi_n_1259);
  xnor csa_tree_sub001036_groupi_g4722__1666(csa_tree_sub001036_groupi_n_1295 ,csa_tree_sub001036_groupi_n_1195 ,csa_tree_sub001036_groupi_n_1217);
  xnor csa_tree_sub001036_groupi_g4723__7410(csa_tree_sub001036_groupi_n_1293 ,csa_tree_sub001036_groupi_n_1123 ,csa_tree_sub001036_groupi_n_1215);
  not csa_tree_sub001036_groupi_g4724(csa_tree_sub001036_groupi_n_1283 ,csa_tree_sub001036_groupi_n_1282);
  or csa_tree_sub001036_groupi_g4725__6417(csa_tree_sub001036_groupi_n_1281 ,csa_tree_sub001036_groupi_n_1148 ,csa_tree_sub001036_groupi_n_1231);
  and csa_tree_sub001036_groupi_g4726__5477(csa_tree_sub001036_groupi_n_1280 ,csa_tree_sub001036_groupi_n_1213 ,csa_tree_sub001036_groupi_n_1239);
  nor csa_tree_sub001036_groupi_g4727__2398(csa_tree_sub001036_groupi_n_1279 ,csa_tree_sub001036_groupi_n_1238 ,csa_tree_sub001036_groupi_n_1251);
  nor csa_tree_sub001036_groupi_g4728__5107(csa_tree_sub001036_groupi_n_1278 ,csa_tree_sub001036_groupi_n_1248 ,csa_tree_sub001036_groupi_n_1229);
  or csa_tree_sub001036_groupi_g4729__6260(csa_tree_sub001036_groupi_n_1277 ,csa_tree_sub001036_groupi_n_156 ,csa_tree_sub001036_groupi_n_1244);
  nor csa_tree_sub001036_groupi_g4730__4319(csa_tree_sub001036_groupi_n_1276 ,csa_tree_sub001036_groupi_n_48 ,csa_tree_sub001036_groupi_n_1245);
  nor csa_tree_sub001036_groupi_g4731__8428(csa_tree_sub001036_groupi_n_1275 ,csa_tree_sub001036_groupi_n_1153 ,csa_tree_sub001036_groupi_n_1224);
  and csa_tree_sub001036_groupi_g4732__5526(csa_tree_sub001036_groupi_n_1274 ,csa_tree_sub001036_groupi_n_1153 ,csa_tree_sub001036_groupi_n_1224);
  or csa_tree_sub001036_groupi_g4733__6783(csa_tree_sub001036_groupi_n_1273 ,csa_tree_sub001036_groupi_n_1249 ,csa_tree_sub001036_groupi_n_1228);
  or csa_tree_sub001036_groupi_g4734__3680(csa_tree_sub001036_groupi_n_1272 ,csa_tree_sub001036_groupi_n_1168 ,csa_tree_sub001036_groupi_n_1235);
  and csa_tree_sub001036_groupi_g4735__1617(csa_tree_sub001036_groupi_n_1271 ,csa_tree_sub001036_groupi_n_1220 ,csa_tree_sub001036_groupi_n_1250);
  or csa_tree_sub001036_groupi_g4736__2802(csa_tree_sub001036_groupi_n_1285 ,csa_tree_sub001036_groupi_n_1185 ,csa_tree_sub001036_groupi_n_1218);
  and csa_tree_sub001036_groupi_g4737__1705(csa_tree_sub001036_groupi_n_1284 ,csa_tree_sub001036_groupi_n_1201 ,csa_tree_sub001036_groupi_n_1241);
  or csa_tree_sub001036_groupi_g4738__5122(csa_tree_sub001036_groupi_n_1282 ,csa_tree_sub001036_groupi_n_1204 ,csa_tree_sub001036_groupi_n_1237);
  not csa_tree_sub001036_groupi_g4739(csa_tree_sub001036_groupi_n_1267 ,csa_tree_sub001036_groupi_n_1266);
  not csa_tree_sub001036_groupi_g4740(csa_tree_sub001036_groupi_n_1265 ,csa_tree_sub001036_groupi_n_1264);
  not csa_tree_sub001036_groupi_g4741(csa_tree_sub001036_groupi_n_1263 ,csa_tree_sub001036_groupi_n_1262);
  and csa_tree_sub001036_groupi_g4742__8246(csa_tree_sub001036_groupi_n_1260 ,csa_tree_sub001036_groupi_n_1148 ,csa_tree_sub001036_groupi_n_1231);
  or csa_tree_sub001036_groupi_g4743__7098(csa_tree_sub001036_groupi_n_1259 ,csa_tree_sub001036_groupi_n_1234 ,csa_tree_sub001036_groupi_n_1236);
  xnor csa_tree_sub001036_groupi_g4744__6131(csa_tree_sub001036_groupi_n_1258 ,csa_tree_sub001036_groupi_n_1210 ,csa_tree_sub001036_groupi_n_1194);
  xnor csa_tree_sub001036_groupi_g4745__1881(csa_tree_sub001036_groupi_n_1257 ,csa_tree_sub001036_groupi_n_1126 ,csa_tree_sub001036_groupi_n_1190);
  xor csa_tree_sub001036_groupi_g4746__5115(csa_tree_sub001036_groupi_n_1256 ,csa_tree_sub001036_groupi_n_1148 ,csa_tree_sub001036_groupi_n_1196);
  xnor csa_tree_sub001036_groupi_g4747__7482(csa_tree_sub001036_groupi_n_1255 ,csa_tree_sub001036_groupi_n_1212 ,csa_tree_sub001036_groupi_n_1097);
  xnor csa_tree_sub001036_groupi_g4748__4733(csa_tree_sub001036_groupi_n_1254 ,csa_tree_sub001036_groupi_n_1125 ,csa_tree_sub001036_groupi_n_1192);
  xnor csa_tree_sub001036_groupi_g4749__6161(csa_tree_sub001036_groupi_n_1270 ,csa_tree_sub001036_groupi_n_1155 ,csa_tree_sub001036_groupi_n_1179);
  xnor csa_tree_sub001036_groupi_g4750__9315(csa_tree_sub001036_groupi_n_1269 ,csa_tree_sub001036_groupi_n_1135 ,csa_tree_sub001036_groupi_n_1181);
  xnor csa_tree_sub001036_groupi_g4751__9945(csa_tree_sub001036_groupi_n_1268 ,csa_tree_sub001036_groupi_n_1157 ,csa_tree_sub001036_groupi_n_1180);
  xnor csa_tree_sub001036_groupi_g4752__2883(csa_tree_sub001036_groupi_n_1266 ,csa_tree_sub001036_groupi_n_1154 ,csa_tree_sub001036_groupi_n_1184);
  xnor csa_tree_sub001036_groupi_g4753__2346(csa_tree_sub001036_groupi_n_1264 ,csa_tree_sub001036_groupi_n_1106 ,csa_tree_sub001036_groupi_n_1182);
  xnor csa_tree_sub001036_groupi_g4754__1666(csa_tree_sub001036_groupi_n_1262 ,csa_tree_sub001036_groupi_n_1152 ,csa_tree_sub001036_groupi_n_1183);
  xnor csa_tree_sub001036_groupi_g4755__7410(csa_tree_sub001036_groupi_n_1261 ,csa_tree_sub001036_groupi_n_1092 ,csa_tree_sub001036_groupi_n_2);
  not csa_tree_sub001036_groupi_g4756(csa_tree_sub001036_groupi_n_1249 ,csa_tree_sub001036_groupi_n_1248);
  not csa_tree_sub001036_groupi_g4757(csa_tree_sub001036_groupi_n_1247 ,csa_tree_sub001036_groupi_n_1246);
  not csa_tree_sub001036_groupi_g4758(csa_tree_sub001036_groupi_n_1244 ,csa_tree_sub001036_groupi_n_1245);
  nor csa_tree_sub001036_groupi_g4759__6417(csa_tree_sub001036_groupi_n_1243 ,csa_tree_sub001036_groupi_n_1127 ,csa_tree_sub001036_groupi_n_1190);
  or csa_tree_sub001036_groupi_g4760__5477(csa_tree_sub001036_groupi_n_1242 ,csa_tree_sub001036_groupi_n_1209 ,csa_tree_sub001036_groupi_n_1194);
  or csa_tree_sub001036_groupi_g4761__2398(csa_tree_sub001036_groupi_n_1241 ,csa_tree_sub001036_groupi_n_1131 ,csa_tree_sub001036_groupi_n_1200);
  nor csa_tree_sub001036_groupi_g4762__5107(csa_tree_sub001036_groupi_n_1240 ,csa_tree_sub001036_groupi_n_1124 ,csa_tree_sub001036_groupi_n_1192);
  or csa_tree_sub001036_groupi_g4763__6260(csa_tree_sub001036_groupi_n_1239 ,csa_tree_sub001036_groupi_n_1125 ,csa_tree_sub001036_groupi_n_1191);
  and csa_tree_sub001036_groupi_g4764__4319(csa_tree_sub001036_groupi_n_1238 ,csa_tree_sub001036_groupi_n_1127 ,csa_tree_sub001036_groupi_n_1190);
  nor csa_tree_sub001036_groupi_g4765__8428(csa_tree_sub001036_groupi_n_1237 ,csa_tree_sub001036_groupi_n_1079 ,csa_tree_sub001036_groupi_n_1203);
  nor csa_tree_sub001036_groupi_g4766__5526(csa_tree_sub001036_groupi_n_1236 ,csa_tree_sub001036_groupi_n_1210 ,csa_tree_sub001036_groupi_n_1193);
  and csa_tree_sub001036_groupi_g4767__6783(csa_tree_sub001036_groupi_n_1253 ,csa_tree_sub001036_groupi_n_1173 ,csa_tree_sub001036_groupi_n_1206);
  and csa_tree_sub001036_groupi_g4768__3680(csa_tree_sub001036_groupi_n_1252 ,csa_tree_sub001036_groupi_n_1164 ,csa_tree_sub001036_groupi_n_1199);
  and csa_tree_sub001036_groupi_g4769__1617(csa_tree_sub001036_groupi_n_1251 ,csa_tree_sub001036_groupi_n_1171 ,csa_tree_sub001036_groupi_n_1205);
  or csa_tree_sub001036_groupi_g4770__2802(csa_tree_sub001036_groupi_n_1250 ,csa_tree_sub001036_groupi_n_1167 ,csa_tree_sub001036_groupi_n_1202);
  or csa_tree_sub001036_groupi_g4771__1705(csa_tree_sub001036_groupi_n_1248 ,csa_tree_sub001036_groupi_n_1176 ,csa_tree_sub001036_groupi_n_1207);
  or csa_tree_sub001036_groupi_g4772__5122(csa_tree_sub001036_groupi_n_1246 ,csa_tree_sub001036_groupi_n_1049 ,csa_tree_sub001036_groupi_n_1188);
  or csa_tree_sub001036_groupi_g4773__8246(csa_tree_sub001036_groupi_n_1245 ,csa_tree_sub001036_groupi_n_1162 ,csa_tree_sub001036_groupi_n_1198);
  not csa_tree_sub001036_groupi_g4775(csa_tree_sub001036_groupi_n_1234 ,csa_tree_sub001036_groupi_n_1233);
  not csa_tree_sub001036_groupi_g4777(csa_tree_sub001036_groupi_n_1231 ,csa_tree_sub001036_groupi_n_1230);
  not csa_tree_sub001036_groupi_g4778(csa_tree_sub001036_groupi_n_1229 ,csa_tree_sub001036_groupi_n_1228);
  not csa_tree_sub001036_groupi_g4779(csa_tree_sub001036_groupi_n_1226 ,csa_tree_sub001036_groupi_n_1225);
  not csa_tree_sub001036_groupi_g4780(csa_tree_sub001036_groupi_n_1224 ,csa_tree_sub001036_groupi_n_1223);
  not csa_tree_sub001036_groupi_g4781(csa_tree_sub001036_groupi_n_1221 ,csa_tree_sub001036_groupi_n_1222);
  or csa_tree_sub001036_groupi_g4782__7098(csa_tree_sub001036_groupi_n_1220 ,csa_tree_sub001036_groupi_n_1212 ,csa_tree_sub001036_groupi_n_1096);
  nor csa_tree_sub001036_groupi_g4783__6131(csa_tree_sub001036_groupi_n_1219 ,csa_tree_sub001036_groupi_n_1211 ,csa_tree_sub001036_groupi_n_1097);
  and csa_tree_sub001036_groupi_g4784__1881(csa_tree_sub001036_groupi_n_1218 ,csa_tree_sub001036_groupi_n_1186 ,csa_tree_sub001036_groupi_n_1195);
  xnor csa_tree_sub001036_groupi_g4785__5115(csa_tree_sub001036_groupi_n_1217 ,csa_tree_sub001036_groupi_n_1150 ,csa_tree_sub001036_groupi_n_1104);
  xnor csa_tree_sub001036_groupi_g4786__7482(csa_tree_sub001036_groupi_n_1216 ,csa_tree_sub001036_groupi_n_1178 ,csa_tree_sub001036_groupi_n_47);
  xnor csa_tree_sub001036_groupi_g4787__4733(csa_tree_sub001036_groupi_n_1215 ,csa_tree_sub001036_groupi_n_1090 ,csa_tree_sub001036_groupi_n_1158);
  xnor csa_tree_sub001036_groupi_g4788__6161(csa_tree_sub001036_groupi_n_1235 ,csa_tree_sub001036_groupi_n_1156 ,csa_tree_sub001036_groupi_n_1083);
  or csa_tree_sub001036_groupi_g4789__9315(csa_tree_sub001036_groupi_n_1233 ,csa_tree_sub001036_groupi_n_1147 ,csa_tree_sub001036_groupi_n_1208);
  xnor csa_tree_sub001036_groupi_g4790__9945(csa_tree_sub001036_groupi_n_1232 ,csa_tree_sub001036_groupi_n_1082 ,csa_tree_sub001036_groupi_n_1136);
  and csa_tree_sub001036_groupi_g4791__2883(csa_tree_sub001036_groupi_n_1230 ,csa_tree_sub001036_groupi_n_1146 ,csa_tree_sub001036_groupi_n_1189);
  xnor csa_tree_sub001036_groupi_g4792__2346(csa_tree_sub001036_groupi_n_1228 ,csa_tree_sub001036_groupi_n_1102 ,csa_tree_sub001036_groupi_n_1139);
  xnor csa_tree_sub001036_groupi_g4793__1666(csa_tree_sub001036_groupi_n_1227 ,csa_tree_sub001036_groupi_n_1098 ,csa_tree_sub001036_groupi_n_1138);
  xnor csa_tree_sub001036_groupi_g4794__7410(csa_tree_sub001036_groupi_n_1225 ,csa_tree_sub001036_groupi_n_1076 ,csa_tree_sub001036_groupi_n_1137);
  xnor csa_tree_sub001036_groupi_g4795__6417(csa_tree_sub001036_groupi_n_1223 ,csa_tree_sub001036_groupi_n_1133 ,csa_tree_sub001036_groupi_n_1140);
  xnor csa_tree_sub001036_groupi_g4796__5477(csa_tree_sub001036_groupi_n_1222 ,csa_tree_sub001036_groupi_n_1077 ,csa_tree_sub001036_groupi_n_1141);
  not csa_tree_sub001036_groupi_g4797(csa_tree_sub001036_groupi_n_1211 ,csa_tree_sub001036_groupi_n_1212);
  not csa_tree_sub001036_groupi_g4798(csa_tree_sub001036_groupi_n_1209 ,csa_tree_sub001036_groupi_n_1210);
  nor csa_tree_sub001036_groupi_g4799__2398(csa_tree_sub001036_groupi_n_1208 ,csa_tree_sub001036_groupi_n_1110 ,csa_tree_sub001036_groupi_n_1177);
  nor csa_tree_sub001036_groupi_g4800__5107(csa_tree_sub001036_groupi_n_1207 ,csa_tree_sub001036_groupi_n_1135 ,csa_tree_sub001036_groupi_n_1175);
  or csa_tree_sub001036_groupi_g4801__6260(csa_tree_sub001036_groupi_n_1206 ,csa_tree_sub001036_groupi_n_1172 ,csa_tree_sub001036_groupi_n_1157);
  or csa_tree_sub001036_groupi_g4802__4319(csa_tree_sub001036_groupi_n_1205 ,csa_tree_sub001036_groupi_n_1080 ,csa_tree_sub001036_groupi_n_1170);
  and csa_tree_sub001036_groupi_g4803__8428(csa_tree_sub001036_groupi_n_1204 ,csa_tree_sub001036_groupi_n_1105 ,csa_tree_sub001036_groupi_n_1154);
  nor csa_tree_sub001036_groupi_g4804__5526(csa_tree_sub001036_groupi_n_1203 ,csa_tree_sub001036_groupi_n_1105 ,csa_tree_sub001036_groupi_n_1154);
  nor csa_tree_sub001036_groupi_g4805__6783(csa_tree_sub001036_groupi_n_1202 ,csa_tree_sub001036_groupi_n_1081 ,csa_tree_sub001036_groupi_n_1166);
  or csa_tree_sub001036_groupi_g4806__3680(csa_tree_sub001036_groupi_n_1201 ,csa_tree_sub001036_groupi_n_1095 ,csa_tree_sub001036_groupi_n_1151);
  nor csa_tree_sub001036_groupi_g4807__1617(csa_tree_sub001036_groupi_n_1200 ,csa_tree_sub001036_groupi_n_1094 ,csa_tree_sub001036_groupi_n_1152);
  or csa_tree_sub001036_groupi_g4808__2802(csa_tree_sub001036_groupi_n_1199 ,csa_tree_sub001036_groupi_n_1158 ,csa_tree_sub001036_groupi_n_1163);
  and csa_tree_sub001036_groupi_g4809__1705(csa_tree_sub001036_groupi_n_1198 ,csa_tree_sub001036_groupi_n_1161 ,csa_tree_sub001036_groupi_n_1155);
  and csa_tree_sub001036_groupi_g4810__5122(csa_tree_sub001036_groupi_n_1197 ,csa_tree_sub001036_groupi_n_57 ,csa_tree_sub001036_groupi_n_1178);
  and csa_tree_sub001036_groupi_g4811__8246(csa_tree_sub001036_groupi_n_1214 ,csa_tree_sub001036_groupi_n_1115 ,csa_tree_sub001036_groupi_n_1160);
  or csa_tree_sub001036_groupi_g4812__7098(csa_tree_sub001036_groupi_n_1213 ,csa_tree_sub001036_groupi_n_1119 ,csa_tree_sub001036_groupi_n_1169);
  or csa_tree_sub001036_groupi_g4813__6131(csa_tree_sub001036_groupi_n_1212 ,csa_tree_sub001036_groupi_n_1112 ,csa_tree_sub001036_groupi_n_1165);
  or csa_tree_sub001036_groupi_g4814__1881(csa_tree_sub001036_groupi_n_1210 ,csa_tree_sub001036_groupi_n_1118 ,csa_tree_sub001036_groupi_n_1159);
  not csa_tree_sub001036_groupi_g4815(csa_tree_sub001036_groupi_n_1193 ,csa_tree_sub001036_groupi_n_1194);
  not csa_tree_sub001036_groupi_g4816(csa_tree_sub001036_groupi_n_1192 ,csa_tree_sub001036_groupi_n_1191);
  or csa_tree_sub001036_groupi_g4817__5115(csa_tree_sub001036_groupi_n_1189 ,csa_tree_sub001036_groupi_n_1132 ,csa_tree_sub001036_groupi_n_1145);
  nor csa_tree_sub001036_groupi_g4818__7482(csa_tree_sub001036_groupi_n_1188 ,csa_tree_sub001036_groupi_n_1050 ,csa_tree_sub001036_groupi_n_1156);
  or csa_tree_sub001036_groupi_g4819__4733(csa_tree_sub001036_groupi_n_1187 ,csa_tree_sub001036_groupi_n_91 ,csa_tree_sub001036_groupi_n_1178);
  or csa_tree_sub001036_groupi_g4820__6161(csa_tree_sub001036_groupi_n_1186 ,csa_tree_sub001036_groupi_n_1103 ,csa_tree_sub001036_groupi_n_1149);
  nor csa_tree_sub001036_groupi_g4821__9315(csa_tree_sub001036_groupi_n_1185 ,csa_tree_sub001036_groupi_n_1104 ,csa_tree_sub001036_groupi_n_1150);
  xnor csa_tree_sub001036_groupi_g4822__9945(csa_tree_sub001036_groupi_n_1184 ,csa_tree_sub001036_groupi_n_1079 ,csa_tree_sub001036_groupi_n_1105);
  xnor csa_tree_sub001036_groupi_g4823__2883(csa_tree_sub001036_groupi_n_1183 ,csa_tree_sub001036_groupi_n_1095 ,csa_tree_sub001036_groupi_n_1131);
  xor csa_tree_sub001036_groupi_g4825__2346(csa_tree_sub001036_groupi_n_1182 ,csa_tree_sub001036_groupi_n_1110 ,csa_tree_sub001036_groupi_n_1033);
  xnor csa_tree_sub001036_groupi_g4826__1666(csa_tree_sub001036_groupi_n_1181 ,csa_tree_sub001036_groupi_n_1053 ,csa_tree_sub001036_groupi_n_1107);
  xnor csa_tree_sub001036_groupi_g4827__7410(csa_tree_sub001036_groupi_n_1180 ,csa_tree_sub001036_groupi_n_1130 ,csa_tree_sub001036_groupi_n_1100);
  xnor csa_tree_sub001036_groupi_g4828__6417(csa_tree_sub001036_groupi_n_1179 ,csa_tree_sub001036_groupi_n_1075 ,csa_tree_sub001036_groupi_n_1109);
  or csa_tree_sub001036_groupi_g4829__5477(csa_tree_sub001036_groupi_n_1196 ,csa_tree_sub001036_groupi_n_1088 ,csa_tree_sub001036_groupi_n_1144);
  or csa_tree_sub001036_groupi_g4830__2398(csa_tree_sub001036_groupi_n_1195 ,csa_tree_sub001036_groupi_n_1114 ,csa_tree_sub001036_groupi_n_1174);
  xnor csa_tree_sub001036_groupi_g4831__5107(csa_tree_sub001036_groupi_n_1194 ,csa_tree_sub001036_groupi_n_1072 ,csa_tree_sub001036_groupi_n_1084);
  xnor csa_tree_sub001036_groupi_g4832__6260(csa_tree_sub001036_groupi_n_1191 ,csa_tree_sub001036_groupi_n_982 ,csa_tree_sub001036_groupi_n_1086);
  xnor csa_tree_sub001036_groupi_g4833__4319(csa_tree_sub001036_groupi_n_1190 ,csa_tree_sub001036_groupi_n_1059 ,csa_tree_sub001036_groupi_n_1085);
  nor csa_tree_sub001036_groupi_g4834__8428(csa_tree_sub001036_groupi_n_1177 ,csa_tree_sub001036_groupi_n_1033 ,csa_tree_sub001036_groupi_n_1106);
  nor csa_tree_sub001036_groupi_g4835__5526(csa_tree_sub001036_groupi_n_1176 ,csa_tree_sub001036_groupi_n_1054 ,csa_tree_sub001036_groupi_n_1107);
  and csa_tree_sub001036_groupi_g4836__6783(csa_tree_sub001036_groupi_n_1175 ,csa_tree_sub001036_groupi_n_1054 ,csa_tree_sub001036_groupi_n_1107);
  and csa_tree_sub001036_groupi_g4837__3680(csa_tree_sub001036_groupi_n_1174 ,csa_tree_sub001036_groupi_n_1077 ,csa_tree_sub001036_groupi_n_1116);
  or csa_tree_sub001036_groupi_g4838__1617(csa_tree_sub001036_groupi_n_1173 ,csa_tree_sub001036_groupi_n_1129 ,csa_tree_sub001036_groupi_n_1100);
  nor csa_tree_sub001036_groupi_g4839__2802(csa_tree_sub001036_groupi_n_1172 ,csa_tree_sub001036_groupi_n_1130 ,csa_tree_sub001036_groupi_n_1099);
  or csa_tree_sub001036_groupi_g4840__1705(csa_tree_sub001036_groupi_n_1171 ,csa_tree_sub001036_groupi_n_1057 ,csa_tree_sub001036_groupi_n_1101);
  nor csa_tree_sub001036_groupi_g4841__5122(csa_tree_sub001036_groupi_n_1170 ,csa_tree_sub001036_groupi_n_1058 ,csa_tree_sub001036_groupi_n_1102);
  and csa_tree_sub001036_groupi_g4842__8246(csa_tree_sub001036_groupi_n_1169 ,csa_tree_sub001036_groupi_n_1037 ,csa_tree_sub001036_groupi_n_1111);
  and csa_tree_sub001036_groupi_g4843__7098(csa_tree_sub001036_groupi_n_1168 ,csa_tree_sub001036_groupi_n_1093 ,csa_tree_sub001036_groupi_n_1128);
  and csa_tree_sub001036_groupi_g4844__6131(csa_tree_sub001036_groupi_n_1167 ,csa_tree_sub001036_groupi_n_1071 ,csa_tree_sub001036_groupi_n_1098);
  nor csa_tree_sub001036_groupi_g4845__1881(csa_tree_sub001036_groupi_n_1166 ,csa_tree_sub001036_groupi_n_1071 ,csa_tree_sub001036_groupi_n_1098);
  nor csa_tree_sub001036_groupi_g4846__5115(csa_tree_sub001036_groupi_n_1165 ,csa_tree_sub001036_groupi_n_1038 ,csa_tree_sub001036_groupi_n_1113);
  or csa_tree_sub001036_groupi_g4847__7482(csa_tree_sub001036_groupi_n_1164 ,csa_tree_sub001036_groupi_n_1122 ,csa_tree_sub001036_groupi_n_1089);
  nor csa_tree_sub001036_groupi_g4848__4733(csa_tree_sub001036_groupi_n_1163 ,csa_tree_sub001036_groupi_n_1123 ,csa_tree_sub001036_groupi_n_1090);
  nor csa_tree_sub001036_groupi_g4849__6161(csa_tree_sub001036_groupi_n_1162 ,csa_tree_sub001036_groupi_n_1075 ,csa_tree_sub001036_groupi_n_1108);
  or csa_tree_sub001036_groupi_g4850__9315(csa_tree_sub001036_groupi_n_1161 ,csa_tree_sub001036_groupi_n_1074 ,csa_tree_sub001036_groupi_n_1109);
  or csa_tree_sub001036_groupi_g4851__9945(csa_tree_sub001036_groupi_n_1160 ,csa_tree_sub001036_groupi_n_1117 ,csa_tree_sub001036_groupi_n_1134);
  and csa_tree_sub001036_groupi_g4852__2883(csa_tree_sub001036_groupi_n_1159 ,csa_tree_sub001036_groupi_n_1082 ,csa_tree_sub001036_groupi_n_1120);
  or csa_tree_sub001036_groupi_g4853__2346(csa_tree_sub001036_groupi_n_1178 ,csa_tree_sub001036_groupi_n_831 ,csa_tree_sub001036_groupi_n_1121);
  not csa_tree_sub001036_groupi_g4854(csa_tree_sub001036_groupi_n_1152 ,csa_tree_sub001036_groupi_n_1151);
  not csa_tree_sub001036_groupi_g4855(csa_tree_sub001036_groupi_n_1149 ,csa_tree_sub001036_groupi_n_1150);
  and csa_tree_sub001036_groupi_g4856__1666(csa_tree_sub001036_groupi_n_1147 ,csa_tree_sub001036_groupi_n_1033 ,csa_tree_sub001036_groupi_n_1106);
  or csa_tree_sub001036_groupi_g4857__7410(csa_tree_sub001036_groupi_n_1146 ,csa_tree_sub001036_groupi_n_1056 ,csa_tree_sub001036_groupi_n_1091);
  nor csa_tree_sub001036_groupi_g4858__6417(csa_tree_sub001036_groupi_n_1145 ,csa_tree_sub001036_groupi_n_1 ,csa_tree_sub001036_groupi_n_1092);
  nor csa_tree_sub001036_groupi_g4859__5477(csa_tree_sub001036_groupi_n_1144 ,csa_tree_sub001036_groupi_n_1036 ,csa_tree_sub001036_groupi_n_1087);
  xnor csa_tree_sub001036_groupi_g4860__2398(out1[1] ,csa_tree_sub001036_groupi_n_645 ,csa_tree_sub001036_groupi_n_1046);
  or csa_tree_sub001036_groupi_g4861__5107(csa_tree_sub001036_groupi_n_1142 ,csa_tree_sub001036_groupi_n_1093 ,csa_tree_sub001036_groupi_n_1128);
  xnor csa_tree_sub001036_groupi_g4862__6260(csa_tree_sub001036_groupi_n_1141 ,csa_tree_sub001036_groupi_n_1052 ,csa_tree_sub001036_groupi_n_1061);
  xnor csa_tree_sub001036_groupi_g4863__4319(csa_tree_sub001036_groupi_n_1140 ,csa_tree_sub001036_groupi_n_1055 ,csa_tree_sub001036_groupi_n_1008);
  xnor csa_tree_sub001036_groupi_g4864__8428(csa_tree_sub001036_groupi_n_1139 ,csa_tree_sub001036_groupi_n_1058 ,csa_tree_sub001036_groupi_n_1080);
  xnor csa_tree_sub001036_groupi_g4865__5526(csa_tree_sub001036_groupi_n_1138 ,csa_tree_sub001036_groupi_n_1071 ,csa_tree_sub001036_groupi_n_1081);
  xnor csa_tree_sub001036_groupi_g4866__6783(csa_tree_sub001036_groupi_n_1137 ,csa_tree_sub001036_groupi_n_1035 ,csa_tree_sub001036_groupi_n_1073);
  xnor csa_tree_sub001036_groupi_g4867__3680(csa_tree_sub001036_groupi_n_1136 ,csa_tree_sub001036_groupi_n_921 ,csa_tree_sub001036_groupi_n_1060);
  xnor csa_tree_sub001036_groupi_g4868__1617(csa_tree_sub001036_groupi_n_1158 ,csa_tree_sub001036_groupi_n_939 ,csa_tree_sub001036_groupi_n_1041);
  xnor csa_tree_sub001036_groupi_g4869__2802(csa_tree_sub001036_groupi_n_1157 ,csa_tree_sub001036_groupi_n_947 ,csa_tree_sub001036_groupi_n_1042);
  xnor csa_tree_sub001036_groupi_g4870__1705(csa_tree_sub001036_groupi_n_1156 ,csa_tree_sub001036_groupi_n_948 ,csa_tree_sub001036_groupi_n_1043);
  xnor csa_tree_sub001036_groupi_g4871__5122(csa_tree_sub001036_groupi_n_1155 ,csa_tree_sub001036_groupi_n_949 ,csa_tree_sub001036_groupi_n_1045);
  xnor csa_tree_sub001036_groupi_g4872__8246(csa_tree_sub001036_groupi_n_1154 ,csa_tree_sub001036_groupi_n_944 ,csa_tree_sub001036_groupi_n_1044);
  xnor csa_tree_sub001036_groupi_g4873__7098(csa_tree_sub001036_groupi_n_1153 ,csa_tree_sub001036_groupi_n_943 ,csa_tree_sub001036_groupi_n_1047);
  xnor csa_tree_sub001036_groupi_g4874__6131(csa_tree_sub001036_groupi_n_1151 ,csa_tree_sub001036_groupi_n_946 ,csa_tree_sub001036_groupi_n_1040);
  xnor csa_tree_sub001036_groupi_g4875__1881(csa_tree_sub001036_groupi_n_1150 ,csa_tree_sub001036_groupi_n_1078 ,csa_tree_sub001036_groupi_n_0);
  xnor csa_tree_sub001036_groupi_g4876__5115(csa_tree_sub001036_groupi_n_1148 ,csa_tree_sub001036_groupi_n_1034 ,csa_tree_sub001036_groupi_n_1039);
  not csa_tree_sub001036_groupi_g4877(csa_tree_sub001036_groupi_n_1134 ,csa_tree_sub001036_groupi_n_1133);
  not csa_tree_sub001036_groupi_g4879(csa_tree_sub001036_groupi_n_1129 ,csa_tree_sub001036_groupi_n_1130);
  not csa_tree_sub001036_groupi_g4880(csa_tree_sub001036_groupi_n_1127 ,csa_tree_sub001036_groupi_n_1126);
  not csa_tree_sub001036_groupi_g4881(csa_tree_sub001036_groupi_n_1124 ,csa_tree_sub001036_groupi_n_1125);
  not csa_tree_sub001036_groupi_g4882(csa_tree_sub001036_groupi_n_1123 ,csa_tree_sub001036_groupi_n_1122);
  and csa_tree_sub001036_groupi_g4883__7482(csa_tree_sub001036_groupi_n_1121 ,csa_tree_sub001036_groupi_n_874 ,csa_tree_sub001036_groupi_n_1078);
  or csa_tree_sub001036_groupi_g4884__4733(csa_tree_sub001036_groupi_n_1120 ,csa_tree_sub001036_groupi_n_921 ,csa_tree_sub001036_groupi_n_1060);
  and csa_tree_sub001036_groupi_g4885__6161(csa_tree_sub001036_groupi_n_1119 ,csa_tree_sub001036_groupi_n_891 ,csa_tree_sub001036_groupi_n_1072);
  and csa_tree_sub001036_groupi_g4886__9315(csa_tree_sub001036_groupi_n_1118 ,csa_tree_sub001036_groupi_n_921 ,csa_tree_sub001036_groupi_n_1060);
  and csa_tree_sub001036_groupi_g4887__9945(csa_tree_sub001036_groupi_n_1117 ,csa_tree_sub001036_groupi_n_1008 ,csa_tree_sub001036_groupi_n_1055);
  or csa_tree_sub001036_groupi_g4888__2883(csa_tree_sub001036_groupi_n_1116 ,csa_tree_sub001036_groupi_n_1052 ,csa_tree_sub001036_groupi_n_1061);
  or csa_tree_sub001036_groupi_g4889__2346(csa_tree_sub001036_groupi_n_1115 ,csa_tree_sub001036_groupi_n_1008 ,csa_tree_sub001036_groupi_n_1055);
  and csa_tree_sub001036_groupi_g4890__1666(csa_tree_sub001036_groupi_n_1114 ,csa_tree_sub001036_groupi_n_1052 ,csa_tree_sub001036_groupi_n_1061);
  nor csa_tree_sub001036_groupi_g4891__7410(csa_tree_sub001036_groupi_n_1113 ,csa_tree_sub001036_groupi_n_880 ,csa_tree_sub001036_groupi_n_1059);
  and csa_tree_sub001036_groupi_g4892__6417(csa_tree_sub001036_groupi_n_1112 ,csa_tree_sub001036_groupi_n_880 ,csa_tree_sub001036_groupi_n_1059);
  or csa_tree_sub001036_groupi_g4893__5477(csa_tree_sub001036_groupi_n_1111 ,csa_tree_sub001036_groupi_n_891 ,csa_tree_sub001036_groupi_n_1072);
  and csa_tree_sub001036_groupi_g4894__2398(csa_tree_sub001036_groupi_n_1135 ,csa_tree_sub001036_groupi_n_1031 ,csa_tree_sub001036_groupi_n_1069);
  or csa_tree_sub001036_groupi_g4895__5107(csa_tree_sub001036_groupi_n_1133 ,csa_tree_sub001036_groupi_n_1003 ,csa_tree_sub001036_groupi_n_1068);
  and csa_tree_sub001036_groupi_g4896__6260(csa_tree_sub001036_groupi_n_1132 ,csa_tree_sub001036_groupi_n_1014 ,csa_tree_sub001036_groupi_n_1065);
  and csa_tree_sub001036_groupi_g4897__4319(csa_tree_sub001036_groupi_n_1131 ,csa_tree_sub001036_groupi_n_1017 ,csa_tree_sub001036_groupi_n_1062);
  or csa_tree_sub001036_groupi_g4898__8428(csa_tree_sub001036_groupi_n_1130 ,csa_tree_sub001036_groupi_n_1028 ,csa_tree_sub001036_groupi_n_1064);
  and csa_tree_sub001036_groupi_g4899__5526(csa_tree_sub001036_groupi_n_1128 ,csa_tree_sub001036_groupi_n_1000 ,csa_tree_sub001036_groupi_n_1051);
  or csa_tree_sub001036_groupi_g4900__6783(csa_tree_sub001036_groupi_n_1126 ,csa_tree_sub001036_groupi_n_1004 ,csa_tree_sub001036_groupi_n_1063);
  or csa_tree_sub001036_groupi_g4901__3680(csa_tree_sub001036_groupi_n_1125 ,csa_tree_sub001036_groupi_n_1018 ,csa_tree_sub001036_groupi_n_1067);
  and csa_tree_sub001036_groupi_g4902__1617(csa_tree_sub001036_groupi_n_1122 ,csa_tree_sub001036_groupi_n_1024 ,csa_tree_sub001036_groupi_n_1066);
  not csa_tree_sub001036_groupi_g4903(csa_tree_sub001036_groupi_n_1108 ,csa_tree_sub001036_groupi_n_1109);
  not csa_tree_sub001036_groupi_g4904(csa_tree_sub001036_groupi_n_1103 ,csa_tree_sub001036_groupi_n_1104);
  not csa_tree_sub001036_groupi_g4905(csa_tree_sub001036_groupi_n_1102 ,csa_tree_sub001036_groupi_n_1101);
  not csa_tree_sub001036_groupi_g4906(csa_tree_sub001036_groupi_n_1100 ,csa_tree_sub001036_groupi_n_1099);
  not csa_tree_sub001036_groupi_g4907(csa_tree_sub001036_groupi_n_1097 ,csa_tree_sub001036_groupi_n_1096);
  not csa_tree_sub001036_groupi_g4908(csa_tree_sub001036_groupi_n_1095 ,csa_tree_sub001036_groupi_n_1094);
  not csa_tree_sub001036_groupi_g4909(csa_tree_sub001036_groupi_n_1091 ,csa_tree_sub001036_groupi_n_1092);
  not csa_tree_sub001036_groupi_g4910(csa_tree_sub001036_groupi_n_1089 ,csa_tree_sub001036_groupi_n_1090);
  and csa_tree_sub001036_groupi_g4911__2802(csa_tree_sub001036_groupi_n_1088 ,csa_tree_sub001036_groupi_n_1073 ,csa_tree_sub001036_groupi_n_1076);
  nor csa_tree_sub001036_groupi_g4912__1705(csa_tree_sub001036_groupi_n_1087 ,csa_tree_sub001036_groupi_n_1073 ,csa_tree_sub001036_groupi_n_1076);
  xnor csa_tree_sub001036_groupi_g4913__5122(csa_tree_sub001036_groupi_n_1086 ,csa_tree_sub001036_groupi_n_937 ,csa_tree_sub001036_groupi_n_1010);
  xnor csa_tree_sub001036_groupi_g4914__8246(csa_tree_sub001036_groupi_n_1085 ,csa_tree_sub001036_groupi_n_880 ,csa_tree_sub001036_groupi_n_1038);
  xor csa_tree_sub001036_groupi_g4915__7098(csa_tree_sub001036_groupi_n_1084 ,csa_tree_sub001036_groupi_n_891 ,csa_tree_sub001036_groupi_n_1037);
  xnor csa_tree_sub001036_groupi_g4916__6131(csa_tree_sub001036_groupi_n_1083 ,csa_tree_sub001036_groupi_n_1009 ,csa_tree_sub001036_groupi_n_983);
  and csa_tree_sub001036_groupi_g4917__1881(csa_tree_sub001036_groupi_n_1110 ,csa_tree_sub001036_groupi_n_996 ,csa_tree_sub001036_groupi_n_1070);
  xnor csa_tree_sub001036_groupi_g4918__5115(csa_tree_sub001036_groupi_n_1109 ,csa_tree_sub001036_groupi_n_849 ,csa_tree_sub001036_groupi_n_985);
  xnor csa_tree_sub001036_groupi_g4919__7482(csa_tree_sub001036_groupi_n_1107 ,csa_tree_sub001036_groupi_n_940 ,csa_tree_sub001036_groupi_n_991);
  xnor csa_tree_sub001036_groupi_g4920__4733(csa_tree_sub001036_groupi_n_1106 ,csa_tree_sub001036_groupi_n_855 ,csa_tree_sub001036_groupi_n_988);
  xnor csa_tree_sub001036_groupi_g4921__6161(csa_tree_sub001036_groupi_n_1105 ,csa_tree_sub001036_groupi_n_861 ,csa_tree_sub001036_groupi_n_994);
  and csa_tree_sub001036_groupi_g4922__9315(csa_tree_sub001036_groupi_n_1104 ,csa_tree_sub001036_groupi_n_999 ,csa_tree_sub001036_groupi_n_1048);
  xnor csa_tree_sub001036_groupi_g4923__9945(csa_tree_sub001036_groupi_n_1101 ,csa_tree_sub001036_groupi_n_896 ,csa_tree_sub001036_groupi_n_993);
  xnor csa_tree_sub001036_groupi_g4924__2883(csa_tree_sub001036_groupi_n_1099 ,csa_tree_sub001036_groupi_n_898 ,csa_tree_sub001036_groupi_n_990);
  xnor csa_tree_sub001036_groupi_g4925__2346(csa_tree_sub001036_groupi_n_1098 ,csa_tree_sub001036_groupi_n_854 ,csa_tree_sub001036_groupi_n_989);
  xnor csa_tree_sub001036_groupi_g4926__1666(csa_tree_sub001036_groupi_n_1096 ,csa_tree_sub001036_groupi_n_942 ,csa_tree_sub001036_groupi_n_992);
  xnor csa_tree_sub001036_groupi_g4927__7410(csa_tree_sub001036_groupi_n_1094 ,csa_tree_sub001036_groupi_n_904 ,csa_tree_sub001036_groupi_n_995);
  xnor csa_tree_sub001036_groupi_g4928__6417(csa_tree_sub001036_groupi_n_1093 ,csa_tree_sub001036_groupi_n_866 ,csa_tree_sub001036_groupi_n_984);
  xnor csa_tree_sub001036_groupi_g4929__5477(csa_tree_sub001036_groupi_n_1092 ,csa_tree_sub001036_groupi_n_860 ,csa_tree_sub001036_groupi_n_987);
  xnor csa_tree_sub001036_groupi_g4930__2398(csa_tree_sub001036_groupi_n_1090 ,csa_tree_sub001036_groupi_n_924 ,csa_tree_sub001036_groupi_n_986);
  not csa_tree_sub001036_groupi_g4931(csa_tree_sub001036_groupi_n_1075 ,csa_tree_sub001036_groupi_n_1074);
  or csa_tree_sub001036_groupi_g4932__5107(csa_tree_sub001036_groupi_n_1070 ,csa_tree_sub001036_groupi_n_950 ,csa_tree_sub001036_groupi_n_1032);
  or csa_tree_sub001036_groupi_g4933__6260(csa_tree_sub001036_groupi_n_1069 ,csa_tree_sub001036_groupi_n_900 ,csa_tree_sub001036_groupi_n_1030);
  and csa_tree_sub001036_groupi_g4934__4319(csa_tree_sub001036_groupi_n_1068 ,csa_tree_sub001036_groupi_n_948 ,csa_tree_sub001036_groupi_n_1002);
  and csa_tree_sub001036_groupi_g4935__8428(csa_tree_sub001036_groupi_n_1067 ,csa_tree_sub001036_groupi_n_947 ,csa_tree_sub001036_groupi_n_1007);
  or csa_tree_sub001036_groupi_g4936__5526(csa_tree_sub001036_groupi_n_1066 ,csa_tree_sub001036_groupi_n_943 ,csa_tree_sub001036_groupi_n_1026);
  or csa_tree_sub001036_groupi_g4937__6783(csa_tree_sub001036_groupi_n_1065 ,csa_tree_sub001036_groupi_n_946 ,csa_tree_sub001036_groupi_n_1013);
  nor csa_tree_sub001036_groupi_g4938__3680(csa_tree_sub001036_groupi_n_1064 ,csa_tree_sub001036_groupi_n_903 ,csa_tree_sub001036_groupi_n_1027);
  and csa_tree_sub001036_groupi_g4939__1617(csa_tree_sub001036_groupi_n_1063 ,csa_tree_sub001036_groupi_n_1010 ,csa_tree_sub001036_groupi_n_1005);
  or csa_tree_sub001036_groupi_g4940__2802(csa_tree_sub001036_groupi_n_1062 ,csa_tree_sub001036_groupi_n_945 ,csa_tree_sub001036_groupi_n_1016);
  or csa_tree_sub001036_groupi_g4941__1705(csa_tree_sub001036_groupi_n_1082 ,csa_tree_sub001036_groupi_n_952 ,csa_tree_sub001036_groupi_n_1001);
  and csa_tree_sub001036_groupi_g4942__5122(csa_tree_sub001036_groupi_n_1081 ,csa_tree_sub001036_groupi_n_966 ,csa_tree_sub001036_groupi_n_1019);
  and csa_tree_sub001036_groupi_g4943__8246(csa_tree_sub001036_groupi_n_1080 ,csa_tree_sub001036_groupi_n_976 ,csa_tree_sub001036_groupi_n_1029);
  and csa_tree_sub001036_groupi_g4944__7098(csa_tree_sub001036_groupi_n_1079 ,csa_tree_sub001036_groupi_n_963 ,csa_tree_sub001036_groupi_n_998);
  or csa_tree_sub001036_groupi_g4945__6131(csa_tree_sub001036_groupi_n_1078 ,csa_tree_sub001036_groupi_n_978 ,csa_tree_sub001036_groupi_n_1023);
  or csa_tree_sub001036_groupi_g4946__1881(csa_tree_sub001036_groupi_n_1077 ,csa_tree_sub001036_groupi_n_977 ,csa_tree_sub001036_groupi_n_1025);
  or csa_tree_sub001036_groupi_g4947__5115(csa_tree_sub001036_groupi_n_1076 ,csa_tree_sub001036_groupi_n_961 ,csa_tree_sub001036_groupi_n_1012);
  or csa_tree_sub001036_groupi_g4948__7482(csa_tree_sub001036_groupi_n_1074 ,csa_tree_sub001036_groupi_n_957 ,csa_tree_sub001036_groupi_n_1006);
  or csa_tree_sub001036_groupi_g4949__4733(csa_tree_sub001036_groupi_n_1073 ,csa_tree_sub001036_groupi_n_969 ,csa_tree_sub001036_groupi_n_1011);
  or csa_tree_sub001036_groupi_g4950__6161(csa_tree_sub001036_groupi_n_1072 ,csa_tree_sub001036_groupi_n_975 ,csa_tree_sub001036_groupi_n_1022);
  or csa_tree_sub001036_groupi_g4951__9315(csa_tree_sub001036_groupi_n_1071 ,csa_tree_sub001036_groupi_n_968 ,csa_tree_sub001036_groupi_n_1020);
  not csa_tree_sub001036_groupi_g4952(csa_tree_sub001036_groupi_n_1057 ,csa_tree_sub001036_groupi_n_1058);
  not csa_tree_sub001036_groupi_g4953(csa_tree_sub001036_groupi_n_1056 ,csa_tree_sub001036_groupi_n_1);
  not csa_tree_sub001036_groupi_g4954(csa_tree_sub001036_groupi_n_1054 ,csa_tree_sub001036_groupi_n_1053);
  or csa_tree_sub001036_groupi_g4955__9945(csa_tree_sub001036_groupi_n_1051 ,csa_tree_sub001036_groupi_n_941 ,csa_tree_sub001036_groupi_n_1015);
  and csa_tree_sub001036_groupi_g4956__2883(csa_tree_sub001036_groupi_n_1050 ,csa_tree_sub001036_groupi_n_983 ,csa_tree_sub001036_groupi_n_1009);
  nor csa_tree_sub001036_groupi_g4957__2346(csa_tree_sub001036_groupi_n_1049 ,csa_tree_sub001036_groupi_n_983 ,csa_tree_sub001036_groupi_n_1009);
  or csa_tree_sub001036_groupi_g4958__1666(csa_tree_sub001036_groupi_n_1048 ,csa_tree_sub001036_groupi_n_1021 ,csa_tree_sub001036_groupi_n_1034);
  xnor csa_tree_sub001036_groupi_g4959__7410(csa_tree_sub001036_groupi_n_1047 ,csa_tree_sub001036_groupi_n_883 ,csa_tree_sub001036_groupi_n_932);
  xnor csa_tree_sub001036_groupi_g4960__6417(csa_tree_sub001036_groupi_n_1046 ,csa_tree_sub001036_groupi_n_941 ,csa_tree_sub001036_groupi_n_928);
  xnor csa_tree_sub001036_groupi_g4961__5477(csa_tree_sub001036_groupi_n_1045 ,csa_tree_sub001036_groupi_n_933 ,csa_tree_sub001036_groupi_n_839);
  xnor csa_tree_sub001036_groupi_g4962__2398(csa_tree_sub001036_groupi_n_1044 ,csa_tree_sub001036_groupi_n_914 ,csa_tree_sub001036_groupi_n_926);
  xnor csa_tree_sub001036_groupi_g4963__5107(csa_tree_sub001036_groupi_n_1043 ,csa_tree_sub001036_groupi_n_844 ,csa_tree_sub001036_groupi_n_920);
  xnor csa_tree_sub001036_groupi_g4964__6260(csa_tree_sub001036_groupi_n_1042 ,csa_tree_sub001036_groupi_n_923 ,csa_tree_sub001036_groupi_n_935);
  xor csa_tree_sub001036_groupi_g4965__4319(csa_tree_sub001036_groupi_n_1041 ,csa_tree_sub001036_groupi_n_930 ,csa_tree_sub001036_groupi_n_900);
  xnor csa_tree_sub001036_groupi_g4966__8428(csa_tree_sub001036_groupi_n_1040 ,csa_tree_sub001036_groupi_n_846 ,csa_tree_sub001036_groupi_n_918);
  xnor csa_tree_sub001036_groupi_g4967__5526(csa_tree_sub001036_groupi_n_1039 ,csa_tree_sub001036_groupi_n_842 ,csa_tree_sub001036_groupi_n_916);
  xnor csa_tree_sub001036_groupi_g4968__6783(csa_tree_sub001036_groupi_n_1061 ,csa_tree_sub001036_groupi_n_881 ,csa_tree_sub001036_groupi_n_906);
  xnor csa_tree_sub001036_groupi_g4969__3680(csa_tree_sub001036_groupi_n_1060 ,csa_tree_sub001036_groupi_n_759 ,csa_tree_sub001036_groupi_n_911);
  xnor csa_tree_sub001036_groupi_g4970__1617(csa_tree_sub001036_groupi_n_1059 ,csa_tree_sub001036_groupi_n_818 ,csa_tree_sub001036_groupi_n_909);
  xnor csa_tree_sub001036_groupi_g4971__2802(csa_tree_sub001036_groupi_n_1058 ,csa_tree_sub001036_groupi_n_822 ,csa_tree_sub001036_groupi_n_908);
  xnor csa_tree_sub001036_groupi_g4973__1705(csa_tree_sub001036_groupi_n_1055 ,csa_tree_sub001036_groupi_n_789 ,csa_tree_sub001036_groupi_n_907);
  xnor csa_tree_sub001036_groupi_g4974__5122(csa_tree_sub001036_groupi_n_1053 ,csa_tree_sub001036_groupi_n_760 ,csa_tree_sub001036_groupi_n_905);
  or csa_tree_sub001036_groupi_g4975__8246(csa_tree_sub001036_groupi_n_1052 ,csa_tree_sub001036_groupi_n_912 ,csa_tree_sub001036_groupi_n_997);
  not csa_tree_sub001036_groupi_g4976(csa_tree_sub001036_groupi_n_1036 ,csa_tree_sub001036_groupi_n_1035);
  and csa_tree_sub001036_groupi_g4977__7098(csa_tree_sub001036_groupi_n_1032 ,csa_tree_sub001036_groupi_n_839 ,csa_tree_sub001036_groupi_n_933);
  or csa_tree_sub001036_groupi_g4978__6131(csa_tree_sub001036_groupi_n_1031 ,csa_tree_sub001036_groupi_n_930 ,csa_tree_sub001036_groupi_n_938);
  nor csa_tree_sub001036_groupi_g4979__1881(csa_tree_sub001036_groupi_n_1030 ,csa_tree_sub001036_groupi_n_929 ,csa_tree_sub001036_groupi_n_939);
  or csa_tree_sub001036_groupi_g4980__5115(csa_tree_sub001036_groupi_n_1029 ,csa_tree_sub001036_groupi_n_899 ,csa_tree_sub001036_groupi_n_974);
  and csa_tree_sub001036_groupi_g4981__7482(csa_tree_sub001036_groupi_n_1028 ,csa_tree_sub001036_groupi_n_893 ,csa_tree_sub001036_groupi_n_924);
  nor csa_tree_sub001036_groupi_g4982__4733(csa_tree_sub001036_groupi_n_1027 ,csa_tree_sub001036_groupi_n_893 ,csa_tree_sub001036_groupi_n_924);
  nor csa_tree_sub001036_groupi_g4983__6161(csa_tree_sub001036_groupi_n_1026 ,csa_tree_sub001036_groupi_n_883 ,csa_tree_sub001036_groupi_n_932);
  and csa_tree_sub001036_groupi_g4984__9315(csa_tree_sub001036_groupi_n_1025 ,csa_tree_sub001036_groupi_n_973 ,csa_tree_sub001036_groupi_n_942);
  or csa_tree_sub001036_groupi_g4985__9945(csa_tree_sub001036_groupi_n_1024 ,csa_tree_sub001036_groupi_n_882 ,csa_tree_sub001036_groupi_n_931);
  nor csa_tree_sub001036_groupi_g4986__2883(csa_tree_sub001036_groupi_n_1023 ,csa_tree_sub001036_groupi_n_827 ,csa_tree_sub001036_groupi_n_951);
  nor csa_tree_sub001036_groupi_g4987__2346(csa_tree_sub001036_groupi_n_1022 ,csa_tree_sub001036_groupi_n_895 ,csa_tree_sub001036_groupi_n_980);
  nor csa_tree_sub001036_groupi_g4988__1666(csa_tree_sub001036_groupi_n_1021 ,csa_tree_sub001036_groupi_n_841 ,csa_tree_sub001036_groupi_n_916);
  nor csa_tree_sub001036_groupi_g4989__7410(csa_tree_sub001036_groupi_n_1020 ,csa_tree_sub001036_groupi_n_867 ,csa_tree_sub001036_groupi_n_967);
  or csa_tree_sub001036_groupi_g4990__6417(csa_tree_sub001036_groupi_n_1019 ,csa_tree_sub001036_groupi_n_897 ,csa_tree_sub001036_groupi_n_965);
  nor csa_tree_sub001036_groupi_g4991__5477(csa_tree_sub001036_groupi_n_1018 ,csa_tree_sub001036_groupi_n_923 ,csa_tree_sub001036_groupi_n_934);
  or csa_tree_sub001036_groupi_g4992__2398(csa_tree_sub001036_groupi_n_1017 ,csa_tree_sub001036_groupi_n_913 ,csa_tree_sub001036_groupi_n_925);
  nor csa_tree_sub001036_groupi_g4993__5107(csa_tree_sub001036_groupi_n_1016 ,csa_tree_sub001036_groupi_n_914 ,csa_tree_sub001036_groupi_n_926);
  nor csa_tree_sub001036_groupi_g4994__6260(csa_tree_sub001036_groupi_n_1015 ,csa_tree_sub001036_groupi_n_644 ,csa_tree_sub001036_groupi_n_928);
  or csa_tree_sub001036_groupi_g4995__4319(csa_tree_sub001036_groupi_n_1014 ,csa_tree_sub001036_groupi_n_845 ,csa_tree_sub001036_groupi_n_917);
  nor csa_tree_sub001036_groupi_g4996__8428(csa_tree_sub001036_groupi_n_1013 ,csa_tree_sub001036_groupi_n_846 ,csa_tree_sub001036_groupi_n_918);
  and csa_tree_sub001036_groupi_g4997__5526(csa_tree_sub001036_groupi_n_1012 ,csa_tree_sub001036_groupi_n_904 ,csa_tree_sub001036_groupi_n_960);
  nor csa_tree_sub001036_groupi_g4998__6783(csa_tree_sub001036_groupi_n_1011 ,csa_tree_sub001036_groupi_n_894 ,csa_tree_sub001036_groupi_n_970);
  and csa_tree_sub001036_groupi_g4999__3680(csa_tree_sub001036_groupi_n_1038 ,csa_tree_sub001036_groupi_n_869 ,csa_tree_sub001036_groupi_n_972);
  or csa_tree_sub001036_groupi_g5000__1617(csa_tree_sub001036_groupi_n_1037 ,csa_tree_sub001036_groupi_n_871 ,csa_tree_sub001036_groupi_n_962);
  or csa_tree_sub001036_groupi_g5001__2802(csa_tree_sub001036_groupi_n_1035 ,csa_tree_sub001036_groupi_n_875 ,csa_tree_sub001036_groupi_n_959);
  and csa_tree_sub001036_groupi_g5002__1705(csa_tree_sub001036_groupi_n_1034 ,csa_tree_sub001036_groupi_n_879 ,csa_tree_sub001036_groupi_n_956);
  or csa_tree_sub001036_groupi_g5003__5122(csa_tree_sub001036_groupi_n_1033 ,csa_tree_sub001036_groupi_n_833 ,csa_tree_sub001036_groupi_n_971);
  or csa_tree_sub001036_groupi_g5004__8246(csa_tree_sub001036_groupi_n_1007 ,csa_tree_sub001036_groupi_n_922 ,csa_tree_sub001036_groupi_n_935);
  nor csa_tree_sub001036_groupi_g5005__7098(csa_tree_sub001036_groupi_n_1006 ,csa_tree_sub001036_groupi_n_866 ,csa_tree_sub001036_groupi_n_955);
  or csa_tree_sub001036_groupi_g5006__6131(csa_tree_sub001036_groupi_n_1005 ,csa_tree_sub001036_groupi_n_981 ,csa_tree_sub001036_groupi_n_936);
  nor csa_tree_sub001036_groupi_g5007__1881(csa_tree_sub001036_groupi_n_1004 ,csa_tree_sub001036_groupi_n_982 ,csa_tree_sub001036_groupi_n_937);
  nor csa_tree_sub001036_groupi_g5008__5115(csa_tree_sub001036_groupi_n_1003 ,csa_tree_sub001036_groupi_n_844 ,csa_tree_sub001036_groupi_n_919);
  or csa_tree_sub001036_groupi_g5009__7482(csa_tree_sub001036_groupi_n_1002 ,csa_tree_sub001036_groupi_n_843 ,csa_tree_sub001036_groupi_n_920);
  nor csa_tree_sub001036_groupi_g5010__4733(csa_tree_sub001036_groupi_n_1001 ,csa_tree_sub001036_groupi_n_865 ,csa_tree_sub001036_groupi_n_958);
  or csa_tree_sub001036_groupi_g5011__6161(csa_tree_sub001036_groupi_n_1000 ,csa_tree_sub001036_groupi_n_645 ,csa_tree_sub001036_groupi_n_927);
  or csa_tree_sub001036_groupi_g5012__9315(csa_tree_sub001036_groupi_n_999 ,csa_tree_sub001036_groupi_n_842 ,csa_tree_sub001036_groupi_n_915);
  or csa_tree_sub001036_groupi_g5013__9945(csa_tree_sub001036_groupi_n_998 ,csa_tree_sub001036_groupi_n_940 ,csa_tree_sub001036_groupi_n_964);
  nor csa_tree_sub001036_groupi_g5014__2883(csa_tree_sub001036_groupi_n_997 ,csa_tree_sub001036_groupi_n_902 ,csa_tree_sub001036_groupi_n_979);
  or csa_tree_sub001036_groupi_g5015__2346(csa_tree_sub001036_groupi_n_996 ,csa_tree_sub001036_groupi_n_839 ,csa_tree_sub001036_groupi_n_933);
  xnor csa_tree_sub001036_groupi_g5016__1666(csa_tree_sub001036_groupi_n_995 ,csa_tree_sub001036_groupi_n_892 ,csa_tree_sub001036_groupi_n_852);
  xnor csa_tree_sub001036_groupi_g5017__7410(csa_tree_sub001036_groupi_n_994 ,csa_tree_sub001036_groupi_n_867 ,csa_tree_sub001036_groupi_n_758);
  xnor csa_tree_sub001036_groupi_g5018__6417(csa_tree_sub001036_groupi_n_993 ,csa_tree_sub001036_groupi_n_888 ,csa_tree_sub001036_groupi_n_890);
  xnor csa_tree_sub001036_groupi_g5019__5477(csa_tree_sub001036_groupi_n_992 ,csa_tree_sub001036_groupi_n_886 ,csa_tree_sub001036_groupi_n_857);
  xnor csa_tree_sub001036_groupi_g5020__2398(csa_tree_sub001036_groupi_n_991 ,csa_tree_sub001036_groupi_n_838 ,csa_tree_sub001036_groupi_n_848);
  xnor csa_tree_sub001036_groupi_g5021__5107(csa_tree_sub001036_groupi_n_990 ,csa_tree_sub001036_groupi_n_859 ,csa_tree_sub001036_groupi_n_885);
  xor csa_tree_sub001036_groupi_g5022__6260(csa_tree_sub001036_groupi_n_989 ,csa_tree_sub001036_groupi_n_853 ,csa_tree_sub001036_groupi_n_894);
  xor csa_tree_sub001036_groupi_g5023__4319(csa_tree_sub001036_groupi_n_988 ,csa_tree_sub001036_groupi_n_895 ,csa_tree_sub001036_groupi_n_856);
  xnor csa_tree_sub001036_groupi_g5024__8428(csa_tree_sub001036_groupi_n_987 ,csa_tree_sub001036_groupi_n_851 ,csa_tree_sub001036_groupi_n_901);
  xor csa_tree_sub001036_groupi_g5025__5526(csa_tree_sub001036_groupi_n_986 ,csa_tree_sub001036_groupi_n_903 ,csa_tree_sub001036_groupi_n_893);
  xnor csa_tree_sub001036_groupi_g5026__6783(csa_tree_sub001036_groupi_n_985 ,csa_tree_sub001036_groupi_n_840 ,csa_tree_sub001036_groupi_n_864);
  xnor csa_tree_sub001036_groupi_g5027__3680(csa_tree_sub001036_groupi_n_984 ,csa_tree_sub001036_groupi_n_825 ,csa_tree_sub001036_groupi_n_850);
  or csa_tree_sub001036_groupi_g5028__1617(csa_tree_sub001036_groupi_n_1010 ,csa_tree_sub001036_groupi_n_873 ,csa_tree_sub001036_groupi_n_953);
  xnor csa_tree_sub001036_groupi_g5029__2802(csa_tree_sub001036_groupi_n_1009 ,csa_tree_sub001036_groupi_n_868 ,csa_tree_sub001036_groupi_n_782);
  and csa_tree_sub001036_groupi_g5030__1705(csa_tree_sub001036_groupi_n_1008 ,csa_tree_sub001036_groupi_n_699 ,csa_tree_sub001036_groupi_n_954);
  not csa_tree_sub001036_groupi_g5031(csa_tree_sub001036_groupi_n_982 ,csa_tree_sub001036_groupi_n_981);
  nor csa_tree_sub001036_groupi_g5032__5122(csa_tree_sub001036_groupi_n_980 ,csa_tree_sub001036_groupi_n_856 ,csa_tree_sub001036_groupi_n_855);
  nor csa_tree_sub001036_groupi_g5033__8246(csa_tree_sub001036_groupi_n_979 ,csa_tree_sub001036_groupi_n_851 ,csa_tree_sub001036_groupi_n_860);
  and csa_tree_sub001036_groupi_g5034__7098(csa_tree_sub001036_groupi_n_978 ,csa_tree_sub001036_groupi_n_819 ,csa_tree_sub001036_groupi_n_881);
  and csa_tree_sub001036_groupi_g5035__6131(csa_tree_sub001036_groupi_n_977 ,csa_tree_sub001036_groupi_n_886 ,csa_tree_sub001036_groupi_n_857);
  or csa_tree_sub001036_groupi_g5036__1881(csa_tree_sub001036_groupi_n_976 ,csa_tree_sub001036_groupi_n_858 ,csa_tree_sub001036_groupi_n_884);
  and csa_tree_sub001036_groupi_g5037__5115(csa_tree_sub001036_groupi_n_975 ,csa_tree_sub001036_groupi_n_856 ,csa_tree_sub001036_groupi_n_855);
  nor csa_tree_sub001036_groupi_g5038__7482(csa_tree_sub001036_groupi_n_974 ,csa_tree_sub001036_groupi_n_859 ,csa_tree_sub001036_groupi_n_885);
  or csa_tree_sub001036_groupi_g5039__4733(csa_tree_sub001036_groupi_n_973 ,csa_tree_sub001036_groupi_n_886 ,csa_tree_sub001036_groupi_n_857);
  or csa_tree_sub001036_groupi_g5040__6161(csa_tree_sub001036_groupi_n_972 ,csa_tree_sub001036_groupi_n_826 ,csa_tree_sub001036_groupi_n_870);
  and csa_tree_sub001036_groupi_g5041__9315(csa_tree_sub001036_groupi_n_971 ,csa_tree_sub001036_groupi_n_792 ,csa_tree_sub001036_groupi_n_872);
  nor csa_tree_sub001036_groupi_g5042__9945(csa_tree_sub001036_groupi_n_970 ,csa_tree_sub001036_groupi_n_854 ,csa_tree_sub001036_groupi_n_853);
  and csa_tree_sub001036_groupi_g5043__2883(csa_tree_sub001036_groupi_n_969 ,csa_tree_sub001036_groupi_n_854 ,csa_tree_sub001036_groupi_n_853);
  nor csa_tree_sub001036_groupi_g5044__2346(csa_tree_sub001036_groupi_n_968 ,csa_tree_sub001036_groupi_n_758 ,csa_tree_sub001036_groupi_n_862);
  and csa_tree_sub001036_groupi_g5045__1666(csa_tree_sub001036_groupi_n_967 ,csa_tree_sub001036_groupi_n_758 ,csa_tree_sub001036_groupi_n_862);
  or csa_tree_sub001036_groupi_g5046__7410(csa_tree_sub001036_groupi_n_966 ,csa_tree_sub001036_groupi_n_888 ,csa_tree_sub001036_groupi_n_889);
  nor csa_tree_sub001036_groupi_g5047__6417(csa_tree_sub001036_groupi_n_965 ,csa_tree_sub001036_groupi_n_887 ,csa_tree_sub001036_groupi_n_890);
  nor csa_tree_sub001036_groupi_g5048__5477(csa_tree_sub001036_groupi_n_964 ,csa_tree_sub001036_groupi_n_838 ,csa_tree_sub001036_groupi_n_848);
  or csa_tree_sub001036_groupi_g5049__2398(csa_tree_sub001036_groupi_n_963 ,csa_tree_sub001036_groupi_n_837 ,csa_tree_sub001036_groupi_n_847);
  nor csa_tree_sub001036_groupi_g5050__5107(csa_tree_sub001036_groupi_n_962 ,csa_tree_sub001036_groupi_n_793 ,csa_tree_sub001036_groupi_n_878);
  and csa_tree_sub001036_groupi_g5051__6260(csa_tree_sub001036_groupi_n_961 ,csa_tree_sub001036_groupi_n_892 ,csa_tree_sub001036_groupi_n_852);
  or csa_tree_sub001036_groupi_g5052__4319(csa_tree_sub001036_groupi_n_960 ,csa_tree_sub001036_groupi_n_892 ,csa_tree_sub001036_groupi_n_852);
  nor csa_tree_sub001036_groupi_g5053__8428(csa_tree_sub001036_groupi_n_959 ,csa_tree_sub001036_groupi_n_830 ,csa_tree_sub001036_groupi_n_877);
  nor csa_tree_sub001036_groupi_g5054__5526(csa_tree_sub001036_groupi_n_958 ,csa_tree_sub001036_groupi_n_840 ,csa_tree_sub001036_groupi_n_849);
  and csa_tree_sub001036_groupi_g5055__6783(csa_tree_sub001036_groupi_n_957 ,csa_tree_sub001036_groupi_n_825 ,csa_tree_sub001036_groupi_n_850);
  or csa_tree_sub001036_groupi_g5056__3680(csa_tree_sub001036_groupi_n_956 ,csa_tree_sub001036_groupi_n_863 ,csa_tree_sub001036_groupi_n_836);
  nor csa_tree_sub001036_groupi_g5057__1617(csa_tree_sub001036_groupi_n_955 ,csa_tree_sub001036_groupi_n_825 ,csa_tree_sub001036_groupi_n_850);
  or csa_tree_sub001036_groupi_g5058__2802(csa_tree_sub001036_groupi_n_954 ,csa_tree_sub001036_groupi_n_693 ,csa_tree_sub001036_groupi_n_868);
  nor csa_tree_sub001036_groupi_g5059__1705(csa_tree_sub001036_groupi_n_953 ,csa_tree_sub001036_groupi_n_794 ,csa_tree_sub001036_groupi_n_834);
  and csa_tree_sub001036_groupi_g5060__5122(csa_tree_sub001036_groupi_n_952 ,csa_tree_sub001036_groupi_n_840 ,csa_tree_sub001036_groupi_n_849);
  nor csa_tree_sub001036_groupi_g5061__8246(csa_tree_sub001036_groupi_n_951 ,csa_tree_sub001036_groupi_n_819 ,csa_tree_sub001036_groupi_n_881);
  and csa_tree_sub001036_groupi_g5062__7098(csa_tree_sub001036_groupi_n_983 ,csa_tree_sub001036_groupi_n_734 ,csa_tree_sub001036_groupi_n_832);
  or csa_tree_sub001036_groupi_g5063__6131(csa_tree_sub001036_groupi_n_981 ,csa_tree_sub001036_groupi_n_704 ,csa_tree_sub001036_groupi_n_835);
  not csa_tree_sub001036_groupi_g5064(csa_tree_sub001036_groupi_n_950 ,csa_tree_sub001036_groupi_n_949);
  not csa_tree_sub001036_groupi_g5065(csa_tree_sub001036_groupi_n_945 ,csa_tree_sub001036_groupi_n_944);
  not csa_tree_sub001036_groupi_g5066(csa_tree_sub001036_groupi_n_939 ,csa_tree_sub001036_groupi_n_938);
  not csa_tree_sub001036_groupi_g5067(csa_tree_sub001036_groupi_n_937 ,csa_tree_sub001036_groupi_n_936);
  not csa_tree_sub001036_groupi_g5068(csa_tree_sub001036_groupi_n_934 ,csa_tree_sub001036_groupi_n_935);
  not csa_tree_sub001036_groupi_g5069(csa_tree_sub001036_groupi_n_931 ,csa_tree_sub001036_groupi_n_932);
  not csa_tree_sub001036_groupi_g5070(csa_tree_sub001036_groupi_n_929 ,csa_tree_sub001036_groupi_n_930);
  not csa_tree_sub001036_groupi_g5071(csa_tree_sub001036_groupi_n_927 ,csa_tree_sub001036_groupi_n_928);
  not csa_tree_sub001036_groupi_g5072(csa_tree_sub001036_groupi_n_925 ,csa_tree_sub001036_groupi_n_926);
  not csa_tree_sub001036_groupi_g5073(csa_tree_sub001036_groupi_n_922 ,csa_tree_sub001036_groupi_n_923);
  not csa_tree_sub001036_groupi_g5074(csa_tree_sub001036_groupi_n_919 ,csa_tree_sub001036_groupi_n_920);
  not csa_tree_sub001036_groupi_g5075(csa_tree_sub001036_groupi_n_917 ,csa_tree_sub001036_groupi_n_918);
  not csa_tree_sub001036_groupi_g5076(csa_tree_sub001036_groupi_n_915 ,csa_tree_sub001036_groupi_n_916);
  not csa_tree_sub001036_groupi_g5077(csa_tree_sub001036_groupi_n_913 ,csa_tree_sub001036_groupi_n_914);
  and csa_tree_sub001036_groupi_g5078__1881(csa_tree_sub001036_groupi_n_912 ,csa_tree_sub001036_groupi_n_851 ,csa_tree_sub001036_groupi_n_860);
  xor csa_tree_sub001036_groupi_g5079__5115(csa_tree_sub001036_groupi_n_911 ,csa_tree_sub001036_groupi_n_793 ,csa_tree_sub001036_groupi_n_820);
  xnor csa_tree_sub001036_groupi_g5080__7482(csa_tree_sub001036_groupi_n_910 ,csa_tree_sub001036_groupi_n_816 ,csa_tree_sub001036_groupi_n_824);
  xor csa_tree_sub001036_groupi_g5081__4733(csa_tree_sub001036_groupi_n_909 ,csa_tree_sub001036_groupi_n_585 ,csa_tree_sub001036_groupi_n_830);
  xor csa_tree_sub001036_groupi_g5082__6161(csa_tree_sub001036_groupi_n_908 ,csa_tree_sub001036_groupi_n_647 ,csa_tree_sub001036_groupi_n_826);
  xnor csa_tree_sub001036_groupi_g5083__9315(csa_tree_sub001036_groupi_n_907 ,csa_tree_sub001036_groupi_n_711 ,csa_tree_sub001036_groupi_n_792);
  xor csa_tree_sub001036_groupi_g5084__9945(csa_tree_sub001036_groupi_n_906 ,csa_tree_sub001036_groupi_n_827 ,csa_tree_sub001036_groupi_n_819);
  xor csa_tree_sub001036_groupi_g5086__2883(csa_tree_sub001036_groupi_n_905 ,csa_tree_sub001036_groupi_n_794 ,csa_tree_sub001036_groupi_n_790);
  xnor csa_tree_sub001036_groupi_g5087__2346(csa_tree_sub001036_groupi_n_949 ,csa_tree_sub001036_groupi_n_656 ,csa_tree_sub001036_groupi_n_776);
  xnor csa_tree_sub001036_groupi_g5088__1666(csa_tree_sub001036_groupi_n_948 ,csa_tree_sub001036_groupi_n_588 ,csa_tree_sub001036_groupi_n_761);
  xnor csa_tree_sub001036_groupi_g5089__7410(csa_tree_sub001036_groupi_n_947 ,csa_tree_sub001036_groupi_n_828 ,csa_tree_sub001036_groupi_n_763);
  xnor csa_tree_sub001036_groupi_g5090__6417(csa_tree_sub001036_groupi_n_946 ,csa_tree_sub001036_groupi_n_498 ,csa_tree_sub001036_groupi_n_769);
  xnor csa_tree_sub001036_groupi_g5091__5477(csa_tree_sub001036_groupi_n_944 ,csa_tree_sub001036_groupi_n_469 ,csa_tree_sub001036_groupi_n_768);
  xnor csa_tree_sub001036_groupi_g5092__2398(csa_tree_sub001036_groupi_n_943 ,csa_tree_sub001036_groupi_n_594 ,csa_tree_sub001036_groupi_n_764);
  xnor csa_tree_sub001036_groupi_g5093__5107(csa_tree_sub001036_groupi_n_942 ,csa_tree_sub001036_groupi_n_829 ,csa_tree_sub001036_groupi_n_771);
  xnor csa_tree_sub001036_groupi_g5094__6260(csa_tree_sub001036_groupi_n_941 ,csa_tree_sub001036_groupi_n_591 ,csa_tree_sub001036_groupi_n_775);
  xnor csa_tree_sub001036_groupi_g5095__4319(csa_tree_sub001036_groupi_n_940 ,csa_tree_sub001036_groupi_n_590 ,csa_tree_sub001036_groupi_n_777);
  xnor csa_tree_sub001036_groupi_g5096__8428(csa_tree_sub001036_groupi_n_938 ,csa_tree_sub001036_groupi_n_540 ,csa_tree_sub001036_groupi_n_774);
  xnor csa_tree_sub001036_groupi_g5097__5526(csa_tree_sub001036_groupi_n_936 ,csa_tree_sub001036_groupi_n_554 ,csa_tree_sub001036_groupi_n_778);
  xnor csa_tree_sub001036_groupi_g5098__6783(csa_tree_sub001036_groupi_n_935 ,csa_tree_sub001036_groupi_n_466 ,csa_tree_sub001036_groupi_n_766);
  xnor csa_tree_sub001036_groupi_g5099__3680(csa_tree_sub001036_groupi_n_933 ,csa_tree_sub001036_groupi_n_595 ,csa_tree_sub001036_groupi_n_784);
  xnor csa_tree_sub001036_groupi_g5100__1617(csa_tree_sub001036_groupi_n_932 ,csa_tree_sub001036_groupi_n_592 ,csa_tree_sub001036_groupi_n_765);
  xnor csa_tree_sub001036_groupi_g5101__2802(csa_tree_sub001036_groupi_n_930 ,csa_tree_sub001036_groupi_n_608 ,csa_tree_sub001036_groupi_n_783);
  xnor csa_tree_sub001036_groupi_g5102__1705(csa_tree_sub001036_groupi_n_928 ,csa_tree_sub001036_groupi_n_791 ,csa_tree_sub001036_groupi_n_779);
  xnor csa_tree_sub001036_groupi_g5103__5122(csa_tree_sub001036_groupi_n_926 ,csa_tree_sub001036_groupi_n_659 ,csa_tree_sub001036_groupi_n_762);
  xnor csa_tree_sub001036_groupi_g5104__8246(csa_tree_sub001036_groupi_n_924 ,csa_tree_sub001036_groupi_n_576 ,csa_tree_sub001036_groupi_n_773);
  xnor csa_tree_sub001036_groupi_g5105__7098(csa_tree_sub001036_groupi_n_923 ,csa_tree_sub001036_groupi_n_562 ,csa_tree_sub001036_groupi_n_781);
  xnor csa_tree_sub001036_groupi_g5106__6131(csa_tree_sub001036_groupi_n_921 ,csa_tree_sub001036_groupi_n_713 ,csa_tree_sub001036_groupi_n_780);
  xnor csa_tree_sub001036_groupi_g5107__1881(csa_tree_sub001036_groupi_n_920 ,csa_tree_sub001036_groupi_n_600 ,csa_tree_sub001036_groupi_n_770);
  xnor csa_tree_sub001036_groupi_g5108__5115(csa_tree_sub001036_groupi_n_918 ,csa_tree_sub001036_groupi_n_657 ,csa_tree_sub001036_groupi_n_767);
  or csa_tree_sub001036_groupi_g5109__7482(csa_tree_sub001036_groupi_n_916 ,csa_tree_sub001036_groupi_n_705 ,csa_tree_sub001036_groupi_n_876);
  xnor csa_tree_sub001036_groupi_g5110__4733(csa_tree_sub001036_groupi_n_914 ,csa_tree_sub001036_groupi_n_460 ,csa_tree_sub001036_groupi_n_772);
  not csa_tree_sub001036_groupi_g5111(csa_tree_sub001036_groupi_n_902 ,csa_tree_sub001036_groupi_n_901);
  not csa_tree_sub001036_groupi_g5112(csa_tree_sub001036_groupi_n_899 ,csa_tree_sub001036_groupi_n_898);
  not csa_tree_sub001036_groupi_g5113(csa_tree_sub001036_groupi_n_897 ,csa_tree_sub001036_groupi_n_896);
  not csa_tree_sub001036_groupi_g5114(csa_tree_sub001036_groupi_n_889 ,csa_tree_sub001036_groupi_n_890);
  not csa_tree_sub001036_groupi_g5115(csa_tree_sub001036_groupi_n_888 ,csa_tree_sub001036_groupi_n_887);
  not csa_tree_sub001036_groupi_g5116(csa_tree_sub001036_groupi_n_884 ,csa_tree_sub001036_groupi_n_885);
  not csa_tree_sub001036_groupi_g5117(csa_tree_sub001036_groupi_n_882 ,csa_tree_sub001036_groupi_n_883);
  or csa_tree_sub001036_groupi_g5118__6161(csa_tree_sub001036_groupi_n_879 ,csa_tree_sub001036_groupi_n_815 ,csa_tree_sub001036_groupi_n_823);
  nor csa_tree_sub001036_groupi_g5119__9315(csa_tree_sub001036_groupi_n_878 ,csa_tree_sub001036_groupi_n_759 ,csa_tree_sub001036_groupi_n_820);
  nor csa_tree_sub001036_groupi_g5120__9945(csa_tree_sub001036_groupi_n_877 ,csa_tree_sub001036_groupi_n_585 ,csa_tree_sub001036_groupi_n_818);
  and csa_tree_sub001036_groupi_g5121__2883(csa_tree_sub001036_groupi_n_876 ,csa_tree_sub001036_groupi_n_829 ,csa_tree_sub001036_groupi_n_724);
  and csa_tree_sub001036_groupi_g5122__2346(csa_tree_sub001036_groupi_n_875 ,csa_tree_sub001036_groupi_n_585 ,csa_tree_sub001036_groupi_n_818);
  or csa_tree_sub001036_groupi_g5123__1666(csa_tree_sub001036_groupi_n_874 ,csa_tree_sub001036_groupi_n_90 ,csa_tree_sub001036_groupi_n_817);
  and csa_tree_sub001036_groupi_g5124__7410(csa_tree_sub001036_groupi_n_873 ,csa_tree_sub001036_groupi_n_760 ,csa_tree_sub001036_groupi_n_790);
  or csa_tree_sub001036_groupi_g5125__6417(csa_tree_sub001036_groupi_n_872 ,csa_tree_sub001036_groupi_n_712 ,csa_tree_sub001036_groupi_n_789);
  and csa_tree_sub001036_groupi_g5126__5477(csa_tree_sub001036_groupi_n_871 ,csa_tree_sub001036_groupi_n_759 ,csa_tree_sub001036_groupi_n_820);
  nor csa_tree_sub001036_groupi_g5127__2398(csa_tree_sub001036_groupi_n_870 ,csa_tree_sub001036_groupi_n_647 ,csa_tree_sub001036_groupi_n_822);
  or csa_tree_sub001036_groupi_g5128__5107(csa_tree_sub001036_groupi_n_869 ,csa_tree_sub001036_groupi_n_646 ,csa_tree_sub001036_groupi_n_821);
  or csa_tree_sub001036_groupi_g5129__6260(csa_tree_sub001036_groupi_n_904 ,csa_tree_sub001036_groupi_n_716 ,csa_tree_sub001036_groupi_n_805);
  and csa_tree_sub001036_groupi_g5130__4319(csa_tree_sub001036_groupi_n_903 ,csa_tree_sub001036_groupi_n_729 ,csa_tree_sub001036_groupi_n_814);
  or csa_tree_sub001036_groupi_g5131__8428(csa_tree_sub001036_groupi_n_901 ,csa_tree_sub001036_groupi_n_755 ,csa_tree_sub001036_groupi_n_798);
  and csa_tree_sub001036_groupi_g5132__5526(csa_tree_sub001036_groupi_n_900 ,csa_tree_sub001036_groupi_n_753 ,csa_tree_sub001036_groupi_n_811);
  or csa_tree_sub001036_groupi_g5133__6783(csa_tree_sub001036_groupi_n_898 ,csa_tree_sub001036_groupi_n_757 ,csa_tree_sub001036_groupi_n_802);
  or csa_tree_sub001036_groupi_g5134__3680(csa_tree_sub001036_groupi_n_896 ,csa_tree_sub001036_groupi_n_750 ,csa_tree_sub001036_groupi_n_810);
  and csa_tree_sub001036_groupi_g5135__1617(csa_tree_sub001036_groupi_n_895 ,csa_tree_sub001036_groupi_n_719 ,csa_tree_sub001036_groupi_n_796);
  and csa_tree_sub001036_groupi_g5136__2802(csa_tree_sub001036_groupi_n_894 ,csa_tree_sub001036_groupi_n_727 ,csa_tree_sub001036_groupi_n_801);
  or csa_tree_sub001036_groupi_g5137__1705(csa_tree_sub001036_groupi_n_893 ,csa_tree_sub001036_groupi_n_731 ,csa_tree_sub001036_groupi_n_800);
  or csa_tree_sub001036_groupi_g5138__5122(csa_tree_sub001036_groupi_n_892 ,csa_tree_sub001036_groupi_n_715 ,csa_tree_sub001036_groupi_n_807);
  or csa_tree_sub001036_groupi_g5139__8246(csa_tree_sub001036_groupi_n_891 ,csa_tree_sub001036_groupi_n_743 ,csa_tree_sub001036_groupi_n_806);
  or csa_tree_sub001036_groupi_g5140__7098(csa_tree_sub001036_groupi_n_890 ,csa_tree_sub001036_groupi_n_746 ,csa_tree_sub001036_groupi_n_808);
  or csa_tree_sub001036_groupi_g5141__6131(csa_tree_sub001036_groupi_n_887 ,csa_tree_sub001036_groupi_n_748 ,csa_tree_sub001036_groupi_n_809);
  or csa_tree_sub001036_groupi_g5142__1881(csa_tree_sub001036_groupi_n_886 ,csa_tree_sub001036_groupi_n_742 ,csa_tree_sub001036_groupi_n_803);
  or csa_tree_sub001036_groupi_g5143__5115(csa_tree_sub001036_groupi_n_885 ,csa_tree_sub001036_groupi_n_737 ,csa_tree_sub001036_groupi_n_804);
  or csa_tree_sub001036_groupi_g5144__7482(csa_tree_sub001036_groupi_n_883 ,csa_tree_sub001036_groupi_n_708 ,csa_tree_sub001036_groupi_n_812);
  or csa_tree_sub001036_groupi_g5145__4733(csa_tree_sub001036_groupi_n_881 ,csa_tree_sub001036_groupi_n_756 ,csa_tree_sub001036_groupi_n_799);
  or csa_tree_sub001036_groupi_g5146__6161(csa_tree_sub001036_groupi_n_880 ,csa_tree_sub001036_groupi_n_721 ,csa_tree_sub001036_groupi_n_795);
  not csa_tree_sub001036_groupi_g5147(csa_tree_sub001036_groupi_n_865 ,csa_tree_sub001036_groupi_n_864);
  not csa_tree_sub001036_groupi_g5149(csa_tree_sub001036_groupi_n_862 ,csa_tree_sub001036_groupi_n_861);
  not csa_tree_sub001036_groupi_g5150(csa_tree_sub001036_groupi_n_858 ,csa_tree_sub001036_groupi_n_859);
  not csa_tree_sub001036_groupi_g5151(csa_tree_sub001036_groupi_n_847 ,csa_tree_sub001036_groupi_n_848);
  not csa_tree_sub001036_groupi_g5152(csa_tree_sub001036_groupi_n_846 ,csa_tree_sub001036_groupi_n_845);
  not csa_tree_sub001036_groupi_g5153(csa_tree_sub001036_groupi_n_844 ,csa_tree_sub001036_groupi_n_843);
  not csa_tree_sub001036_groupi_g5154(csa_tree_sub001036_groupi_n_842 ,csa_tree_sub001036_groupi_n_841);
  not csa_tree_sub001036_groupi_g5155(csa_tree_sub001036_groupi_n_837 ,csa_tree_sub001036_groupi_n_838);
  nor csa_tree_sub001036_groupi_g5156__9315(csa_tree_sub001036_groupi_n_836 ,csa_tree_sub001036_groupi_n_816 ,csa_tree_sub001036_groupi_n_824);
  and csa_tree_sub001036_groupi_g5157__9945(csa_tree_sub001036_groupi_n_835 ,csa_tree_sub001036_groupi_n_720 ,csa_tree_sub001036_groupi_n_828);
  nor csa_tree_sub001036_groupi_g5158__2883(csa_tree_sub001036_groupi_n_834 ,csa_tree_sub001036_groupi_n_760 ,csa_tree_sub001036_groupi_n_790);
  and csa_tree_sub001036_groupi_g5159__2346(csa_tree_sub001036_groupi_n_833 ,csa_tree_sub001036_groupi_n_712 ,csa_tree_sub001036_groupi_n_789);
  or csa_tree_sub001036_groupi_g5160__1666(csa_tree_sub001036_groupi_n_832 ,csa_tree_sub001036_groupi_n_689 ,csa_tree_sub001036_groupi_n_791);
  and csa_tree_sub001036_groupi_g5161__7410(csa_tree_sub001036_groupi_n_831 ,csa_tree_sub001036_groupi_n_90 ,csa_tree_sub001036_groupi_n_817);
  xnor csa_tree_sub001036_groupi_g5162__6417(csa_tree_sub001036_groupi_n_868 ,csa_tree_sub001036_groupi_n_515 ,csa_tree_sub001036_groupi_n_682);
  xnor csa_tree_sub001036_groupi_g5163__5477(csa_tree_sub001036_groupi_n_867 ,csa_tree_sub001036_groupi_n_535 ,csa_tree_sub001036_groupi_n_677);
  and csa_tree_sub001036_groupi_g5164__2398(csa_tree_sub001036_groupi_n_866 ,csa_tree_sub001036_groupi_n_701 ,csa_tree_sub001036_groupi_n_813);
  or csa_tree_sub001036_groupi_g5165__5107(csa_tree_sub001036_groupi_n_864 ,csa_tree_sub001036_groupi_n_688 ,csa_tree_sub001036_groupi_n_787);
  and csa_tree_sub001036_groupi_g5166__6260(csa_tree_sub001036_groupi_n_863 ,csa_tree_sub001036_groupi_n_698 ,csa_tree_sub001036_groupi_n_797);
  xnor csa_tree_sub001036_groupi_g5167__4319(csa_tree_sub001036_groupi_n_861 ,csa_tree_sub001036_groupi_n_491 ,csa_tree_sub001036_groupi_n_678);
  xnor csa_tree_sub001036_groupi_g5168__8428(csa_tree_sub001036_groupi_n_860 ,csa_tree_sub001036_groupi_n_484 ,csa_tree_sub001036_groupi_n_679);
  xnor csa_tree_sub001036_groupi_g5169__5526(csa_tree_sub001036_groupi_n_859 ,csa_tree_sub001036_groupi_n_529 ,csa_tree_sub001036_groupi_n_676);
  xnor csa_tree_sub001036_groupi_g5170__6783(csa_tree_sub001036_groupi_n_857 ,csa_tree_sub001036_groupi_n_650 ,csa_tree_sub001036_groupi_n_674);
  xnor csa_tree_sub001036_groupi_g5171__3680(csa_tree_sub001036_groupi_n_856 ,csa_tree_sub001036_groupi_n_536 ,csa_tree_sub001036_groupi_n_675);
  xnor csa_tree_sub001036_groupi_g5172__1617(csa_tree_sub001036_groupi_n_855 ,csa_tree_sub001036_groupi_n_516 ,csa_tree_sub001036_groupi_n_673);
  xnor csa_tree_sub001036_groupi_g5173__2802(csa_tree_sub001036_groupi_n_854 ,csa_tree_sub001036_groupi_n_527 ,csa_tree_sub001036_groupi_n_672);
  xnor csa_tree_sub001036_groupi_g5174__1705(csa_tree_sub001036_groupi_n_853 ,csa_tree_sub001036_groupi_n_485 ,csa_tree_sub001036_groupi_n_671);
  xnor csa_tree_sub001036_groupi_g5175__5122(csa_tree_sub001036_groupi_n_852 ,csa_tree_sub001036_groupi_n_597 ,csa_tree_sub001036_groupi_n_670);
  xnor csa_tree_sub001036_groupi_g5176__8246(csa_tree_sub001036_groupi_n_851 ,csa_tree_sub001036_groupi_n_545 ,csa_tree_sub001036_groupi_n_666);
  xnor csa_tree_sub001036_groupi_g5177__7098(csa_tree_sub001036_groupi_n_850 ,csa_tree_sub001036_groupi_n_567 ,csa_tree_sub001036_groupi_n_669);
  xnor csa_tree_sub001036_groupi_g5178__6131(csa_tree_sub001036_groupi_n_849 ,csa_tree_sub001036_groupi_n_490 ,csa_tree_sub001036_groupi_n_668);
  xnor csa_tree_sub001036_groupi_g5179__1881(csa_tree_sub001036_groupi_n_848 ,csa_tree_sub001036_groupi_n_471 ,csa_tree_sub001036_groupi_n_667);
  xnor csa_tree_sub001036_groupi_g5180__5115(csa_tree_sub001036_groupi_n_845 ,csa_tree_sub001036_groupi_n_561 ,csa_tree_sub001036_groupi_n_681);
  xnor csa_tree_sub001036_groupi_g5181__7482(csa_tree_sub001036_groupi_n_843 ,csa_tree_sub001036_groupi_n_663 ,csa_tree_sub001036_groupi_n_680);
  xnor csa_tree_sub001036_groupi_g5182__4733(csa_tree_sub001036_groupi_n_841 ,csa_tree_sub001036_groupi_n_665 ,csa_tree_sub001036_groupi_n_504);
  or csa_tree_sub001036_groupi_g5183__6161(csa_tree_sub001036_groupi_n_840 ,csa_tree_sub001036_groupi_n_695 ,csa_tree_sub001036_groupi_n_785);
  xnor csa_tree_sub001036_groupi_g5184__9315(csa_tree_sub001036_groupi_n_839 ,csa_tree_sub001036_groupi_n_480 ,csa_tree_sub001036_groupi_n_683);
  or csa_tree_sub001036_groupi_g5185__9945(csa_tree_sub001036_groupi_n_838 ,csa_tree_sub001036_groupi_n_697 ,csa_tree_sub001036_groupi_n_786);
  not csa_tree_sub001036_groupi_g5186(csa_tree_sub001036_groupi_n_823 ,csa_tree_sub001036_groupi_n_824);
  not csa_tree_sub001036_groupi_g5187(csa_tree_sub001036_groupi_n_821 ,csa_tree_sub001036_groupi_n_822);
  not csa_tree_sub001036_groupi_g5188(csa_tree_sub001036_groupi_n_815 ,csa_tree_sub001036_groupi_n_816);
  or csa_tree_sub001036_groupi_g5189__2883(csa_tree_sub001036_groupi_n_814 ,csa_tree_sub001036_groupi_n_664 ,csa_tree_sub001036_groupi_n_728);
  or csa_tree_sub001036_groupi_g5190__2346(csa_tree_sub001036_groupi_n_813 ,csa_tree_sub001036_groupi_n_591 ,csa_tree_sub001036_groupi_n_744);
  nor csa_tree_sub001036_groupi_g5191__1666(csa_tree_sub001036_groupi_n_812 ,csa_tree_sub001036_groupi_n_602 ,csa_tree_sub001036_groupi_n_718);
  or csa_tree_sub001036_groupi_g5192__7410(csa_tree_sub001036_groupi_n_811 ,csa_tree_sub001036_groupi_n_594 ,csa_tree_sub001036_groupi_n_751);
  nor csa_tree_sub001036_groupi_g5193__6417(csa_tree_sub001036_groupi_n_810 ,csa_tree_sub001036_groupi_n_605 ,csa_tree_sub001036_groupi_n_749);
  nor csa_tree_sub001036_groupi_g5194__5477(csa_tree_sub001036_groupi_n_809 ,csa_tree_sub001036_groupi_n_593 ,csa_tree_sub001036_groupi_n_747);
  nor csa_tree_sub001036_groupi_g5195__2398(csa_tree_sub001036_groupi_n_808 ,csa_tree_sub001036_groupi_n_603 ,csa_tree_sub001036_groupi_n_745);
  nor csa_tree_sub001036_groupi_g5196__5107(csa_tree_sub001036_groupi_n_807 ,csa_tree_sub001036_groupi_n_604 ,csa_tree_sub001036_groupi_n_710);
  nor csa_tree_sub001036_groupi_g5197__6260(csa_tree_sub001036_groupi_n_806 ,csa_tree_sub001036_groupi_n_713 ,csa_tree_sub001036_groupi_n_735);
  nor csa_tree_sub001036_groupi_g5198__4319(csa_tree_sub001036_groupi_n_805 ,csa_tree_sub001036_groupi_n_607 ,csa_tree_sub001036_groupi_n_707);
  nor csa_tree_sub001036_groupi_g5199__8428(csa_tree_sub001036_groupi_n_804 ,csa_tree_sub001036_groupi_n_606 ,csa_tree_sub001036_groupi_n_736);
  nor csa_tree_sub001036_groupi_g5200__5526(csa_tree_sub001036_groupi_n_803 ,csa_tree_sub001036_groupi_n_498 ,csa_tree_sub001036_groupi_n_726);
  nor csa_tree_sub001036_groupi_g5201__6783(csa_tree_sub001036_groupi_n_802 ,csa_tree_sub001036_groupi_n_540 ,csa_tree_sub001036_groupi_n_733);
  or csa_tree_sub001036_groupi_g5202__3680(csa_tree_sub001036_groupi_n_801 ,csa_tree_sub001036_groupi_n_601 ,csa_tree_sub001036_groupi_n_739);
  and csa_tree_sub001036_groupi_g5203__1617(csa_tree_sub001036_groupi_n_800 ,csa_tree_sub001036_groupi_n_592 ,csa_tree_sub001036_groupi_n_730);
  nor csa_tree_sub001036_groupi_g5204__2802(csa_tree_sub001036_groupi_n_799 ,csa_tree_sub001036_groupi_n_533 ,csa_tree_sub001036_groupi_n_725);
  nor csa_tree_sub001036_groupi_g5205__1705(csa_tree_sub001036_groupi_n_798 ,csa_tree_sub001036_groupi_n_662 ,csa_tree_sub001036_groupi_n_752);
  or csa_tree_sub001036_groupi_g5206__5122(csa_tree_sub001036_groupi_n_797 ,csa_tree_sub001036_groupi_n_489 ,csa_tree_sub001036_groupi_n_687);
  or csa_tree_sub001036_groupi_g5207__8246(csa_tree_sub001036_groupi_n_796 ,csa_tree_sub001036_groupi_n_596 ,csa_tree_sub001036_groupi_n_691);
  and csa_tree_sub001036_groupi_g5208__7098(csa_tree_sub001036_groupi_n_795 ,csa_tree_sub001036_groupi_n_598 ,csa_tree_sub001036_groupi_n_692);
  and csa_tree_sub001036_groupi_g5209__6131(csa_tree_sub001036_groupi_n_830 ,csa_tree_sub001036_groupi_n_615 ,csa_tree_sub001036_groupi_n_722);
  or csa_tree_sub001036_groupi_g5210__1881(csa_tree_sub001036_groupi_n_829 ,csa_tree_sub001036_groupi_n_641 ,csa_tree_sub001036_groupi_n_740);
  or csa_tree_sub001036_groupi_g5211__5115(csa_tree_sub001036_groupi_n_828 ,csa_tree_sub001036_groupi_n_621 ,csa_tree_sub001036_groupi_n_706);
  and csa_tree_sub001036_groupi_g5212__7482(csa_tree_sub001036_groupi_n_827 ,csa_tree_sub001036_groupi_n_629 ,csa_tree_sub001036_groupi_n_754);
  and csa_tree_sub001036_groupi_g5213__4733(csa_tree_sub001036_groupi_n_826 ,csa_tree_sub001036_groupi_n_638 ,csa_tree_sub001036_groupi_n_738);
  or csa_tree_sub001036_groupi_g5214__6161(csa_tree_sub001036_groupi_n_825 ,csa_tree_sub001036_groupi_n_502 ,csa_tree_sub001036_groupi_n_702);
  or csa_tree_sub001036_groupi_g5215__9315(csa_tree_sub001036_groupi_n_824 ,csa_tree_sub001036_groupi_n_628 ,csa_tree_sub001036_groupi_n_732);
  or csa_tree_sub001036_groupi_g5216__9945(csa_tree_sub001036_groupi_n_822 ,csa_tree_sub001036_groupi_n_640 ,csa_tree_sub001036_groupi_n_741);
  or csa_tree_sub001036_groupi_g5217__2883(csa_tree_sub001036_groupi_n_820 ,csa_tree_sub001036_groupi_n_631 ,csa_tree_sub001036_groupi_n_714);
  or csa_tree_sub001036_groupi_g5218__2346(csa_tree_sub001036_groupi_n_819 ,csa_tree_sub001036_groupi_n_636 ,csa_tree_sub001036_groupi_n_700);
  or csa_tree_sub001036_groupi_g5219__1666(csa_tree_sub001036_groupi_n_818 ,csa_tree_sub001036_groupi_n_633 ,csa_tree_sub001036_groupi_n_723);
  or csa_tree_sub001036_groupi_g5220__7410(csa_tree_sub001036_groupi_n_817 ,csa_tree_sub001036_groupi_n_642 ,csa_tree_sub001036_groupi_n_709);
  or csa_tree_sub001036_groupi_g5221__6417(csa_tree_sub001036_groupi_n_816 ,csa_tree_sub001036_groupi_n_616 ,csa_tree_sub001036_groupi_n_717);
  xor csa_tree_sub001036_groupi_g5222__5477(out1[0] ,csa_tree_sub001036_groupi_n_548 ,csa_tree_sub001036_groupi_n_138);
  and csa_tree_sub001036_groupi_g5223__2398(csa_tree_sub001036_groupi_n_787 ,csa_tree_sub001036_groupi_n_600 ,csa_tree_sub001036_groupi_n_686);
  and csa_tree_sub001036_groupi_g5224__5107(csa_tree_sub001036_groupi_n_786 ,csa_tree_sub001036_groupi_n_608 ,csa_tree_sub001036_groupi_n_694);
  nor csa_tree_sub001036_groupi_g5225__6260(csa_tree_sub001036_groupi_n_785 ,csa_tree_sub001036_groupi_n_496 ,csa_tree_sub001036_groupi_n_690);
  xnor csa_tree_sub001036_groupi_g5226__4319(csa_tree_sub001036_groupi_n_784 ,csa_tree_sub001036_groupi_n_468 ,csa_tree_sub001036_groupi_n_577);
  xnor csa_tree_sub001036_groupi_g5227__8428(csa_tree_sub001036_groupi_n_783 ,csa_tree_sub001036_groupi_n_526 ,csa_tree_sub001036_groupi_n_557);
  xnor csa_tree_sub001036_groupi_g5228__5526(csa_tree_sub001036_groupi_n_782 ,csa_tree_sub001036_groupi_n_555 ,csa_tree_sub001036_groupi_n_551);
  xnor csa_tree_sub001036_groupi_g5229__6783(csa_tree_sub001036_groupi_n_781 ,csa_tree_sub001036_groupi_n_457 ,csa_tree_sub001036_groupi_n_593);
  xnor csa_tree_sub001036_groupi_g5230__3680(csa_tree_sub001036_groupi_n_780 ,csa_tree_sub001036_groupi_n_563 ,csa_tree_sub001036_groupi_n_648);
  xnor csa_tree_sub001036_groupi_g5231__1617(csa_tree_sub001036_groupi_n_779 ,csa_tree_sub001036_groupi_n_552 ,csa_tree_sub001036_groupi_n_579);
  xnor csa_tree_sub001036_groupi_g5232__2802(csa_tree_sub001036_groupi_n_778 ,csa_tree_sub001036_groupi_n_465 ,csa_tree_sub001036_groupi_n_598);
  xnor csa_tree_sub001036_groupi_g5233__1705(csa_tree_sub001036_groupi_n_777 ,csa_tree_sub001036_groupi_n_519 ,csa_tree_sub001036_groupi_n_605);
  xor csa_tree_sub001036_groupi_g5234__5122(csa_tree_sub001036_groupi_n_776 ,csa_tree_sub001036_groupi_n_664 ,csa_tree_sub001036_groupi_n_582);
  xnor csa_tree_sub001036_groupi_g5235__8246(csa_tree_sub001036_groupi_n_775 ,csa_tree_sub001036_groupi_n_569 ,csa_tree_sub001036_groupi_n_574);
  xnor csa_tree_sub001036_groupi_g5236__7098(csa_tree_sub001036_groupi_n_774 ,csa_tree_sub001036_groupi_n_653 ,csa_tree_sub001036_groupi_n_660);
  xor csa_tree_sub001036_groupi_g5237__6131(csa_tree_sub001036_groupi_n_773 ,csa_tree_sub001036_groupi_n_606 ,csa_tree_sub001036_groupi_n_572);
  xor csa_tree_sub001036_groupi_g5238__1881(csa_tree_sub001036_groupi_n_772 ,csa_tree_sub001036_groupi_n_604 ,csa_tree_sub001036_groupi_n_586);
  xnor csa_tree_sub001036_groupi_g5239__5115(csa_tree_sub001036_groupi_n_771 ,csa_tree_sub001036_groupi_n_570 ,csa_tree_sub001036_groupi_n_661);
  xnor csa_tree_sub001036_groupi_g5240__7482(csa_tree_sub001036_groupi_n_770 ,csa_tree_sub001036_groupi_n_456 ,csa_tree_sub001036_groupi_n_583);
  xnor csa_tree_sub001036_groupi_g5241__4733(csa_tree_sub001036_groupi_n_769 ,csa_tree_sub001036_groupi_n_550 ,csa_tree_sub001036_groupi_n_571);
  xor csa_tree_sub001036_groupi_g5242__6161(csa_tree_sub001036_groupi_n_768 ,csa_tree_sub001036_groupi_n_607 ,csa_tree_sub001036_groupi_n_564);
  xor csa_tree_sub001036_groupi_g5243__9315(csa_tree_sub001036_groupi_n_767 ,csa_tree_sub001036_groupi_n_662 ,csa_tree_sub001036_groupi_n_654);
  xor csa_tree_sub001036_groupi_g5244__9945(csa_tree_sub001036_groupi_n_766 ,csa_tree_sub001036_groupi_n_603 ,csa_tree_sub001036_groupi_n_584);
  xnor csa_tree_sub001036_groupi_g5245__2883(csa_tree_sub001036_groupi_n_765 ,csa_tree_sub001036_groupi_n_520 ,csa_tree_sub001036_groupi_n_575);
  xnor csa_tree_sub001036_groupi_g5246__2346(csa_tree_sub001036_groupi_n_764 ,csa_tree_sub001036_groupi_n_522 ,csa_tree_sub001036_groupi_n_652);
  xnor csa_tree_sub001036_groupi_g5247__1666(csa_tree_sub001036_groupi_n_763 ,csa_tree_sub001036_groupi_n_559 ,csa_tree_sub001036_groupi_n_587);
  xor csa_tree_sub001036_groupi_g5248__7410(csa_tree_sub001036_groupi_n_762 ,csa_tree_sub001036_groupi_n_601 ,csa_tree_sub001036_groupi_n_566);
  xor csa_tree_sub001036_groupi_g5249__6417(csa_tree_sub001036_groupi_n_761 ,csa_tree_sub001036_groupi_n_602 ,csa_tree_sub001036_groupi_n_589);
  and csa_tree_sub001036_groupi_g5250__5477(csa_tree_sub001036_groupi_n_794 ,csa_tree_sub001036_groupi_n_643 ,csa_tree_sub001036_groupi_n_696);
  and csa_tree_sub001036_groupi_g5251__2398(csa_tree_sub001036_groupi_n_793 ,csa_tree_sub001036_groupi_n_626 ,csa_tree_sub001036_groupi_n_703);
  or csa_tree_sub001036_groupi_g5252__5107(csa_tree_sub001036_groupi_n_792 ,csa_tree_sub001036_groupi_n_622 ,csa_tree_sub001036_groupi_n_684);
  xnor csa_tree_sub001036_groupi_g5253__6260(csa_tree_sub001036_groupi_n_791 ,csa_tree_sub001036_groupi_n_599 ,csa_tree_sub001036_groupi_n_549);
  xnor csa_tree_sub001036_groupi_g5254__4319(csa_tree_sub001036_groupi_n_790 ,csa_tree_sub001036_groupi_n_538 ,csa_tree_sub001036_groupi_n_547);
  or csa_tree_sub001036_groupi_g5255__8428(csa_tree_sub001036_groupi_n_789 ,csa_tree_sub001036_groupi_n_634 ,csa_tree_sub001036_groupi_n_685);
  and csa_tree_sub001036_groupi_g5256__5526(csa_tree_sub001036_groupi_n_757 ,csa_tree_sub001036_groupi_n_653 ,csa_tree_sub001036_groupi_n_660);
  and csa_tree_sub001036_groupi_g5257__6783(csa_tree_sub001036_groupi_n_756 ,csa_tree_sub001036_groupi_n_486 ,csa_tree_sub001036_groupi_n_650);
  and csa_tree_sub001036_groupi_g5258__3680(csa_tree_sub001036_groupi_n_755 ,csa_tree_sub001036_groupi_n_654 ,csa_tree_sub001036_groupi_n_657);
  or csa_tree_sub001036_groupi_g5259__1617(csa_tree_sub001036_groupi_n_754 ,csa_tree_sub001036_groupi_n_499 ,csa_tree_sub001036_groupi_n_625);
  or csa_tree_sub001036_groupi_g5260__2802(csa_tree_sub001036_groupi_n_753 ,csa_tree_sub001036_groupi_n_521 ,csa_tree_sub001036_groupi_n_651);
  nor csa_tree_sub001036_groupi_g5261__1705(csa_tree_sub001036_groupi_n_752 ,csa_tree_sub001036_groupi_n_654 ,csa_tree_sub001036_groupi_n_657);
  nor csa_tree_sub001036_groupi_g5262__5122(csa_tree_sub001036_groupi_n_751 ,csa_tree_sub001036_groupi_n_522 ,csa_tree_sub001036_groupi_n_652);
  and csa_tree_sub001036_groupi_g5263__8246(csa_tree_sub001036_groupi_n_750 ,csa_tree_sub001036_groupi_n_519 ,csa_tree_sub001036_groupi_n_590);
  nor csa_tree_sub001036_groupi_g5264__7098(csa_tree_sub001036_groupi_n_749 ,csa_tree_sub001036_groupi_n_519 ,csa_tree_sub001036_groupi_n_590);
  and csa_tree_sub001036_groupi_g5265__6131(csa_tree_sub001036_groupi_n_748 ,csa_tree_sub001036_groupi_n_457 ,csa_tree_sub001036_groupi_n_562);
  nor csa_tree_sub001036_groupi_g5266__1881(csa_tree_sub001036_groupi_n_747 ,csa_tree_sub001036_groupi_n_457 ,csa_tree_sub001036_groupi_n_562);
  and csa_tree_sub001036_groupi_g5267__5115(csa_tree_sub001036_groupi_n_746 ,csa_tree_sub001036_groupi_n_466 ,csa_tree_sub001036_groupi_n_584);
  nor csa_tree_sub001036_groupi_g5268__7482(csa_tree_sub001036_groupi_n_745 ,csa_tree_sub001036_groupi_n_466 ,csa_tree_sub001036_groupi_n_584);
  nor csa_tree_sub001036_groupi_g5269__4733(csa_tree_sub001036_groupi_n_744 ,csa_tree_sub001036_groupi_n_569 ,csa_tree_sub001036_groupi_n_574);
  nor csa_tree_sub001036_groupi_g5270__6161(csa_tree_sub001036_groupi_n_743 ,csa_tree_sub001036_groupi_n_563 ,csa_tree_sub001036_groupi_n_649);
  and csa_tree_sub001036_groupi_g5271__9315(csa_tree_sub001036_groupi_n_742 ,csa_tree_sub001036_groupi_n_550 ,csa_tree_sub001036_groupi_n_571);
  nor csa_tree_sub001036_groupi_g5272__9945(csa_tree_sub001036_groupi_n_741 ,csa_tree_sub001036_groupi_n_532 ,csa_tree_sub001036_groupi_n_639);
  nor csa_tree_sub001036_groupi_g5273__2883(csa_tree_sub001036_groupi_n_740 ,csa_tree_sub001036_groupi_n_534 ,csa_tree_sub001036_groupi_n_635);
  nor csa_tree_sub001036_groupi_g5274__2346(csa_tree_sub001036_groupi_n_739 ,csa_tree_sub001036_groupi_n_566 ,csa_tree_sub001036_groupi_n_659);
  or csa_tree_sub001036_groupi_g5275__1666(csa_tree_sub001036_groupi_n_738 ,csa_tree_sub001036_groupi_n_487 ,csa_tree_sub001036_groupi_n_637);
  and csa_tree_sub001036_groupi_g5276__7410(csa_tree_sub001036_groupi_n_737 ,csa_tree_sub001036_groupi_n_576 ,csa_tree_sub001036_groupi_n_572);
  nor csa_tree_sub001036_groupi_g5277__6417(csa_tree_sub001036_groupi_n_736 ,csa_tree_sub001036_groupi_n_576 ,csa_tree_sub001036_groupi_n_572);
  and csa_tree_sub001036_groupi_g5278__5477(csa_tree_sub001036_groupi_n_735 ,csa_tree_sub001036_groupi_n_563 ,csa_tree_sub001036_groupi_n_649);
  or csa_tree_sub001036_groupi_g5279__2398(csa_tree_sub001036_groupi_n_734 ,csa_tree_sub001036_groupi_n_580 ,csa_tree_sub001036_groupi_n_552);
  nor csa_tree_sub001036_groupi_g5280__5107(csa_tree_sub001036_groupi_n_733 ,csa_tree_sub001036_groupi_n_653 ,csa_tree_sub001036_groupi_n_660);
  and csa_tree_sub001036_groupi_g5281__6260(csa_tree_sub001036_groupi_n_732 ,csa_tree_sub001036_groupi_n_619 ,csa_tree_sub001036_groupi_n_597);
  and csa_tree_sub001036_groupi_g5282__4319(csa_tree_sub001036_groupi_n_731 ,csa_tree_sub001036_groupi_n_520 ,csa_tree_sub001036_groupi_n_575);
  or csa_tree_sub001036_groupi_g5283__8428(csa_tree_sub001036_groupi_n_730 ,csa_tree_sub001036_groupi_n_520 ,csa_tree_sub001036_groupi_n_575);
  or csa_tree_sub001036_groupi_g5284__5526(csa_tree_sub001036_groupi_n_729 ,csa_tree_sub001036_groupi_n_655 ,csa_tree_sub001036_groupi_n_581);
  nor csa_tree_sub001036_groupi_g5285__6783(csa_tree_sub001036_groupi_n_728 ,csa_tree_sub001036_groupi_n_656 ,csa_tree_sub001036_groupi_n_582);
  or csa_tree_sub001036_groupi_g5286__3680(csa_tree_sub001036_groupi_n_727 ,csa_tree_sub001036_groupi_n_565 ,csa_tree_sub001036_groupi_n_658);
  nor csa_tree_sub001036_groupi_g5287__1617(csa_tree_sub001036_groupi_n_726 ,csa_tree_sub001036_groupi_n_550 ,csa_tree_sub001036_groupi_n_571);
  nor csa_tree_sub001036_groupi_g5288__2802(csa_tree_sub001036_groupi_n_725 ,csa_tree_sub001036_groupi_n_486 ,csa_tree_sub001036_groupi_n_650);
  or csa_tree_sub001036_groupi_g5289__1705(csa_tree_sub001036_groupi_n_724 ,csa_tree_sub001036_groupi_n_570 ,csa_tree_sub001036_groupi_n_661);
  and csa_tree_sub001036_groupi_g5290__5122(csa_tree_sub001036_groupi_n_723 ,csa_tree_sub001036_groupi_n_535 ,csa_tree_sub001036_groupi_n_617);
  or csa_tree_sub001036_groupi_g5291__8246(csa_tree_sub001036_groupi_n_722 ,csa_tree_sub001036_groupi_n_492 ,csa_tree_sub001036_groupi_n_610);
  nor csa_tree_sub001036_groupi_g5292__7098(csa_tree_sub001036_groupi_n_721 ,csa_tree_sub001036_groupi_n_465 ,csa_tree_sub001036_groupi_n_554);
  or csa_tree_sub001036_groupi_g5293__6131(csa_tree_sub001036_groupi_n_720 ,csa_tree_sub001036_groupi_n_155 ,csa_tree_sub001036_groupi_n_558);
  or csa_tree_sub001036_groupi_g5294__1881(csa_tree_sub001036_groupi_n_719 ,csa_tree_sub001036_groupi_n_468 ,csa_tree_sub001036_groupi_n_578);
  nor csa_tree_sub001036_groupi_g5295__5115(csa_tree_sub001036_groupi_n_718 ,csa_tree_sub001036_groupi_n_589 ,csa_tree_sub001036_groupi_n_588);
  nor csa_tree_sub001036_groupi_g5296__7482(csa_tree_sub001036_groupi_n_717 ,csa_tree_sub001036_groupi_n_488 ,csa_tree_sub001036_groupi_n_624);
  and csa_tree_sub001036_groupi_g5297__4733(csa_tree_sub001036_groupi_n_716 ,csa_tree_sub001036_groupi_n_469 ,csa_tree_sub001036_groupi_n_564);
  and csa_tree_sub001036_groupi_g5298__6161(csa_tree_sub001036_groupi_n_715 ,csa_tree_sub001036_groupi_n_460 ,csa_tree_sub001036_groupi_n_586);
  and csa_tree_sub001036_groupi_g5299__9315(csa_tree_sub001036_groupi_n_714 ,csa_tree_sub001036_groupi_n_490 ,csa_tree_sub001036_groupi_n_627);
  or csa_tree_sub001036_groupi_g5300__9945(csa_tree_sub001036_groupi_n_760 ,csa_tree_sub001036_groupi_n_314 ,csa_tree_sub001036_groupi_n_630);
  or csa_tree_sub001036_groupi_g5301__2883(csa_tree_sub001036_groupi_n_759 ,csa_tree_sub001036_groupi_n_315 ,csa_tree_sub001036_groupi_n_632);
  and csa_tree_sub001036_groupi_g5302__2346(csa_tree_sub001036_groupi_n_758 ,csa_tree_sub001036_groupi_n_500 ,csa_tree_sub001036_groupi_n_618);
  not csa_tree_sub001036_groupi_g5303(csa_tree_sub001036_groupi_n_712 ,csa_tree_sub001036_groupi_n_711);
  nor csa_tree_sub001036_groupi_g5304__1666(csa_tree_sub001036_groupi_n_710 ,csa_tree_sub001036_groupi_n_460 ,csa_tree_sub001036_groupi_n_586);
  nor csa_tree_sub001036_groupi_g5305__7410(csa_tree_sub001036_groupi_n_709 ,csa_tree_sub001036_groupi_n_544 ,csa_tree_sub001036_groupi_n_614);
  and csa_tree_sub001036_groupi_g5306__6417(csa_tree_sub001036_groupi_n_708 ,csa_tree_sub001036_groupi_n_589 ,csa_tree_sub001036_groupi_n_588);
  nor csa_tree_sub001036_groupi_g5307__5477(csa_tree_sub001036_groupi_n_707 ,csa_tree_sub001036_groupi_n_469 ,csa_tree_sub001036_groupi_n_564);
  nor csa_tree_sub001036_groupi_g5308__2398(csa_tree_sub001036_groupi_n_706 ,csa_tree_sub001036_groupi_n_542 ,csa_tree_sub001036_groupi_n_620);
  and csa_tree_sub001036_groupi_g5309__5107(csa_tree_sub001036_groupi_n_705 ,csa_tree_sub001036_groupi_n_570 ,csa_tree_sub001036_groupi_n_661);
  nor csa_tree_sub001036_groupi_g5310__6260(csa_tree_sub001036_groupi_n_704 ,csa_tree_sub001036_groupi_n_49 ,csa_tree_sub001036_groupi_n_559);
  or csa_tree_sub001036_groupi_g5311__4319(csa_tree_sub001036_groupi_n_703 ,csa_tree_sub001036_groupi_n_494 ,csa_tree_sub001036_groupi_n_623);
  and csa_tree_sub001036_groupi_g5312__8428(csa_tree_sub001036_groupi_n_702 ,csa_tree_sub001036_groupi_n_458 ,csa_tree_sub001036_groupi_n_599);
  or csa_tree_sub001036_groupi_g5313__5526(csa_tree_sub001036_groupi_n_701 ,csa_tree_sub001036_groupi_n_568 ,csa_tree_sub001036_groupi_n_573);
  and csa_tree_sub001036_groupi_g5314__6783(csa_tree_sub001036_groupi_n_700 ,csa_tree_sub001036_groupi_n_545 ,csa_tree_sub001036_groupi_n_611);
  or csa_tree_sub001036_groupi_g5315__3680(csa_tree_sub001036_groupi_n_699 ,csa_tree_sub001036_groupi_n_551 ,csa_tree_sub001036_groupi_n_555);
  or csa_tree_sub001036_groupi_g5316__1617(csa_tree_sub001036_groupi_n_698 ,csa_tree_sub001036_groupi_n_472 ,csa_tree_sub001036_groupi_n_560);
  nor csa_tree_sub001036_groupi_g5317__2802(csa_tree_sub001036_groupi_n_697 ,csa_tree_sub001036_groupi_n_526 ,csa_tree_sub001036_groupi_n_556);
  or csa_tree_sub001036_groupi_g5318__1705(csa_tree_sub001036_groupi_n_696 ,csa_tree_sub001036_groupi_n_537 ,csa_tree_sub001036_groupi_n_613);
  and csa_tree_sub001036_groupi_g5319__5122(csa_tree_sub001036_groupi_n_695 ,csa_tree_sub001036_groupi_n_478 ,csa_tree_sub001036_groupi_n_567);
  or csa_tree_sub001036_groupi_g5320__8246(csa_tree_sub001036_groupi_n_694 ,csa_tree_sub001036_groupi_n_525 ,csa_tree_sub001036_groupi_n_557);
  and csa_tree_sub001036_groupi_g5321__7098(csa_tree_sub001036_groupi_n_693 ,csa_tree_sub001036_groupi_n_551 ,csa_tree_sub001036_groupi_n_555);
  or csa_tree_sub001036_groupi_g5322__6131(csa_tree_sub001036_groupi_n_692 ,csa_tree_sub001036_groupi_n_464 ,csa_tree_sub001036_groupi_n_553);
  and csa_tree_sub001036_groupi_g5323__1881(csa_tree_sub001036_groupi_n_691 ,csa_tree_sub001036_groupi_n_468 ,csa_tree_sub001036_groupi_n_578);
  nor csa_tree_sub001036_groupi_g5324__5115(csa_tree_sub001036_groupi_n_690 ,csa_tree_sub001036_groupi_n_478 ,csa_tree_sub001036_groupi_n_567);
  and csa_tree_sub001036_groupi_g5325__7482(csa_tree_sub001036_groupi_n_689 ,csa_tree_sub001036_groupi_n_580 ,csa_tree_sub001036_groupi_n_552);
  and csa_tree_sub001036_groupi_g5326__4733(csa_tree_sub001036_groupi_n_688 ,csa_tree_sub001036_groupi_n_456 ,csa_tree_sub001036_groupi_n_583);
  nor csa_tree_sub001036_groupi_g5327__6161(csa_tree_sub001036_groupi_n_687 ,csa_tree_sub001036_groupi_n_473 ,csa_tree_sub001036_groupi_n_561);
  or csa_tree_sub001036_groupi_g5328__9315(csa_tree_sub001036_groupi_n_686 ,csa_tree_sub001036_groupi_n_456 ,csa_tree_sub001036_groupi_n_583);
  and csa_tree_sub001036_groupi_g5329__9945(csa_tree_sub001036_groupi_n_685 ,csa_tree_sub001036_groupi_n_612 ,csa_tree_sub001036_groupi_n_663);
  and csa_tree_sub001036_groupi_g5330__2883(csa_tree_sub001036_groupi_n_684 ,csa_tree_sub001036_groupi_n_546 ,csa_tree_sub001036_groupi_n_609);
  xnor csa_tree_sub001036_groupi_g5331__2346(csa_tree_sub001036_groupi_n_683 ,csa_tree_sub001036_groupi_n_493 ,csa_tree_sub001036_groupi_n_323);
  xnor csa_tree_sub001036_groupi_g5332__1666(csa_tree_sub001036_groupi_n_682 ,csa_tree_sub001036_groupi_n_257 ,csa_tree_sub001036_groupi_n_546);
  xnor csa_tree_sub001036_groupi_g5333__7410(csa_tree_sub001036_groupi_n_681 ,csa_tree_sub001036_groupi_n_489 ,csa_tree_sub001036_groupi_n_473);
  xnor csa_tree_sub001036_groupi_g5334__6417(csa_tree_sub001036_groupi_n_680 ,csa_tree_sub001036_groupi_n_467 ,csa_tree_sub001036_groupi_n_475);
  xor csa_tree_sub001036_groupi_g5335__5477(csa_tree_sub001036_groupi_n_679 ,csa_tree_sub001036_groupi_n_499 ,csa_tree_sub001036_groupi_n_463);
  xnor csa_tree_sub001036_groupi_g5336__2398(csa_tree_sub001036_groupi_n_678 ,csa_tree_sub001036_groupi_n_507 ,csa_tree_sub001036_groupi_n_513);
  xnor csa_tree_sub001036_groupi_g5337__5107(csa_tree_sub001036_groupi_n_677 ,csa_tree_sub001036_groupi_n_523 ,csa_tree_sub001036_groupi_n_253);
  xor csa_tree_sub001036_groupi_g5338__6260(csa_tree_sub001036_groupi_n_676 ,csa_tree_sub001036_groupi_n_532 ,csa_tree_sub001036_groupi_n_528);
  xnor csa_tree_sub001036_groupi_g5339__4319(csa_tree_sub001036_groupi_n_675 ,csa_tree_sub001036_groupi_n_531 ,csa_tree_sub001036_groupi_n_518);
  xor csa_tree_sub001036_groupi_g5340__8428(csa_tree_sub001036_groupi_n_674 ,csa_tree_sub001036_groupi_n_533 ,csa_tree_sub001036_groupi_n_486);
  xnor csa_tree_sub001036_groupi_g5341__5526(csa_tree_sub001036_groupi_n_673 ,csa_tree_sub001036_groupi_n_510 ,csa_tree_sub001036_groupi_n_541);
  xor csa_tree_sub001036_groupi_g5342__6783(csa_tree_sub001036_groupi_n_672 ,csa_tree_sub001036_groupi_n_534 ,csa_tree_sub001036_groupi_n_45);
  xor csa_tree_sub001036_groupi_g5343__3680(csa_tree_sub001036_groupi_n_671 ,csa_tree_sub001036_groupi_n_488 ,csa_tree_sub001036_groupi_n_511);
  xnor csa_tree_sub001036_groupi_g5344__1617(csa_tree_sub001036_groupi_n_670 ,csa_tree_sub001036_groupi_n_482 ,csa_tree_sub001036_groupi_n_481);
  xor csa_tree_sub001036_groupi_g5345__2802(csa_tree_sub001036_groupi_n_669 ,csa_tree_sub001036_groupi_n_496 ,csa_tree_sub001036_groupi_n_478);
  xnor csa_tree_sub001036_groupi_g5346__1705(csa_tree_sub001036_groupi_n_668 ,csa_tree_sub001036_groupi_n_476 ,csa_tree_sub001036_groupi_n_477);
  xor csa_tree_sub001036_groupi_g5347__5122(csa_tree_sub001036_groupi_n_667 ,csa_tree_sub001036_groupi_n_487 ,csa_tree_sub001036_groupi_n_509);
  xnor csa_tree_sub001036_groupi_g5348__8246(csa_tree_sub001036_groupi_n_666 ,csa_tree_sub001036_groupi_n_461 ,csa_tree_sub001036_groupi_n_474);
  xnor csa_tree_sub001036_groupi_g5349__7098(csa_tree_sub001036_groupi_n_665 ,csa_tree_sub001036_groupi_n_524 ,csa_tree_sub001036_groupi_n_543);
  xnor csa_tree_sub001036_groupi_g5350__6131(csa_tree_sub001036_groupi_n_713 ,csa_tree_sub001036_groupi_n_495 ,csa_tree_sub001036_groupi_n_383);
  xnor csa_tree_sub001036_groupi_g5351__1881(csa_tree_sub001036_groupi_n_711 ,csa_tree_sub001036_groupi_n_497 ,csa_tree_sub001036_groupi_n_384);
  not csa_tree_sub001036_groupi_g5352(csa_tree_sub001036_groupi_n_658 ,csa_tree_sub001036_groupi_n_659);
  not csa_tree_sub001036_groupi_g5353(csa_tree_sub001036_groupi_n_655 ,csa_tree_sub001036_groupi_n_656);
  not csa_tree_sub001036_groupi_g5354(csa_tree_sub001036_groupi_n_651 ,csa_tree_sub001036_groupi_n_652);
  not csa_tree_sub001036_groupi_g5355(csa_tree_sub001036_groupi_n_649 ,csa_tree_sub001036_groupi_n_648);
  not csa_tree_sub001036_groupi_g5356(csa_tree_sub001036_groupi_n_646 ,csa_tree_sub001036_groupi_n_647);
  not csa_tree_sub001036_groupi_g5357(csa_tree_sub001036_groupi_n_644 ,csa_tree_sub001036_groupi_n_645);
  or csa_tree_sub001036_groupi_g5358__5115(csa_tree_sub001036_groupi_n_643 ,csa_tree_sub001036_groupi_n_530 ,csa_tree_sub001036_groupi_n_517);
  and csa_tree_sub001036_groupi_g5359__7482(csa_tree_sub001036_groupi_n_642 ,csa_tree_sub001036_groupi_n_524 ,csa_tree_sub001036_groupi_n_91);
  and csa_tree_sub001036_groupi_g5360__4733(csa_tree_sub001036_groupi_n_641 ,csa_tree_sub001036_groupi_n_26 ,csa_tree_sub001036_groupi_n_527);
  and csa_tree_sub001036_groupi_g5361__6161(csa_tree_sub001036_groupi_n_640 ,csa_tree_sub001036_groupi_n_529 ,csa_tree_sub001036_groupi_n_528);
  nor csa_tree_sub001036_groupi_g5362__9315(csa_tree_sub001036_groupi_n_639 ,csa_tree_sub001036_groupi_n_529 ,csa_tree_sub001036_groupi_n_528);
  or csa_tree_sub001036_groupi_g5363__9945(csa_tree_sub001036_groupi_n_638 ,csa_tree_sub001036_groupi_n_470 ,csa_tree_sub001036_groupi_n_508);
  nor csa_tree_sub001036_groupi_g5364__2883(csa_tree_sub001036_groupi_n_637 ,csa_tree_sub001036_groupi_n_471 ,csa_tree_sub001036_groupi_n_509);
  and csa_tree_sub001036_groupi_g5365__2346(csa_tree_sub001036_groupi_n_636 ,csa_tree_sub001036_groupi_n_461 ,csa_tree_sub001036_groupi_n_474);
  nor csa_tree_sub001036_groupi_g5366__1666(csa_tree_sub001036_groupi_n_635 ,csa_tree_sub001036_groupi_n_144 ,csa_tree_sub001036_groupi_n_527);
  and csa_tree_sub001036_groupi_g5367__7410(csa_tree_sub001036_groupi_n_634 ,csa_tree_sub001036_groupi_n_467 ,csa_tree_sub001036_groupi_n_475);
  and csa_tree_sub001036_groupi_g5368__6417(csa_tree_sub001036_groupi_n_633 ,csa_tree_sub001036_groupi_n_252 ,csa_tree_sub001036_groupi_n_523);
  and csa_tree_sub001036_groupi_g5369__5477(csa_tree_sub001036_groupi_n_632 ,csa_tree_sub001036_groupi_n_313 ,csa_tree_sub001036_groupi_n_497);
  and csa_tree_sub001036_groupi_g5370__2398(csa_tree_sub001036_groupi_n_631 ,csa_tree_sub001036_groupi_n_476 ,csa_tree_sub001036_groupi_n_477);
  and csa_tree_sub001036_groupi_g5371__5107(csa_tree_sub001036_groupi_n_630 ,csa_tree_sub001036_groupi_n_316 ,csa_tree_sub001036_groupi_n_495);
  or csa_tree_sub001036_groupi_g5372__6260(csa_tree_sub001036_groupi_n_629 ,csa_tree_sub001036_groupi_n_462 ,csa_tree_sub001036_groupi_n_483);
  and csa_tree_sub001036_groupi_g5373__4319(csa_tree_sub001036_groupi_n_628 ,csa_tree_sub001036_groupi_n_482 ,csa_tree_sub001036_groupi_n_481);
  or csa_tree_sub001036_groupi_g5374__8428(csa_tree_sub001036_groupi_n_627 ,csa_tree_sub001036_groupi_n_476 ,csa_tree_sub001036_groupi_n_477);
  or csa_tree_sub001036_groupi_g5375__5526(csa_tree_sub001036_groupi_n_626 ,csa_tree_sub001036_groupi_n_58 ,csa_tree_sub001036_groupi_n_479);
  nor csa_tree_sub001036_groupi_g5376__6783(csa_tree_sub001036_groupi_n_625 ,csa_tree_sub001036_groupi_n_463 ,csa_tree_sub001036_groupi_n_484);
  nor csa_tree_sub001036_groupi_g5377__3680(csa_tree_sub001036_groupi_n_624 ,csa_tree_sub001036_groupi_n_485 ,csa_tree_sub001036_groupi_n_511);
  nor csa_tree_sub001036_groupi_g5378__1617(csa_tree_sub001036_groupi_n_623 ,csa_tree_sub001036_groupi_n_154 ,csa_tree_sub001036_groupi_n_480);
  nor csa_tree_sub001036_groupi_g5379__2802(csa_tree_sub001036_groupi_n_622 ,csa_tree_sub001036_groupi_n_257 ,csa_tree_sub001036_groupi_n_514);
  and csa_tree_sub001036_groupi_g5380__1705(csa_tree_sub001036_groupi_n_621 ,csa_tree_sub001036_groupi_n_510 ,csa_tree_sub001036_groupi_n_516);
  nor csa_tree_sub001036_groupi_g5381__5122(csa_tree_sub001036_groupi_n_620 ,csa_tree_sub001036_groupi_n_510 ,csa_tree_sub001036_groupi_n_516);
  or csa_tree_sub001036_groupi_g5382__8246(csa_tree_sub001036_groupi_n_619 ,csa_tree_sub001036_groupi_n_482 ,csa_tree_sub001036_groupi_n_481);
  or csa_tree_sub001036_groupi_g5383__7098(csa_tree_sub001036_groupi_n_618 ,csa_tree_sub001036_groupi_n_539 ,csa_tree_sub001036_groupi_n_501);
  or csa_tree_sub001036_groupi_g5384__6131(csa_tree_sub001036_groupi_n_617 ,csa_tree_sub001036_groupi_n_252 ,csa_tree_sub001036_groupi_n_523);
  and csa_tree_sub001036_groupi_g5385__1881(csa_tree_sub001036_groupi_n_616 ,csa_tree_sub001036_groupi_n_485 ,csa_tree_sub001036_groupi_n_511);
  or csa_tree_sub001036_groupi_g5386__5115(csa_tree_sub001036_groupi_n_615 ,csa_tree_sub001036_groupi_n_506 ,csa_tree_sub001036_groupi_n_512);
  nor csa_tree_sub001036_groupi_g5387__7482(csa_tree_sub001036_groupi_n_614 ,csa_tree_sub001036_groupi_n_57 ,csa_tree_sub001036_groupi_n_524);
  nor csa_tree_sub001036_groupi_g5388__4733(csa_tree_sub001036_groupi_n_613 ,csa_tree_sub001036_groupi_n_531 ,csa_tree_sub001036_groupi_n_518);
  or csa_tree_sub001036_groupi_g5389__6161(csa_tree_sub001036_groupi_n_612 ,csa_tree_sub001036_groupi_n_467 ,csa_tree_sub001036_groupi_n_475);
  or csa_tree_sub001036_groupi_g5390__9315(csa_tree_sub001036_groupi_n_611 ,csa_tree_sub001036_groupi_n_461 ,csa_tree_sub001036_groupi_n_474);
  nor csa_tree_sub001036_groupi_g5391__9945(csa_tree_sub001036_groupi_n_610 ,csa_tree_sub001036_groupi_n_507 ,csa_tree_sub001036_groupi_n_513);
  or csa_tree_sub001036_groupi_g5392__2883(csa_tree_sub001036_groupi_n_609 ,csa_tree_sub001036_groupi_n_256 ,csa_tree_sub001036_groupi_n_515);
  xor csa_tree_sub001036_groupi_g5393__2346(csa_tree_sub001036_groupi_n_664 ,csa_tree_sub001036_groupi_n_346 ,in11[2]);
  xnor csa_tree_sub001036_groupi_g5394__1666(csa_tree_sub001036_groupi_n_663 ,csa_tree_sub001036_groupi_n_354 ,in25[0]);
  xor csa_tree_sub001036_groupi_g5395__7410(csa_tree_sub001036_groupi_n_662 ,csa_tree_sub001036_groupi_n_361 ,in27[5]);
  xnor csa_tree_sub001036_groupi_g5396__6417(csa_tree_sub001036_groupi_n_661 ,csa_tree_sub001036_groupi_n_363 ,in30[6]);
  xnor csa_tree_sub001036_groupi_g5397__5477(csa_tree_sub001036_groupi_n_660 ,csa_tree_sub001036_groupi_n_326 ,in26[2]);
  xnor csa_tree_sub001036_groupi_g5398__2398(csa_tree_sub001036_groupi_n_659 ,csa_tree_sub001036_groupi_n_336 ,in7[5]);
  xnor csa_tree_sub001036_groupi_g5399__5107(csa_tree_sub001036_groupi_n_657 ,csa_tree_sub001036_groupi_n_364 ,in8[6]);
  xnor csa_tree_sub001036_groupi_g5400__6260(csa_tree_sub001036_groupi_n_656 ,csa_tree_sub001036_groupi_n_368 ,in10[2]);
  xnor csa_tree_sub001036_groupi_g5401__4319(csa_tree_sub001036_groupi_n_654 ,csa_tree_sub001036_groupi_n_366 ,in12[6]);
  xnor csa_tree_sub001036_groupi_g5402__8428(csa_tree_sub001036_groupi_n_653 ,csa_tree_sub001036_groupi_n_371 ,in11[3]);
  xnor csa_tree_sub001036_groupi_g5403__5526(csa_tree_sub001036_groupi_n_652 ,csa_tree_sub001036_groupi_n_374 ,csa_tree_sub001036_groupi_n_112);
  xnor csa_tree_sub001036_groupi_g5404__6783(csa_tree_sub001036_groupi_n_650 ,csa_tree_sub001036_groupi_n_351 ,in29[6]);
  xnor csa_tree_sub001036_groupi_g5405__3680(csa_tree_sub001036_groupi_n_648 ,csa_tree_sub001036_groupi_n_387 ,csa_tree_sub001036_groupi_n_85);
  xnor csa_tree_sub001036_groupi_g5406__1617(csa_tree_sub001036_groupi_n_647 ,csa_tree_sub001036_groupi_n_386 ,csa_tree_sub001036_groupi_n_145);
  and csa_tree_sub001036_groupi_g5407__2802(csa_tree_sub001036_groupi_n_645 ,csa_tree_sub001036_groupi_n_295 ,csa_tree_sub001036_groupi_n_459);
  not csa_tree_sub001036_groupi_g5408(csa_tree_sub001036_groupi_n_596 ,csa_tree_sub001036_groupi_n_595);
  not csa_tree_sub001036_groupi_g5410(csa_tree_sub001036_groupi_n_581 ,csa_tree_sub001036_groupi_n_582);
  not csa_tree_sub001036_groupi_g5411(csa_tree_sub001036_groupi_n_580 ,csa_tree_sub001036_groupi_n_579);
  not csa_tree_sub001036_groupi_g5412(csa_tree_sub001036_groupi_n_578 ,csa_tree_sub001036_groupi_n_577);
  not csa_tree_sub001036_groupi_g5413(csa_tree_sub001036_groupi_n_573 ,csa_tree_sub001036_groupi_n_574);
  not csa_tree_sub001036_groupi_g5414(csa_tree_sub001036_groupi_n_568 ,csa_tree_sub001036_groupi_n_569);
  not csa_tree_sub001036_groupi_g5415(csa_tree_sub001036_groupi_n_565 ,csa_tree_sub001036_groupi_n_566);
  not csa_tree_sub001036_groupi_g5416(csa_tree_sub001036_groupi_n_560 ,csa_tree_sub001036_groupi_n_561);
  not csa_tree_sub001036_groupi_g5417(csa_tree_sub001036_groupi_n_558 ,csa_tree_sub001036_groupi_n_559);
  not csa_tree_sub001036_groupi_g5418(csa_tree_sub001036_groupi_n_556 ,csa_tree_sub001036_groupi_n_557);
  not csa_tree_sub001036_groupi_g5419(csa_tree_sub001036_groupi_n_553 ,csa_tree_sub001036_groupi_n_554);
  xnor csa_tree_sub001036_groupi_g5420__1705(csa_tree_sub001036_groupi_n_549 ,csa_tree_sub001036_groupi_n_255 ,csa_tree_sub001036_groupi_n_391);
  xnor csa_tree_sub001036_groupi_g5421__5122(csa_tree_sub001036_groupi_n_548 ,csa_tree_sub001036_groupi_n_392 ,csa_tree_sub001036_groupi_n_106);
  xnor csa_tree_sub001036_groupi_g5422__8246(csa_tree_sub001036_groupi_n_547 ,csa_tree_sub001036_groupi_n_389 ,csa_tree_sub001036_groupi_n_142);
  xnor csa_tree_sub001036_groupi_g5423__7098(csa_tree_sub001036_groupi_n_608 ,csa_tree_sub001036_groupi_n_359 ,in10[3]);
  xor csa_tree_sub001036_groupi_g5424__6131(csa_tree_sub001036_groupi_n_607 ,csa_tree_sub001036_groupi_n_352 ,in30[4]);
  xor csa_tree_sub001036_groupi_g5425__1881(csa_tree_sub001036_groupi_n_606 ,csa_tree_sub001036_groupi_n_348 ,in30[2]);
  xor csa_tree_sub001036_groupi_g5426__5115(csa_tree_sub001036_groupi_n_605 ,csa_tree_sub001036_groupi_n_370 ,in25[3]);
  xor csa_tree_sub001036_groupi_g5427__7482(csa_tree_sub001036_groupi_n_604 ,csa_tree_sub001036_groupi_n_335 ,in26[4]);
  xor csa_tree_sub001036_groupi_g5428__4733(csa_tree_sub001036_groupi_n_603 ,csa_tree_sub001036_groupi_n_330 ,in15[4]);
  xor csa_tree_sub001036_groupi_g5429__6161(csa_tree_sub001036_groupi_n_602 ,csa_tree_sub001036_groupi_n_339 ,in15[1]);
  xor csa_tree_sub001036_groupi_g5430__9315(csa_tree_sub001036_groupi_n_601 ,csa_tree_sub001036_groupi_n_343 ,in8[5]);
  xnor csa_tree_sub001036_groupi_g5431__9945(csa_tree_sub001036_groupi_n_600 ,csa_tree_sub001036_groupi_n_355 ,in13[1]);
  xnor csa_tree_sub001036_groupi_g5432__2883(csa_tree_sub001036_groupi_n_599 ,csa_tree_sub001036_groupi_n_328 ,in11[0]);
  xnor csa_tree_sub001036_groupi_g5433__2346(csa_tree_sub001036_groupi_n_598 ,csa_tree_sub001036_groupi_n_258 ,csa_tree_sub001036_groupi_n_376);
  xnor csa_tree_sub001036_groupi_g5434__1666(csa_tree_sub001036_groupi_n_597 ,csa_tree_sub001036_groupi_n_341 ,in26[5]);
  xnor csa_tree_sub001036_groupi_g5435__7410(csa_tree_sub001036_groupi_n_595 ,csa_tree_sub001036_groupi_n_360 ,in28[1]);
  xnor csa_tree_sub001036_groupi_g5436__6417(csa_tree_sub001036_groupi_n_594 ,csa_tree_sub001036_groupi_n_393 ,csa_tree_sub001036_groupi_n_39);
  xnor csa_tree_sub001036_groupi_g5437__5477(csa_tree_sub001036_groupi_n_593 ,csa_tree_sub001036_groupi_n_345 ,csa_tree_sub001036_groupi_n_88);
  xnor csa_tree_sub001036_groupi_g5438__2398(csa_tree_sub001036_groupi_n_592 ,csa_tree_sub001036_groupi_n_356 ,in8[2]);
  xnor csa_tree_sub001036_groupi_g5439__5107(csa_tree_sub001036_groupi_n_591 ,csa_tree_sub001036_groupi_n_379 ,csa_tree_sub001036_groupi_n_105);
  xnor csa_tree_sub001036_groupi_g5440__6260(csa_tree_sub001036_groupi_n_590 ,csa_tree_sub001036_groupi_n_367 ,in13[4]);
  xnor csa_tree_sub001036_groupi_g5441__4319(csa_tree_sub001036_groupi_n_589 ,csa_tree_sub001036_groupi_n_332 ,in27[0]);
  xnor csa_tree_sub001036_groupi_g5442__8428(csa_tree_sub001036_groupi_n_588 ,csa_tree_sub001036_groupi_n_378 ,csa_tree_sub001036_groupi_n_117);
  xnor csa_tree_sub001036_groupi_g5443__5526(csa_tree_sub001036_groupi_n_587 ,csa_tree_sub001036_groupi_n_377 ,csa_tree_sub001036_groupi_n_37);
  xnor csa_tree_sub001036_groupi_g5444__6783(csa_tree_sub001036_groupi_n_586 ,csa_tree_sub001036_groupi_n_337 ,in11[5]);
  xnor csa_tree_sub001036_groupi_g5445__3680(csa_tree_sub001036_groupi_n_585 ,csa_tree_sub001036_groupi_n_373 ,csa_tree_sub001036_groupi_n_72);
  xnor csa_tree_sub001036_groupi_g5446__1617(csa_tree_sub001036_groupi_n_584 ,csa_tree_sub001036_groupi_n_349 ,in9[4]);
  xnor csa_tree_sub001036_groupi_g5447__2802(csa_tree_sub001036_groupi_n_583 ,csa_tree_sub001036_groupi_n_333 ,in24[0]);
  xnor csa_tree_sub001036_groupi_g5448__1705(csa_tree_sub001036_groupi_n_582 ,csa_tree_sub001036_groupi_n_369 ,in30[1]);
  xnor csa_tree_sub001036_groupi_g5449__5122(csa_tree_sub001036_groupi_n_579 ,csa_tree_sub001036_groupi_n_372 ,csa_tree_sub001036_groupi_n_61);
  xnor csa_tree_sub001036_groupi_g5450__8246(csa_tree_sub001036_groupi_n_577 ,csa_tree_sub001036_groupi_n_350 ,in7[2]);
  xnor csa_tree_sub001036_groupi_g5451__7098(csa_tree_sub001036_groupi_n_576 ,csa_tree_sub001036_groupi_n_358 ,in28[2]);
  xnor csa_tree_sub001036_groupi_g5452__6131(csa_tree_sub001036_groupi_n_575 ,csa_tree_sub001036_groupi_n_353 ,in26[1]);
  xnor csa_tree_sub001036_groupi_g5453__1881(csa_tree_sub001036_groupi_n_574 ,csa_tree_sub001036_groupi_n_334 ,in9[0]);
  xnor csa_tree_sub001036_groupi_g5454__5115(csa_tree_sub001036_groupi_n_572 ,csa_tree_sub001036_groupi_n_357 ,in8[3]);
  xnor csa_tree_sub001036_groupi_g5455__7482(csa_tree_sub001036_groupi_n_571 ,csa_tree_sub001036_groupi_n_338 ,in28[5]);
  xnor csa_tree_sub001036_groupi_g5456__4733(csa_tree_sub001036_groupi_n_570 ,csa_tree_sub001036_groupi_n_331 ,in24[6]);
  xnor csa_tree_sub001036_groupi_g5457__6161(csa_tree_sub001036_groupi_n_569 ,csa_tree_sub001036_groupi_n_327 ,in10[0]);
  xnor csa_tree_sub001036_groupi_g5458__9315(csa_tree_sub001036_groupi_n_567 ,csa_tree_sub001036_groupi_n_362 ,in9[1]);
  xnor csa_tree_sub001036_groupi_g5459__9945(csa_tree_sub001036_groupi_n_566 ,csa_tree_sub001036_groupi_n_365 ,in10[5]);
  xnor csa_tree_sub001036_groupi_g5460__2883(csa_tree_sub001036_groupi_n_564 ,csa_tree_sub001036_groupi_n_340 ,in28[4]);
  xnor csa_tree_sub001036_groupi_g5461__2346(csa_tree_sub001036_groupi_n_563 ,csa_tree_sub001036_groupi_n_388 ,csa_tree_sub001036_groupi_n_103);
  xnor csa_tree_sub001036_groupi_g5462__1666(csa_tree_sub001036_groupi_n_562 ,csa_tree_sub001036_groupi_n_342 ,in27[3]);
  xnor csa_tree_sub001036_groupi_g5463__7410(csa_tree_sub001036_groupi_n_561 ,csa_tree_sub001036_groupi_n_344 ,in23[5]);
  xnor csa_tree_sub001036_groupi_g5464__6417(csa_tree_sub001036_groupi_n_559 ,csa_tree_sub001036_groupi_n_381 ,csa_tree_sub001036_groupi_n_84);
  xnor csa_tree_sub001036_groupi_g5465__5477(csa_tree_sub001036_groupi_n_557 ,csa_tree_sub001036_groupi_n_347 ,in7[3]);
  xnor csa_tree_sub001036_groupi_g5466__2398(csa_tree_sub001036_groupi_n_555 ,csa_tree_sub001036_groupi_n_380 ,csa_tree_sub001036_groupi_n_35);
  xnor csa_tree_sub001036_groupi_g5467__5107(csa_tree_sub001036_groupi_n_554 ,csa_tree_sub001036_groupi_n_382 ,csa_tree_sub001036_groupi_n_43);
  xnor csa_tree_sub001036_groupi_g5468__6260(csa_tree_sub001036_groupi_n_552 ,csa_tree_sub001036_groupi_n_385 ,csa_tree_sub001036_groupi_n_76);
  xnor csa_tree_sub001036_groupi_g5469__4319(csa_tree_sub001036_groupi_n_551 ,csa_tree_sub001036_groupi_n_375 ,csa_tree_sub001036_groupi_n_109);
  xnor csa_tree_sub001036_groupi_g5470__8428(csa_tree_sub001036_groupi_n_550 ,csa_tree_sub001036_groupi_n_329 ,in18[6]);
  not csa_tree_sub001036_groupi_g5471(csa_tree_sub001036_groupi_n_544 ,csa_tree_sub001036_groupi_n_543);
  not csa_tree_sub001036_groupi_g5472(csa_tree_sub001036_groupi_n_542 ,csa_tree_sub001036_groupi_n_541);
  not csa_tree_sub001036_groupi_g5473(csa_tree_sub001036_groupi_n_539 ,csa_tree_sub001036_groupi_n_538);
  not csa_tree_sub001036_groupi_g5474(csa_tree_sub001036_groupi_n_537 ,csa_tree_sub001036_groupi_n_536);
  not csa_tree_sub001036_groupi_g5475(csa_tree_sub001036_groupi_n_530 ,csa_tree_sub001036_groupi_n_531);
  not csa_tree_sub001036_groupi_g5476(csa_tree_sub001036_groupi_n_525 ,csa_tree_sub001036_groupi_n_526);
  not csa_tree_sub001036_groupi_g5477(csa_tree_sub001036_groupi_n_521 ,csa_tree_sub001036_groupi_n_522);
  not csa_tree_sub001036_groupi_g5478(csa_tree_sub001036_groupi_n_517 ,csa_tree_sub001036_groupi_n_518);
  not csa_tree_sub001036_groupi_g5479(csa_tree_sub001036_groupi_n_514 ,csa_tree_sub001036_groupi_n_515);
  not csa_tree_sub001036_groupi_g5480(csa_tree_sub001036_groupi_n_512 ,csa_tree_sub001036_groupi_n_513);
  not csa_tree_sub001036_groupi_g5481(csa_tree_sub001036_groupi_n_508 ,csa_tree_sub001036_groupi_n_509);
  not csa_tree_sub001036_groupi_g5482(csa_tree_sub001036_groupi_n_506 ,csa_tree_sub001036_groupi_n_507);
  not csa_tree_sub001036_groupi_g5483(csa_tree_sub001036_groupi_n_504 ,csa_tree_sub001036_groupi_n_47);
  not csa_tree_sub001036_groupi_g5484(csa_tree_sub001036_groupi_n_503 ,csa_tree_sub001036_groupi_n_505);
  nor csa_tree_sub001036_groupi_g5485__5526(csa_tree_sub001036_groupi_n_502 ,csa_tree_sub001036_groupi_n_254 ,csa_tree_sub001036_groupi_n_391);
  and csa_tree_sub001036_groupi_g5486__6783(csa_tree_sub001036_groupi_n_501 ,csa_tree_sub001036_groupi_n_38 ,csa_tree_sub001036_groupi_n_389);
  or csa_tree_sub001036_groupi_g5487__3680(csa_tree_sub001036_groupi_n_500 ,csa_tree_sub001036_groupi_n_32 ,csa_tree_sub001036_groupi_n_389);
  or csa_tree_sub001036_groupi_g5488__1617(csa_tree_sub001036_groupi_n_546 ,csa_tree_sub001036_groupi_n_217 ,csa_tree_sub001036_groupi_n_426);
  or csa_tree_sub001036_groupi_g5489__2802(csa_tree_sub001036_groupi_n_545 ,csa_tree_sub001036_groupi_n_200 ,csa_tree_sub001036_groupi_n_413);
  or csa_tree_sub001036_groupi_g5490__1705(csa_tree_sub001036_groupi_n_543 ,csa_tree_sub001036_groupi_n_216 ,csa_tree_sub001036_groupi_n_428);
  or csa_tree_sub001036_groupi_g5491__5122(csa_tree_sub001036_groupi_n_541 ,csa_tree_sub001036_groupi_n_286 ,csa_tree_sub001036_groupi_n_418);
  and csa_tree_sub001036_groupi_g5492__8246(csa_tree_sub001036_groupi_n_540 ,csa_tree_sub001036_groupi_n_213 ,csa_tree_sub001036_groupi_n_406);
  or csa_tree_sub001036_groupi_g5493__7098(csa_tree_sub001036_groupi_n_538 ,csa_tree_sub001036_groupi_n_239 ,csa_tree_sub001036_groupi_n_449);
  or csa_tree_sub001036_groupi_g5494__6131(csa_tree_sub001036_groupi_n_536 ,csa_tree_sub001036_groupi_n_218 ,csa_tree_sub001036_groupi_n_438);
  or csa_tree_sub001036_groupi_g5495__1881(csa_tree_sub001036_groupi_n_535 ,csa_tree_sub001036_groupi_n_263 ,csa_tree_sub001036_groupi_n_447);
  and csa_tree_sub001036_groupi_g5496__5115(csa_tree_sub001036_groupi_n_534 ,csa_tree_sub001036_groupi_n_265 ,csa_tree_sub001036_groupi_n_436);
  and csa_tree_sub001036_groupi_g5497__7482(csa_tree_sub001036_groupi_n_533 ,csa_tree_sub001036_groupi_n_238 ,csa_tree_sub001036_groupi_n_434);
  and csa_tree_sub001036_groupi_g5498__4733(csa_tree_sub001036_groupi_n_532 ,csa_tree_sub001036_groupi_n_273 ,csa_tree_sub001036_groupi_n_441);
  or csa_tree_sub001036_groupi_g5499__6161(csa_tree_sub001036_groupi_n_531 ,csa_tree_sub001036_groupi_n_247 ,csa_tree_sub001036_groupi_n_443);
  or csa_tree_sub001036_groupi_g5500__9315(csa_tree_sub001036_groupi_n_529 ,csa_tree_sub001036_groupi_n_241 ,csa_tree_sub001036_groupi_n_429);
  or csa_tree_sub001036_groupi_g5501__9945(csa_tree_sub001036_groupi_n_528 ,csa_tree_sub001036_groupi_n_219 ,csa_tree_sub001036_groupi_n_442);
  or csa_tree_sub001036_groupi_g5502__2883(csa_tree_sub001036_groupi_n_527 ,csa_tree_sub001036_groupi_n_193 ,csa_tree_sub001036_groupi_n_440);
  and csa_tree_sub001036_groupi_g5503__2346(csa_tree_sub001036_groupi_n_526 ,csa_tree_sub001036_groupi_n_304 ,csa_tree_sub001036_groupi_n_407);
  or csa_tree_sub001036_groupi_g5504__1666(csa_tree_sub001036_groupi_n_524 ,csa_tree_sub001036_groupi_n_196 ,csa_tree_sub001036_groupi_n_455);
  or csa_tree_sub001036_groupi_g5505__7410(csa_tree_sub001036_groupi_n_523 ,csa_tree_sub001036_groupi_n_276 ,csa_tree_sub001036_groupi_n_445);
  or csa_tree_sub001036_groupi_g5506__6417(csa_tree_sub001036_groupi_n_522 ,csa_tree_sub001036_groupi_n_320 ,csa_tree_sub001036_groupi_n_446);
  or csa_tree_sub001036_groupi_g5507__5477(csa_tree_sub001036_groupi_n_520 ,csa_tree_sub001036_groupi_n_302 ,csa_tree_sub001036_groupi_n_405);
  or csa_tree_sub001036_groupi_g5508__2398(csa_tree_sub001036_groupi_n_519 ,csa_tree_sub001036_groupi_n_325 ,csa_tree_sub001036_groupi_n_396);
  or csa_tree_sub001036_groupi_g5509__5107(csa_tree_sub001036_groupi_n_518 ,csa_tree_sub001036_groupi_n_243 ,csa_tree_sub001036_groupi_n_435);
  or csa_tree_sub001036_groupi_g5510__6260(csa_tree_sub001036_groupi_n_516 ,csa_tree_sub001036_groupi_n_259 ,csa_tree_sub001036_groupi_n_433);
  or csa_tree_sub001036_groupi_g5511__4319(csa_tree_sub001036_groupi_n_515 ,csa_tree_sub001036_groupi_n_292 ,csa_tree_sub001036_groupi_n_454);
  or csa_tree_sub001036_groupi_g5512__8428(csa_tree_sub001036_groupi_n_513 ,csa_tree_sub001036_groupi_n_191 ,csa_tree_sub001036_groupi_n_451);
  or csa_tree_sub001036_groupi_g5513__5526(csa_tree_sub001036_groupi_n_511 ,csa_tree_sub001036_groupi_n_288 ,csa_tree_sub001036_groupi_n_419);
  or csa_tree_sub001036_groupi_g5514__6783(csa_tree_sub001036_groupi_n_510 ,csa_tree_sub001036_groupi_n_207 ,csa_tree_sub001036_groupi_n_432);
  or csa_tree_sub001036_groupi_g5515__3680(csa_tree_sub001036_groupi_n_509 ,csa_tree_sub001036_groupi_n_192 ,csa_tree_sub001036_groupi_n_421);
  or csa_tree_sub001036_groupi_g5516__1617(csa_tree_sub001036_groupi_n_507 ,csa_tree_sub001036_groupi_n_277 ,csa_tree_sub001036_groupi_n_450);
  or csa_tree_sub001036_groupi_g5517__2802(csa_tree_sub001036_groupi_n_505 ,csa_tree_sub001036_groupi_n_189 ,csa_tree_sub001036_groupi_n_444);
  not csa_tree_sub001036_groupi_g5518(csa_tree_sub001036_groupi_n_494 ,csa_tree_sub001036_groupi_n_493);
  not csa_tree_sub001036_groupi_g5519(csa_tree_sub001036_groupi_n_492 ,csa_tree_sub001036_groupi_n_491);
  not csa_tree_sub001036_groupi_g5520(csa_tree_sub001036_groupi_n_483 ,csa_tree_sub001036_groupi_n_484);
  not csa_tree_sub001036_groupi_g5521(csa_tree_sub001036_groupi_n_479 ,csa_tree_sub001036_groupi_n_480);
  not csa_tree_sub001036_groupi_g5522(csa_tree_sub001036_groupi_n_473 ,csa_tree_sub001036_groupi_n_472);
  not csa_tree_sub001036_groupi_g5523(csa_tree_sub001036_groupi_n_470 ,csa_tree_sub001036_groupi_n_471);
  not csa_tree_sub001036_groupi_g5524(csa_tree_sub001036_groupi_n_465 ,csa_tree_sub001036_groupi_n_464);
  not csa_tree_sub001036_groupi_g5525(csa_tree_sub001036_groupi_n_462 ,csa_tree_sub001036_groupi_n_463);
  or csa_tree_sub001036_groupi_g5526__1705(csa_tree_sub001036_groupi_n_459 ,csa_tree_sub001036_groupi_n_290 ,csa_tree_sub001036_groupi_n_392);
  or csa_tree_sub001036_groupi_g5527__5122(csa_tree_sub001036_groupi_n_458 ,csa_tree_sub001036_groupi_n_255 ,csa_tree_sub001036_groupi_n_390);
  and csa_tree_sub001036_groupi_g5528__8246(csa_tree_sub001036_groupi_n_499 ,csa_tree_sub001036_groupi_n_230 ,csa_tree_sub001036_groupi_n_414);
  and csa_tree_sub001036_groupi_g5529__7098(csa_tree_sub001036_groupi_n_498 ,csa_tree_sub001036_groupi_n_309 ,csa_tree_sub001036_groupi_n_403);
  or csa_tree_sub001036_groupi_g5530__6131(csa_tree_sub001036_groupi_n_497 ,csa_tree_sub001036_groupi_n_250 ,csa_tree_sub001036_groupi_n_416);
  and csa_tree_sub001036_groupi_g5531__1881(csa_tree_sub001036_groupi_n_496 ,csa_tree_sub001036_groupi_n_283 ,csa_tree_sub001036_groupi_n_411);
  or csa_tree_sub001036_groupi_g5532__5115(csa_tree_sub001036_groupi_n_495 ,csa_tree_sub001036_groupi_n_214 ,csa_tree_sub001036_groupi_n_439);
  or csa_tree_sub001036_groupi_g5533__7482(csa_tree_sub001036_groupi_n_493 ,csa_tree_sub001036_groupi_n_284 ,csa_tree_sub001036_groupi_n_425);
  or csa_tree_sub001036_groupi_g5534__4733(csa_tree_sub001036_groupi_n_491 ,csa_tree_sub001036_groupi_n_232 ,csa_tree_sub001036_groupi_n_453);
  or csa_tree_sub001036_groupi_g5535__6161(csa_tree_sub001036_groupi_n_490 ,csa_tree_sub001036_groupi_n_297 ,csa_tree_sub001036_groupi_n_427);
  and csa_tree_sub001036_groupi_g5536__9315(csa_tree_sub001036_groupi_n_489 ,csa_tree_sub001036_groupi_n_202 ,csa_tree_sub001036_groupi_n_400);
  and csa_tree_sub001036_groupi_g5537__9945(csa_tree_sub001036_groupi_n_488 ,csa_tree_sub001036_groupi_n_287 ,csa_tree_sub001036_groupi_n_452);
  and csa_tree_sub001036_groupi_g5538__2883(csa_tree_sub001036_groupi_n_487 ,csa_tree_sub001036_groupi_n_266 ,csa_tree_sub001036_groupi_n_409);
  or csa_tree_sub001036_groupi_g5539__2346(csa_tree_sub001036_groupi_n_486 ,csa_tree_sub001036_groupi_n_220 ,csa_tree_sub001036_groupi_n_448);
  or csa_tree_sub001036_groupi_g5540__1666(csa_tree_sub001036_groupi_n_485 ,csa_tree_sub001036_groupi_n_228 ,csa_tree_sub001036_groupi_n_430);
  or csa_tree_sub001036_groupi_g5541__7410(csa_tree_sub001036_groupi_n_484 ,csa_tree_sub001036_groupi_n_201 ,csa_tree_sub001036_groupi_n_431);
  or csa_tree_sub001036_groupi_g5542__6417(csa_tree_sub001036_groupi_n_482 ,csa_tree_sub001036_groupi_n_322 ,csa_tree_sub001036_groupi_n_408);
  or csa_tree_sub001036_groupi_g5543__5477(csa_tree_sub001036_groupi_n_481 ,csa_tree_sub001036_groupi_n_296 ,csa_tree_sub001036_groupi_n_394);
  or csa_tree_sub001036_groupi_g5544__2398(csa_tree_sub001036_groupi_n_480 ,csa_tree_sub001036_groupi_n_209 ,csa_tree_sub001036_groupi_n_415);
  or csa_tree_sub001036_groupi_g5545__5107(csa_tree_sub001036_groupi_n_478 ,csa_tree_sub001036_groupi_n_289 ,csa_tree_sub001036_groupi_n_412);
  or csa_tree_sub001036_groupi_g5546__6260(csa_tree_sub001036_groupi_n_477 ,csa_tree_sub001036_groupi_n_280 ,csa_tree_sub001036_groupi_n_420);
  or csa_tree_sub001036_groupi_g5547__4319(csa_tree_sub001036_groupi_n_476 ,csa_tree_sub001036_groupi_n_188 ,csa_tree_sub001036_groupi_n_422);
  or csa_tree_sub001036_groupi_g5548__8428(csa_tree_sub001036_groupi_n_475 ,csa_tree_sub001036_groupi_n_306 ,csa_tree_sub001036_groupi_n_397);
  or csa_tree_sub001036_groupi_g5549__5526(csa_tree_sub001036_groupi_n_474 ,csa_tree_sub001036_groupi_n_237 ,csa_tree_sub001036_groupi_n_437);
  and csa_tree_sub001036_groupi_g5550__6783(csa_tree_sub001036_groupi_n_472 ,csa_tree_sub001036_groupi_n_215 ,csa_tree_sub001036_groupi_n_402);
  or csa_tree_sub001036_groupi_g5551__3680(csa_tree_sub001036_groupi_n_471 ,csa_tree_sub001036_groupi_n_211 ,csa_tree_sub001036_groupi_n_410);
  or csa_tree_sub001036_groupi_g5552__1617(csa_tree_sub001036_groupi_n_469 ,csa_tree_sub001036_groupi_n_319 ,csa_tree_sub001036_groupi_n_417);
  and csa_tree_sub001036_groupi_g5553__2802(csa_tree_sub001036_groupi_n_468 ,csa_tree_sub001036_groupi_n_301 ,csa_tree_sub001036_groupi_n_401);
  or csa_tree_sub001036_groupi_g5554__1705(csa_tree_sub001036_groupi_n_467 ,csa_tree_sub001036_groupi_n_190 ,csa_tree_sub001036_groupi_n_404);
  or csa_tree_sub001036_groupi_g5555__5122(csa_tree_sub001036_groupi_n_466 ,csa_tree_sub001036_groupi_n_308 ,csa_tree_sub001036_groupi_n_395);
  or csa_tree_sub001036_groupi_g5556__8246(csa_tree_sub001036_groupi_n_464 ,csa_tree_sub001036_groupi_n_324 ,csa_tree_sub001036_groupi_n_399);
  or csa_tree_sub001036_groupi_g5557__7098(csa_tree_sub001036_groupi_n_463 ,csa_tree_sub001036_groupi_n_223 ,csa_tree_sub001036_groupi_n_424);
  or csa_tree_sub001036_groupi_g5558__6131(csa_tree_sub001036_groupi_n_461 ,csa_tree_sub001036_groupi_n_222 ,csa_tree_sub001036_groupi_n_423);
  or csa_tree_sub001036_groupi_g5559__1881(csa_tree_sub001036_groupi_n_460 ,csa_tree_sub001036_groupi_n_307 ,csa_tree_sub001036_groupi_n_398);
  and csa_tree_sub001036_groupi_g5560__5115(csa_tree_sub001036_groupi_n_455 ,in26[6] ,csa_tree_sub001036_groupi_n_226);
  and csa_tree_sub001036_groupi_g5561__7482(csa_tree_sub001036_groupi_n_454 ,in9[0] ,csa_tree_sub001036_groupi_n_251);
  and csa_tree_sub001036_groupi_g5562__4733(csa_tree_sub001036_groupi_n_453 ,in18[4] ,csa_tree_sub001036_groupi_n_282);
  or csa_tree_sub001036_groupi_g5563__6161(csa_tree_sub001036_groupi_n_452 ,csa_tree_sub001036_groupi_n_182 ,csa_tree_sub001036_groupi_n_210);
  and csa_tree_sub001036_groupi_g5564__9315(csa_tree_sub001036_groupi_n_451 ,in31[3] ,csa_tree_sub001036_groupi_n_294);
  and csa_tree_sub001036_groupi_g5565__9945(csa_tree_sub001036_groupi_n_450 ,in17[4] ,csa_tree_sub001036_groupi_n_249);
  and csa_tree_sub001036_groupi_g5566__2883(csa_tree_sub001036_groupi_n_449 ,in15[3] ,csa_tree_sub001036_groupi_n_278);
  and csa_tree_sub001036_groupi_g5567__2346(csa_tree_sub001036_groupi_n_448 ,csa_tree_sub001036_groupi_n_73 ,csa_tree_sub001036_groupi_n_225);
  and csa_tree_sub001036_groupi_g5568__1666(csa_tree_sub001036_groupi_n_447 ,in12[4] ,csa_tree_sub001036_groupi_n_281);
  and csa_tree_sub001036_groupi_g5569__7410(csa_tree_sub001036_groupi_n_446 ,csa_tree_sub001036_groupi_n_35 ,csa_tree_sub001036_groupi_n_318);
  and csa_tree_sub001036_groupi_g5570__6417(csa_tree_sub001036_groupi_n_445 ,in29[3] ,csa_tree_sub001036_groupi_n_274);
  and csa_tree_sub001036_groupi_g5571__5477(csa_tree_sub001036_groupi_n_444 ,in23[6] ,csa_tree_sub001036_groupi_n_199);
  and csa_tree_sub001036_groupi_g5572__2398(csa_tree_sub001036_groupi_n_443 ,in11[2] ,csa_tree_sub001036_groupi_n_208);
  and csa_tree_sub001036_groupi_g5573__5107(csa_tree_sub001036_groupi_n_442 ,in14[3] ,csa_tree_sub001036_groupi_n_197);
  or csa_tree_sub001036_groupi_g5574__6260(csa_tree_sub001036_groupi_n_441 ,csa_tree_sub001036_groupi_n_170 ,csa_tree_sub001036_groupi_n_293);
  and csa_tree_sub001036_groupi_g5575__4319(csa_tree_sub001036_groupi_n_440 ,in27[4] ,csa_tree_sub001036_groupi_n_272);
  and csa_tree_sub001036_groupi_g5576__8428(csa_tree_sub001036_groupi_n_439 ,in15[2] ,csa_tree_sub001036_groupi_n_240);
  and csa_tree_sub001036_groupi_g5577__5526(csa_tree_sub001036_groupi_n_438 ,in8[2] ,csa_tree_sub001036_groupi_n_279);
  and csa_tree_sub001036_groupi_g5578__6783(csa_tree_sub001036_groupi_n_437 ,in9[6] ,csa_tree_sub001036_groupi_n_275);
  or csa_tree_sub001036_groupi_g5579__3680(csa_tree_sub001036_groupi_n_436 ,csa_tree_sub001036_groupi_n_183 ,csa_tree_sub001036_groupi_n_245);
  and csa_tree_sub001036_groupi_g5580__1617(csa_tree_sub001036_groupi_n_435 ,in12[2] ,csa_tree_sub001036_groupi_n_270);
  or csa_tree_sub001036_groupi_g5581__2802(csa_tree_sub001036_groupi_n_434 ,csa_tree_sub001036_groupi_n_169 ,csa_tree_sub001036_groupi_n_291);
  and csa_tree_sub001036_groupi_g5582__1705(csa_tree_sub001036_groupi_n_433 ,in14[2] ,csa_tree_sub001036_groupi_n_233);
  and csa_tree_sub001036_groupi_g5583__5122(csa_tree_sub001036_groupi_n_432 ,in9[2] ,csa_tree_sub001036_groupi_n_298);
  and csa_tree_sub001036_groupi_g5584__8246(csa_tree_sub001036_groupi_n_431 ,in11[6] ,csa_tree_sub001036_groupi_n_268);
  and csa_tree_sub001036_groupi_g5585__7098(csa_tree_sub001036_groupi_n_430 ,in29[4] ,csa_tree_sub001036_groupi_n_242);
  and csa_tree_sub001036_groupi_g5586__6131(csa_tree_sub001036_groupi_n_429 ,in13[3] ,csa_tree_sub001036_groupi_n_205);
  and csa_tree_sub001036_groupi_g5587__1881(csa_tree_sub001036_groupi_n_428 ,in28[6] ,csa_tree_sub001036_groupi_n_234);
  and csa_tree_sub001036_groupi_g5588__5115(csa_tree_sub001036_groupi_n_427 ,in25[0] ,csa_tree_sub001036_groupi_n_285);
  and csa_tree_sub001036_groupi_g5589__7482(csa_tree_sub001036_groupi_n_426 ,in11[0] ,csa_tree_sub001036_groupi_n_261);
  and csa_tree_sub001036_groupi_g5590__4733(csa_tree_sub001036_groupi_n_425 ,in15[1] ,csa_tree_sub001036_groupi_n_212);
  and csa_tree_sub001036_groupi_g5591__6161(csa_tree_sub001036_groupi_n_424 ,in26[5] ,csa_tree_sub001036_groupi_n_227);
  and csa_tree_sub001036_groupi_g5592(csa_tree_sub001036_groupi_n_423 ,in7[6] ,csa_tree_sub001036_groupi_n_221);
  and csa_tree_sub001036_groupi_g5593(csa_tree_sub001036_groupi_n_422 ,in24[0] ,csa_tree_sub001036_groupi_n_203);
  and csa_tree_sub001036_groupi_g5594(csa_tree_sub001036_groupi_n_421 ,in27[2] ,csa_tree_sub001036_groupi_n_260);
  and csa_tree_sub001036_groupi_g5595(csa_tree_sub001036_groupi_n_420 ,in27[0] ,csa_tree_sub001036_groupi_n_198);
  and csa_tree_sub001036_groupi_g5596(csa_tree_sub001036_groupi_n_419 ,in16[5] ,csa_tree_sub001036_groupi_n_248);
  and csa_tree_sub001036_groupi_g5597(csa_tree_sub001036_groupi_n_418 ,in24[1] ,csa_tree_sub001036_groupi_n_231);
  and csa_tree_sub001036_groupi_g5598(csa_tree_sub001036_groupi_n_417 ,in10[4] ,csa_tree_sub001036_groupi_n_317);
  and csa_tree_sub001036_groupi_g5599(csa_tree_sub001036_groupi_n_416 ,in9[1] ,csa_tree_sub001036_groupi_n_264);
  and csa_tree_sub001036_groupi_g5600(csa_tree_sub001036_groupi_n_415 ,in13[1] ,csa_tree_sub001036_groupi_n_271);
  or csa_tree_sub001036_groupi_g5601(csa_tree_sub001036_groupi_n_414 ,csa_tree_sub001036_groupi_n_180 ,csa_tree_sub001036_groupi_n_267);
  and csa_tree_sub001036_groupi_g5602(csa_tree_sub001036_groupi_n_413 ,in14[6] ,csa_tree_sub001036_groupi_n_194);
  and csa_tree_sub001036_groupi_g5603(csa_tree_sub001036_groupi_n_412 ,csa_tree_sub001036_groupi_n_105 ,csa_tree_sub001036_groupi_n_321);
  or csa_tree_sub001036_groupi_g5604(csa_tree_sub001036_groupi_n_411 ,csa_tree_sub001036_groupi_n_168 ,csa_tree_sub001036_groupi_n_195);
  and csa_tree_sub001036_groupi_g5605(csa_tree_sub001036_groupi_n_410 ,in9[3] ,csa_tree_sub001036_groupi_n_204);
  or csa_tree_sub001036_groupi_g5606(csa_tree_sub001036_groupi_n_409 ,csa_tree_sub001036_groupi_n_179 ,csa_tree_sub001036_groupi_n_236);
  and csa_tree_sub001036_groupi_g5607(csa_tree_sub001036_groupi_n_408 ,in15[5] ,csa_tree_sub001036_groupi_n_246);
  or csa_tree_sub001036_groupi_g5608(csa_tree_sub001036_groupi_n_407 ,csa_tree_sub001036_groupi_n_18 ,csa_tree_sub001036_groupi_n_311);
  or csa_tree_sub001036_groupi_g5609(csa_tree_sub001036_groupi_n_406 ,csa_tree_sub001036_groupi_n_78 ,csa_tree_sub001036_groupi_n_229);
  and csa_tree_sub001036_groupi_g5610(csa_tree_sub001036_groupi_n_405 ,csa_tree_sub001036_groupi_n_20 ,csa_tree_sub001036_groupi_n_303);
  and csa_tree_sub001036_groupi_g5611(csa_tree_sub001036_groupi_n_404 ,csa_tree_sub001036_groupi_n_60 ,csa_tree_sub001036_groupi_n_224);
  or csa_tree_sub001036_groupi_g5612(csa_tree_sub001036_groupi_n_403 ,csa_tree_sub001036_groupi_n_258 ,csa_tree_sub001036_groupi_n_305);
  or csa_tree_sub001036_groupi_g5613(csa_tree_sub001036_groupi_n_402 ,csa_tree_sub001036_groupi_n_72 ,csa_tree_sub001036_groupi_n_235);
  or csa_tree_sub001036_groupi_g5614(csa_tree_sub001036_groupi_n_401 ,csa_tree_sub001036_groupi_n_39 ,csa_tree_sub001036_groupi_n_310);
  or csa_tree_sub001036_groupi_g5615(csa_tree_sub001036_groupi_n_400 ,csa_tree_sub001036_groupi_n_165 ,csa_tree_sub001036_groupi_n_262);
  nor csa_tree_sub001036_groupi_g5616(csa_tree_sub001036_groupi_n_399 ,csa_tree_sub001036_groupi_n_82 ,csa_tree_sub001036_groupi_n_325);
  and csa_tree_sub001036_groupi_g5617(csa_tree_sub001036_groupi_n_398 ,csa_tree_sub001036_groupi_n_14 ,csa_tree_sub001036_groupi_n_300);
  and csa_tree_sub001036_groupi_g5618(csa_tree_sub001036_groupi_n_397 ,csa_tree_sub001036_groupi_n_75 ,csa_tree_sub001036_groupi_n_312);
  nor csa_tree_sub001036_groupi_g5619(csa_tree_sub001036_groupi_n_396 ,csa_tree_sub001036_groupi_n_175 ,csa_tree_sub001036_groupi_n_324);
  and csa_tree_sub001036_groupi_g5620(csa_tree_sub001036_groupi_n_395 ,csa_tree_sub001036_groupi_n_13 ,csa_tree_sub001036_groupi_n_299);
  and csa_tree_sub001036_groupi_g5621(csa_tree_sub001036_groupi_n_394 ,in13[5] ,csa_tree_sub001036_groupi_n_206);
  xnor csa_tree_sub001036_groupi_g5622(csa_tree_sub001036_groupi_n_393 ,csa_tree_sub001036_groupi_n_17 ,csa_tree_sub001036_groupi_n_79);
  or csa_tree_sub001036_groupi_g5623(csa_tree_sub001036_groupi_n_457 ,csa_tree_sub001036_groupi_n_269 ,csa_tree_sub001036_groupi_n_253);
  or csa_tree_sub001036_groupi_g5624(csa_tree_sub001036_groupi_n_456 ,csa_tree_sub001036_groupi_n_244 ,csa_tree_sub001036_groupi_n_323);
  not csa_tree_sub001036_groupi_g5625(csa_tree_sub001036_groupi_n_390 ,csa_tree_sub001036_groupi_n_391);
  xnor csa_tree_sub001036_groupi_g5626(csa_tree_sub001036_groupi_n_388 ,csa_tree_sub001036_groupi_n_13 ,csa_tree_sub001036_groupi_n_123);
  xnor csa_tree_sub001036_groupi_g5627(csa_tree_sub001036_groupi_n_387 ,csa_tree_sub001036_groupi_n_67 ,csa_tree_sub001036_groupi_n_79);
  xnor csa_tree_sub001036_groupi_g5628(csa_tree_sub001036_groupi_n_386 ,csa_tree_sub001036_groupi_n_28 ,csa_tree_sub001036_groupi_n_81);
  xnor csa_tree_sub001036_groupi_g5629(csa_tree_sub001036_groupi_n_385 ,csa_tree_sub001036_groupi_n_22 ,csa_tree_sub001036_groupi_n_41);
  xnor csa_tree_sub001036_groupi_g5630(csa_tree_sub001036_groupi_n_384 ,csa_tree_sub001036_groupi_n_96 ,csa_tree_sub001036_groupi_n_70);
  xnor csa_tree_sub001036_groupi_g5631(csa_tree_sub001036_groupi_n_383 ,csa_tree_sub001036_groupi_n_14 ,csa_tree_sub001036_groupi_n_115);
  xnor csa_tree_sub001036_groupi_g5632(csa_tree_sub001036_groupi_n_382 ,csa_tree_sub001036_groupi_n_32 ,csa_tree_sub001036_groupi_n_73);
  xnor csa_tree_sub001036_groupi_g5633(csa_tree_sub001036_groupi_n_381 ,csa_tree_sub001036_groupi_n_81 ,csa_tree_sub001036_groupi_n_67);
  xnor csa_tree_sub001036_groupi_g5634(csa_tree_sub001036_groupi_n_380 ,csa_tree_sub001036_groupi_n_69 ,in10[1]);
  xnor csa_tree_sub001036_groupi_g5635(csa_tree_sub001036_groupi_n_379 ,csa_tree_sub001036_groupi_n_64 ,in12[0]);
  xnor csa_tree_sub001036_groupi_g5636(csa_tree_sub001036_groupi_n_378 ,csa_tree_sub001036_groupi_n_17 ,csa_tree_sub001036_groupi_n_126);
  xnor csa_tree_sub001036_groupi_g5637(csa_tree_sub001036_groupi_n_377 ,csa_tree_sub001036_groupi_n_93 ,csa_tree_sub001036_groupi_n_129);
  xnor csa_tree_sub001036_groupi_g5638(csa_tree_sub001036_groupi_n_376 ,csa_tree_sub001036_groupi_n_12 ,csa_tree_sub001036_groupi_n_87);
  xnor csa_tree_sub001036_groupi_g5639(csa_tree_sub001036_groupi_n_375 ,csa_tree_sub001036_groupi_n_30 ,csa_tree_sub001036_groupi_n_64);
  xnor csa_tree_sub001036_groupi_g5640(csa_tree_sub001036_groupi_n_374 ,csa_tree_sub001036_groupi_n_34 ,csa_tree_sub001036_groupi_n_115);
  xnor csa_tree_sub001036_groupi_g5641(csa_tree_sub001036_groupi_n_373 ,csa_tree_sub001036_groupi_n_12 ,csa_tree_sub001036_groupi_n_136);
  xnor csa_tree_sub001036_groupi_g5642(csa_tree_sub001036_groupi_n_372 ,csa_tree_sub001036_groupi_n_20 ,csa_tree_sub001036_groupi_n_120);
  xnor csa_tree_sub001036_groupi_g5643(csa_tree_sub001036_groupi_n_371 ,in25[2] ,in29[2]);
  xnor csa_tree_sub001036_groupi_g5644(csa_tree_sub001036_groupi_n_370 ,in26[3] ,in29[3]);
  xnor csa_tree_sub001036_groupi_g5645(csa_tree_sub001036_groupi_n_369 ,in27[1] ,in12[2]);
  xnor csa_tree_sub001036_groupi_g5646(csa_tree_sub001036_groupi_n_368 ,in23[1] ,in24[1]);
  xnor csa_tree_sub001036_groupi_g5647(csa_tree_sub001036_groupi_n_367 ,in17[4] ,in11[4]);
  xnor csa_tree_sub001036_groupi_g5648(csa_tree_sub001036_groupi_n_366 ,in9[6] ,in24[5]);
  xnor csa_tree_sub001036_groupi_g5649(csa_tree_sub001036_groupi_n_365 ,in23[4] ,in24[4]);
  xnor csa_tree_sub001036_groupi_g5650(csa_tree_sub001036_groupi_n_364 ,in7[6] ,in10[6]);
  xnor csa_tree_sub001036_groupi_g5651(csa_tree_sub001036_groupi_n_363 ,in27[6] ,in28[6]);
  xnor csa_tree_sub001036_groupi_g5652(csa_tree_sub001036_groupi_n_362 ,in18[1] ,in7[1]);
  xnor csa_tree_sub001036_groupi_g5653(csa_tree_sub001036_groupi_n_361 ,in13[6] ,in15[6]);
  xnor csa_tree_sub001036_groupi_g5654(csa_tree_sub001036_groupi_n_360 ,in9[2] ,in18[2]);
  xnor csa_tree_sub001036_groupi_g5655(csa_tree_sub001036_groupi_n_359 ,in23[2] ,in24[2]);
  xnor csa_tree_sub001036_groupi_g5656(csa_tree_sub001036_groupi_n_358 ,in9[3] ,in18[3]);
  xnor csa_tree_sub001036_groupi_g5657(csa_tree_sub001036_groupi_n_357 ,in17[3] ,in13[3]);
  xnor csa_tree_sub001036_groupi_g5658(csa_tree_sub001036_groupi_n_356 ,in17[2] ,in13[2]);
  xnor csa_tree_sub001036_groupi_g5659(csa_tree_sub001036_groupi_n_355 ,in17[1] ,in11[1]);
  xnor csa_tree_sub001036_groupi_g5660(csa_tree_sub001036_groupi_n_354 ,in26[0] ,in29[0]);
  xnor csa_tree_sub001036_groupi_g5661(csa_tree_sub001036_groupi_n_353 ,in14[2] ,in16[2]);
  xnor csa_tree_sub001036_groupi_g5662(csa_tree_sub001036_groupi_n_352 ,in27[4] ,in12[5]);
  xnor csa_tree_sub001036_groupi_g5663(csa_tree_sub001036_groupi_n_351 ,in23[6] ,in31[6]);
  xnor csa_tree_sub001036_groupi_g5664(csa_tree_sub001036_groupi_n_350 ,in31[1] ,in15[2]);
  xnor csa_tree_sub001036_groupi_g5665(csa_tree_sub001036_groupi_n_349 ,in18[4] ,in7[4]);
  xnor csa_tree_sub001036_groupi_g5666(csa_tree_sub001036_groupi_n_348 ,in27[2] ,in12[3]);
  xnor csa_tree_sub001036_groupi_g5667(csa_tree_sub001036_groupi_n_347 ,in31[2] ,in15[3]);
  xnor csa_tree_sub001036_groupi_g5668(csa_tree_sub001036_groupi_n_346 ,in25[1] ,in29[1]);
  xnor csa_tree_sub001036_groupi_g5669(csa_tree_sub001036_groupi_n_345 ,in24[3] ,in10[4]);
  xnor csa_tree_sub001036_groupi_g5670(csa_tree_sub001036_groupi_n_344 ,in14[6] ,in16[6]);
  xnor csa_tree_sub001036_groupi_g5671(csa_tree_sub001036_groupi_n_343 ,in17[5] ,in13[5]);
  xnor csa_tree_sub001036_groupi_g5672(csa_tree_sub001036_groupi_n_342 ,in28[3] ,in12[4]);
  xnor csa_tree_sub001036_groupi_g5673(csa_tree_sub001036_groupi_n_341 ,in25[5] ,in29[5]);
  xnor csa_tree_sub001036_groupi_g5674(csa_tree_sub001036_groupi_n_340 ,in9[5] ,in18[5]);
  xnor csa_tree_sub001036_groupi_g5675(csa_tree_sub001036_groupi_n_339 ,in31[0] ,in8[1]);
  xnor csa_tree_sub001036_groupi_g5676(csa_tree_sub001036_groupi_n_338 ,in30[5] ,in11[6]);
  xnor csa_tree_sub001036_groupi_g5677(csa_tree_sub001036_groupi_n_337 ,in25[4] ,in29[4]);
  xnor csa_tree_sub001036_groupi_g5678(csa_tree_sub001036_groupi_n_336 ,in31[4] ,in15[5]);
  xnor csa_tree_sub001036_groupi_g5679(csa_tree_sub001036_groupi_n_335 ,in14[5] ,in16[5]);
  xnor csa_tree_sub001036_groupi_g5680(csa_tree_sub001036_groupi_n_334 ,in8[0] ,in13[0]);
  xnor csa_tree_sub001036_groupi_g5681(csa_tree_sub001036_groupi_n_333 ,in23[0] ,in30[0]);
  xnor csa_tree_sub001036_groupi_g5682(csa_tree_sub001036_groupi_n_332 ,in28[0] ,in12[1]);
  xnor csa_tree_sub001036_groupi_g5683(csa_tree_sub001036_groupi_n_331 ,in25[6] ,in26[6]);
  xnor csa_tree_sub001036_groupi_g5684(csa_tree_sub001036_groupi_n_330 ,in31[3] ,in8[4]);
  xnor csa_tree_sub001036_groupi_g5685(csa_tree_sub001036_groupi_n_329 ,in31[5] ,in17[6]);
  xnor csa_tree_sub001036_groupi_g5686(csa_tree_sub001036_groupi_n_328 ,in7[0] ,in15[0]);
  xnor csa_tree_sub001036_groupi_g5687(csa_tree_sub001036_groupi_n_327 ,in17[0] ,in18[0]);
  xnor csa_tree_sub001036_groupi_g5688(csa_tree_sub001036_groupi_n_326 ,in14[3] ,in16[3]);
  xnor csa_tree_sub001036_groupi_g5689(csa_tree_sub001036_groupi_n_392 ,csa_tree_sub001036_groupi_n_61 ,csa_tree_sub001036_groupi_n_75);
  xnor csa_tree_sub001036_groupi_g5690(csa_tree_sub001036_groupi_n_391 ,in14[0] ,in16[0]);
  xnor csa_tree_sub001036_groupi_g5691(csa_tree_sub001036_groupi_n_389 ,in14[4] ,in16[4]);
  and csa_tree_sub001036_groupi_g5693(csa_tree_sub001036_groupi_n_322 ,in31[4] ,in7[5]);
  or csa_tree_sub001036_groupi_g5694(csa_tree_sub001036_groupi_n_321 ,csa_tree_sub001036_groupi_n_53 ,in12[0]);
  and csa_tree_sub001036_groupi_g5695(csa_tree_sub001036_groupi_n_320 ,in10[1] ,csa_tree_sub001036_groupi_n_55);
  and csa_tree_sub001036_groupi_g5696(csa_tree_sub001036_groupi_n_319 ,in24[3] ,csa_tree_sub001036_groupi_n_173);
  or csa_tree_sub001036_groupi_g5697(csa_tree_sub001036_groupi_n_318 ,csa_tree_sub001036_groupi_n_55 ,in10[1]);
  or csa_tree_sub001036_groupi_g5698(csa_tree_sub001036_groupi_n_317 ,csa_tree_sub001036_groupi_n_51 ,in24[3]);
  or csa_tree_sub001036_groupi_g5699(csa_tree_sub001036_groupi_n_316 ,csa_tree_sub001036_groupi_n_153 ,csa_tree_sub001036_groupi_n_18);
  nor csa_tree_sub001036_groupi_g5700(csa_tree_sub001036_groupi_n_315 ,csa_tree_sub001036_groupi_n_172 ,csa_tree_sub001036_groupi_n_96);
  nor csa_tree_sub001036_groupi_g5701(csa_tree_sub001036_groupi_n_314 ,csa_tree_sub001036_groupi_n_149 ,csa_tree_sub001036_groupi_n_93);
  or csa_tree_sub001036_groupi_g5702(csa_tree_sub001036_groupi_n_313 ,csa_tree_sub001036_groupi_n_150 ,csa_tree_sub001036_groupi_n_70);
  or csa_tree_sub001036_groupi_g5703(csa_tree_sub001036_groupi_n_312 ,csa_tree_sub001036_groupi_n_161 ,csa_tree_sub001036_groupi_n_15);
  nor csa_tree_sub001036_groupi_g5704(csa_tree_sub001036_groupi_n_311 ,csa_tree_sub001036_groupi_n_162 ,csa_tree_sub001036_groupi_n_111);
  nor csa_tree_sub001036_groupi_g5705(csa_tree_sub001036_groupi_n_310 ,csa_tree_sub001036_groupi_n_157 ,csa_tree_sub001036_groupi_n_126);
  or csa_tree_sub001036_groupi_g5706(csa_tree_sub001036_groupi_n_309 ,csa_tree_sub001036_groupi_n_51 ,csa_tree_sub001036_groupi_n_132);
  nor csa_tree_sub001036_groupi_g5707(csa_tree_sub001036_groupi_n_308 ,csa_tree_sub001036_groupi_n_162 ,csa_tree_sub001036_groupi_n_123);
  nor csa_tree_sub001036_groupi_g5708(csa_tree_sub001036_groupi_n_307 ,csa_tree_sub001036_groupi_n_158 ,csa_tree_sub001036_groupi_n_129);
  nor csa_tree_sub001036_groupi_g5709(csa_tree_sub001036_groupi_n_306 ,csa_tree_sub001036_groupi_n_146 ,csa_tree_sub001036_groupi_n_41);
  nor csa_tree_sub001036_groupi_g5710(csa_tree_sub001036_groupi_n_305 ,csa_tree_sub001036_groupi_n_152 ,csa_tree_sub001036_groupi_n_87);
  or csa_tree_sub001036_groupi_g5711(csa_tree_sub001036_groupi_n_304 ,csa_tree_sub001036_groupi_n_163 ,csa_tree_sub001036_groupi_n_34);
  or csa_tree_sub001036_groupi_g5712(csa_tree_sub001036_groupi_n_303 ,csa_tree_sub001036_groupi_n_163 ,csa_tree_sub001036_groupi_n_63);
  nor csa_tree_sub001036_groupi_g5713(csa_tree_sub001036_groupi_n_302 ,csa_tree_sub001036_groupi_n_160 ,csa_tree_sub001036_groupi_n_30);
  or csa_tree_sub001036_groupi_g5714(csa_tree_sub001036_groupi_n_301 ,csa_tree_sub001036_groupi_n_161 ,csa_tree_sub001036_groupi_n_99);
  or csa_tree_sub001036_groupi_g5715(csa_tree_sub001036_groupi_n_300 ,csa_tree_sub001036_groupi_n_159 ,csa_tree_sub001036_groupi_n_37);
  or csa_tree_sub001036_groupi_g5716(csa_tree_sub001036_groupi_n_299 ,csa_tree_sub001036_groupi_n_158 ,csa_tree_sub001036_groupi_n_102);
  or csa_tree_sub001036_groupi_g5717(csa_tree_sub001036_groupi_n_298 ,in28[1] ,in18[2]);
  and csa_tree_sub001036_groupi_g5718(csa_tree_sub001036_groupi_n_297 ,in26[0] ,in29[0]);
  and csa_tree_sub001036_groupi_g5719(csa_tree_sub001036_groupi_n_296 ,in17[5] ,in8[5]);
  or csa_tree_sub001036_groupi_g5720(csa_tree_sub001036_groupi_n_295 ,csa_tree_sub001036_groupi_n_22 ,csa_tree_sub001036_groupi_n_24);
  or csa_tree_sub001036_groupi_g5721(csa_tree_sub001036_groupi_n_294 ,in8[4] ,in15[4]);
  nor csa_tree_sub001036_groupi_g5722(csa_tree_sub001036_groupi_n_293 ,in29[2] ,in11[3]);
  and csa_tree_sub001036_groupi_g5723(csa_tree_sub001036_groupi_n_292 ,in8[0] ,in13[0]);
  nor csa_tree_sub001036_groupi_g5724(csa_tree_sub001036_groupi_n_291 ,in31[5] ,in18[6]);
  and csa_tree_sub001036_groupi_g5725(csa_tree_sub001036_groupi_n_290 ,csa_tree_sub001036_groupi_n_15 ,csa_tree_sub001036_groupi_n_24);
  and csa_tree_sub001036_groupi_g5726(csa_tree_sub001036_groupi_n_289 ,in12[0] ,csa_tree_sub001036_groupi_n_53);
  and csa_tree_sub001036_groupi_g5727(csa_tree_sub001036_groupi_n_288 ,in26[4] ,in14[5]);
  nand csa_tree_sub001036_groupi_g5728(csa_tree_sub001036_groupi_n_287 ,in23[4] ,in10[5]);
  and csa_tree_sub001036_groupi_g5729(csa_tree_sub001036_groupi_n_286 ,in23[1] ,in10[2]);
  or csa_tree_sub001036_groupi_g5730(csa_tree_sub001036_groupi_n_285 ,in26[0] ,in29[0]);
  and csa_tree_sub001036_groupi_g5731(csa_tree_sub001036_groupi_n_284 ,in31[0] ,in8[1]);
  nand csa_tree_sub001036_groupi_g5732(csa_tree_sub001036_groupi_n_283 ,in17[0] ,in18[0]);
  or csa_tree_sub001036_groupi_g5733(csa_tree_sub001036_groupi_n_282 ,in9[4] ,in7[4]);
  or csa_tree_sub001036_groupi_g5734(csa_tree_sub001036_groupi_n_281 ,in27[3] ,in28[3]);
  and csa_tree_sub001036_groupi_g5735(csa_tree_sub001036_groupi_n_280 ,in28[0] ,in12[1]);
  or csa_tree_sub001036_groupi_g5736(csa_tree_sub001036_groupi_n_279 ,in17[2] ,in13[2]);
  or csa_tree_sub001036_groupi_g5737(csa_tree_sub001036_groupi_n_278 ,in31[2] ,in7[3]);
  and csa_tree_sub001036_groupi_g5738(csa_tree_sub001036_groupi_n_277 ,in11[4] ,in13[4]);
  and csa_tree_sub001036_groupi_g5739(csa_tree_sub001036_groupi_n_276 ,in25[3] ,in26[3]);
  or csa_tree_sub001036_groupi_g5740(csa_tree_sub001036_groupi_n_275 ,in24[5] ,in12[6]);
  or csa_tree_sub001036_groupi_g5741(csa_tree_sub001036_groupi_n_274 ,in25[3] ,in26[3]);
  nand csa_tree_sub001036_groupi_g5742(csa_tree_sub001036_groupi_n_273 ,in29[2] ,in11[3]);
  or csa_tree_sub001036_groupi_g5743(csa_tree_sub001036_groupi_n_272 ,in30[4] ,in12[5]);
  or csa_tree_sub001036_groupi_g5744(csa_tree_sub001036_groupi_n_271 ,in17[1] ,in11[1]);
  or csa_tree_sub001036_groupi_g5745(csa_tree_sub001036_groupi_n_270 ,in27[1] ,in30[1]);
  and csa_tree_sub001036_groupi_g5746(csa_tree_sub001036_groupi_n_269 ,in23[3] ,in30[3]);
  or csa_tree_sub001036_groupi_g5747(csa_tree_sub001036_groupi_n_268 ,in28[5] ,in30[5]);
  nor csa_tree_sub001036_groupi_g5748(csa_tree_sub001036_groupi_n_267 ,in27[5] ,in13[6]);
  nand csa_tree_sub001036_groupi_g5749(csa_tree_sub001036_groupi_n_266 ,in23[2] ,in10[3]);
  nand csa_tree_sub001036_groupi_g5750(csa_tree_sub001036_groupi_n_265 ,in28[4] ,in18[5]);
  or csa_tree_sub001036_groupi_g5751(csa_tree_sub001036_groupi_n_264 ,in18[1] ,in7[1]);
  and csa_tree_sub001036_groupi_g5752(csa_tree_sub001036_groupi_n_263 ,in27[3] ,in28[3]);
  and csa_tree_sub001036_groupi_g5753(csa_tree_sub001036_groupi_n_262 ,csa_tree_sub001036_groupi_n_26 ,csa_tree_sub001036_groupi_n_28);
  or csa_tree_sub001036_groupi_g5754(csa_tree_sub001036_groupi_n_261 ,in7[0] ,in15[0]);
  or csa_tree_sub001036_groupi_g5755(csa_tree_sub001036_groupi_n_260 ,in30[2] ,in12[3]);
  and csa_tree_sub001036_groupi_g5756(csa_tree_sub001036_groupi_n_259 ,in26[1] ,in16[2]);
  and csa_tree_sub001036_groupi_g5757(csa_tree_sub001036_groupi_n_325 ,csa_tree_sub001036_groupi_n_166 ,csa_tree_sub001036_groupi_n_176);
  and csa_tree_sub001036_groupi_g5758(csa_tree_sub001036_groupi_n_324 ,csa_tree_sub001036_groupi_n_84 ,csa_tree_sub001036_groupi_n_66);
  and csa_tree_sub001036_groupi_g5759(csa_tree_sub001036_groupi_n_323 ,csa_tree_sub001036_groupi_n_186 ,csa_tree_sub001036_groupi_n_185);
  not csa_tree_sub001036_groupi_g5760(csa_tree_sub001036_groupi_n_256 ,csa_tree_sub001036_groupi_n_257);
  not csa_tree_sub001036_groupi_g5761(csa_tree_sub001036_groupi_n_254 ,csa_tree_sub001036_groupi_n_255);
  not csa_tree_sub001036_groupi_g5762(csa_tree_sub001036_groupi_n_252 ,csa_tree_sub001036_groupi_n_253);
  or csa_tree_sub001036_groupi_g5763(csa_tree_sub001036_groupi_n_251 ,in8[0] ,in13[0]);
  and csa_tree_sub001036_groupi_g5764(csa_tree_sub001036_groupi_n_250 ,in18[1] ,in7[1]);
  or csa_tree_sub001036_groupi_g5765(csa_tree_sub001036_groupi_n_249 ,in11[4] ,in13[4]);
  or csa_tree_sub001036_groupi_g5766(csa_tree_sub001036_groupi_n_248 ,in26[4] ,in14[5]);
  and csa_tree_sub001036_groupi_g5767(csa_tree_sub001036_groupi_n_247 ,in25[1] ,in29[1]);
  or csa_tree_sub001036_groupi_g5768(csa_tree_sub001036_groupi_n_246 ,in31[4] ,in7[5]);
  nor csa_tree_sub001036_groupi_g5769(csa_tree_sub001036_groupi_n_245 ,in28[4] ,in18[5]);
  nor csa_tree_sub001036_groupi_g5770(csa_tree_sub001036_groupi_n_244 ,csa_tree_sub001036_groupi_n_186 ,csa_tree_sub001036_groupi_n_185);
  and csa_tree_sub001036_groupi_g5771(csa_tree_sub001036_groupi_n_243 ,in27[1] ,in30[1]);
  or csa_tree_sub001036_groupi_g5772(csa_tree_sub001036_groupi_n_242 ,in25[4] ,in11[5]);
  and csa_tree_sub001036_groupi_g5773(csa_tree_sub001036_groupi_n_241 ,in17[3] ,in8[3]);
  or csa_tree_sub001036_groupi_g5774(csa_tree_sub001036_groupi_n_240 ,in31[1] ,in7[2]);
  and csa_tree_sub001036_groupi_g5775(csa_tree_sub001036_groupi_n_239 ,in31[2] ,in7[3]);
  nand csa_tree_sub001036_groupi_g5776(csa_tree_sub001036_groupi_n_238 ,in31[5] ,in18[6]);
  and csa_tree_sub001036_groupi_g5777(csa_tree_sub001036_groupi_n_237 ,in24[5] ,in12[6]);
  nor csa_tree_sub001036_groupi_g5778(csa_tree_sub001036_groupi_n_236 ,in23[2] ,in10[3]);
  nor csa_tree_sub001036_groupi_g5779(csa_tree_sub001036_groupi_n_235 ,csa_tree_sub001036_groupi_n_141 ,csa_tree_sub001036_groupi_n_43);
  or csa_tree_sub001036_groupi_g5780(csa_tree_sub001036_groupi_n_234 ,in27[6] ,in30[6]);
  or csa_tree_sub001036_groupi_g5781(csa_tree_sub001036_groupi_n_233 ,in26[1] ,in16[2]);
  and csa_tree_sub001036_groupi_g5782(csa_tree_sub001036_groupi_n_232 ,in9[4] ,in7[4]);
  or csa_tree_sub001036_groupi_g5783(csa_tree_sub001036_groupi_n_231 ,in23[1] ,in10[2]);
  nand csa_tree_sub001036_groupi_g5784(csa_tree_sub001036_groupi_n_230 ,in27[5] ,in13[6]);
  nor csa_tree_sub001036_groupi_g5785(csa_tree_sub001036_groupi_n_229 ,csa_tree_sub001036_groupi_n_99 ,csa_tree_sub001036_groupi_n_117);
  and csa_tree_sub001036_groupi_g5786(csa_tree_sub001036_groupi_n_228 ,in25[4] ,in11[5]);
  or csa_tree_sub001036_groupi_g5787(csa_tree_sub001036_groupi_n_227 ,in25[5] ,in29[5]);
  or csa_tree_sub001036_groupi_g5788(csa_tree_sub001036_groupi_n_226 ,in24[6] ,in25[6]);
  or csa_tree_sub001036_groupi_g5789(csa_tree_sub001036_groupi_n_225 ,csa_tree_sub001036_groupi_n_9 ,csa_tree_sub001036_groupi_n_135);
  or csa_tree_sub001036_groupi_g5790(csa_tree_sub001036_groupi_n_224 ,csa_tree_sub001036_groupi_n_164 ,csa_tree_sub001036_groupi_n_148);
  and csa_tree_sub001036_groupi_g5791(csa_tree_sub001036_groupi_n_223 ,in25[5] ,in29[5]);
  and csa_tree_sub001036_groupi_g5792(csa_tree_sub001036_groupi_n_222 ,in8[6] ,in10[6]);
  or csa_tree_sub001036_groupi_g5793(csa_tree_sub001036_groupi_n_221 ,in8[6] ,in10[6]);
  and csa_tree_sub001036_groupi_g5794(csa_tree_sub001036_groupi_n_220 ,csa_tree_sub001036_groupi_n_9 ,csa_tree_sub001036_groupi_n_11);
  and csa_tree_sub001036_groupi_g5795(csa_tree_sub001036_groupi_n_219 ,in26[2] ,in16[3]);
  and csa_tree_sub001036_groupi_g5796(csa_tree_sub001036_groupi_n_218 ,in17[2] ,in13[2]);
  and csa_tree_sub001036_groupi_g5797(csa_tree_sub001036_groupi_n_217 ,in7[0] ,in15[0]);
  and csa_tree_sub001036_groupi_g5798(csa_tree_sub001036_groupi_n_216 ,in27[6] ,in30[6]);
  or csa_tree_sub001036_groupi_g5799(csa_tree_sub001036_groupi_n_215 ,csa_tree_sub001036_groupi_n_147 ,csa_tree_sub001036_groupi_n_159);
  and csa_tree_sub001036_groupi_g5800(csa_tree_sub001036_groupi_n_214 ,in31[1] ,in7[2]);
  or csa_tree_sub001036_groupi_g5801(csa_tree_sub001036_groupi_n_213 ,csa_tree_sub001036_groupi_n_157 ,csa_tree_sub001036_groupi_n_151);
  or csa_tree_sub001036_groupi_g5802(csa_tree_sub001036_groupi_n_212 ,in31[0] ,in8[1]);
  and csa_tree_sub001036_groupi_g5803(csa_tree_sub001036_groupi_n_211 ,in28[2] ,in18[3]);
  nor csa_tree_sub001036_groupi_g5804(csa_tree_sub001036_groupi_n_210 ,in23[4] ,in10[5]);
  and csa_tree_sub001036_groupi_g5805(csa_tree_sub001036_groupi_n_209 ,in17[1] ,in11[1]);
  or csa_tree_sub001036_groupi_g5806(csa_tree_sub001036_groupi_n_208 ,in25[1] ,in29[1]);
  and csa_tree_sub001036_groupi_g5807(csa_tree_sub001036_groupi_n_207 ,in28[1] ,in18[2]);
  or csa_tree_sub001036_groupi_g5808(csa_tree_sub001036_groupi_n_206 ,in17[5] ,in8[5]);
  or csa_tree_sub001036_groupi_g5809(csa_tree_sub001036_groupi_n_205 ,in17[3] ,in8[3]);
  or csa_tree_sub001036_groupi_g5810(csa_tree_sub001036_groupi_n_204 ,in28[2] ,in18[3]);
  or csa_tree_sub001036_groupi_g5811(csa_tree_sub001036_groupi_n_203 ,in23[0] ,in30[0]);
  or csa_tree_sub001036_groupi_g5812(csa_tree_sub001036_groupi_n_202 ,csa_tree_sub001036_groupi_n_45 ,csa_tree_sub001036_groupi_n_11);
  and csa_tree_sub001036_groupi_g5813(csa_tree_sub001036_groupi_n_201 ,in28[5] ,in30[5]);
  and csa_tree_sub001036_groupi_g5814(csa_tree_sub001036_groupi_n_200 ,in23[5] ,in16[6]);
  or csa_tree_sub001036_groupi_g5815(csa_tree_sub001036_groupi_n_199 ,in29[6] ,in31[6]);
  or csa_tree_sub001036_groupi_g5816(csa_tree_sub001036_groupi_n_198 ,in28[0] ,in12[1]);
  or csa_tree_sub001036_groupi_g5817(csa_tree_sub001036_groupi_n_197 ,in26[2] ,in16[3]);
  and csa_tree_sub001036_groupi_g5818(csa_tree_sub001036_groupi_n_196 ,in24[6] ,in25[6]);
  nor csa_tree_sub001036_groupi_g5819(csa_tree_sub001036_groupi_n_195 ,in17[0] ,in18[0]);
  or csa_tree_sub001036_groupi_g5820(csa_tree_sub001036_groupi_n_194 ,in23[5] ,in16[6]);
  and csa_tree_sub001036_groupi_g5821(csa_tree_sub001036_groupi_n_193 ,in30[4] ,in12[5]);
  and csa_tree_sub001036_groupi_g5822(csa_tree_sub001036_groupi_n_192 ,in30[2] ,in12[3]);
  and csa_tree_sub001036_groupi_g5823(csa_tree_sub001036_groupi_n_191 ,in8[4] ,in15[4]);
  nor csa_tree_sub001036_groupi_g5824(csa_tree_sub001036_groupi_n_190 ,csa_tree_sub001036_groupi_n_108 ,csa_tree_sub001036_groupi_n_120);
  and csa_tree_sub001036_groupi_g5825(csa_tree_sub001036_groupi_n_189 ,in29[6] ,in31[6]);
  and csa_tree_sub001036_groupi_g5826(csa_tree_sub001036_groupi_n_188 ,in23[0] ,in30[0]);
  or csa_tree_sub001036_groupi_g5827(csa_tree_sub001036_groupi_n_258 ,csa_tree_sub001036_groupi_n_178 ,csa_tree_sub001036_groupi_n_181);
  or csa_tree_sub001036_groupi_g5828(csa_tree_sub001036_groupi_n_257 ,csa_tree_sub001036_groupi_n_177 ,csa_tree_sub001036_groupi_n_184);
  and csa_tree_sub001036_groupi_g5829(csa_tree_sub001036_groupi_n_255 ,csa_tree_sub001036_groupi_n_167 ,csa_tree_sub001036_groupi_n_174);
  and csa_tree_sub001036_groupi_g5830(csa_tree_sub001036_groupi_n_253 ,csa_tree_sub001036_groupi_n_171 ,csa_tree_sub001036_groupi_n_187);
  not csa_tree_sub001036_groupi_g5831(csa_tree_sub001036_groupi_n_187 ,in30[3]);
  not csa_tree_sub001036_groupi_g5832(csa_tree_sub001036_groupi_n_186 ,in14[1]);
  not csa_tree_sub001036_groupi_g5833(csa_tree_sub001036_groupi_n_185 ,in16[1]);
  not csa_tree_sub001036_groupi_g5834(csa_tree_sub001036_groupi_n_184 ,in16[0]);
  not csa_tree_sub001036_groupi_g5835(csa_tree_sub001036_groupi_n_183 ,in9[5]);
  not csa_tree_sub001036_groupi_g5836(csa_tree_sub001036_groupi_n_182 ,in24[4]);
  not csa_tree_sub001036_groupi_g5837(csa_tree_sub001036_groupi_n_181 ,in16[4]);
  not csa_tree_sub001036_groupi_g5838(csa_tree_sub001036_groupi_n_180 ,in15[6]);
  not csa_tree_sub001036_groupi_g5839(csa_tree_sub001036_groupi_n_179 ,in24[2]);
  not csa_tree_sub001036_groupi_g5840(csa_tree_sub001036_groupi_n_178 ,in14[4]);
  not csa_tree_sub001036_groupi_g5841(csa_tree_sub001036_groupi_n_177 ,in14[0]);
  not csa_tree_sub001036_groupi_g5842(csa_tree_sub001036_groupi_n_176 ,csa_tree_sub001036_groupi_n_66);
  not csa_tree_sub001036_groupi_g5843(csa_tree_sub001036_groupi_n_175 ,csa_tree_sub001036_groupi_n_78);
  not csa_tree_sub001036_groupi_g5844(csa_tree_sub001036_groupi_n_174 ,csa_tree_sub001036_groupi_n_76);
  not csa_tree_sub001036_groupi_g5847(csa_tree_sub001036_groupi_n_173 ,csa_tree_sub001036_groupi_n_88);
  not csa_tree_sub001036_groupi_g5848(csa_tree_sub001036_groupi_n_172 ,csa_tree_sub001036_groupi_n_69);
  not csa_tree_sub001036_groupi_g5849(csa_tree_sub001036_groupi_n_171 ,in23[3]);
  not csa_tree_sub001036_groupi_g5850(csa_tree_sub001036_groupi_n_170 ,in25[2]);
  not csa_tree_sub001036_groupi_g5851(csa_tree_sub001036_groupi_n_169 ,in17[6]);
  not csa_tree_sub001036_groupi_g5852(csa_tree_sub001036_groupi_n_168 ,in10[0]);
  not csa_tree_sub001036_groupi_g5853(csa_tree_sub001036_groupi_n_167 ,csa_tree_sub001036_groupi_n_60);
  not csa_tree_sub001036_groupi_g5854(csa_tree_sub001036_groupi_n_166 ,csa_tree_sub001036_groupi_n_85);
  not csa_tree_sub001036_groupi_g5855(csa_tree_sub001036_groupi_n_165 ,csa_tree_sub001036_groupi_n_82);
  not csa_tree_sub001036_groupi_g5859(csa_tree_sub001036_groupi_n_164 ,csa_tree_sub001036_groupi_n_109);
  not csa_tree_sub001036_groupi_g5861(csa_tree_sub001036_groupi_n_163 ,csa_tree_sub001036_groupi_n_112);
  not csa_tree_sub001036_groupi_g5862(csa_tree_sub001036_groupi_n_162 ,csa_tree_sub001036_groupi_n_102);
  not csa_tree_sub001036_groupi_g5863(csa_tree_sub001036_groupi_n_161 ,csa_tree_sub001036_groupi_n_127);
  not csa_tree_sub001036_groupi_g5864(csa_tree_sub001036_groupi_n_160 ,csa_tree_sub001036_groupi_n_63);
  not csa_tree_sub001036_groupi_g5865(csa_tree_sub001036_groupi_n_159 ,csa_tree_sub001036_groupi_n_130);
  not csa_tree_sub001036_groupi_g5868(csa_tree_sub001036_groupi_n_158 ,csa_tree_sub001036_groupi_n_124);
  not csa_tree_sub001036_groupi_g5869(csa_tree_sub001036_groupi_n_157 ,csa_tree_sub001036_groupi_n_100);
  not csa_tree_sub001036_groupi_drc_bufs(csa_tree_sub001036_groupi_n_145 ,csa_tree_sub001036_groupi_n_143);
  not csa_tree_sub001036_groupi_drc_bufs5870(csa_tree_sub001036_groupi_n_144 ,csa_tree_sub001036_groupi_n_143);
  not csa_tree_sub001036_groupi_drc_bufs5871(csa_tree_sub001036_groupi_n_143 ,n_127);
  not csa_tree_sub001036_groupi_drc_bufs5873(csa_tree_sub001036_groupi_n_142 ,csa_tree_sub001036_groupi_n_140);
  not csa_tree_sub001036_groupi_drc_bufs5874(csa_tree_sub001036_groupi_n_141 ,csa_tree_sub001036_groupi_n_140);
  not csa_tree_sub001036_groupi_drc_bufs5875(csa_tree_sub001036_groupi_n_140 ,n_140);
  not csa_tree_sub001036_groupi_drc_bufs5877(csa_tree_sub001036_groupi_n_139 ,csa_tree_sub001036_groupi_n_137);
  not csa_tree_sub001036_groupi_drc_bufs5878(csa_tree_sub001036_groupi_n_138 ,csa_tree_sub001036_groupi_n_137);
  not csa_tree_sub001036_groupi_drc_bufs5879(csa_tree_sub001036_groupi_n_137 ,n_121);
  not csa_tree_sub001036_groupi_drc_bufs5881(csa_tree_sub001036_groupi_n_136 ,csa_tree_sub001036_groupi_n_134);
  not csa_tree_sub001036_groupi_drc_bufs5882(csa_tree_sub001036_groupi_n_135 ,csa_tree_sub001036_groupi_n_134);
  not csa_tree_sub001036_groupi_drc_bufs5883(csa_tree_sub001036_groupi_n_134 ,n_120);
  not csa_tree_sub001036_groupi_drc_bufs5885(csa_tree_sub001036_groupi_n_133 ,csa_tree_sub001036_groupi_n_131);
  not csa_tree_sub001036_groupi_drc_bufs5886(csa_tree_sub001036_groupi_n_132 ,csa_tree_sub001036_groupi_n_131);
  not csa_tree_sub001036_groupi_drc_bufs5887(csa_tree_sub001036_groupi_n_131 ,n_141);
  not csa_tree_sub001036_groupi_drc_bufs5893(csa_tree_sub001036_groupi_n_130 ,csa_tree_sub001036_groupi_n_128);
  not csa_tree_sub001036_groupi_drc_bufs5894(csa_tree_sub001036_groupi_n_129 ,csa_tree_sub001036_groupi_n_128);
  not csa_tree_sub001036_groupi_drc_bufs5895(csa_tree_sub001036_groupi_n_128 ,n_133);
  not csa_tree_sub001036_groupi_drc_bufs5897(csa_tree_sub001036_groupi_n_127 ,csa_tree_sub001036_groupi_n_125);
  not csa_tree_sub001036_groupi_drc_bufs5898(csa_tree_sub001036_groupi_n_126 ,csa_tree_sub001036_groupi_n_125);
  not csa_tree_sub001036_groupi_drc_bufs5899(csa_tree_sub001036_groupi_n_125 ,n_115);
  not csa_tree_sub001036_groupi_drc_bufs5901(csa_tree_sub001036_groupi_n_124 ,csa_tree_sub001036_groupi_n_122);
  not csa_tree_sub001036_groupi_drc_bufs5902(csa_tree_sub001036_groupi_n_123 ,csa_tree_sub001036_groupi_n_122);
  not csa_tree_sub001036_groupi_drc_bufs5903(csa_tree_sub001036_groupi_n_122 ,n_132);
  not csa_tree_sub001036_groupi_drc_bufs5905(csa_tree_sub001036_groupi_n_121 ,csa_tree_sub001036_groupi_n_119);
  not csa_tree_sub001036_groupi_drc_bufs5906(csa_tree_sub001036_groupi_n_120 ,csa_tree_sub001036_groupi_n_119);
  not csa_tree_sub001036_groupi_drc_bufs5907(csa_tree_sub001036_groupi_n_119 ,n_122);
  not csa_tree_sub001036_groupi_drc_bufs5909(csa_tree_sub001036_groupi_n_118 ,csa_tree_sub001036_groupi_n_116);
  not csa_tree_sub001036_groupi_drc_bufs5910(csa_tree_sub001036_groupi_n_117 ,csa_tree_sub001036_groupi_n_116);
  not csa_tree_sub001036_groupi_drc_bufs5911(csa_tree_sub001036_groupi_n_116 ,n_116);
  not csa_tree_sub001036_groupi_drc_bufs5913(csa_tree_sub001036_groupi_n_115 ,csa_tree_sub001036_groupi_n_113);
  not csa_tree_sub001036_groupi_drc_bufs5914(csa_tree_sub001036_groupi_n_114 ,csa_tree_sub001036_groupi_n_113);
  not csa_tree_sub001036_groupi_drc_bufs5915(csa_tree_sub001036_groupi_n_113 ,n_124);
  not csa_tree_sub001036_groupi_drc_bufs5917(csa_tree_sub001036_groupi_n_112 ,csa_tree_sub001036_groupi_n_110);
  not csa_tree_sub001036_groupi_drc_bufs5918(csa_tree_sub001036_groupi_n_111 ,csa_tree_sub001036_groupi_n_110);
  not csa_tree_sub001036_groupi_drc_bufs5919(csa_tree_sub001036_groupi_n_110 ,n_137);
  not csa_tree_sub001036_groupi_drc_bufs5921(csa_tree_sub001036_groupi_n_109 ,csa_tree_sub001036_groupi_n_107);
  not csa_tree_sub001036_groupi_drc_bufs5922(csa_tree_sub001036_groupi_n_108 ,csa_tree_sub001036_groupi_n_107);
  not csa_tree_sub001036_groupi_drc_bufs5923(csa_tree_sub001036_groupi_n_107 ,n_129);
  not csa_tree_sub001036_groupi_drc_bufs5925(csa_tree_sub001036_groupi_n_106 ,csa_tree_sub001036_groupi_n_104);
  not csa_tree_sub001036_groupi_drc_bufs5926(csa_tree_sub001036_groupi_n_105 ,csa_tree_sub001036_groupi_n_104);
  not csa_tree_sub001036_groupi_drc_bufs5927(csa_tree_sub001036_groupi_n_104 ,n_114);
  not csa_tree_sub001036_groupi_drc_bufs5929(csa_tree_sub001036_groupi_n_103 ,csa_tree_sub001036_groupi_n_101);
  not csa_tree_sub001036_groupi_drc_bufs5930(csa_tree_sub001036_groupi_n_102 ,csa_tree_sub001036_groupi_n_101);
  not csa_tree_sub001036_groupi_drc_bufs5931(csa_tree_sub001036_groupi_n_101 ,n_131);
  not csa_tree_sub001036_groupi_drc_bufs5933(csa_tree_sub001036_groupi_n_100 ,csa_tree_sub001036_groupi_n_98);
  not csa_tree_sub001036_groupi_drc_bufs5934(csa_tree_sub001036_groupi_n_99 ,csa_tree_sub001036_groupi_n_98);
  not csa_tree_sub001036_groupi_drc_bufs5935(csa_tree_sub001036_groupi_n_98 ,n_130);
  not csa_tree_sub001036_groupi_drc_bufs5937(csa_tree_sub001036_groupi_n_97 ,csa_tree_sub001036_groupi_n_95);
  not csa_tree_sub001036_groupi_drc_bufs5938(csa_tree_sub001036_groupi_n_96 ,csa_tree_sub001036_groupi_n_95);
  not csa_tree_sub001036_groupi_drc_bufs5939(csa_tree_sub001036_groupi_n_95 ,n_138);
  not csa_tree_sub001036_groupi_drc_bufs5941(csa_tree_sub001036_groupi_n_94 ,csa_tree_sub001036_groupi_n_92);
  not csa_tree_sub001036_groupi_drc_bufs5942(csa_tree_sub001036_groupi_n_93 ,csa_tree_sub001036_groupi_n_92);
  not csa_tree_sub001036_groupi_drc_bufs5943(csa_tree_sub001036_groupi_n_92 ,n_139);
  not csa_tree_sub001036_groupi_drc_bufs5945(csa_tree_sub001036_groupi_n_91 ,csa_tree_sub001036_groupi_n_89);
  not csa_tree_sub001036_groupi_drc_bufs5946(csa_tree_sub001036_groupi_n_90 ,csa_tree_sub001036_groupi_n_89);
  not csa_tree_sub001036_groupi_drc_bufs5947(csa_tree_sub001036_groupi_n_89 ,csa_tree_sub001036_groupi_n_503);
  not csa_tree_sub001036_groupi_drc_bufs5949(csa_tree_sub001036_groupi_n_88 ,csa_tree_sub001036_groupi_n_86);
  not csa_tree_sub001036_groupi_drc_bufs5950(csa_tree_sub001036_groupi_n_87 ,csa_tree_sub001036_groupi_n_86);
  not csa_tree_sub001036_groupi_drc_bufs5951(csa_tree_sub001036_groupi_n_86 ,n_126);
  not csa_tree_sub001036_groupi_drc_bufs5953(csa_tree_sub001036_groupi_n_85 ,csa_tree_sub001036_groupi_n_83);
  not csa_tree_sub001036_groupi_drc_bufs5954(csa_tree_sub001036_groupi_n_84 ,csa_tree_sub001036_groupi_n_83);
  not csa_tree_sub001036_groupi_drc_bufs5955(csa_tree_sub001036_groupi_n_83 ,n_125);
  not csa_tree_sub001036_groupi_drc_bufs5957(csa_tree_sub001036_groupi_n_82 ,csa_tree_sub001036_groupi_n_80);
  not csa_tree_sub001036_groupi_drc_bufs5958(csa_tree_sub001036_groupi_n_81 ,csa_tree_sub001036_groupi_n_80);
  not csa_tree_sub001036_groupi_drc_bufs5959(csa_tree_sub001036_groupi_n_80 ,n_119);
  not csa_tree_sub001036_groupi_drc_bufs5961(csa_tree_sub001036_groupi_n_79 ,csa_tree_sub001036_groupi_n_77);
  not csa_tree_sub001036_groupi_drc_bufs5962(csa_tree_sub001036_groupi_n_78 ,csa_tree_sub001036_groupi_n_77);
  not csa_tree_sub001036_groupi_drc_bufs5963(csa_tree_sub001036_groupi_n_77 ,n_117);
  not csa_tree_sub001036_groupi_drc_bufs5965(csa_tree_sub001036_groupi_n_76 ,csa_tree_sub001036_groupi_n_74);
  not csa_tree_sub001036_groupi_drc_bufs5966(csa_tree_sub001036_groupi_n_75 ,csa_tree_sub001036_groupi_n_74);
  not csa_tree_sub001036_groupi_drc_bufs5967(csa_tree_sub001036_groupi_n_74 ,n_128);
  not csa_tree_sub001036_groupi_drc_bufs5969(csa_tree_sub001036_groupi_n_73 ,csa_tree_sub001036_groupi_n_71);
  not csa_tree_sub001036_groupi_drc_bufs5970(csa_tree_sub001036_groupi_n_72 ,csa_tree_sub001036_groupi_n_71);
  not csa_tree_sub001036_groupi_drc_bufs5971(csa_tree_sub001036_groupi_n_71 ,n_134);
  not csa_tree_sub001036_groupi_drc_bufs5973(csa_tree_sub001036_groupi_n_70 ,csa_tree_sub001036_groupi_n_68);
  not csa_tree_sub001036_groupi_drc_bufs5974(csa_tree_sub001036_groupi_n_69 ,csa_tree_sub001036_groupi_n_68);
  not csa_tree_sub001036_groupi_drc_bufs5975(csa_tree_sub001036_groupi_n_68 ,n_123);
  not csa_tree_sub001036_groupi_drc_bufs5977(csa_tree_sub001036_groupi_n_67 ,csa_tree_sub001036_groupi_n_65);
  not csa_tree_sub001036_groupi_drc_bufs5978(csa_tree_sub001036_groupi_n_66 ,csa_tree_sub001036_groupi_n_65);
  not csa_tree_sub001036_groupi_drc_bufs5979(csa_tree_sub001036_groupi_n_65 ,n_118);
  not csa_tree_sub001036_groupi_drc_bufs5981(csa_tree_sub001036_groupi_n_64 ,csa_tree_sub001036_groupi_n_62);
  not csa_tree_sub001036_groupi_drc_bufs5982(csa_tree_sub001036_groupi_n_63 ,csa_tree_sub001036_groupi_n_62);
  not csa_tree_sub001036_groupi_drc_bufs5983(csa_tree_sub001036_groupi_n_62 ,n_136);
  not csa_tree_sub001036_groupi_drc_bufs5985(csa_tree_sub001036_groupi_n_61 ,csa_tree_sub001036_groupi_n_59);
  not csa_tree_sub001036_groupi_drc_bufs5986(csa_tree_sub001036_groupi_n_60 ,csa_tree_sub001036_groupi_n_59);
  not csa_tree_sub001036_groupi_drc_bufs5987(csa_tree_sub001036_groupi_n_59 ,n_135);
  not csa_tree_sub001036_groupi_drc_bufs5990(csa_tree_sub001036_groupi_n_58 ,csa_tree_sub001036_groupi_n_154);
  not csa_tree_sub001036_groupi_drc_bufs5991(csa_tree_sub001036_groupi_n_154 ,csa_tree_sub001036_groupi_n_323);
  not csa_tree_sub001036_groupi_drc_bufs5993(csa_tree_sub001036_groupi_n_57 ,csa_tree_sub001036_groupi_n_56);
  not csa_tree_sub001036_groupi_drc_bufs5995(csa_tree_sub001036_groupi_n_56 ,csa_tree_sub001036_groupi_n_504);
  not csa_tree_sub001036_groupi_drc_bufs5998(csa_tree_sub001036_groupi_n_55 ,csa_tree_sub001036_groupi_n_54);
  not csa_tree_sub001036_groupi_drc_bufs5999(csa_tree_sub001036_groupi_n_54 ,csa_tree_sub001036_groupi_n_172);
  not csa_tree_sub001036_groupi_drc_bufs6002(csa_tree_sub001036_groupi_n_53 ,csa_tree_sub001036_groupi_n_52);
  not csa_tree_sub001036_groupi_drc_bufs6003(csa_tree_sub001036_groupi_n_52 ,csa_tree_sub001036_groupi_n_160);
  not csa_tree_sub001036_groupi_drc_bufs6005(csa_tree_sub001036_groupi_n_51 ,csa_tree_sub001036_groupi_n_50);
  not csa_tree_sub001036_groupi_drc_bufs6007(csa_tree_sub001036_groupi_n_50 ,csa_tree_sub001036_groupi_n_173);
  not csa_tree_sub001036_groupi_drc_bufs6017(csa_tree_sub001036_groupi_n_49 ,csa_tree_sub001036_groupi_n_155);
  not csa_tree_sub001036_groupi_drc_bufs6018(csa_tree_sub001036_groupi_n_155 ,csa_tree_sub001036_groupi_n_587);
  not csa_tree_sub001036_groupi_drc_bufs6021(csa_tree_sub001036_groupi_n_48 ,csa_tree_sub001036_groupi_n_156);
  not csa_tree_sub001036_groupi_drc_bufs6022(csa_tree_sub001036_groupi_n_156 ,csa_tree_sub001036_groupi_n_1232);
  not csa_tree_sub001036_groupi_drc_bufs6024(csa_tree_sub001036_groupi_n_47 ,csa_tree_sub001036_groupi_n_46);
  not csa_tree_sub001036_groupi_drc_bufs6026(csa_tree_sub001036_groupi_n_46 ,csa_tree_sub001036_groupi_n_505);
  not csa_tree_sub001036_groupi_drc_bufs6028(csa_tree_sub001036_groupi_n_45 ,csa_tree_sub001036_groupi_n_44);
  not csa_tree_sub001036_groupi_drc_bufs6030(csa_tree_sub001036_groupi_n_44 ,csa_tree_sub001036_groupi_n_145);
  not csa_tree_sub001036_groupi_drc_bufs6032(csa_tree_sub001036_groupi_n_43 ,csa_tree_sub001036_groupi_n_42);
  not csa_tree_sub001036_groupi_drc_bufs6034(csa_tree_sub001036_groupi_n_42 ,csa_tree_sub001036_groupi_n_130);
  not csa_tree_sub001036_groupi_drc_bufs6036(csa_tree_sub001036_groupi_n_41 ,csa_tree_sub001036_groupi_n_40);
  not csa_tree_sub001036_groupi_drc_bufs6038(csa_tree_sub001036_groupi_n_40 ,csa_tree_sub001036_groupi_n_127);
  not csa_tree_sub001036_groupi_drc_bufs6040(csa_tree_sub001036_groupi_n_39 ,csa_tree_sub001036_groupi_n_151);
  not csa_tree_sub001036_groupi_drc_bufs6042(csa_tree_sub001036_groupi_n_151 ,csa_tree_sub001036_groupi_n_118);
  not csa_tree_sub001036_groupi_drc_bufs6044(csa_tree_sub001036_groupi_n_38 ,csa_tree_sub001036_groupi_n_147);
  not csa_tree_sub001036_groupi_drc_bufs6046(csa_tree_sub001036_groupi_n_147 ,csa_tree_sub001036_groupi_n_142);
  not csa_tree_sub001036_groupi_drc_bufs6048(csa_tree_sub001036_groupi_n_37 ,csa_tree_sub001036_groupi_n_36);
  not csa_tree_sub001036_groupi_drc_bufs6050(csa_tree_sub001036_groupi_n_36 ,csa_tree_sub001036_groupi_n_124);
  not csa_tree_sub001036_groupi_drc_bufs6052(csa_tree_sub001036_groupi_n_35 ,csa_tree_sub001036_groupi_n_148);
  not csa_tree_sub001036_groupi_drc_bufs6054(csa_tree_sub001036_groupi_n_148 ,csa_tree_sub001036_groupi_n_121);
  not csa_tree_sub001036_groupi_drc_bufs6057(csa_tree_sub001036_groupi_n_34 ,csa_tree_sub001036_groupi_n_33);
  not csa_tree_sub001036_groupi_drc_bufs6058(csa_tree_sub001036_groupi_n_33 ,csa_tree_sub001036_groupi_n_103);
  not csa_tree_sub001036_groupi_drc_bufs6061(csa_tree_sub001036_groupi_n_32 ,csa_tree_sub001036_groupi_n_31);
  not csa_tree_sub001036_groupi_drc_bufs6062(csa_tree_sub001036_groupi_n_31 ,csa_tree_sub001036_groupi_n_141);
  not csa_tree_sub001036_groupi_drc_bufs6064(csa_tree_sub001036_groupi_n_30 ,csa_tree_sub001036_groupi_n_29);
  not csa_tree_sub001036_groupi_drc_bufs6066(csa_tree_sub001036_groupi_n_29 ,csa_tree_sub001036_groupi_n_111);
  not csa_tree_sub001036_groupi_drc_bufs6069(csa_tree_sub001036_groupi_n_28 ,csa_tree_sub001036_groupi_n_27);
  not csa_tree_sub001036_groupi_drc_bufs6070(csa_tree_sub001036_groupi_n_27 ,csa_tree_sub001036_groupi_n_136);
  not csa_tree_sub001036_groupi_drc_bufs6073(csa_tree_sub001036_groupi_n_26 ,csa_tree_sub001036_groupi_n_25);
  not csa_tree_sub001036_groupi_drc_bufs6074(csa_tree_sub001036_groupi_n_25 ,csa_tree_sub001036_groupi_n_144);
  not csa_tree_sub001036_groupi_drc_bufs6077(csa_tree_sub001036_groupi_n_24 ,csa_tree_sub001036_groupi_n_23);
  not csa_tree_sub001036_groupi_drc_bufs6078(csa_tree_sub001036_groupi_n_23 ,csa_tree_sub001036_groupi_n_106);
  not csa_tree_sub001036_groupi_drc_bufs6081(csa_tree_sub001036_groupi_n_22 ,csa_tree_sub001036_groupi_n_21);
  not csa_tree_sub001036_groupi_drc_bufs6082(csa_tree_sub001036_groupi_n_21 ,csa_tree_sub001036_groupi_n_138);
  not csa_tree_sub001036_groupi_drc_bufs6085(csa_tree_sub001036_groupi_n_20 ,csa_tree_sub001036_groupi_n_19);
  not csa_tree_sub001036_groupi_drc_bufs6086(csa_tree_sub001036_groupi_n_19 ,csa_tree_sub001036_groupi_n_108);
  not csa_tree_sub001036_groupi_drc_bufs6089(csa_tree_sub001036_groupi_n_18 ,csa_tree_sub001036_groupi_n_149);
  not csa_tree_sub001036_groupi_drc_bufs6090(csa_tree_sub001036_groupi_n_149 ,csa_tree_sub001036_groupi_n_114);
  not csa_tree_sub001036_groupi_drc_bufs6093(csa_tree_sub001036_groupi_n_17 ,csa_tree_sub001036_groupi_n_16);
  not csa_tree_sub001036_groupi_drc_bufs6094(csa_tree_sub001036_groupi_n_16 ,csa_tree_sub001036_groupi_n_100);
  not csa_tree_sub001036_groupi_drc_bufs6097(csa_tree_sub001036_groupi_n_15 ,csa_tree_sub001036_groupi_n_146);
  not csa_tree_sub001036_groupi_drc_bufs6098(csa_tree_sub001036_groupi_n_146 ,csa_tree_sub001036_groupi_n_139);
  not csa_tree_sub001036_groupi_drc_bufs6101(csa_tree_sub001036_groupi_n_14 ,csa_tree_sub001036_groupi_n_153);
  not csa_tree_sub001036_groupi_drc_bufs6102(csa_tree_sub001036_groupi_n_153 ,csa_tree_sub001036_groupi_n_94);
  not csa_tree_sub001036_groupi_drc_bufs6105(csa_tree_sub001036_groupi_n_13 ,csa_tree_sub001036_groupi_n_150);
  not csa_tree_sub001036_groupi_drc_bufs6106(csa_tree_sub001036_groupi_n_150 ,csa_tree_sub001036_groupi_n_97);
  not csa_tree_sub001036_groupi_drc_bufs6109(csa_tree_sub001036_groupi_n_12 ,csa_tree_sub001036_groupi_n_152);
  not csa_tree_sub001036_groupi_drc_bufs6110(csa_tree_sub001036_groupi_n_152 ,csa_tree_sub001036_groupi_n_133);
  not csa_tree_sub001036_groupi_drc_bufs6112(csa_tree_sub001036_groupi_n_11 ,csa_tree_sub001036_groupi_n_10);
  not csa_tree_sub001036_groupi_drc_bufs6114(csa_tree_sub001036_groupi_n_10 ,csa_tree_sub001036_groupi_n_135);
  not csa_tree_sub001036_groupi_drc_bufs6116(csa_tree_sub001036_groupi_n_9 ,csa_tree_sub001036_groupi_n_8);
  not csa_tree_sub001036_groupi_drc_bufs6118(csa_tree_sub001036_groupi_n_8 ,csa_tree_sub001036_groupi_n_132);
  xor csa_tree_sub001036_groupi_g2(out1[10] ,csa_tree_sub001036_groupi_n_1472 ,csa_tree_sub001036_groupi_n_1453);
  xor csa_tree_sub001036_groupi_g6120(out1[9] ,csa_tree_sub001036_groupi_n_1470 ,csa_tree_sub001036_groupi_n_1461);
  xor csa_tree_sub001036_groupi_g6121(csa_tree_sub001036_groupi_n_5 ,csa_tree_sub001036_groupi_n_1346 ,csa_tree_sub001036_groupi_n_1361);
  xor csa_tree_sub001036_groupi_g6122(csa_tree_sub001036_groupi_n_4 ,csa_tree_sub001036_groupi_n_1338 ,csa_tree_sub001036_groupi_n_1363);
  xor csa_tree_sub001036_groupi_g6123(csa_tree_sub001036_groupi_n_3 ,csa_tree_sub001036_groupi_n_1093 ,csa_tree_sub001036_groupi_n_1235);
  xor csa_tree_sub001036_groupi_g6124(csa_tree_sub001036_groupi_n_2 ,csa_tree_sub001036_groupi_n_1056 ,csa_tree_sub001036_groupi_n_1132);
  xor csa_tree_sub001036_groupi_g6125(csa_tree_sub001036_groupi_n_1 ,csa_tree_sub001036_groupi_n_863 ,csa_tree_sub001036_groupi_n_910);
  xor csa_tree_sub001036_groupi_g6126(csa_tree_sub001036_groupi_n_0 ,csa_tree_sub001036_groupi_n_817 ,csa_tree_sub001036_groupi_n_46);
endmodule
