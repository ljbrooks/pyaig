module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, out1);
  input [3:0] in1;
  input [25:0] in2, in4;
  input in3, in5, in6, in7, in8, in9, in10, in12;
  input [6:0] in11;
  input [2:0] in13, in14, in15, in16, in17;
  output [25:0] out1;
  wire [3:0] in1;
  wire [25:0] in2, in4;
  wire in3, in5, in6, in7, in8, in9, in10, in12;
  wire [6:0] in11;
  wire [2:0] in13, in14, in15, in16, in17;
  wire [25:0] out1;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__139, w__140, w__141, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__157, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__171, w__172, w__173, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662;
  not g__1(w__278 ,w__279);
  not g__2(w__359 ,in3);
  or g__3(w__350 ,w__252 ,w__277);
  and g__4(w__277 ,in15[0] ,w__272);
  or g__5(w__276 ,w__261 ,w__271);
  or g__6(w__275 ,w__262 ,w__269);
  or g__7(w__346 ,w__270 ,w__268);
  and g__8(w__274 ,in15[2] ,w__272);
  and g__9(w__273 ,in15[1] ,w__272);
  or g__10(w__271 ,w__265 ,w__259);
  and g__11(w__272 ,w__243 ,w__263);
  or g__12(w__270 ,w__248 ,w__260);
  or g__13(w__269 ,w__266 ,w__264);
  or g__14(w__268 ,w__255 ,w__267);
  and g__15(w__267 ,in16[0] ,w__256);
  and g__16(w__266 ,in16[2] ,w__256);
  and g__17(w__265 ,in16[1] ,w__256);
  and g__18(w__264 ,in17[2] ,w__258);
  not g__19(w__279 ,w__263);
  or g__20(w__262 ,w__247 ,w__254);
  or g__21(w__261 ,w__246 ,w__257);
  and g__22(w__260 ,in17[0] ,w__258);
  and g__23(w__259 ,in17[1] ,w__258);
  and g__24(w__263 ,w__242 ,w__280);
  and g__25(w__257 ,in14[1] ,w__253);
  or g__26(w__280 ,in10 ,w__250);
  and g__27(w__258 ,w__244 ,w__249);
  and g__28(w__349 ,in1[3] ,w__252);
  and g__29(w__255 ,in14[0] ,w__253);
  and g__30(w__254 ,in14[2] ,w__253);
  and g__31(w__256 ,in9 ,w__245);
  not g__32(w__251 ,w__252);
  or g__33(w__250 ,in8 ,in9);
  nor g__34(w__249 ,in7 ,in9);
  and g__35(w__253 ,in8 ,w__243);
  and g__36(w__252 ,in7 ,w__242);
  and g__37(w__248 ,in1[0] ,in7);
  and g__38(w__247 ,in1[2] ,in7);
  and g__39(w__246 ,in1[1] ,in7);
  nor g__40(w__245 ,in7 ,in8);
  not g__41(w__244 ,in8);
  not g__42(w__243 ,in7);
  not g__43(w__242 ,in6);
  buf g__44(w__348 ,w__275);
  buf g__45(w__347 ,w__276);
  buf g__46(w__352 ,w__274);
  buf g__47(w__351 ,w__273);
  buf g__48(w__662 ,w__251);
  or g__49(w__241 ,w__223 ,w__238);
  or g__50(w__240 ,w__214 ,w__229);
  or g__51(w__239 ,w__224 ,w__232);
  or g__52(w__238 ,w__213 ,w__234);
  or g__53(w__337 ,w__231 ,w__227);
  or g__54(w__237 ,w__216 ,w__228);
  or g__55(w__335 ,w__235 ,w__236);
  or g__56(w__334 ,w__230 ,w__233);
  or g__57(w__236 ,w__215 ,w__222);
  and g__58(w__235 ,in11[1] ,w__226);
  and g__59(w__234 ,in11[2] ,w__203);
  or g__60(w__233 ,w__212 ,w__221);
  and g__61(w__232 ,in11[4] ,w__206);
  and g__62(w__231 ,in11[3] ,w__203);
  and g__63(w__230 ,in11[0] ,w__206);
  and g__64(w__229 ,in11[6] ,w__205);
  and g__65(w__228 ,in11[5] ,w__205);
  or g__66(w__227 ,w__211 ,w__225);
  or g__67(w__224 ,w__219 ,w__218);
  and g__68(w__226 ,w__209 ,w__217);
  and g__69(w__223 ,w__343 ,w__220);
  and g__70(w__222 ,w__342 ,w__208);
  and g__71(w__221 ,w__341 ,w__208);
  and g__72(w__219 ,in6 ,w__356);
  nor g__73(w__217 ,in7 ,w__280);
  and g__74(w__216 ,in6 ,w__357);
  or g__75(w__220 ,w__210 ,w__278);
  and g__76(w__215 ,in6 ,w__353);
  and g__77(w__214 ,in6 ,w__358);
  and g__78(w__213 ,in6 ,w__354);
  and g__79(w__212 ,in1[0] ,in6);
  and g__80(w__211 ,in6 ,w__355);
  not g__81(w__210 ,w__662);
  not g__82(w__209 ,in6);
  not g__83(w__208 ,w__207);
  not g__84(w__207 ,w__220);
  buf g__85(w__336 ,w__241);
  buf g__86(w__338 ,w__239);
  buf g__87(w__340 ,w__240);
  buf g__88(w__339 ,w__237);
  not g__89(w__206 ,w__204);
  not g__90(w__205 ,w__204);
  not g__91(w__204 ,w__226);
  not g__92(w__203 ,w__202);
  not g__93(w__202 ,w__226);
  buf g__94(w__494 ,w__407);
  buf g__95(w__493 ,w__419);
  buf g__96(w__492 ,w__418);
  buf g__97(w__491 ,w__417);
  buf g__98(w__490 ,w__416);
  buf g__99(w__489 ,w__415);
  buf g__100(w__488 ,w__414);
  buf g__101(w__487 ,w__413);
  buf g__102(w__486 ,w__412);
  buf g__103(w__485 ,w__411);
  buf g__104(w__484 ,in2[24]);
  buf g__105(w__483 ,w__409);
  buf g__106(w__482 ,w__408);
  buf g__107(w__481 ,w__420);
  buf g__108(w__480 ,w__406);
  buf g__109(w__479 ,w__405);
  buf g__110(w__478 ,w__424);
  buf g__111(w__477 ,w__425);
  buf g__112(w__476 ,w__426);
  buf g__113(w__475 ,w__428);
  buf g__114(w__474 ,w__429);
  buf g__115(w__473 ,w__423);
  buf g__116(w__472 ,w__427);
  buf g__117(w__471 ,w__410);
  buf g__118(w__470 ,w__422);
  buf g__119(w__469 ,w__421);
  or g__120(w__468 ,w__400 ,w__441);
  or g__121(w__467 ,w__399 ,w__437);
  or g__122(w__466 ,w__402 ,w__449);
  or g__123(w__465 ,w__397 ,w__431);
  or g__124(w__455 ,w__398 ,w__434);
  or g__125(w__454 ,w__396 ,w__445);
  or g__126(w__453 ,w__401 ,w__403);
  and g__127(w__452 ,w__483 ,w__363);
  and g__128(w__451 ,w__493 ,w__380);
  and g__129(w__450 ,w__494 ,w__377);
  and g__130(w__449 ,w__475 ,w__365);
  and g__131(w__448 ,w__481 ,w__361);
  and g__132(w__447 ,w__486 ,w__371);
  and g__133(w__446 ,w__469 ,w__365);
  and g__134(w__445 ,w__474 ,w__375);
  and g__135(w__444 ,w__470 ,w__375);
  and g__136(w__333 ,w__484 ,w__378);
  and g__137(w__443 ,w__482 ,w__380);
  and g__138(w__442 ,w__487 ,w__371);
  and g__139(w__441 ,w__473 ,w__369);
  and g__140(w__440 ,w__479 ,w__374);
  and g__141(w__439 ,w__488 ,w__363);
  and g__142(w__438 ,w__485 ,w__374);
  and g__143(w__437 ,w__478 ,w__372);
  and g__144(w__436 ,w__489 ,w__369);
  and g__145(w__435 ,w__480 ,w__368);
  and g__146(w__434 ,w__477 ,w__366);
  and g__147(w__433 ,w__490 ,w__381);
  and g__148(w__432 ,w__491 ,w__368);
  and g__149(w__431 ,w__476 ,w__372);
  and g__150(w__430 ,w__471 ,w__366);
  and g__151(w__404 ,w__492 ,w__361);
  and g__152(w__403 ,w__472 ,w__377);
  and g__153(w__402 ,w__385 ,w__335);
  and g__154(w__401 ,w__383 ,w__336);
  and g__155(w__400 ,w__393 ,w__340);
  and g__156(w__399 ,w__383 ,w__339);
  and g__157(w__398 ,w__386 ,w__338);
  and g__158(w__397 ,w__386 ,w__337);
  and g__159(w__396 ,w__385 ,w__334);
  not g__160(w__395 ,w__389);
  not g__161(w__394 ,w__388);
  not g__162(w__393 ,w__391);
  not g__163(w__392 ,w__391);
  not g__164(w__391 ,w__388);
  not g__165(w__390 ,w__389);
  not g__166(w__389 ,w__387);
  not g__167(w__388 ,w__387);
  not g__168(w__387 ,w__359);
  not g__169(w__386 ,w__384);
  not g__170(w__385 ,w__384);
  not g__171(w__384 ,w__392);
  not g__172(w__383 ,w__382);
  not g__173(w__382 ,w__393);
  buf g__174(w__308 ,w__454);
  buf g__175(w__313 ,w__467);
  buf g__176(w__310 ,w__453);
  buf g__177(w__309 ,w__466);
  buf g__178(w__311 ,w__465);
  buf g__179(w__314 ,w__468);
  buf g__180(w__312 ,w__455);
  buf g__181(w__319 ,w__404);
  buf g__182(w__329 ,w__443);
  buf g__183(w__328 ,w__452);
  buf g__184(w__323 ,w__439);
  buf g__185(w__318 ,w__451);
  buf g__186(w__330 ,w__450);
  buf g__187(w__321 ,w__433);
  buf g__188(w__317 ,w__448);
  buf g__189(w__320 ,w__432);
  buf g__190(w__324 ,w__442);
  buf g__191(w__327 ,w__430);
  buf g__192(w__331 ,w__435);
  buf g__193(w__326 ,w__438);
  buf g__194(w__322 ,w__436);
  buf g__195(w__316 ,w__446);
  buf g__196(w__332 ,w__440);
  buf g__197(w__325 ,w__447);
  buf g__198(w__315 ,w__444);
  not g__199(w__381 ,w__379);
  not g__200(w__380 ,w__379);
  not g__201(w__379 ,w__390);
  not g__202(w__378 ,w__376);
  not g__203(w__377 ,w__376);
  not g__204(w__376 ,w__390);
  not g__205(w__375 ,w__373);
  not g__206(w__374 ,w__373);
  not g__207(w__373 ,w__394);
  not g__208(w__372 ,w__370);
  not g__209(w__371 ,w__370);
  not g__210(w__370 ,w__395);
  not g__211(w__369 ,w__367);
  not g__212(w__368 ,w__367);
  not g__213(w__367 ,w__395);
  not g__214(w__366 ,w__364);
  not g__215(w__365 ,w__364);
  not g__216(w__364 ,w__394);
  not g__217(w__363 ,w__362);
  not g__218(w__362 ,w__381);
  not g__219(w__361 ,w__360);
  not g__220(w__360 ,w__378);
  buf g__221(w__658 ,in2[11]);
  buf g__222(w__657 ,in2[23]);
  buf g__223(w__656 ,in2[22]);
  buf g__224(w__655 ,in2[21]);
  buf g__225(w__654 ,in2[20]);
  buf g__226(w__653 ,in2[19]);
  buf g__227(w__652 ,in2[18]);
  buf g__228(w__651 ,in2[17]);
  buf g__229(w__650 ,in2[16]);
  buf g__230(w__649 ,in2[15]);
  buf g__231(w__648 ,in2[14]);
  buf g__232(w__647 ,in2[13]);
  buf g__233(w__646 ,in2[12]);
  buf g__234(w__645 ,w__456);
  buf g__235(w__644 ,in2[10]);
  buf g__236(w__643 ,in2[9]);
  buf g__237(w__642 ,in2[8]);
  buf g__238(w__641 ,in2[7]);
  buf g__239(w__640 ,w__457);
  buf g__240(w__639 ,w__458);
  buf g__241(w__638 ,w__459);
  buf g__242(w__637 ,w__460);
  buf g__243(w__636 ,w__461);
  buf g__244(w__635 ,w__462);
  buf g__245(w__634 ,w__463);
  buf g__246(w__633 ,w__464);
  or g__247(w__307 ,w__573 ,w__595);
  or g__248(w__632 ,w__578 ,w__599);
  or g__249(w__631 ,w__580 ,w__605);
  or g__250(w__630 ,w__579 ,w__604);
  or g__251(w__629 ,w__576 ,w__601);
  or g__252(w__628 ,w__577 ,w__603);
  or g__253(w__627 ,w__575 ,w__602);
  or g__254(w__626 ,w__567 ,w__594);
  or g__255(w__625 ,w__571 ,w__598);
  or g__256(w__624 ,w__572 ,w__600);
  or g__257(w__623 ,w__570 ,w__597);
  or g__258(w__622 ,w__566 ,w__592);
  or g__259(w__621 ,w__568 ,w__608);
  or g__260(w__620 ,w__581 ,w__596);
  or g__261(w__619 ,w__557 ,w__588);
  or g__262(w__618 ,w__565 ,w__593);
  or g__263(w__617 ,w__564 ,w__591);
  or g__264(w__616 ,w__561 ,w__583);
  or g__265(w__615 ,w__563 ,w__590);
  or g__266(w__614 ,w__562 ,w__589);
  or g__267(w__613 ,w__559 ,w__585);
  or g__268(w__612 ,w__560 ,w__587);
  or g__269(w__611 ,w__558 ,w__586);
  or g__270(w__610 ,w__574 ,w__606);
  or g__271(w__609 ,w__582 ,w__584);
  or g__272(w__282 ,w__569 ,w__607);
  and g__273(w__608 ,w__640 ,w__504);
  and g__274(w__607 ,w__633 ,w__510);
  and g__275(w__606 ,w__646 ,w__498);
  and g__276(w__605 ,w__652 ,w__524);
  and g__277(w__604 ,w__658 ,w__521);
  and g__278(w__603 ,w__644 ,w__500);
  and g__279(w__602 ,w__643 ,w__496);
  and g__280(w__601 ,w__651 ,w__532);
  and g__281(w__600 ,w__642 ,w__501);
  and g__282(w__599 ,w__655 ,w__529);
  and g__283(w__598 ,w__650 ,w__542);
  and g__284(w__597 ,w__641 ,w__504);
  and g__285(w__596 ,w__657 ,w__503);
  and g__286(w__595 ,w__645 ,w__510);
  and g__287(w__594 ,w__654 ,w__532);
  and g__288(w__593 ,w__639 ,w__529);
  and g__289(w__592 ,w__649 ,w__496);
  and g__290(w__591 ,w__638 ,w__531);
  and g__291(w__590 ,w__648 ,w__501);
  and g__292(w__589 ,w__637 ,w__503);
  and g__293(w__588 ,w__656 ,w__528);
  and g__294(w__587 ,w__636 ,w__498);
  and g__295(w__586 ,w__635 ,w__528);
  and g__296(w__585 ,w__647 ,w__509);
  and g__297(w__584 ,w__634 ,w__500);
  and g__298(w__583 ,w__653 ,w__531);
  and g__299(w__582 ,in4[1] ,w__534);
  and g__300(w__581 ,in4[24] ,w__538);
  and g__301(w__580 ,in4[19] ,w__534);
  and g__302(w__579 ,in4[12] ,w__513);
  and g__303(w__578 ,in4[22] ,w__507);
  and g__304(w__577 ,in4[11] ,w__506);
  and g__305(w__576 ,in4[18] ,w__538);
  and g__306(w__575 ,in4[10] ,w__513);
  and g__307(w__574 ,in4[13] ,w__541);
  and g__308(w__573 ,in4[25] ,w__518);
  and g__309(w__572 ,in4[9] ,w__515);
  and g__310(w__571 ,in4[17] ,w__518);
  and g__311(w__570 ,in4[8] ,w__515);
  and g__312(w__569 ,in4[0] ,w__535);
  and g__313(w__568 ,in4[7] ,w__535);
  and g__314(w__567 ,in4[21] ,w__512);
  and g__315(w__566 ,in4[16] ,w__537);
  and g__316(w__565 ,in4[6] ,w__540);
  and g__317(w__564 ,in4[5] ,w__516);
  and g__318(w__563 ,in4[15] ,w__537);
  and g__319(w__562 ,in4[4] ,w__540);
  and g__320(w__561 ,in4[20] ,w__507);
  and g__321(w__560 ,in4[3] ,w__519);
  and g__322(w__559 ,in4[14] ,w__541);
  and g__323(w__558 ,in4[2] ,w__516);
  and g__324(w__557 ,in4[23] ,w__519);
  not g__325(w__556 ,w__526);
  not g__326(w__555 ,w__526);
  not g__327(w__554 ,w__545);
  not g__328(w__553 ,w__544);
  not g__329(w__552 ,w__544);
  not g__330(w__551 ,w__550);
  not g__331(w__550 ,w__548);
  not g__332(w__549 ,w__548);
  not g__333(w__548 ,w__545);
  not g__334(w__545 ,w__543);
  not g__335(w__544 ,w__543);
  not g__336(w__543 ,w__359);
  not g__337(w__542 ,w__546);
  not g__338(w__546 ,w__552);
  not g__339(w__541 ,w__539);
  not g__340(w__540 ,w__539);
  not g__341(w__539 ,w__546);
  not g__342(w__538 ,w__536);
  not g__343(w__537 ,w__536);
  not g__344(w__536 ,w__555);
  not g__345(w__535 ,w__533);
  not g__346(w__534 ,w__533);
  not g__347(w__533 ,w__547);
  not g__348(w__532 ,w__530);
  not g__349(w__531 ,w__530);
  not g__350(w__530 ,w__551);
  not g__351(w__529 ,w__527);
  not g__352(w__528 ,w__527);
  not g__353(w__527 ,w__551);
  not g__354(w__526 ,w__547);
  not g__355(w__547 ,w__554);
  buf g__356(w__283 ,w__609);
  buf g__357(w__295 ,w__610);
  buf g__358(w__284 ,w__611);
  buf g__359(w__285 ,w__612);
  buf g__360(w__296 ,w__613);
  buf g__361(w__286 ,w__614);
  buf g__362(w__297 ,w__615);
  buf g__363(w__299 ,w__625);
  buf g__364(w__302 ,w__616);
  buf g__365(w__294 ,w__630);
  buf g__366(w__287 ,w__617);
  buf g__367(w__304 ,w__632);
  buf g__368(w__301 ,w__631);
  buf g__369(w__298 ,w__622);
  buf g__370(w__290 ,w__623);
  buf g__371(w__291 ,w__624);
  buf g__372(w__292 ,w__627);
  buf g__373(w__303 ,w__626);
  buf g__374(w__305 ,w__619);
  buf g__375(w__288 ,w__618);
  buf g__376(w__300 ,w__629);
  buf g__377(w__306 ,w__620);
  buf g__378(w__293 ,w__628);
  buf g__379(w__289 ,w__621);
  not g__380(w__525 ,w__523);
  not g__381(w__524 ,w__523);
  not g__382(w__523 ,w__553);
  not g__383(w__522 ,w__520);
  not g__384(w__521 ,w__520);
  not g__385(w__520 ,w__553);
  not g__386(w__519 ,w__517);
  not g__387(w__518 ,w__517);
  not g__388(w__517 ,w__549);
  not g__389(w__516 ,w__514);
  not g__390(w__515 ,w__514);
  not g__391(w__514 ,w__549);
  not g__392(w__513 ,w__511);
  not g__393(w__512 ,w__511);
  not g__394(w__511 ,w__556);
  not g__395(w__510 ,w__508);
  not g__396(w__509 ,w__508);
  not g__397(w__508 ,w__552);
  not g__398(w__507 ,w__505);
  not g__399(w__506 ,w__505);
  not g__400(w__505 ,w__556);
  not g__401(w__504 ,w__502);
  not g__402(w__503 ,w__502);
  not g__403(w__502 ,w__525);
  not g__404(w__501 ,w__499);
  not g__405(w__500 ,w__499);
  not g__406(w__499 ,w__522);
  not g__407(w__498 ,w__497);
  not g__408(w__497 ,w__521);
  not g__409(w__496 ,w__495);
  not g__410(w__495 ,w__524);
  buf g__411(w__661 ,in1[0]);
  not g__412(w__660 ,w__359);
  and g__413(w__659 ,w__661 ,w__660);
  buf g__414(w__281 ,w__659);
  xnor g__415(w__344 ,w__18 ,w__349);
  nor g__416(w__19 ,w__18 ,w__4);
  and g__417(w__18 ,w__11 ,w__17);
  xnor g__418(w__343 ,w__15 ,w__13);
  or g__419(w__17 ,w__9 ,w__16);
  xor g__420(w__342 ,w__6 ,w__12);
  not g__421(w__16 ,w__15);
  or g__422(w__15 ,w__8 ,w__14);
  nor g__423(w__14 ,w__6 ,w__10);
  and g__424(w__341 ,w__6 ,w__7);
  xnor g__425(w__13 ,w__352 ,w__348);
  xnor g__426(w__12 ,w__351 ,w__347);
  or g__427(w__11 ,w__1 ,w__5);
  nor g__428(w__10 ,w__351 ,w__347);
  nor g__429(w__9 ,w__352 ,w__348);
  and g__430(w__8 ,w__351 ,w__347);
  or g__431(w__7 ,w__350 ,w__346);
  or g__432(w__6 ,w__3 ,w__2);
  not g__433(w__5 ,w__348);
  not g__434(w__4 ,w__349);
  not g__435(w__3 ,w__350);
  not g__436(w__2 ,w__346);
  not g__437(w__1 ,w__352);
  buf g__438(w__345 ,w__19);
  xnor g__439(w__357 ,w__51 ,in13[2]);
  nor g__440(w__53 ,w__51 ,w__21);
  and g__441(w__356 ,w__51 ,w__52);
  or g__442(w__52 ,w__36 ,w__49);
  or g__443(w__51 ,w__37 ,w__50);
  xnor g__444(w__355 ,w__46 ,w__47);
  not g__445(w__50 ,w__49);
  or g__446(w__49 ,w__45 ,w__48);
  and g__447(w__48 ,w__46 ,w__44);
  xnor g__448(w__354 ,w__30 ,w__42);
  xnor g__449(w__47 ,w__28 ,w__41);
  or g__450(w__46 ,w__39 ,w__43);
  nor g__451(w__45 ,w__28 ,w__41);
  or g__452(w__44 ,w__27 ,w__40);
  nor g__453(w__43 ,w__30 ,w__38);
  xnor g__454(w__42 ,w__33 ,in1[2]);
  not g__455(w__41 ,w__40);
  xnor g__456(w__40 ,w__34 ,w__24);
  nor g__457(w__39 ,w__26 ,w__33);
  and g__458(w__38 ,w__26 ,w__33);
  not g__459(w__37 ,w__36);
  or g__460(w__36 ,w__31 ,w__35);
  and g__461(w__35 ,in1[3] ,w__32);
  and g__462(w__353 ,w__30 ,w__29);
  xnor g__463(w__34 ,in13[1] ,in1[3]);
  xnor g__464(w__33 ,in13[1] ,in13[0]);
  or g__465(w__32 ,w__21 ,in13[1]);
  and g__466(w__31 ,in13[1] ,w__24);
  or g__467(w__30 ,w__25 ,w__23);
  or g__468(w__29 ,in13[0] ,in1[1]);
  not g__469(w__27 ,w__28);
  or g__470(w__28 ,w__22 ,w__25);
  not g__471(w__26 ,in1[2]);
  not g__472(w__25 ,in13[0]);
  not g__473(w__24 ,in13[2]);
  not g__474(w__23 ,in1[1]);
  not g__475(w__22 ,in13[1]);
  not g__476(w__21 ,w__20);
  not g__477(w__20 ,w__24);
  buf g__478(w__358 ,w__53);
  xnor g__479(w__428 ,w__71 ,in2[0]);
  xor g__480(w__426 ,w__70 ,w__56);
  xor g__481(w__427 ,w__72 ,w__336);
  or g__482(w__462 ,w__62 ,w__75);
  or g__483(w__425 ,w__54 ,w__73);
  or g__484(w__461 ,w__64 ,w__74);
  nor g__485(w__75 ,w__464 ,w__63);
  and g__486(w__74 ,in2[2] ,w__69);
  and g__487(w__73 ,in2[3] ,w__65);
  xnor g__488(w__423 ,w__340 ,in2[6]);
  xnor g__489(w__459 ,w__339 ,in2[5]);
  xnor g__490(w__460 ,w__338 ,in2[4]);
  xnor g__491(w__72 ,in1[2] ,in2[2]);
  xnor g__492(w__71 ,in1[1] ,in2[1]);
  xnor g__493(w__70 ,in1[3] ,in2[3]);
  or g__494(w__69 ,w__58 ,in1[2]);
  nor g__495(w__68 ,w__339 ,w__59);
  nor g__496(w__67 ,w__340 ,w__61);
  nor g__497(w__66 ,w__338 ,w__60);
  or g__498(w__65 ,w__57 ,in1[3]);
  and g__499(w__64 ,in1[2] ,w__58);
  nor g__500(w__63 ,in1[1] ,in2[1]);
  and g__501(w__62 ,in1[1] ,in2[1]);
  not g__502(w__456 ,in2[25]);
  not g__503(w__429 ,w__334);
  not g__504(w__408 ,in2[21]);
  not g__505(w__406 ,in2[23]);
  not g__506(w__412 ,in2[17]);
  not g__507(w__421 ,in2[8]);
  not g__508(w__415 ,in2[14]);
  not g__509(w__61 ,in2[6]);
  not g__510(w__409 ,in2[20]);
  not g__511(w__457 ,in2[7]);
  not g__512(w__417 ,in2[12]);
  not g__513(w__60 ,in2[4]);
  not g__514(w__410 ,in2[19]);
  not g__515(w__463 ,w__335);
  not g__516(w__418 ,in2[11]);
  not g__517(w__420 ,in2[9]);
  not g__518(w__419 ,in2[10]);
  not g__519(w__405 ,in2[24]);
  not g__520(w__414 ,in2[15]);
  not g__521(w__407 ,in2[22]);
  not g__522(w__413 ,in2[16]);
  not g__523(w__59 ,in2[5]);
  not g__524(w__416 ,in2[13]);
  not g__525(w__411 ,in2[18]);
  not g__526(w__58 ,w__336);
  not g__527(w__57 ,w__56);
  not g__528(w__464 ,in2[0]);
  not g__529(w__56 ,w__55);
  not g__530(w__55 ,w__337);
  buf g__531(w__424 ,w__66);
  buf g__532(w__422 ,w__67);
  buf g__533(w__458 ,w__68);
  and g__534(w__54 ,in1[3] ,w__55);
  xnor g__535(out1[25] ,w__136 ,w__201);
  or g__536(w__201 ,w__94 ,w__200);
  xnor g__537(out1[24] ,w__199 ,w__143);
  and g__538(w__200 ,w__77 ,w__199);
  or g__539(w__199 ,w__76 ,w__198);
  xnor g__540(out1[23] ,w__197 ,w__142);
  and g__541(w__198 ,w__96 ,w__197);
  or g__542(w__197 ,w__101 ,w__196);
  xnor g__543(out1[22] ,w__195 ,w__141);
  and g__544(w__196 ,w__91 ,w__195);
  or g__545(w__195 ,w__117 ,w__194);
  xnor g__546(out1[21] ,w__193 ,w__126);
  and g__547(w__194 ,w__100 ,w__193);
  or g__548(w__193 ,w__121 ,w__192);
  xnor g__549(out1[20] ,w__191 ,w__138);
  and g__550(w__192 ,w__98 ,w__191);
  or g__551(w__191 ,w__105 ,w__190);
  xnor g__552(out1[19] ,w__189 ,w__137);
  and g__553(w__190 ,w__99 ,w__189);
  or g__554(w__189 ,w__124 ,w__188);
  xnor g__555(out1[18] ,w__187 ,w__135);
  and g__556(w__188 ,w__92 ,w__187);
  or g__557(w__187 ,w__89 ,w__186);
  xnor g__558(out1[17] ,w__185 ,w__134);
  and g__559(w__186 ,w__83 ,w__185);
  or g__560(w__185 ,w__86 ,w__184);
  xnor g__561(out1[16] ,w__183 ,w__133);
  and g__562(w__184 ,w__79 ,w__183);
  or g__563(w__183 ,w__80 ,w__182);
  xnor g__564(out1[15] ,w__181 ,w__132);
  and g__565(w__182 ,w__82 ,w__181);
  or g__566(w__181 ,w__90 ,w__180);
  xnor g__567(out1[14] ,w__179 ,w__131);
  and g__568(w__180 ,w__95 ,w__179);
  or g__569(w__179 ,w__88 ,w__178);
  xnor g__570(out1[13] ,w__177 ,w__130);
  and g__571(w__178 ,w__78 ,w__177);
  or g__572(w__177 ,w__103 ,w__176);
  xnor g__573(out1[12] ,w__175 ,w__129);
  and g__574(w__176 ,w__113 ,w__175);
  or g__575(w__175 ,w__107 ,w__174);
  xnor g__576(out1[11] ,w__173 ,w__128);
  and g__577(w__174 ,w__116 ,w__173);
  or g__578(w__173 ,w__119 ,w__172);
  xnor g__579(out1[10] ,w__171 ,w__127);
  and g__580(w__172 ,w__110 ,w__171);
  or g__581(w__171 ,w__109 ,w__170);
  xnor g__582(out1[9] ,w__169 ,w__139);
  and g__583(w__170 ,w__115 ,w__169);
  or g__584(w__169 ,w__120 ,w__168);
  xnor g__585(out1[8] ,w__167 ,w__140);
  and g__586(w__168 ,w__87 ,w__167);
  or g__587(w__167 ,w__118 ,w__166);
  xnor g__588(out1[7] ,w__165 ,w__145);
  and g__589(w__166 ,w__93 ,w__165);
  or g__590(w__165 ,w__85 ,w__164);
  xnor g__591(out1[6] ,w__163 ,w__150);
  and g__592(w__164 ,w__84 ,w__163);
  or g__593(w__163 ,w__125 ,w__162);
  xnor g__594(out1[5] ,w__161 ,w__149);
  and g__595(w__162 ,w__81 ,w__161);
  or g__596(w__161 ,w__108 ,w__160);
  xnor g__597(out1[4] ,w__159 ,w__148);
  and g__598(w__160 ,w__112 ,w__159);
  or g__599(w__159 ,w__114 ,w__158);
  xnor g__600(out1[3] ,w__157 ,w__147);
  and g__601(w__158 ,w__123 ,w__157);
  or g__602(w__157 ,w__97 ,w__156);
  xnor g__603(out1[2] ,w__155 ,w__146);
  and g__604(w__156 ,w__106 ,w__155);
  or g__605(w__155 ,w__111 ,w__154);
  xnor g__606(out1[1] ,w__153 ,w__151);
  and g__607(w__154 ,w__122 ,w__153);
  xnor g__608(out1[0] ,w__144 ,w__281);
  or g__609(w__153 ,w__102 ,w__152);
  and g__610(w__152 ,w__282 ,w__104);
  xnor g__611(w__151 ,w__309 ,w__283);
  xnor g__612(w__150 ,w__314 ,w__288);
  xnor g__613(w__149 ,w__313 ,w__287);
  xnor g__614(w__148 ,w__312 ,w__286);
  xnor g__615(w__147 ,w__311 ,w__285);
  xnor g__616(w__146 ,w__310 ,w__284);
  xnor g__617(w__145 ,w__315 ,w__289);
  xnor g__618(w__144 ,w__308 ,w__282);
  xnor g__619(w__143 ,w__332 ,w__306);
  xnor g__620(w__142 ,w__331 ,w__305);
  xnor g__621(w__141 ,w__330 ,w__304);
  xnor g__622(w__140 ,w__316 ,w__290);
  xnor g__623(w__139 ,w__317 ,w__291);
  xnor g__624(w__138 ,w__328 ,w__302);
  xnor g__625(w__137 ,w__327 ,w__301);
  xnor g__626(w__136 ,w__333 ,w__307);
  xnor g__627(w__135 ,w__326 ,w__300);
  xnor g__628(w__134 ,w__325 ,w__299);
  xnor g__629(w__133 ,w__324 ,w__298);
  xnor g__630(w__132 ,w__323 ,w__297);
  xnor g__631(w__131 ,w__322 ,w__296);
  xnor g__632(w__130 ,w__321 ,w__295);
  xnor g__633(w__129 ,w__320 ,w__294);
  xnor g__634(w__128 ,w__319 ,w__293);
  xnor g__635(w__127 ,w__318 ,w__292);
  xnor g__636(w__126 ,w__329 ,w__303);
  and g__637(w__125 ,w__313 ,w__287);
  and g__638(w__124 ,w__326 ,w__300);
  or g__639(w__123 ,w__311 ,w__285);
  or g__640(w__122 ,w__309 ,w__283);
  and g__641(w__121 ,w__328 ,w__302);
  and g__642(w__120 ,w__316 ,w__290);
  and g__643(w__119 ,w__318 ,w__292);
  and g__644(w__118 ,w__315 ,w__289);
  and g__645(w__117 ,w__329 ,w__303);
  or g__646(w__116 ,w__319 ,w__293);
  or g__647(w__115 ,w__317 ,w__291);
  and g__648(w__114 ,w__311 ,w__285);
  or g__649(w__113 ,w__320 ,w__294);
  or g__650(w__112 ,w__312 ,w__286);
  and g__651(w__111 ,w__309 ,w__283);
  or g__652(w__110 ,w__318 ,w__292);
  and g__653(w__109 ,w__317 ,w__291);
  and g__654(w__108 ,w__312 ,w__286);
  and g__655(w__107 ,w__319 ,w__293);
  or g__656(w__106 ,w__310 ,w__284);
  and g__657(w__105 ,w__327 ,w__301);
  or g__658(w__104 ,w__308 ,w__281);
  and g__659(w__103 ,w__320 ,w__294);
  and g__660(w__102 ,w__308 ,w__281);
  and g__661(w__101 ,w__330 ,w__304);
  or g__662(w__100 ,w__329 ,w__303);
  or g__663(w__99 ,w__327 ,w__301);
  or g__664(w__98 ,w__328 ,w__302);
  and g__665(w__97 ,w__310 ,w__284);
  or g__666(w__96 ,w__331 ,w__305);
  or g__667(w__95 ,w__322 ,w__296);
  and g__668(w__94 ,w__332 ,w__306);
  or g__669(w__93 ,w__315 ,w__289);
  or g__670(w__92 ,w__326 ,w__300);
  or g__671(w__91 ,w__330 ,w__304);
  and g__672(w__90 ,w__322 ,w__296);
  and g__673(w__89 ,w__325 ,w__299);
  and g__674(w__88 ,w__321 ,w__295);
  or g__675(w__87 ,w__316 ,w__290);
  and g__676(w__86 ,w__324 ,w__298);
  and g__677(w__85 ,w__314 ,w__288);
  or g__678(w__84 ,w__314 ,w__288);
  or g__679(w__83 ,w__325 ,w__299);
  or g__680(w__82 ,w__323 ,w__297);
  or g__681(w__81 ,w__313 ,w__287);
  and g__682(w__80 ,w__323 ,w__297);
  or g__683(w__79 ,w__324 ,w__298);
  or g__684(w__78 ,w__321 ,w__295);
  or g__685(w__77 ,w__332 ,w__306);
  and g__686(w__76 ,w__331 ,w__305);
  buf g__687(w__225 ,w__344);
  buf g__688(w__218 ,w__345);
endmodule
