module top(in1, in2, in3, in4, in5, out1, out2);
  input [25:0] in1, in5;
  input in2, in3, in4;
  output [25:0] out1, out2;
  wire [25:0] in1, in5;
  wire in2, in3, in4;
  wire [25:0] out1, out2;
  wire add_12_21_n_0, add_12_21_n_1, add_12_21_n_2, add_12_21_n_3, add_12_21_n_4, add_12_21_n_5, add_12_21_n_6, add_12_21_n_7;
  wire add_12_21_n_8, add_12_21_n_9, add_12_21_n_10, add_12_21_n_11, add_12_21_n_12, add_12_21_n_13, add_12_21_n_14, add_12_21_n_15;
  wire add_12_21_n_16, add_12_21_n_17, add_12_21_n_18, add_12_21_n_19, add_12_21_n_20, add_12_21_n_21, add_12_21_n_22, add_12_21_n_23;
  wire add_12_21_n_24, add_12_21_n_25, add_12_21_n_26, add_12_21_n_27, add_12_21_n_28, add_12_21_n_29, add_12_21_n_30, add_12_21_n_31;
  wire add_12_21_n_32, add_12_21_n_33, add_12_21_n_34, add_12_21_n_35, add_12_21_n_36, add_12_21_n_37, add_12_21_n_38, add_12_21_n_39;
  wire add_12_21_n_40, add_12_21_n_41, add_12_21_n_42, add_12_21_n_43, add_12_21_n_44, add_12_21_n_45, add_12_21_n_46, add_12_21_n_47;
  wire add_12_21_n_48, add_12_21_n_49, add_12_21_n_50, add_12_21_n_51, add_12_21_n_52, add_12_21_n_53, add_12_21_n_54, add_12_21_n_55;
  wire add_12_21_n_56, add_12_21_n_57, add_12_21_n_58, add_12_21_n_59, add_12_21_n_60, add_12_21_n_61, add_12_21_n_62, add_12_21_n_63;
  wire add_12_21_n_64, add_12_21_n_65, add_12_21_n_66, add_12_21_n_67, add_12_21_n_68, add_12_21_n_69, add_12_21_n_70, add_12_21_n_71;
  wire add_12_21_n_72, add_12_21_n_73, add_12_21_n_74, add_12_21_n_75, add_12_21_n_76, add_12_21_n_78, add_12_21_n_79, add_12_21_n_81;
  wire add_12_21_n_83, add_12_21_n_84, add_12_21_n_86, add_12_21_n_87, add_12_21_n_89, add_12_21_n_90, add_12_21_n_92, add_12_21_n_93;
  wire add_12_21_n_95, add_12_21_n_96, add_12_21_n_98, add_12_21_n_99, add_12_21_n_101, add_12_21_n_102, add_12_21_n_104, add_12_21_n_105;
  wire add_12_21_n_107, add_12_21_n_108, add_12_21_n_110, add_12_21_n_111, add_12_21_n_113, add_12_21_n_114, add_12_21_n_116, add_12_21_n_117;
  wire add_12_21_n_119, add_12_21_n_120, add_12_21_n_122, add_12_21_n_123, add_12_21_n_125, add_12_21_n_126, add_12_21_n_128, add_12_21_n_129;
  wire add_12_21_n_131, add_12_21_n_132, add_12_21_n_134, add_12_21_n_135, add_12_21_n_137, add_12_21_n_138, add_12_21_n_140, add_12_21_n_141;
  wire add_12_21_n_143, add_12_21_n_144, add_12_21_n_146, add_12_21_n_147, add_12_21_n_149, inc_add_11_21_n_2, inc_add_11_21_n_3, inc_add_11_21_n_4;
  wire inc_add_11_21_n_5, inc_add_11_21_n_6, inc_add_11_21_n_7, inc_add_11_21_n_8, inc_add_11_21_n_9, inc_add_11_21_n_10, inc_add_11_21_n_11, inc_add_11_21_n_12;
  wire inc_add_11_21_n_13, inc_add_11_21_n_14, inc_add_11_21_n_15, inc_add_11_21_n_16, inc_add_11_21_n_17, inc_add_11_21_n_18, inc_add_11_21_n_19, inc_add_11_21_n_20;
  wire inc_add_11_21_n_21, inc_add_11_21_n_22, inc_add_11_21_n_23, inc_add_11_21_n_24, inc_add_11_21_n_25, inc_add_11_21_n_26, inc_add_11_21_n_27, inc_add_11_21_n_28;
  wire inc_add_11_21_n_29, inc_add_11_21_n_30, inc_add_11_21_n_31, inc_add_11_21_n_32, inc_add_11_21_n_34, inc_add_11_21_n_35, inc_add_11_21_n_36, inc_add_11_21_n_38;
  wire inc_add_11_21_n_39, inc_add_11_21_n_40, inc_add_11_21_n_41, inc_add_11_21_n_42, inc_add_11_21_n_43, inc_add_11_21_n_44, inc_add_11_21_n_45, inc_add_11_21_n_47;
  wire inc_add_11_21_n_48, inc_add_11_21_n_51, inc_add_11_21_n_52, inc_add_11_21_n_54, inc_add_11_21_n_55, inc_add_11_21_n_56, inc_add_11_21_n_57, inc_add_11_21_n_58;
  wire inc_add_11_21_n_60, inc_add_11_21_n_61, inc_add_11_21_n_62, inc_add_11_21_n_66, inc_add_11_21_n_67, inc_add_11_21_n_71, inc_add_11_21_n_72, inc_add_11_21_n_74;
  wire inc_add_11_21_n_75, inc_add_11_21_n_76, inc_add_11_21_n_77, inc_add_11_21_n_78, inc_add_11_21_n_80, inc_add_11_21_n_81, inc_add_11_21_n_82, inc_add_11_21_n_83;
  wire inc_add_11_21_n_87, inc_add_11_21_n_88, inc_add_11_21_n_92, inc_add_11_21_n_94, n_0, n_1, n_2, n_3;
  wire n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11;
  wire n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19;
  wire n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27;
  wire n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35;
  wire n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  and g63__2398(n_50 ,out1[25] ,n_0);
  or g64__5107(n_24 ,in3 ,out1[24]);
  or g65__6260(n_23 ,in3 ,out1[22]);
  or g66__4319(n_22 ,in3 ,out1[18]);
  or g67__8428(n_21 ,in3 ,out1[10]);
  or g68__5526(n_20 ,in3 ,out1[9]);
  or g69__6783(n_19 ,in3 ,out1[17]);
  or g70__3680(n_18 ,in3 ,out1[8]);
  or g71__1617(n_17 ,in3 ,out1[7]);
  or g72__2802(n_16 ,in3 ,out1[21]);
  or g73__1705(n_15 ,in3 ,out1[16]);
  or g74__5122(n_14 ,in3 ,out1[6]);
  or g75__8246(n_13 ,in3 ,out1[5]);
  or g76__7098(n_12 ,in3 ,out1[15]);
  or g77__6131(n_11 ,in3 ,out1[4]);
  or g78__1881(n_10 ,in3 ,out1[3]);
  or g79__5115(n_9 ,in3 ,out1[23]);
  or g80__7482(n_8 ,in3 ,out1[20]);
  or g81__4733(n_7 ,in3 ,out1[14]);
  or g82__6161(n_6 ,in3 ,out1[2]);
  or g83__9315(n_5 ,in3 ,out1[1]);
  or g84__9945(n_4 ,in3 ,out1[13]);
  or g85__2883(n_25 ,in3 ,out1[0]);
  or g86__2346(n_3 ,in3 ,out1[19]);
  or g87__1666(n_2 ,in3 ,out1[12]);
  or g88__7410(n_1 ,in3 ,out1[11]);
  not g89(n_0 ,in3);
  buf drc_bufs(n_26 ,n_5);
  buf drc_bufs90(n_36 ,n_1);
  buf drc_bufs91(n_37 ,n_2);
  buf drc_bufs92(n_44 ,n_3);
  buf drc_bufs93(n_38 ,n_4);
  buf drc_bufs94(n_41 ,n_15);
  buf drc_bufs95(n_27 ,n_6);
  buf drc_bufs96(n_39 ,n_7);
  buf drc_bufs97(n_45 ,n_8);
  buf drc_bufs98(n_49 ,n_24);
  buf drc_bufs99(n_28 ,n_10);
  buf drc_bufs100(n_29 ,n_11);
  buf drc_bufs101(n_40 ,n_12);
  buf drc_bufs102(n_30 ,n_13);
  buf drc_bufs103(n_31 ,n_14);
  buf drc_bufs104(n_34 ,n_20);
  buf drc_bufs105(n_46 ,n_16);
  buf drc_bufs106(n_32 ,n_17);
  buf drc_bufs107(n_33 ,n_18);
  buf drc_bufs108(n_42 ,n_19);
  buf drc_bufs109(n_35 ,n_21);
  buf drc_bufs110(n_48 ,n_9);
  buf drc_bufs111(n_43 ,n_22);
  buf drc_bufs112(n_47 ,n_23);
  xnor add_12_21_g534__6417(out2[25] ,add_12_21_n_63 ,add_12_21_n_149);
  or add_12_21_g535__5477(add_12_21_n_149 ,add_12_21_n_14 ,add_12_21_n_147);
  xnor add_12_21_g536__2398(out2[24] ,add_12_21_n_146 ,add_12_21_n_70);
  and add_12_21_g537__5107(add_12_21_n_147 ,add_12_21_n_47 ,add_12_21_n_146);
  or add_12_21_g538__6260(add_12_21_n_146 ,add_12_21_n_27 ,add_12_21_n_144);
  xnor add_12_21_g539__4319(out2[23] ,add_12_21_n_143 ,add_12_21_n_69);
  and add_12_21_g540__8428(add_12_21_n_144 ,add_12_21_n_36 ,add_12_21_n_143);
  or add_12_21_g541__5526(add_12_21_n_143 ,add_12_21_n_40 ,add_12_21_n_141);
  xnor add_12_21_g542__6783(out2[22] ,add_12_21_n_140 ,add_12_21_n_68);
  and add_12_21_g543__3680(add_12_21_n_141 ,add_12_21_n_17 ,add_12_21_n_140);
  or add_12_21_g544__1617(add_12_21_n_140 ,add_12_21_n_15 ,add_12_21_n_138);
  xnor add_12_21_g545__2802(out2[21] ,add_12_21_n_137 ,add_12_21_n_67);
  and add_12_21_g546__1705(add_12_21_n_138 ,add_12_21_n_11 ,add_12_21_n_137);
  or add_12_21_g547__5122(add_12_21_n_137 ,add_12_21_n_21 ,add_12_21_n_135);
  xnor add_12_21_g548__8246(out2[20] ,add_12_21_n_134 ,add_12_21_n_52);
  and add_12_21_g549__7098(add_12_21_n_135 ,add_12_21_n_26 ,add_12_21_n_134);
  or add_12_21_g550__6131(add_12_21_n_134 ,add_12_21_n_22 ,add_12_21_n_132);
  xnor add_12_21_g551__1881(out2[19] ,add_12_21_n_131 ,add_12_21_n_64);
  and add_12_21_g552__5115(add_12_21_n_132 ,add_12_21_n_31 ,add_12_21_n_131);
  or add_12_21_g553__7482(add_12_21_n_131 ,add_12_21_n_25 ,add_12_21_n_129);
  xnor add_12_21_g554__4733(out2[18] ,add_12_21_n_128 ,add_12_21_n_62);
  and add_12_21_g555__6161(add_12_21_n_129 ,add_12_21_n_30 ,add_12_21_n_128);
  or add_12_21_g556__9315(add_12_21_n_128 ,add_12_21_n_42 ,add_12_21_n_126);
  xnor add_12_21_g557__9945(out2[17] ,add_12_21_n_125 ,add_12_21_n_61);
  and add_12_21_g558__2883(add_12_21_n_126 ,add_12_21_n_8 ,add_12_21_n_125);
  or add_12_21_g559__2346(add_12_21_n_125 ,add_12_21_n_4 ,add_12_21_n_123);
  xnor add_12_21_g560__1666(out2[16] ,add_12_21_n_122 ,add_12_21_n_60);
  and add_12_21_g561__7410(add_12_21_n_123 ,add_12_21_n_43 ,add_12_21_n_122);
  or add_12_21_g562__6417(add_12_21_n_122 ,add_12_21_n_6 ,add_12_21_n_120);
  xnor add_12_21_g563__5477(out2[15] ,add_12_21_n_119 ,add_12_21_n_59);
  and add_12_21_g564__2398(add_12_21_n_120 ,add_12_21_n_45 ,add_12_21_n_119);
  or add_12_21_g565__5107(add_12_21_n_119 ,add_12_21_n_29 ,add_12_21_n_117);
  xnor add_12_21_g566__6260(out2[14] ,add_12_21_n_116 ,add_12_21_n_58);
  and add_12_21_g567__4319(add_12_21_n_117 ,add_12_21_n_28 ,add_12_21_n_116);
  or add_12_21_g568__8428(add_12_21_n_116 ,add_12_21_n_50 ,add_12_21_n_114);
  xnor add_12_21_g569__5526(out2[13] ,add_12_21_n_113 ,add_12_21_n_57);
  and add_12_21_g570__6783(add_12_21_n_114 ,add_12_21_n_33 ,add_12_21_n_113);
  or add_12_21_g571__3680(add_12_21_n_113 ,add_12_21_n_32 ,add_12_21_n_111);
  xnor add_12_21_g572__1617(out2[12] ,add_12_21_n_110 ,add_12_21_n_56);
  and add_12_21_g573__2802(add_12_21_n_111 ,add_12_21_n_24 ,add_12_21_n_110);
  or add_12_21_g574__1705(add_12_21_n_110 ,add_12_21_n_41 ,add_12_21_n_108);
  xnor add_12_21_g575__5122(out2[11] ,add_12_21_n_107 ,add_12_21_n_55);
  and add_12_21_g576__8246(add_12_21_n_108 ,add_12_21_n_37 ,add_12_21_n_107);
  or add_12_21_g577__7098(add_12_21_n_107 ,add_12_21_n_23 ,add_12_21_n_105);
  xnor add_12_21_g578__6131(out2[10] ,add_12_21_n_104 ,add_12_21_n_54);
  and add_12_21_g579__1881(add_12_21_n_105 ,add_12_21_n_19 ,add_12_21_n_104);
  or add_12_21_g580__5115(add_12_21_n_104 ,add_12_21_n_38 ,add_12_21_n_102);
  xnor add_12_21_g581__7482(out2[9] ,add_12_21_n_101 ,add_12_21_n_53);
  and add_12_21_g582__4733(add_12_21_n_102 ,add_12_21_n_9 ,add_12_21_n_101);
  or add_12_21_g583__6161(add_12_21_n_101 ,add_12_21_n_3 ,add_12_21_n_99);
  xnor add_12_21_g584__9315(out2[8] ,add_12_21_n_98 ,add_12_21_n_65);
  and add_12_21_g585__9945(add_12_21_n_99 ,add_12_21_n_46 ,add_12_21_n_98);
  or add_12_21_g586__2883(add_12_21_n_98 ,add_12_21_n_5 ,add_12_21_n_96);
  xnor add_12_21_g587__2346(out2[7] ,add_12_21_n_95 ,add_12_21_n_66);
  and add_12_21_g588__1666(add_12_21_n_96 ,add_12_21_n_49 ,add_12_21_n_95);
  or add_12_21_g589__7410(add_12_21_n_95 ,add_12_21_n_16 ,add_12_21_n_93);
  xnor add_12_21_g590__6417(out2[6] ,add_12_21_n_92 ,add_12_21_n_71);
  and add_12_21_g591__5477(add_12_21_n_93 ,add_12_21_n_2 ,add_12_21_n_92);
  or add_12_21_g592__2398(add_12_21_n_92 ,add_12_21_n_12 ,add_12_21_n_90);
  xnor add_12_21_g593__5107(out2[5] ,add_12_21_n_89 ,add_12_21_n_75);
  and add_12_21_g594__6260(add_12_21_n_90 ,add_12_21_n_10 ,add_12_21_n_89);
  or add_12_21_g595__4319(add_12_21_n_89 ,add_12_21_n_13 ,add_12_21_n_87);
  xnor add_12_21_g596__8428(out2[4] ,add_12_21_n_86 ,add_12_21_n_74);
  and add_12_21_g597__5526(add_12_21_n_87 ,add_12_21_n_20 ,add_12_21_n_86);
  or add_12_21_g598__6783(add_12_21_n_86 ,add_12_21_n_48 ,add_12_21_n_84);
  xnor add_12_21_g599__3680(out2[3] ,add_12_21_n_83 ,add_12_21_n_73);
  and add_12_21_g600__1617(add_12_21_n_84 ,add_12_21_n_39 ,add_12_21_n_83);
  or add_12_21_g601__2802(add_12_21_n_83 ,add_12_21_n_44 ,add_12_21_n_81);
  xnor add_12_21_g602__1705(out2[2] ,add_12_21_n_79 ,add_12_21_n_72);
  and add_12_21_g603__5122(add_12_21_n_81 ,add_12_21_n_35 ,add_12_21_n_79);
  xor add_12_21_g604__8246(out2[1] ,add_12_21_n_51 ,add_12_21_n_76);
  or add_12_21_g605__7098(add_12_21_n_79 ,add_12_21_n_7 ,add_12_21_n_78);
  nor add_12_21_g606__6131(add_12_21_n_78 ,add_12_21_n_51 ,add_12_21_n_18);
  and add_12_21_g607__1881(out2[0] ,add_12_21_n_51 ,add_12_21_n_34);
  xnor add_12_21_g608__5115(add_12_21_n_76 ,n_26 ,in5[1]);
  xnor add_12_21_g609__7482(add_12_21_n_75 ,n_30 ,in5[5]);
  xnor add_12_21_g610__4733(add_12_21_n_74 ,n_29 ,in5[4]);
  xnor add_12_21_g611__6161(add_12_21_n_73 ,n_28 ,in5[3]);
  xnor add_12_21_g612__9315(add_12_21_n_72 ,n_27 ,in5[2]);
  xnor add_12_21_g613__9945(add_12_21_n_71 ,n_31 ,in5[6]);
  xnor add_12_21_g614__2883(add_12_21_n_70 ,n_49 ,in5[24]);
  xnor add_12_21_g615__2346(add_12_21_n_69 ,n_48 ,in5[23]);
  xnor add_12_21_g616__1666(add_12_21_n_68 ,n_47 ,in5[22]);
  xnor add_12_21_g617__7410(add_12_21_n_67 ,n_46 ,in5[21]);
  xnor add_12_21_g618__6417(add_12_21_n_66 ,n_32 ,in5[7]);
  xnor add_12_21_g619__5477(add_12_21_n_65 ,n_33 ,in5[8]);
  xnor add_12_21_g620__2398(add_12_21_n_64 ,n_44 ,in5[19]);
  xnor add_12_21_g621__5107(add_12_21_n_63 ,n_50 ,in5[25]);
  xnor add_12_21_g622__6260(add_12_21_n_62 ,n_43 ,in5[18]);
  xnor add_12_21_g623__4319(add_12_21_n_61 ,n_42 ,in5[17]);
  xnor add_12_21_g624__8428(add_12_21_n_60 ,n_41 ,in5[16]);
  xnor add_12_21_g625__5526(add_12_21_n_59 ,n_40 ,in5[15]);
  xnor add_12_21_g626__6783(add_12_21_n_58 ,n_39 ,in5[14]);
  xnor add_12_21_g627__3680(add_12_21_n_57 ,n_38 ,in5[13]);
  xnor add_12_21_g628__1617(add_12_21_n_56 ,n_37 ,in5[12]);
  xnor add_12_21_g629__2802(add_12_21_n_55 ,n_36 ,in5[11]);
  xnor add_12_21_g630__1705(add_12_21_n_54 ,n_35 ,in5[10]);
  xnor add_12_21_g631__5122(add_12_21_n_53 ,n_34 ,in5[9]);
  xnor add_12_21_g632__8246(add_12_21_n_52 ,n_45 ,in5[20]);
  and add_12_21_g633__7098(add_12_21_n_50 ,in5[13] ,n_38);
  or add_12_21_g634__6131(add_12_21_n_49 ,in5[7] ,n_32);
  and add_12_21_g635__1881(add_12_21_n_48 ,in5[3] ,n_28);
  or add_12_21_g636__5115(add_12_21_n_47 ,in5[24] ,n_49);
  or add_12_21_g637__7482(add_12_21_n_46 ,in5[8] ,n_33);
  or add_12_21_g638__4733(add_12_21_n_45 ,in5[15] ,n_40);
  and add_12_21_g639__6161(add_12_21_n_44 ,in5[2] ,n_27);
  or add_12_21_g640__9315(add_12_21_n_43 ,in5[16] ,n_41);
  and add_12_21_g641__9945(add_12_21_n_42 ,in5[17] ,n_42);
  and add_12_21_g642__2883(add_12_21_n_41 ,in5[11] ,n_36);
  and add_12_21_g643__2346(add_12_21_n_40 ,in5[22] ,n_47);
  or add_12_21_g644__1666(add_12_21_n_39 ,in5[3] ,n_28);
  and add_12_21_g645__7410(add_12_21_n_38 ,in5[9] ,n_34);
  or add_12_21_g646__6417(add_12_21_n_37 ,in5[11] ,n_36);
  or add_12_21_g647__5477(add_12_21_n_36 ,in5[23] ,n_48);
  or add_12_21_g648__2398(add_12_21_n_35 ,in5[2] ,n_27);
  or add_12_21_g649__5107(add_12_21_n_34 ,in5[0] ,n_25);
  or add_12_21_g650__6260(add_12_21_n_33 ,in5[13] ,n_38);
  and add_12_21_g651__4319(add_12_21_n_32 ,in5[12] ,n_37);
  or add_12_21_g652__8428(add_12_21_n_31 ,in5[19] ,n_44);
  or add_12_21_g653__5526(add_12_21_n_30 ,in5[18] ,n_43);
  and add_12_21_g654__6783(add_12_21_n_29 ,in5[14] ,n_39);
  or add_12_21_g655__3680(add_12_21_n_28 ,in5[14] ,n_39);
  and add_12_21_g656__1617(add_12_21_n_27 ,in5[23] ,n_48);
  or add_12_21_g657__2802(add_12_21_n_51 ,add_12_21_n_1 ,add_12_21_n_0);
  or add_12_21_g658__1705(add_12_21_n_26 ,in5[20] ,n_45);
  and add_12_21_g659__5122(add_12_21_n_25 ,in5[18] ,n_43);
  or add_12_21_g660__8246(add_12_21_n_24 ,in5[12] ,n_37);
  and add_12_21_g661__7098(add_12_21_n_23 ,in5[10] ,n_35);
  and add_12_21_g662__6131(add_12_21_n_22 ,in5[19] ,n_44);
  and add_12_21_g663__1881(add_12_21_n_21 ,in5[20] ,n_45);
  or add_12_21_g664__5115(add_12_21_n_20 ,in5[4] ,n_29);
  or add_12_21_g665__7482(add_12_21_n_19 ,in5[10] ,n_35);
  nor add_12_21_g666__4733(add_12_21_n_18 ,in5[1] ,n_26);
  or add_12_21_g667__6161(add_12_21_n_17 ,in5[22] ,n_47);
  and add_12_21_g668__9315(add_12_21_n_16 ,in5[6] ,n_31);
  and add_12_21_g669__9945(add_12_21_n_15 ,in5[21] ,n_46);
  and add_12_21_g670__2883(add_12_21_n_14 ,in5[24] ,n_49);
  and add_12_21_g671__2346(add_12_21_n_13 ,in5[4] ,n_29);
  and add_12_21_g672__1666(add_12_21_n_12 ,in5[5] ,n_30);
  or add_12_21_g673__7410(add_12_21_n_11 ,in5[21] ,n_46);
  or add_12_21_g674__6417(add_12_21_n_10 ,in5[5] ,n_30);
  or add_12_21_g675__5477(add_12_21_n_9 ,in5[9] ,n_34);
  or add_12_21_g676__2398(add_12_21_n_8 ,in5[17] ,n_42);
  and add_12_21_g677__5107(add_12_21_n_7 ,in5[1] ,n_26);
  and add_12_21_g678__6260(add_12_21_n_6 ,in5[15] ,n_40);
  and add_12_21_g679__4319(add_12_21_n_5 ,in5[7] ,n_32);
  and add_12_21_g680__8428(add_12_21_n_4 ,in5[16] ,n_41);
  and add_12_21_g681__5526(add_12_21_n_3 ,in5[8] ,n_33);
  or add_12_21_g682__6783(add_12_21_n_2 ,in5[6] ,n_31);
  not add_12_21_g683(add_12_21_n_1 ,in5[0]);
  not add_12_21_g684(add_12_21_n_0 ,n_25);
  xnor inc_add_11_21_g309__3680(out1[25] ,inc_add_11_21_n_94 ,in1[25]);
  xnor inc_add_11_21_g310__1617(out1[24] ,inc_add_11_21_n_92 ,in1[24]);
  or inc_add_11_21_g311__2802(inc_add_11_21_n_94 ,inc_add_11_21_n_20 ,inc_add_11_21_n_92);
  xnor inc_add_11_21_g312__1705(out1[23] ,inc_add_11_21_n_88 ,in1[23]);
  or inc_add_11_21_g313__5122(inc_add_11_21_n_92 ,inc_add_11_21_n_5 ,inc_add_11_21_n_88);
  and inc_add_11_21_g314__8246(out1[22] ,inc_add_11_21_n_87 ,inc_add_11_21_n_88);
  xnor inc_add_11_21_g315__7098(out1[19] ,inc_add_11_21_n_82 ,in1[19]);
  xnor inc_add_11_21_g316__6131(out1[21] ,inc_add_11_21_n_83 ,in1[21]);
  or inc_add_11_21_g317__1881(inc_add_11_21_n_88 ,inc_add_11_21_n_13 ,inc_add_11_21_n_81);
  or inc_add_11_21_g318__5115(inc_add_11_21_n_87 ,in1[22] ,inc_add_11_21_n_80);
  xor inc_add_11_21_g319__7482(out1[20] ,inc_add_11_21_n_75 ,in1[20]);
  xor inc_add_11_21_g320__4733(out1[18] ,inc_add_11_21_n_76 ,in1[18]);
  xnor inc_add_11_21_g321__6161(out1[17] ,inc_add_11_21_n_78 ,in1[17]);
  or inc_add_11_21_g322__9315(inc_add_11_21_n_83 ,inc_add_11_21_n_7 ,inc_add_11_21_n_74);
  or inc_add_11_21_g323__9945(inc_add_11_21_n_82 ,inc_add_11_21_n_8 ,inc_add_11_21_n_77);
  not inc_add_11_21_g324(inc_add_11_21_n_81 ,inc_add_11_21_n_80);
  and inc_add_11_21_g325__2883(inc_add_11_21_n_80 ,inc_add_11_21_n_23 ,inc_add_11_21_n_75);
  xnor inc_add_11_21_g326__2346(out1[16] ,inc_add_11_21_n_72 ,in1[16]);
  or inc_add_11_21_g327__1666(inc_add_11_21_n_78 ,inc_add_11_21_n_2 ,inc_add_11_21_n_72);
  not inc_add_11_21_g328(inc_add_11_21_n_77 ,inc_add_11_21_n_76);
  and inc_add_11_21_g329__7410(inc_add_11_21_n_76 ,inc_add_11_21_n_26 ,inc_add_11_21_n_71);
  not inc_add_11_21_g330(inc_add_11_21_n_74 ,inc_add_11_21_n_75);
  and inc_add_11_21_g331__6417(inc_add_11_21_n_75 ,inc_add_11_21_n_40 ,inc_add_11_21_n_71);
  xnor inc_add_11_21_g332__5477(out1[15] ,inc_add_11_21_n_67 ,in1[15]);
  not inc_add_11_21_g333(inc_add_11_21_n_71 ,inc_add_11_21_n_72);
  or inc_add_11_21_g334__2398(inc_add_11_21_n_72 ,inc_add_11_21_n_10 ,inc_add_11_21_n_66);
  xnor inc_add_11_21_g335__5107(out1[14] ,inc_add_11_21_n_60 ,in1[14]);
  xnor inc_add_11_21_g336__6260(out1[13] ,inc_add_11_21_n_62 ,in1[13]);
  xnor inc_add_11_21_g337__4319(out1[11] ,inc_add_11_21_n_61 ,in1[11]);
  or inc_add_11_21_g338__8428(inc_add_11_21_n_67 ,inc_add_11_21_n_10 ,inc_add_11_21_n_60);
  or inc_add_11_21_g339__5526(inc_add_11_21_n_66 ,inc_add_11_21_n_3 ,inc_add_11_21_n_60);
  xor inc_add_11_21_g340__6783(out1[12] ,inc_add_11_21_n_54 ,in1[12]);
  xor inc_add_11_21_g341__3680(out1[10] ,inc_add_11_21_n_56 ,in1[10]);
  xnor inc_add_11_21_g342__1617(out1[9] ,inc_add_11_21_n_58 ,in1[9]);
  or inc_add_11_21_g343__2802(inc_add_11_21_n_62 ,inc_add_11_21_n_11 ,inc_add_11_21_n_55);
  or inc_add_11_21_g344__1705(inc_add_11_21_n_61 ,inc_add_11_21_n_6 ,inc_add_11_21_n_57);
  or inc_add_11_21_g345__5122(inc_add_11_21_n_60 ,inc_add_11_21_n_27 ,inc_add_11_21_n_55);
  xnor inc_add_11_21_g346__8246(out1[8] ,inc_add_11_21_n_52 ,in1[8]);
  or inc_add_11_21_g347__7098(inc_add_11_21_n_58 ,inc_add_11_21_n_4 ,inc_add_11_21_n_52);
  not inc_add_11_21_g348(inc_add_11_21_n_57 ,inc_add_11_21_n_56);
  and inc_add_11_21_g349__6131(inc_add_11_21_n_56 ,inc_add_11_21_n_29 ,inc_add_11_21_n_51);
  not inc_add_11_21_g350(inc_add_11_21_n_55 ,inc_add_11_21_n_54);
  and inc_add_11_21_g351__1881(inc_add_11_21_n_54 ,inc_add_11_21_n_38 ,inc_add_11_21_n_51);
  xnor inc_add_11_21_g352__5115(out1[7] ,inc_add_11_21_n_48 ,in1[7]);
  not inc_add_11_21_g353(inc_add_11_21_n_51 ,inc_add_11_21_n_52);
  or inc_add_11_21_g354__7482(inc_add_11_21_n_52 ,inc_add_11_21_n_9 ,inc_add_11_21_n_47);
  xnor inc_add_11_21_g355__4733(out1[6] ,inc_add_11_21_n_43 ,inc_add_11_21_n_9);
  xnor inc_add_11_21_g356__6161(out1[5] ,inc_add_11_21_n_45 ,in1[5]);
  or inc_add_11_21_g357__9315(inc_add_11_21_n_48 ,inc_add_11_21_n_9 ,inc_add_11_21_n_44);
  or inc_add_11_21_g358__9945(inc_add_11_21_n_47 ,inc_add_11_21_n_17 ,inc_add_11_21_n_44);
  xnor inc_add_11_21_g359__2883(out1[4] ,inc_add_11_21_n_42 ,in1[4]);
  or inc_add_11_21_g360__2346(inc_add_11_21_n_45 ,inc_add_11_21_n_12 ,inc_add_11_21_n_42);
  not inc_add_11_21_g361(inc_add_11_21_n_44 ,inc_add_11_21_n_43);
  and inc_add_11_21_g362__1666(inc_add_11_21_n_43 ,inc_add_11_21_n_24 ,inc_add_11_21_n_41);
  not inc_add_11_21_g364(inc_add_11_21_n_42 ,inc_add_11_21_n_41);
  and inc_add_11_21_g365__7410(inc_add_11_21_n_41 ,in1[3] ,inc_add_11_21_n_39);
  nor inc_add_11_21_g367__6417(inc_add_11_21_n_40 ,inc_add_11_21_n_8 ,inc_add_11_21_n_35);
  and inc_add_11_21_g369__5477(inc_add_11_21_n_39 ,in1[2] ,inc_add_11_21_n_34);
  nor inc_add_11_21_g370__2398(inc_add_11_21_n_38 ,inc_add_11_21_n_6 ,inc_add_11_21_n_36);
  xnor inc_add_11_21_g371__5107(out1[1] ,inc_add_11_21_n_32 ,in1[1]);
  or inc_add_11_21_g372__6260(inc_add_11_21_n_36 ,inc_add_11_21_n_14 ,inc_add_11_21_n_28);
  or inc_add_11_21_g373__4319(inc_add_11_21_n_35 ,inc_add_11_21_n_16 ,inc_add_11_21_n_25);
  and inc_add_11_21_g375__8428(inc_add_11_21_n_34 ,in1[1] ,inc_add_11_21_n_31);
  and inc_add_11_21_g376__5526(out1[0] ,inc_add_11_21_n_32 ,inc_add_11_21_n_30);
  not inc_add_11_21_g377(inc_add_11_21_n_31 ,inc_add_11_21_n_32);
  or inc_add_11_21_g378__6783(inc_add_11_21_n_32 ,inc_add_11_21_n_22 ,inc_add_11_21_n_21);
  or inc_add_11_21_g379__3680(inc_add_11_21_n_30 ,in1[0] ,in2);
  not inc_add_11_21_g380(inc_add_11_21_n_29 ,inc_add_11_21_n_28);
  or inc_add_11_21_g381__1617(inc_add_11_21_n_28 ,inc_add_11_21_n_18 ,inc_add_11_21_n_4);
  or inc_add_11_21_g382__2802(inc_add_11_21_n_27 ,inc_add_11_21_n_15 ,inc_add_11_21_n_11);
  not inc_add_11_21_g383(inc_add_11_21_n_26 ,inc_add_11_21_n_25);
  or inc_add_11_21_g384__1705(inc_add_11_21_n_25 ,inc_add_11_21_n_19 ,inc_add_11_21_n_2);
  and inc_add_11_21_g385__5122(inc_add_11_21_n_24 ,in1[5] ,in1[4]);
  and inc_add_11_21_g386__8246(inc_add_11_21_n_23 ,in1[21] ,in1[20]);
  not inc_add_11_21_g387(inc_add_11_21_n_22 ,in1[0]);
  not inc_add_11_21_g388(inc_add_11_21_n_21 ,in2);
  not inc_add_11_21_g389(inc_add_11_21_n_20 ,in1[24]);
  not inc_add_11_21_g390(inc_add_11_21_n_19 ,in1[17]);
  not inc_add_11_21_g391(inc_add_11_21_n_18 ,in1[9]);
  not inc_add_11_21_g392(inc_add_11_21_n_17 ,in1[7]);
  not inc_add_11_21_g393(inc_add_11_21_n_16 ,in1[19]);
  not inc_add_11_21_g394(inc_add_11_21_n_15 ,in1[13]);
  not inc_add_11_21_g395(inc_add_11_21_n_14 ,in1[11]);
  not inc_add_11_21_g396(inc_add_11_21_n_13 ,in1[22]);
  not inc_add_11_21_g397(inc_add_11_21_n_12 ,in1[4]);
  not inc_add_11_21_g398(inc_add_11_21_n_11 ,in1[12]);
  not inc_add_11_21_g399(inc_add_11_21_n_10 ,in1[14]);
  not inc_add_11_21_g400(inc_add_11_21_n_9 ,in1[6]);
  not inc_add_11_21_g401(inc_add_11_21_n_8 ,in1[18]);
  not inc_add_11_21_g402(inc_add_11_21_n_7 ,in1[20]);
  not inc_add_11_21_g403(inc_add_11_21_n_6 ,in1[10]);
  not inc_add_11_21_g404(inc_add_11_21_n_5 ,in1[23]);
  not inc_add_11_21_g405(inc_add_11_21_n_4 ,in1[8]);
  not inc_add_11_21_g406(inc_add_11_21_n_3 ,in1[15]);
  not inc_add_11_21_g407(inc_add_11_21_n_2 ,in1[16]);
  xor inc_add_11_21_g2__7098(out1[3] ,inc_add_11_21_n_39 ,in1[3]);
  xor inc_add_11_21_g408__6131(out1[2] ,inc_add_11_21_n_34 ,in1[2]);
endmodule
