module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, out1, out2);
  input [6:0] in1, in2;
  input [15:0] in3, in9, in31;
  input [14:0] in4;
  input in5, in6, in28, in29;
  input [8:0] in7, in12, in16, in20, in24;
  input [12:0] in8, in13, in17, in21, in25;
  input [4:0] in10, in11, in14, in15, in18, in19, in22, in23, in26, in27;
  input [11:0] in30;
  input [3:0] in32, in33;
  output [15:0] out1, out2;
  wire [6:0] in1, in2;
  wire [15:0] in3, in9, in31;
  wire [14:0] in4;
  wire in5, in6, in28, in29;
  wire [8:0] in7, in12, in16, in20, in24;
  wire [12:0] in8, in13, in17, in21, in25;
  wire [4:0] in10, in11, in14, in15, in18, in19, in22, in23, in26, in27;
  wire [11:0] in30;
  wire [3:0] in32, in33;
  wire [15:0] out1, out2;
  wire add_115_23_pad_n_8, add_115_23_pad_n_9, add_115_23_pad_n_10, add_115_23_pad_n_11, add_115_23_pad_n_12, add_115_23_pad_n_13, add_115_23_pad_n_14, add_115_23_pad_n_15;
  wire add_115_23_pad_n_16, add_115_23_pad_n_17, add_115_23_pad_n_18, add_115_23_pad_n_19, add_115_23_pad_n_20, add_115_23_pad_n_21, add_115_23_pad_n_22, add_115_23_pad_n_23;
  wire add_115_23_pad_n_24, add_115_23_pad_n_25, add_115_23_pad_n_26, add_115_23_pad_n_27, add_115_23_pad_n_28, add_115_23_pad_n_29, add_115_23_pad_n_30, add_115_23_pad_n_31;
  wire add_115_23_pad_n_32, add_115_23_pad_n_33, add_115_23_pad_n_34, add_115_23_pad_n_35, add_115_23_pad_n_36, add_115_23_pad_n_37, add_115_23_pad_n_38, add_115_23_pad_n_39;
  wire add_115_23_pad_n_40, add_115_23_pad_n_41, add_115_23_pad_n_42, add_115_23_pad_n_43, add_115_23_pad_n_44, add_115_23_pad_n_45, add_115_23_pad_n_46, add_115_23_pad_n_47;
  wire add_115_23_pad_n_48, add_115_23_pad_n_49, add_115_23_pad_n_50, add_115_23_pad_n_51, add_115_23_pad_n_52, add_115_23_pad_n_53, add_115_23_pad_n_54, add_115_23_pad_n_55;
  wire add_115_23_pad_n_56, add_115_23_pad_n_57, add_115_23_pad_n_58, add_115_23_pad_n_59, add_115_23_pad_n_60, add_115_23_pad_n_62, add_115_23_pad_n_63, add_115_23_pad_n_65;
  wire add_115_23_pad_n_67, add_115_23_pad_n_68, add_115_23_pad_n_70, add_115_23_pad_n_71, add_115_23_pad_n_73, add_115_23_pad_n_74, add_115_23_pad_n_75, add_115_23_pad_n_77;
  wire add_115_23_pad_n_78, add_115_23_pad_n_79, add_115_23_pad_n_80, add_115_23_pad_n_81, add_115_23_pad_n_82, add_115_23_pad_n_83, add_115_23_pad_n_84, add_115_23_pad_n_85;
  wire add_115_23_pad_n_86, add_115_23_pad_n_87, add_115_23_pad_n_88, add_115_23_pad_n_89, add_115_23_pad_n_90, add_115_23_pad_n_91, add_115_23_pad_n_92, add_115_23_pad_n_94;
  wire add_115_23_pad_n_96, csa_tree_add_83_21_pad_groupi_n_0, csa_tree_add_83_21_pad_groupi_n_1, csa_tree_add_83_21_pad_groupi_n_3, csa_tree_add_83_21_pad_groupi_n_4, csa_tree_add_83_21_pad_groupi_n_5, csa_tree_add_83_21_pad_groupi_n_6, csa_tree_add_83_21_pad_groupi_n_12;
  wire csa_tree_add_83_21_pad_groupi_n_13, csa_tree_add_83_21_pad_groupi_n_14, csa_tree_add_83_21_pad_groupi_n_15, csa_tree_add_83_21_pad_groupi_n_16, csa_tree_add_83_21_pad_groupi_n_17, csa_tree_add_83_21_pad_groupi_n_18, csa_tree_add_83_21_pad_groupi_n_19, csa_tree_add_83_21_pad_groupi_n_20;
  wire csa_tree_add_83_21_pad_groupi_n_21, csa_tree_add_83_21_pad_groupi_n_22, csa_tree_add_83_21_pad_groupi_n_23, csa_tree_add_83_21_pad_groupi_n_24, csa_tree_add_83_21_pad_groupi_n_25, csa_tree_add_83_21_pad_groupi_n_26, csa_tree_add_83_21_pad_groupi_n_27, csa_tree_add_83_21_pad_groupi_n_28;
  wire csa_tree_add_83_21_pad_groupi_n_29, csa_tree_add_83_21_pad_groupi_n_30, csa_tree_add_83_21_pad_groupi_n_31, csa_tree_add_83_21_pad_groupi_n_32, csa_tree_add_83_21_pad_groupi_n_33, csa_tree_add_83_21_pad_groupi_n_34, csa_tree_add_83_21_pad_groupi_n_35, csa_tree_add_83_21_pad_groupi_n_36;
  wire csa_tree_add_83_21_pad_groupi_n_37, csa_tree_add_83_21_pad_groupi_n_38, csa_tree_add_83_21_pad_groupi_n_39, csa_tree_add_83_21_pad_groupi_n_40, csa_tree_add_83_21_pad_groupi_n_41, csa_tree_add_83_21_pad_groupi_n_42, csa_tree_add_83_21_pad_groupi_n_43, csa_tree_add_83_21_pad_groupi_n_45;
  wire csa_tree_add_83_21_pad_groupi_n_46, csa_tree_add_83_21_pad_groupi_n_47, csa_tree_add_83_21_pad_groupi_n_48, csa_tree_add_83_21_pad_groupi_n_50, csa_tree_add_83_21_pad_groupi_n_51, csa_tree_add_83_21_pad_groupi_n_52, csa_tree_add_83_21_pad_groupi_n_53, csa_tree_add_83_21_pad_groupi_n_54;
  wire csa_tree_add_83_21_pad_groupi_n_55, csa_tree_add_83_21_pad_groupi_n_56, csa_tree_add_83_21_pad_groupi_n_57, csa_tree_add_83_21_pad_groupi_n_58, csa_tree_add_83_21_pad_groupi_n_59, csa_tree_add_83_21_pad_groupi_n_60, csa_tree_add_83_21_pad_groupi_n_61, csa_tree_add_83_21_pad_groupi_n_62;
  wire csa_tree_add_83_21_pad_groupi_n_64, csa_tree_add_83_21_pad_groupi_n_65, csa_tree_add_83_21_pad_groupi_n_66, csa_tree_add_83_21_pad_groupi_n_67, csa_tree_add_83_21_pad_groupi_n_68, csa_tree_add_83_21_pad_groupi_n_69, csa_tree_add_83_21_pad_groupi_n_70, csa_tree_add_83_21_pad_groupi_n_71;
  wire csa_tree_add_83_21_pad_groupi_n_72, csa_tree_add_83_21_pad_groupi_n_73, csa_tree_add_83_21_pad_groupi_n_74, csa_tree_add_83_21_pad_groupi_n_75, csa_tree_add_83_21_pad_groupi_n_76, csa_tree_add_83_21_pad_groupi_n_77, csa_tree_add_83_21_pad_groupi_n_78, csa_tree_add_83_21_pad_groupi_n_79;
  wire csa_tree_add_83_21_pad_groupi_n_80, csa_tree_add_83_21_pad_groupi_n_82, csa_tree_add_83_21_pad_groupi_n_83, csa_tree_add_83_21_pad_groupi_n_84, csa_tree_add_83_21_pad_groupi_n_85, csa_tree_add_83_21_pad_groupi_n_86, csa_tree_add_83_21_pad_groupi_n_87, csa_tree_add_83_21_pad_groupi_n_88;
  wire csa_tree_add_83_21_pad_groupi_n_89, csa_tree_add_83_21_pad_groupi_n_90, csa_tree_add_83_21_pad_groupi_n_91, csa_tree_add_83_21_pad_groupi_n_92, csa_tree_add_83_21_pad_groupi_n_93, csa_tree_add_83_21_pad_groupi_n_94, csa_tree_add_83_21_pad_groupi_n_95, csa_tree_add_83_21_pad_groupi_n_96;
  wire csa_tree_add_83_21_pad_groupi_n_97, csa_tree_add_83_21_pad_groupi_n_98, csa_tree_add_83_21_pad_groupi_n_99, csa_tree_add_83_21_pad_groupi_n_100, csa_tree_add_83_21_pad_groupi_n_101, csa_tree_add_83_21_pad_groupi_n_102, csa_tree_add_83_21_pad_groupi_n_103, csa_tree_add_83_21_pad_groupi_n_104;
  wire csa_tree_add_83_21_pad_groupi_n_105, csa_tree_add_83_21_pad_groupi_n_106, csa_tree_add_83_21_pad_groupi_n_107, csa_tree_add_83_21_pad_groupi_n_108, csa_tree_add_83_21_pad_groupi_n_109, csa_tree_add_83_21_pad_groupi_n_110, csa_tree_add_83_21_pad_groupi_n_111, csa_tree_add_83_21_pad_groupi_n_112;
  wire csa_tree_add_83_21_pad_groupi_n_113, csa_tree_add_83_21_pad_groupi_n_114, csa_tree_add_83_21_pad_groupi_n_115, csa_tree_add_83_21_pad_groupi_n_116, csa_tree_add_83_21_pad_groupi_n_117, csa_tree_add_83_21_pad_groupi_n_118, csa_tree_add_83_21_pad_groupi_n_119, csa_tree_add_83_21_pad_groupi_n_120;
  wire csa_tree_add_83_21_pad_groupi_n_121, csa_tree_add_83_21_pad_groupi_n_122, csa_tree_add_83_21_pad_groupi_n_123, csa_tree_add_83_21_pad_groupi_n_124, csa_tree_add_83_21_pad_groupi_n_125, csa_tree_add_83_21_pad_groupi_n_126, csa_tree_add_83_21_pad_groupi_n_127, csa_tree_add_83_21_pad_groupi_n_128;
  wire csa_tree_add_83_21_pad_groupi_n_129, csa_tree_add_83_21_pad_groupi_n_130, csa_tree_add_83_21_pad_groupi_n_131, csa_tree_add_83_21_pad_groupi_n_132, csa_tree_add_83_21_pad_groupi_n_133, csa_tree_add_83_21_pad_groupi_n_134, csa_tree_add_83_21_pad_groupi_n_135, csa_tree_add_83_21_pad_groupi_n_136;
  wire csa_tree_add_83_21_pad_groupi_n_137, csa_tree_add_83_21_pad_groupi_n_138, csa_tree_add_83_21_pad_groupi_n_139, csa_tree_add_83_21_pad_groupi_n_140, csa_tree_add_83_21_pad_groupi_n_141, csa_tree_add_83_21_pad_groupi_n_142, csa_tree_add_83_21_pad_groupi_n_143, csa_tree_add_83_21_pad_groupi_n_144;
  wire csa_tree_add_83_21_pad_groupi_n_145, csa_tree_add_83_21_pad_groupi_n_146, csa_tree_add_83_21_pad_groupi_n_147, csa_tree_add_83_21_pad_groupi_n_148, csa_tree_add_83_21_pad_groupi_n_149, csa_tree_add_83_21_pad_groupi_n_150, csa_tree_add_83_21_pad_groupi_n_151, csa_tree_add_83_21_pad_groupi_n_152;
  wire csa_tree_add_83_21_pad_groupi_n_153, csa_tree_add_83_21_pad_groupi_n_154, csa_tree_add_83_21_pad_groupi_n_155, csa_tree_add_83_21_pad_groupi_n_158, csa_tree_add_83_21_pad_groupi_n_159, csa_tree_add_83_21_pad_groupi_n_160, csa_tree_add_83_21_pad_groupi_n_161, csa_tree_add_83_21_pad_groupi_n_162;
  wire csa_tree_add_83_21_pad_groupi_n_163, csa_tree_add_83_21_pad_groupi_n_164, csa_tree_add_83_21_pad_groupi_n_165, csa_tree_add_83_21_pad_groupi_n_166, csa_tree_add_83_21_pad_groupi_n_167, csa_tree_add_83_21_pad_groupi_n_168, csa_tree_add_83_21_pad_groupi_n_169, csa_tree_add_83_21_pad_groupi_n_170;
  wire csa_tree_add_83_21_pad_groupi_n_171, csa_tree_add_83_21_pad_groupi_n_172, csa_tree_add_83_21_pad_groupi_n_173, csa_tree_add_83_21_pad_groupi_n_174, csa_tree_add_83_21_pad_groupi_n_175, csa_tree_add_83_21_pad_groupi_n_176, csa_tree_add_83_21_pad_groupi_n_177, csa_tree_add_83_21_pad_groupi_n_178;
  wire csa_tree_add_83_21_pad_groupi_n_179, csa_tree_add_83_21_pad_groupi_n_180, csa_tree_add_83_21_pad_groupi_n_181, csa_tree_add_83_21_pad_groupi_n_182, csa_tree_add_83_21_pad_groupi_n_183, csa_tree_add_83_21_pad_groupi_n_184, csa_tree_add_83_21_pad_groupi_n_185, csa_tree_add_83_21_pad_groupi_n_186;
  wire csa_tree_add_83_21_pad_groupi_n_187, csa_tree_add_83_21_pad_groupi_n_188, csa_tree_add_83_21_pad_groupi_n_189, csa_tree_add_83_21_pad_groupi_n_190, csa_tree_add_83_21_pad_groupi_n_191, csa_tree_add_83_21_pad_groupi_n_192, csa_tree_add_83_21_pad_groupi_n_193, csa_tree_add_83_21_pad_groupi_n_194;
  wire csa_tree_add_83_21_pad_groupi_n_195, csa_tree_add_83_21_pad_groupi_n_196, csa_tree_add_83_21_pad_groupi_n_197, csa_tree_add_83_21_pad_groupi_n_198, csa_tree_add_83_21_pad_groupi_n_200, csa_tree_add_83_21_pad_groupi_n_201, csa_tree_add_83_21_pad_groupi_n_202, csa_tree_add_83_21_pad_groupi_n_203;
  wire csa_tree_add_83_21_pad_groupi_n_204, csa_tree_add_83_21_pad_groupi_n_205, csa_tree_add_83_21_pad_groupi_n_206, csa_tree_add_83_21_pad_groupi_n_207, csa_tree_add_83_21_pad_groupi_n_208, csa_tree_add_83_21_pad_groupi_n_209, csa_tree_add_83_21_pad_groupi_n_210, csa_tree_add_83_21_pad_groupi_n_211;
  wire csa_tree_add_83_21_pad_groupi_n_212, csa_tree_add_83_21_pad_groupi_n_213, csa_tree_add_83_21_pad_groupi_n_214, csa_tree_add_83_21_pad_groupi_n_215, csa_tree_add_83_21_pad_groupi_n_216, csa_tree_add_83_21_pad_groupi_n_217, csa_tree_add_83_21_pad_groupi_n_218, csa_tree_add_83_21_pad_groupi_n_219;
  wire csa_tree_add_83_21_pad_groupi_n_220, csa_tree_add_83_21_pad_groupi_n_221, csa_tree_add_83_21_pad_groupi_n_222, csa_tree_add_83_21_pad_groupi_n_223, csa_tree_add_83_21_pad_groupi_n_224, csa_tree_add_83_21_pad_groupi_n_225, csa_tree_add_83_21_pad_groupi_n_226, csa_tree_add_83_21_pad_groupi_n_227;
  wire csa_tree_add_83_21_pad_groupi_n_228, csa_tree_add_83_21_pad_groupi_n_229, csa_tree_add_83_21_pad_groupi_n_230, csa_tree_add_83_21_pad_groupi_n_231, csa_tree_add_83_21_pad_groupi_n_232, csa_tree_add_83_21_pad_groupi_n_233, csa_tree_add_83_21_pad_groupi_n_234, csa_tree_add_83_21_pad_groupi_n_235;
  wire csa_tree_add_83_21_pad_groupi_n_236, csa_tree_add_83_21_pad_groupi_n_237, csa_tree_add_83_21_pad_groupi_n_238, csa_tree_add_83_21_pad_groupi_n_239, csa_tree_add_83_21_pad_groupi_n_240, csa_tree_add_83_21_pad_groupi_n_241, csa_tree_add_83_21_pad_groupi_n_242, csa_tree_add_83_21_pad_groupi_n_243;
  wire csa_tree_add_83_21_pad_groupi_n_244, csa_tree_add_83_21_pad_groupi_n_245, csa_tree_add_83_21_pad_groupi_n_246, csa_tree_add_83_21_pad_groupi_n_247, csa_tree_add_83_21_pad_groupi_n_248, csa_tree_add_83_21_pad_groupi_n_249, csa_tree_add_83_21_pad_groupi_n_250, csa_tree_add_83_21_pad_groupi_n_251;
  wire csa_tree_add_83_21_pad_groupi_n_252, csa_tree_add_83_21_pad_groupi_n_253, csa_tree_add_83_21_pad_groupi_n_254, csa_tree_add_83_21_pad_groupi_n_255, csa_tree_add_83_21_pad_groupi_n_256, csa_tree_add_83_21_pad_groupi_n_257, csa_tree_add_83_21_pad_groupi_n_258, csa_tree_add_83_21_pad_groupi_n_259;
  wire csa_tree_add_83_21_pad_groupi_n_260, csa_tree_add_83_21_pad_groupi_n_261, csa_tree_add_83_21_pad_groupi_n_262, csa_tree_add_83_21_pad_groupi_n_263, csa_tree_add_83_21_pad_groupi_n_264, csa_tree_add_83_21_pad_groupi_n_265, csa_tree_add_83_21_pad_groupi_n_266, csa_tree_add_83_21_pad_groupi_n_267;
  wire csa_tree_add_83_21_pad_groupi_n_268, csa_tree_add_83_21_pad_groupi_n_269, csa_tree_add_83_21_pad_groupi_n_270, csa_tree_add_83_21_pad_groupi_n_271, csa_tree_add_83_21_pad_groupi_n_272, csa_tree_add_83_21_pad_groupi_n_273, csa_tree_add_83_21_pad_groupi_n_274, csa_tree_add_83_21_pad_groupi_n_275;
  wire csa_tree_add_83_21_pad_groupi_n_276, csa_tree_add_83_21_pad_groupi_n_277, csa_tree_add_83_21_pad_groupi_n_278, csa_tree_add_83_21_pad_groupi_n_279, csa_tree_add_83_21_pad_groupi_n_280, csa_tree_add_83_21_pad_groupi_n_281, csa_tree_add_83_21_pad_groupi_n_282, csa_tree_add_83_21_pad_groupi_n_283;
  wire csa_tree_add_83_21_pad_groupi_n_284, csa_tree_add_83_21_pad_groupi_n_285, csa_tree_add_83_21_pad_groupi_n_286, csa_tree_add_83_21_pad_groupi_n_287, csa_tree_add_83_21_pad_groupi_n_288, csa_tree_add_83_21_pad_groupi_n_289, csa_tree_add_83_21_pad_groupi_n_290, csa_tree_add_83_21_pad_groupi_n_291;
  wire csa_tree_add_83_21_pad_groupi_n_292, csa_tree_add_83_21_pad_groupi_n_293, csa_tree_add_83_21_pad_groupi_n_294, csa_tree_add_83_21_pad_groupi_n_295, csa_tree_add_83_21_pad_groupi_n_296, csa_tree_add_83_21_pad_groupi_n_297, csa_tree_add_83_21_pad_groupi_n_298, csa_tree_add_83_21_pad_groupi_n_299;
  wire csa_tree_add_83_21_pad_groupi_n_300, csa_tree_add_83_21_pad_groupi_n_301, csa_tree_add_83_21_pad_groupi_n_302, csa_tree_add_83_21_pad_groupi_n_303, csa_tree_add_83_21_pad_groupi_n_304, csa_tree_add_83_21_pad_groupi_n_305, csa_tree_add_83_21_pad_groupi_n_306, csa_tree_add_83_21_pad_groupi_n_307;
  wire csa_tree_add_83_21_pad_groupi_n_308, csa_tree_add_83_21_pad_groupi_n_309, csa_tree_add_83_21_pad_groupi_n_310, csa_tree_add_83_21_pad_groupi_n_311, csa_tree_add_83_21_pad_groupi_n_312, csa_tree_add_83_21_pad_groupi_n_313, csa_tree_add_83_21_pad_groupi_n_314, csa_tree_add_83_21_pad_groupi_n_315;
  wire csa_tree_add_83_21_pad_groupi_n_316, csa_tree_add_83_21_pad_groupi_n_317, csa_tree_add_83_21_pad_groupi_n_318, csa_tree_add_83_21_pad_groupi_n_319, csa_tree_add_83_21_pad_groupi_n_320, csa_tree_add_83_21_pad_groupi_n_321, csa_tree_add_83_21_pad_groupi_n_322, csa_tree_add_83_21_pad_groupi_n_323;
  wire csa_tree_add_83_21_pad_groupi_n_324, csa_tree_add_83_21_pad_groupi_n_325, csa_tree_add_83_21_pad_groupi_n_326, csa_tree_add_83_21_pad_groupi_n_327, csa_tree_add_83_21_pad_groupi_n_328, csa_tree_add_83_21_pad_groupi_n_329, csa_tree_add_83_21_pad_groupi_n_330, csa_tree_add_83_21_pad_groupi_n_331;
  wire csa_tree_add_83_21_pad_groupi_n_332, csa_tree_add_83_21_pad_groupi_n_333, csa_tree_add_83_21_pad_groupi_n_334, csa_tree_add_83_21_pad_groupi_n_335, csa_tree_add_83_21_pad_groupi_n_336, csa_tree_add_83_21_pad_groupi_n_337, csa_tree_add_83_21_pad_groupi_n_338, csa_tree_add_83_21_pad_groupi_n_339;
  wire csa_tree_add_83_21_pad_groupi_n_340, csa_tree_add_83_21_pad_groupi_n_341, csa_tree_add_83_21_pad_groupi_n_342, csa_tree_add_83_21_pad_groupi_n_343, csa_tree_add_83_21_pad_groupi_n_344, csa_tree_add_83_21_pad_groupi_n_345, csa_tree_add_83_21_pad_groupi_n_346, csa_tree_add_83_21_pad_groupi_n_347;
  wire csa_tree_add_83_21_pad_groupi_n_348, csa_tree_add_83_21_pad_groupi_n_349, csa_tree_add_83_21_pad_groupi_n_350, csa_tree_add_83_21_pad_groupi_n_351, csa_tree_add_83_21_pad_groupi_n_352, csa_tree_add_83_21_pad_groupi_n_353, csa_tree_add_83_21_pad_groupi_n_354, csa_tree_add_83_21_pad_groupi_n_355;
  wire csa_tree_add_83_21_pad_groupi_n_356, csa_tree_add_83_21_pad_groupi_n_357, csa_tree_add_83_21_pad_groupi_n_358, csa_tree_add_83_21_pad_groupi_n_359, csa_tree_add_83_21_pad_groupi_n_361, csa_tree_add_83_21_pad_groupi_n_362, csa_tree_add_83_21_pad_groupi_n_363, csa_tree_add_83_21_pad_groupi_n_364;
  wire csa_tree_add_83_21_pad_groupi_n_365, csa_tree_add_83_21_pad_groupi_n_366, csa_tree_add_83_21_pad_groupi_n_367, csa_tree_add_83_21_pad_groupi_n_368, csa_tree_add_83_21_pad_groupi_n_369, csa_tree_add_83_21_pad_groupi_n_370, csa_tree_add_83_21_pad_groupi_n_371, csa_tree_add_83_21_pad_groupi_n_372;
  wire csa_tree_add_83_21_pad_groupi_n_373, csa_tree_add_83_21_pad_groupi_n_374, csa_tree_add_83_21_pad_groupi_n_375, csa_tree_add_83_21_pad_groupi_n_376, csa_tree_add_83_21_pad_groupi_n_377, csa_tree_add_83_21_pad_groupi_n_378, csa_tree_add_83_21_pad_groupi_n_379, csa_tree_add_83_21_pad_groupi_n_380;
  wire csa_tree_add_83_21_pad_groupi_n_381, csa_tree_add_83_21_pad_groupi_n_382, csa_tree_add_83_21_pad_groupi_n_383, csa_tree_add_83_21_pad_groupi_n_384, csa_tree_add_83_21_pad_groupi_n_385, csa_tree_add_83_21_pad_groupi_n_386, csa_tree_add_83_21_pad_groupi_n_387, csa_tree_add_83_21_pad_groupi_n_388;
  wire csa_tree_add_83_21_pad_groupi_n_389, csa_tree_add_83_21_pad_groupi_n_390, csa_tree_add_83_21_pad_groupi_n_391, csa_tree_add_83_21_pad_groupi_n_392, csa_tree_add_83_21_pad_groupi_n_393, csa_tree_add_83_21_pad_groupi_n_394, csa_tree_add_83_21_pad_groupi_n_395, csa_tree_add_83_21_pad_groupi_n_396;
  wire csa_tree_add_83_21_pad_groupi_n_397, csa_tree_add_83_21_pad_groupi_n_398, csa_tree_add_83_21_pad_groupi_n_399, csa_tree_add_83_21_pad_groupi_n_401, csa_tree_add_83_21_pad_groupi_n_402, csa_tree_add_83_21_pad_groupi_n_403, csa_tree_add_83_21_pad_groupi_n_404, csa_tree_add_83_21_pad_groupi_n_406;
  wire csa_tree_add_83_21_pad_groupi_n_409, csa_tree_add_83_21_pad_groupi_n_410, csa_tree_add_83_21_pad_groupi_n_411, csa_tree_add_83_21_pad_groupi_n_412, csa_tree_add_83_21_pad_groupi_n_413, csa_tree_add_83_21_pad_groupi_n_414, csa_tree_add_83_21_pad_groupi_n_415, csa_tree_add_83_21_pad_groupi_n_416;
  wire csa_tree_add_83_21_pad_groupi_n_417, csa_tree_add_83_21_pad_groupi_n_418, csa_tree_add_83_21_pad_groupi_n_419, csa_tree_add_83_21_pad_groupi_n_420, csa_tree_add_83_21_pad_groupi_n_421, csa_tree_add_83_21_pad_groupi_n_422, csa_tree_add_83_21_pad_groupi_n_423, csa_tree_add_83_21_pad_groupi_n_424;
  wire csa_tree_add_83_21_pad_groupi_n_425, csa_tree_add_83_21_pad_groupi_n_426, csa_tree_add_83_21_pad_groupi_n_427, csa_tree_add_83_21_pad_groupi_n_428, csa_tree_add_83_21_pad_groupi_n_429, csa_tree_add_83_21_pad_groupi_n_430, csa_tree_add_83_21_pad_groupi_n_431, csa_tree_add_83_21_pad_groupi_n_432;
  wire csa_tree_add_83_21_pad_groupi_n_433, csa_tree_add_83_21_pad_groupi_n_434, csa_tree_add_83_21_pad_groupi_n_435, csa_tree_add_83_21_pad_groupi_n_438, csa_tree_add_83_21_pad_groupi_n_439, csa_tree_add_83_21_pad_groupi_n_445, csa_tree_add_83_21_pad_groupi_n_455, csa_tree_add_83_21_pad_groupi_n_456;
  wire csa_tree_add_83_21_pad_groupi_n_457, csa_tree_add_83_21_pad_groupi_n_458, csa_tree_add_83_21_pad_groupi_n_459, csa_tree_add_83_21_pad_groupi_n_460, csa_tree_add_83_21_pad_groupi_n_461, csa_tree_add_83_21_pad_groupi_n_462, csa_tree_add_83_21_pad_groupi_n_463, csa_tree_add_83_21_pad_groupi_n_464;
  wire csa_tree_add_83_21_pad_groupi_n_465, csa_tree_add_83_21_pad_groupi_n_466, csa_tree_add_83_21_pad_groupi_n_467, csa_tree_add_83_21_pad_groupi_n_468, csa_tree_add_83_21_pad_groupi_n_469, csa_tree_add_83_21_pad_groupi_n_470, csa_tree_add_83_21_pad_groupi_n_471, csa_tree_add_83_21_pad_groupi_n_472;
  wire csa_tree_add_83_21_pad_groupi_n_473, csa_tree_add_83_21_pad_groupi_n_474, csa_tree_add_83_21_pad_groupi_n_475, csa_tree_add_83_21_pad_groupi_n_476, csa_tree_add_83_21_pad_groupi_n_477, csa_tree_add_83_21_pad_groupi_n_478, csa_tree_add_83_21_pad_groupi_n_479, csa_tree_add_83_21_pad_groupi_n_480;
  wire csa_tree_add_83_21_pad_groupi_n_481, csa_tree_add_83_21_pad_groupi_n_482, csa_tree_add_83_21_pad_groupi_n_483, csa_tree_add_83_21_pad_groupi_n_484, csa_tree_add_83_21_pad_groupi_n_485, csa_tree_add_83_21_pad_groupi_n_486, csa_tree_add_83_21_pad_groupi_n_487, csa_tree_add_83_21_pad_groupi_n_488;
  wire csa_tree_add_83_21_pad_groupi_n_489, csa_tree_add_83_21_pad_groupi_n_490, csa_tree_add_83_21_pad_groupi_n_491, csa_tree_add_83_21_pad_groupi_n_492, csa_tree_add_83_21_pad_groupi_n_493, csa_tree_add_83_21_pad_groupi_n_494, csa_tree_add_83_21_pad_groupi_n_495, csa_tree_add_83_21_pad_groupi_n_496;
  wire csa_tree_add_83_21_pad_groupi_n_497, csa_tree_add_83_21_pad_groupi_n_498, csa_tree_add_83_21_pad_groupi_n_499, csa_tree_add_83_21_pad_groupi_n_500, csa_tree_add_83_21_pad_groupi_n_501, csa_tree_add_83_21_pad_groupi_n_502, csa_tree_add_83_21_pad_groupi_n_503, csa_tree_add_83_21_pad_groupi_n_504;
  wire csa_tree_add_83_21_pad_groupi_n_505, csa_tree_add_83_21_pad_groupi_n_506, csa_tree_add_83_21_pad_groupi_n_507, csa_tree_add_83_21_pad_groupi_n_508, csa_tree_add_83_21_pad_groupi_n_509, csa_tree_add_83_21_pad_groupi_n_510, csa_tree_add_83_21_pad_groupi_n_511, csa_tree_add_83_21_pad_groupi_n_512;
  wire csa_tree_add_83_21_pad_groupi_n_513, csa_tree_add_83_21_pad_groupi_n_514, csa_tree_add_83_21_pad_groupi_n_515, csa_tree_add_83_21_pad_groupi_n_516, csa_tree_add_83_21_pad_groupi_n_517, csa_tree_add_83_21_pad_groupi_n_518, csa_tree_add_83_21_pad_groupi_n_519, csa_tree_add_83_21_pad_groupi_n_520;
  wire csa_tree_add_83_21_pad_groupi_n_521, csa_tree_add_83_21_pad_groupi_n_522, csa_tree_add_83_21_pad_groupi_n_523, csa_tree_add_83_21_pad_groupi_n_524, csa_tree_add_83_21_pad_groupi_n_525, csa_tree_add_83_21_pad_groupi_n_526, csa_tree_add_83_21_pad_groupi_n_527, csa_tree_add_83_21_pad_groupi_n_528;
  wire csa_tree_add_83_21_pad_groupi_n_529, csa_tree_add_83_21_pad_groupi_n_530, csa_tree_add_83_21_pad_groupi_n_531, csa_tree_add_83_21_pad_groupi_n_532, csa_tree_add_83_21_pad_groupi_n_533, csa_tree_add_83_21_pad_groupi_n_534, csa_tree_add_83_21_pad_groupi_n_535, csa_tree_add_83_21_pad_groupi_n_536;
  wire csa_tree_add_83_21_pad_groupi_n_537, csa_tree_add_83_21_pad_groupi_n_538, csa_tree_add_83_21_pad_groupi_n_539, csa_tree_add_83_21_pad_groupi_n_540, csa_tree_add_83_21_pad_groupi_n_541, csa_tree_add_83_21_pad_groupi_n_542, csa_tree_add_83_21_pad_groupi_n_543, csa_tree_add_83_21_pad_groupi_n_544;
  wire csa_tree_add_83_21_pad_groupi_n_545, csa_tree_add_83_21_pad_groupi_n_546, csa_tree_add_83_21_pad_groupi_n_547, csa_tree_add_83_21_pad_groupi_n_548, csa_tree_add_83_21_pad_groupi_n_549, csa_tree_add_83_21_pad_groupi_n_550, csa_tree_add_83_21_pad_groupi_n_551, csa_tree_add_83_21_pad_groupi_n_552;
  wire csa_tree_add_83_21_pad_groupi_n_553, csa_tree_add_83_21_pad_groupi_n_554, csa_tree_add_83_21_pad_groupi_n_555, csa_tree_add_83_21_pad_groupi_n_556, csa_tree_add_83_21_pad_groupi_n_557, csa_tree_add_83_21_pad_groupi_n_559, csa_tree_add_83_21_pad_groupi_n_561, csa_tree_add_83_21_pad_groupi_n_562;
  wire csa_tree_add_83_21_pad_groupi_n_563, csa_tree_add_83_21_pad_groupi_n_564, csa_tree_add_83_21_pad_groupi_n_565, csa_tree_add_83_21_pad_groupi_n_566, csa_tree_add_83_21_pad_groupi_n_567, csa_tree_add_83_21_pad_groupi_n_568, csa_tree_add_83_21_pad_groupi_n_569, csa_tree_add_83_21_pad_groupi_n_570;
  wire csa_tree_add_83_21_pad_groupi_n_572, csa_tree_add_83_21_pad_groupi_n_573, csa_tree_add_83_21_pad_groupi_n_574, csa_tree_add_83_21_pad_groupi_n_575, csa_tree_add_83_21_pad_groupi_n_576, csa_tree_add_83_21_pad_groupi_n_577, csa_tree_add_83_21_pad_groupi_n_578, csa_tree_add_83_21_pad_groupi_n_579;
  wire csa_tree_add_83_21_pad_groupi_n_580, csa_tree_add_83_21_pad_groupi_n_581, csa_tree_add_83_21_pad_groupi_n_582, csa_tree_add_83_21_pad_groupi_n_583, csa_tree_add_83_21_pad_groupi_n_584, csa_tree_add_83_21_pad_groupi_n_586, csa_tree_add_83_21_pad_groupi_n_587, csa_tree_add_83_21_pad_groupi_n_588;
  wire csa_tree_add_83_21_pad_groupi_n_589, csa_tree_add_83_21_pad_groupi_n_590, csa_tree_add_83_21_pad_groupi_n_591, csa_tree_add_83_21_pad_groupi_n_592, csa_tree_add_83_21_pad_groupi_n_593, csa_tree_add_83_21_pad_groupi_n_594, csa_tree_add_83_21_pad_groupi_n_595, csa_tree_add_83_21_pad_groupi_n_598;
  wire csa_tree_add_83_21_pad_groupi_n_599, csa_tree_add_83_21_pad_groupi_n_600, csa_tree_add_83_21_pad_groupi_n_601, csa_tree_add_83_21_pad_groupi_n_602, csa_tree_add_83_21_pad_groupi_n_603, csa_tree_add_83_21_pad_groupi_n_604, csa_tree_add_83_21_pad_groupi_n_605, csa_tree_add_83_21_pad_groupi_n_606;
  wire csa_tree_add_83_21_pad_groupi_n_607, csa_tree_add_83_21_pad_groupi_n_608, csa_tree_add_83_21_pad_groupi_n_609, csa_tree_add_83_21_pad_groupi_n_610, csa_tree_add_83_21_pad_groupi_n_611, csa_tree_add_83_21_pad_groupi_n_612, csa_tree_add_83_21_pad_groupi_n_613, csa_tree_add_83_21_pad_groupi_n_614;
  wire csa_tree_add_83_21_pad_groupi_n_615, csa_tree_add_83_21_pad_groupi_n_616, csa_tree_add_83_21_pad_groupi_n_617, csa_tree_add_83_21_pad_groupi_n_618, csa_tree_add_83_21_pad_groupi_n_619, csa_tree_add_83_21_pad_groupi_n_620, csa_tree_add_83_21_pad_groupi_n_621, csa_tree_add_83_21_pad_groupi_n_622;
  wire csa_tree_add_83_21_pad_groupi_n_623, csa_tree_add_83_21_pad_groupi_n_624, csa_tree_add_83_21_pad_groupi_n_625, csa_tree_add_83_21_pad_groupi_n_626, csa_tree_add_83_21_pad_groupi_n_627, csa_tree_add_83_21_pad_groupi_n_628, csa_tree_add_83_21_pad_groupi_n_629, csa_tree_add_83_21_pad_groupi_n_630;
  wire csa_tree_add_83_21_pad_groupi_n_631, csa_tree_add_83_21_pad_groupi_n_633, csa_tree_add_83_21_pad_groupi_n_634, csa_tree_add_83_21_pad_groupi_n_635, csa_tree_add_83_21_pad_groupi_n_637, csa_tree_add_83_21_pad_groupi_n_638, csa_tree_add_83_21_pad_groupi_n_639, csa_tree_add_83_21_pad_groupi_n_640;
  wire csa_tree_add_83_21_pad_groupi_n_641, csa_tree_add_83_21_pad_groupi_n_642, csa_tree_add_83_21_pad_groupi_n_643, csa_tree_add_83_21_pad_groupi_n_644, csa_tree_add_83_21_pad_groupi_n_645, csa_tree_add_83_21_pad_groupi_n_646, csa_tree_add_83_21_pad_groupi_n_647, csa_tree_add_83_21_pad_groupi_n_648;
  wire csa_tree_add_83_21_pad_groupi_n_649, csa_tree_add_83_21_pad_groupi_n_650, csa_tree_add_83_21_pad_groupi_n_651, csa_tree_add_83_21_pad_groupi_n_652, csa_tree_add_83_21_pad_groupi_n_653, csa_tree_add_83_21_pad_groupi_n_654, csa_tree_add_83_21_pad_groupi_n_655, csa_tree_add_83_21_pad_groupi_n_656;
  wire csa_tree_add_83_21_pad_groupi_n_657, csa_tree_add_83_21_pad_groupi_n_658, csa_tree_add_83_21_pad_groupi_n_659, csa_tree_add_83_21_pad_groupi_n_660, csa_tree_add_83_21_pad_groupi_n_661, csa_tree_add_83_21_pad_groupi_n_662, csa_tree_add_83_21_pad_groupi_n_663, csa_tree_add_83_21_pad_groupi_n_664;
  wire csa_tree_add_83_21_pad_groupi_n_665, csa_tree_add_83_21_pad_groupi_n_666, csa_tree_add_83_21_pad_groupi_n_667, csa_tree_add_83_21_pad_groupi_n_668, csa_tree_add_83_21_pad_groupi_n_669, csa_tree_add_83_21_pad_groupi_n_670, csa_tree_add_83_21_pad_groupi_n_671, csa_tree_add_83_21_pad_groupi_n_672;
  wire csa_tree_add_83_21_pad_groupi_n_673, csa_tree_add_83_21_pad_groupi_n_674, csa_tree_add_83_21_pad_groupi_n_675, csa_tree_add_83_21_pad_groupi_n_676, csa_tree_add_83_21_pad_groupi_n_677, csa_tree_add_83_21_pad_groupi_n_678, csa_tree_add_83_21_pad_groupi_n_679, csa_tree_add_83_21_pad_groupi_n_680;
  wire csa_tree_add_83_21_pad_groupi_n_681, csa_tree_add_83_21_pad_groupi_n_682, csa_tree_add_83_21_pad_groupi_n_683, csa_tree_add_83_21_pad_groupi_n_684, csa_tree_add_83_21_pad_groupi_n_685, csa_tree_add_83_21_pad_groupi_n_686, csa_tree_add_83_21_pad_groupi_n_688, csa_tree_add_83_21_pad_groupi_n_689;
  wire csa_tree_add_83_21_pad_groupi_n_690, csa_tree_add_83_21_pad_groupi_n_691, csa_tree_add_83_21_pad_groupi_n_692, csa_tree_add_83_21_pad_groupi_n_693, csa_tree_add_83_21_pad_groupi_n_694, csa_tree_add_83_21_pad_groupi_n_695, csa_tree_add_83_21_pad_groupi_n_696, csa_tree_add_83_21_pad_groupi_n_697;
  wire csa_tree_add_83_21_pad_groupi_n_698, csa_tree_add_83_21_pad_groupi_n_699, csa_tree_add_83_21_pad_groupi_n_700, csa_tree_add_83_21_pad_groupi_n_702, csa_tree_add_83_21_pad_groupi_n_703, csa_tree_add_83_21_pad_groupi_n_704, csa_tree_add_83_21_pad_groupi_n_705, csa_tree_add_83_21_pad_groupi_n_706;
  wire csa_tree_add_83_21_pad_groupi_n_707, csa_tree_add_83_21_pad_groupi_n_708, csa_tree_add_83_21_pad_groupi_n_709, csa_tree_add_83_21_pad_groupi_n_710, csa_tree_add_83_21_pad_groupi_n_711, csa_tree_add_83_21_pad_groupi_n_712, csa_tree_add_83_21_pad_groupi_n_713, csa_tree_add_83_21_pad_groupi_n_714;
  wire csa_tree_add_83_21_pad_groupi_n_715, csa_tree_add_83_21_pad_groupi_n_716, csa_tree_add_83_21_pad_groupi_n_717, csa_tree_add_83_21_pad_groupi_n_718, csa_tree_add_83_21_pad_groupi_n_719, csa_tree_add_83_21_pad_groupi_n_720, csa_tree_add_83_21_pad_groupi_n_721, csa_tree_add_83_21_pad_groupi_n_722;
  wire csa_tree_add_83_21_pad_groupi_n_723, csa_tree_add_83_21_pad_groupi_n_724, csa_tree_add_83_21_pad_groupi_n_725, csa_tree_add_83_21_pad_groupi_n_726, csa_tree_add_83_21_pad_groupi_n_727, csa_tree_add_83_21_pad_groupi_n_728, csa_tree_add_83_21_pad_groupi_n_729, csa_tree_add_83_21_pad_groupi_n_730;
  wire csa_tree_add_83_21_pad_groupi_n_731, csa_tree_add_83_21_pad_groupi_n_732, csa_tree_add_83_21_pad_groupi_n_733, csa_tree_add_83_21_pad_groupi_n_734, csa_tree_add_83_21_pad_groupi_n_735, csa_tree_add_83_21_pad_groupi_n_736, csa_tree_add_83_21_pad_groupi_n_737, csa_tree_add_83_21_pad_groupi_n_738;
  wire csa_tree_add_83_21_pad_groupi_n_739, csa_tree_add_83_21_pad_groupi_n_740, csa_tree_add_83_21_pad_groupi_n_741, csa_tree_add_83_21_pad_groupi_n_742, csa_tree_add_83_21_pad_groupi_n_743, csa_tree_add_83_21_pad_groupi_n_744, csa_tree_add_83_21_pad_groupi_n_745, csa_tree_add_83_21_pad_groupi_n_746;
  wire csa_tree_add_83_21_pad_groupi_n_747, csa_tree_add_83_21_pad_groupi_n_748, csa_tree_add_83_21_pad_groupi_n_749, csa_tree_add_83_21_pad_groupi_n_750, csa_tree_add_83_21_pad_groupi_n_751, csa_tree_add_83_21_pad_groupi_n_752, csa_tree_add_83_21_pad_groupi_n_753, csa_tree_add_83_21_pad_groupi_n_754;
  wire csa_tree_add_83_21_pad_groupi_n_755, csa_tree_add_83_21_pad_groupi_n_756, csa_tree_add_83_21_pad_groupi_n_757, csa_tree_add_83_21_pad_groupi_n_758, csa_tree_add_83_21_pad_groupi_n_759, csa_tree_add_83_21_pad_groupi_n_760, csa_tree_add_83_21_pad_groupi_n_761, csa_tree_add_83_21_pad_groupi_n_762;
  wire csa_tree_add_83_21_pad_groupi_n_763, csa_tree_add_83_21_pad_groupi_n_764, csa_tree_add_83_21_pad_groupi_n_765, csa_tree_add_83_21_pad_groupi_n_766, csa_tree_add_83_21_pad_groupi_n_767, csa_tree_add_83_21_pad_groupi_n_768, csa_tree_add_83_21_pad_groupi_n_769, csa_tree_add_83_21_pad_groupi_n_770;
  wire csa_tree_add_83_21_pad_groupi_n_771, csa_tree_add_83_21_pad_groupi_n_772, csa_tree_add_83_21_pad_groupi_n_773, csa_tree_add_83_21_pad_groupi_n_774, csa_tree_add_83_21_pad_groupi_n_775, csa_tree_add_83_21_pad_groupi_n_776, csa_tree_add_83_21_pad_groupi_n_777, csa_tree_add_83_21_pad_groupi_n_778;
  wire csa_tree_add_83_21_pad_groupi_n_779, csa_tree_add_83_21_pad_groupi_n_780, csa_tree_add_83_21_pad_groupi_n_781, csa_tree_add_83_21_pad_groupi_n_782, csa_tree_add_83_21_pad_groupi_n_783, csa_tree_add_83_21_pad_groupi_n_784, csa_tree_add_83_21_pad_groupi_n_785, csa_tree_add_83_21_pad_groupi_n_786;
  wire csa_tree_add_83_21_pad_groupi_n_787, csa_tree_add_83_21_pad_groupi_n_788, csa_tree_add_83_21_pad_groupi_n_789, csa_tree_add_83_21_pad_groupi_n_790, csa_tree_add_83_21_pad_groupi_n_791, csa_tree_add_83_21_pad_groupi_n_792, csa_tree_add_83_21_pad_groupi_n_793, csa_tree_add_83_21_pad_groupi_n_794;
  wire csa_tree_add_83_21_pad_groupi_n_795, csa_tree_add_83_21_pad_groupi_n_796, csa_tree_add_83_21_pad_groupi_n_797, csa_tree_add_83_21_pad_groupi_n_798, csa_tree_add_83_21_pad_groupi_n_799, csa_tree_add_83_21_pad_groupi_n_800, csa_tree_add_83_21_pad_groupi_n_801, csa_tree_add_83_21_pad_groupi_n_802;
  wire csa_tree_add_83_21_pad_groupi_n_803, csa_tree_add_83_21_pad_groupi_n_804, csa_tree_add_83_21_pad_groupi_n_805, csa_tree_add_83_21_pad_groupi_n_806, csa_tree_add_83_21_pad_groupi_n_807, csa_tree_add_83_21_pad_groupi_n_808, csa_tree_add_83_21_pad_groupi_n_809, csa_tree_add_83_21_pad_groupi_n_810;
  wire csa_tree_add_83_21_pad_groupi_n_811, csa_tree_add_83_21_pad_groupi_n_812, csa_tree_add_83_21_pad_groupi_n_813, csa_tree_add_83_21_pad_groupi_n_814, csa_tree_add_83_21_pad_groupi_n_815, csa_tree_add_83_21_pad_groupi_n_816, csa_tree_add_83_21_pad_groupi_n_817, csa_tree_add_83_21_pad_groupi_n_818;
  wire csa_tree_add_83_21_pad_groupi_n_819, csa_tree_add_83_21_pad_groupi_n_820, csa_tree_add_83_21_pad_groupi_n_821, csa_tree_add_83_21_pad_groupi_n_822, csa_tree_add_83_21_pad_groupi_n_823, csa_tree_add_83_21_pad_groupi_n_824, csa_tree_add_83_21_pad_groupi_n_825, csa_tree_add_83_21_pad_groupi_n_826;
  wire csa_tree_add_83_21_pad_groupi_n_827, csa_tree_add_83_21_pad_groupi_n_828, csa_tree_add_83_21_pad_groupi_n_829, csa_tree_add_83_21_pad_groupi_n_830, csa_tree_add_83_21_pad_groupi_n_831, csa_tree_add_83_21_pad_groupi_n_832, csa_tree_add_83_21_pad_groupi_n_833, csa_tree_add_83_21_pad_groupi_n_834;
  wire csa_tree_add_83_21_pad_groupi_n_835, csa_tree_add_83_21_pad_groupi_n_836, csa_tree_add_83_21_pad_groupi_n_837, csa_tree_add_83_21_pad_groupi_n_838, csa_tree_add_83_21_pad_groupi_n_839, csa_tree_add_83_21_pad_groupi_n_840, csa_tree_add_83_21_pad_groupi_n_841, csa_tree_add_83_21_pad_groupi_n_842;
  wire csa_tree_add_83_21_pad_groupi_n_843, csa_tree_add_83_21_pad_groupi_n_844, csa_tree_add_83_21_pad_groupi_n_845, csa_tree_add_83_21_pad_groupi_n_846, csa_tree_add_83_21_pad_groupi_n_847, csa_tree_add_83_21_pad_groupi_n_848, csa_tree_add_83_21_pad_groupi_n_849, csa_tree_add_83_21_pad_groupi_n_851;
  wire csa_tree_add_83_21_pad_groupi_n_852, csa_tree_add_83_21_pad_groupi_n_853, csa_tree_add_83_21_pad_groupi_n_854, csa_tree_add_83_21_pad_groupi_n_855, csa_tree_add_83_21_pad_groupi_n_856, csa_tree_add_83_21_pad_groupi_n_857, csa_tree_add_83_21_pad_groupi_n_858, csa_tree_add_83_21_pad_groupi_n_859;
  wire csa_tree_add_83_21_pad_groupi_n_860, csa_tree_add_83_21_pad_groupi_n_861, csa_tree_add_83_21_pad_groupi_n_862, csa_tree_add_83_21_pad_groupi_n_863, csa_tree_add_83_21_pad_groupi_n_864, csa_tree_add_83_21_pad_groupi_n_865, csa_tree_add_83_21_pad_groupi_n_866, csa_tree_add_83_21_pad_groupi_n_867;
  wire csa_tree_add_83_21_pad_groupi_n_868, csa_tree_add_83_21_pad_groupi_n_869, csa_tree_add_83_21_pad_groupi_n_870, csa_tree_add_83_21_pad_groupi_n_871, csa_tree_add_83_21_pad_groupi_n_872, csa_tree_add_83_21_pad_groupi_n_873, csa_tree_add_83_21_pad_groupi_n_874, csa_tree_add_83_21_pad_groupi_n_875;
  wire csa_tree_add_83_21_pad_groupi_n_876, csa_tree_add_83_21_pad_groupi_n_877, csa_tree_add_83_21_pad_groupi_n_878, csa_tree_add_83_21_pad_groupi_n_879, csa_tree_add_83_21_pad_groupi_n_880, csa_tree_add_83_21_pad_groupi_n_881, csa_tree_add_83_21_pad_groupi_n_882, csa_tree_add_83_21_pad_groupi_n_883;
  wire csa_tree_add_83_21_pad_groupi_n_884, csa_tree_add_83_21_pad_groupi_n_885, csa_tree_add_83_21_pad_groupi_n_886, csa_tree_add_83_21_pad_groupi_n_887, csa_tree_add_83_21_pad_groupi_n_888, csa_tree_add_83_21_pad_groupi_n_889, csa_tree_add_83_21_pad_groupi_n_890, csa_tree_add_83_21_pad_groupi_n_891;
  wire csa_tree_add_83_21_pad_groupi_n_892, csa_tree_add_83_21_pad_groupi_n_893, csa_tree_add_83_21_pad_groupi_n_894, csa_tree_add_83_21_pad_groupi_n_895, csa_tree_add_83_21_pad_groupi_n_896, csa_tree_add_83_21_pad_groupi_n_897, csa_tree_add_83_21_pad_groupi_n_898, csa_tree_add_83_21_pad_groupi_n_899;
  wire csa_tree_add_83_21_pad_groupi_n_900, csa_tree_add_83_21_pad_groupi_n_901, csa_tree_add_83_21_pad_groupi_n_902, csa_tree_add_83_21_pad_groupi_n_903, csa_tree_add_83_21_pad_groupi_n_904, csa_tree_add_83_21_pad_groupi_n_905, csa_tree_add_83_21_pad_groupi_n_906, csa_tree_add_83_21_pad_groupi_n_907;
  wire csa_tree_add_83_21_pad_groupi_n_908, csa_tree_add_83_21_pad_groupi_n_909, csa_tree_add_83_21_pad_groupi_n_910, csa_tree_add_83_21_pad_groupi_n_911, csa_tree_add_83_21_pad_groupi_n_912, csa_tree_add_83_21_pad_groupi_n_913, csa_tree_add_83_21_pad_groupi_n_914, csa_tree_add_83_21_pad_groupi_n_915;
  wire csa_tree_add_83_21_pad_groupi_n_916, csa_tree_add_83_21_pad_groupi_n_917, csa_tree_add_83_21_pad_groupi_n_918, csa_tree_add_83_21_pad_groupi_n_919, csa_tree_add_83_21_pad_groupi_n_920, csa_tree_add_83_21_pad_groupi_n_921, csa_tree_add_83_21_pad_groupi_n_922, csa_tree_add_83_21_pad_groupi_n_923;
  wire csa_tree_add_83_21_pad_groupi_n_924, csa_tree_add_83_21_pad_groupi_n_925, csa_tree_add_83_21_pad_groupi_n_926, csa_tree_add_83_21_pad_groupi_n_927, csa_tree_add_83_21_pad_groupi_n_928, csa_tree_add_83_21_pad_groupi_n_929, csa_tree_add_83_21_pad_groupi_n_930, csa_tree_add_83_21_pad_groupi_n_931;
  wire csa_tree_add_83_21_pad_groupi_n_932, csa_tree_add_83_21_pad_groupi_n_933, csa_tree_add_83_21_pad_groupi_n_934, csa_tree_add_83_21_pad_groupi_n_935, csa_tree_add_83_21_pad_groupi_n_936, csa_tree_add_83_21_pad_groupi_n_937, csa_tree_add_83_21_pad_groupi_n_938, csa_tree_add_83_21_pad_groupi_n_939;
  wire csa_tree_add_83_21_pad_groupi_n_940, csa_tree_add_83_21_pad_groupi_n_941, csa_tree_add_83_21_pad_groupi_n_942, csa_tree_add_83_21_pad_groupi_n_943, csa_tree_add_83_21_pad_groupi_n_944, csa_tree_add_83_21_pad_groupi_n_945, csa_tree_add_83_21_pad_groupi_n_946, csa_tree_add_83_21_pad_groupi_n_947;
  wire csa_tree_add_83_21_pad_groupi_n_948, csa_tree_add_83_21_pad_groupi_n_949, csa_tree_add_83_21_pad_groupi_n_950, csa_tree_add_83_21_pad_groupi_n_951, csa_tree_add_83_21_pad_groupi_n_952, csa_tree_add_83_21_pad_groupi_n_953, csa_tree_add_83_21_pad_groupi_n_954, csa_tree_add_83_21_pad_groupi_n_955;
  wire csa_tree_add_83_21_pad_groupi_n_956, csa_tree_add_83_21_pad_groupi_n_957, csa_tree_add_83_21_pad_groupi_n_958, csa_tree_add_83_21_pad_groupi_n_959, csa_tree_add_83_21_pad_groupi_n_960, csa_tree_add_83_21_pad_groupi_n_961, csa_tree_add_83_21_pad_groupi_n_962, csa_tree_add_83_21_pad_groupi_n_963;
  wire csa_tree_add_83_21_pad_groupi_n_964, csa_tree_add_83_21_pad_groupi_n_965, csa_tree_add_83_21_pad_groupi_n_966, csa_tree_add_83_21_pad_groupi_n_967, csa_tree_add_83_21_pad_groupi_n_968, csa_tree_add_83_21_pad_groupi_n_969, csa_tree_add_83_21_pad_groupi_n_970, csa_tree_add_83_21_pad_groupi_n_971;
  wire csa_tree_add_83_21_pad_groupi_n_972, csa_tree_add_83_21_pad_groupi_n_973, csa_tree_add_83_21_pad_groupi_n_974, csa_tree_add_83_21_pad_groupi_n_975, csa_tree_add_83_21_pad_groupi_n_976, csa_tree_add_83_21_pad_groupi_n_977, csa_tree_add_83_21_pad_groupi_n_978, csa_tree_add_83_21_pad_groupi_n_979;
  wire csa_tree_add_83_21_pad_groupi_n_980, csa_tree_add_83_21_pad_groupi_n_981, csa_tree_add_83_21_pad_groupi_n_982, csa_tree_add_83_21_pad_groupi_n_983, csa_tree_add_83_21_pad_groupi_n_984, csa_tree_add_83_21_pad_groupi_n_985, csa_tree_add_83_21_pad_groupi_n_986, csa_tree_add_83_21_pad_groupi_n_987;
  wire csa_tree_add_83_21_pad_groupi_n_988, csa_tree_add_83_21_pad_groupi_n_989, csa_tree_add_83_21_pad_groupi_n_990, csa_tree_add_83_21_pad_groupi_n_991, csa_tree_add_83_21_pad_groupi_n_992, csa_tree_add_83_21_pad_groupi_n_993, csa_tree_add_83_21_pad_groupi_n_994, csa_tree_add_83_21_pad_groupi_n_995;
  wire csa_tree_add_83_21_pad_groupi_n_996, csa_tree_add_83_21_pad_groupi_n_997, csa_tree_add_83_21_pad_groupi_n_998, csa_tree_add_83_21_pad_groupi_n_999, csa_tree_add_83_21_pad_groupi_n_1000, csa_tree_add_83_21_pad_groupi_n_1001, csa_tree_add_83_21_pad_groupi_n_1002, csa_tree_add_83_21_pad_groupi_n_1003;
  wire csa_tree_add_83_21_pad_groupi_n_1004, csa_tree_add_83_21_pad_groupi_n_1005, csa_tree_add_83_21_pad_groupi_n_1006, csa_tree_add_83_21_pad_groupi_n_1007, csa_tree_add_83_21_pad_groupi_n_1008, csa_tree_add_83_21_pad_groupi_n_1009, csa_tree_add_83_21_pad_groupi_n_1010, csa_tree_add_83_21_pad_groupi_n_1011;
  wire csa_tree_add_83_21_pad_groupi_n_1012, csa_tree_add_83_21_pad_groupi_n_1013, csa_tree_add_83_21_pad_groupi_n_1014, csa_tree_add_83_21_pad_groupi_n_1015, csa_tree_add_83_21_pad_groupi_n_1016, csa_tree_add_83_21_pad_groupi_n_1017, csa_tree_add_83_21_pad_groupi_n_1018, csa_tree_add_83_21_pad_groupi_n_1019;
  wire csa_tree_add_83_21_pad_groupi_n_1020, csa_tree_add_83_21_pad_groupi_n_1021, csa_tree_add_83_21_pad_groupi_n_1022, csa_tree_add_83_21_pad_groupi_n_1023, csa_tree_add_83_21_pad_groupi_n_1024, csa_tree_add_83_21_pad_groupi_n_1025, csa_tree_add_83_21_pad_groupi_n_1026, csa_tree_add_83_21_pad_groupi_n_1027;
  wire csa_tree_add_83_21_pad_groupi_n_1028, csa_tree_add_83_21_pad_groupi_n_1029, csa_tree_add_83_21_pad_groupi_n_1030, csa_tree_add_83_21_pad_groupi_n_1031, csa_tree_add_83_21_pad_groupi_n_1032, csa_tree_add_83_21_pad_groupi_n_1033, csa_tree_add_83_21_pad_groupi_n_1034, csa_tree_add_83_21_pad_groupi_n_1035;
  wire csa_tree_add_83_21_pad_groupi_n_1036, csa_tree_add_83_21_pad_groupi_n_1037, csa_tree_add_83_21_pad_groupi_n_1038, csa_tree_add_83_21_pad_groupi_n_1039, csa_tree_add_83_21_pad_groupi_n_1040, csa_tree_add_83_21_pad_groupi_n_1041, csa_tree_add_83_21_pad_groupi_n_1042, csa_tree_add_83_21_pad_groupi_n_1043;
  wire csa_tree_add_83_21_pad_groupi_n_1044, csa_tree_add_83_21_pad_groupi_n_1045, csa_tree_add_83_21_pad_groupi_n_1046, csa_tree_add_83_21_pad_groupi_n_1047, csa_tree_add_83_21_pad_groupi_n_1048, csa_tree_add_83_21_pad_groupi_n_1049, csa_tree_add_83_21_pad_groupi_n_1050, csa_tree_add_83_21_pad_groupi_n_1051;
  wire csa_tree_add_83_21_pad_groupi_n_1052, csa_tree_add_83_21_pad_groupi_n_1053, csa_tree_add_83_21_pad_groupi_n_1054, csa_tree_add_83_21_pad_groupi_n_1055, csa_tree_add_83_21_pad_groupi_n_1056, csa_tree_add_83_21_pad_groupi_n_1057, csa_tree_add_83_21_pad_groupi_n_1058, csa_tree_add_83_21_pad_groupi_n_1059;
  wire csa_tree_add_83_21_pad_groupi_n_1060, csa_tree_add_83_21_pad_groupi_n_1061, csa_tree_add_83_21_pad_groupi_n_1062, csa_tree_add_83_21_pad_groupi_n_1063, csa_tree_add_83_21_pad_groupi_n_1064, csa_tree_add_83_21_pad_groupi_n_1065, csa_tree_add_83_21_pad_groupi_n_1066, csa_tree_add_83_21_pad_groupi_n_1067;
  wire csa_tree_add_83_21_pad_groupi_n_1068, csa_tree_add_83_21_pad_groupi_n_1069, csa_tree_add_83_21_pad_groupi_n_1070, csa_tree_add_83_21_pad_groupi_n_1071, csa_tree_add_83_21_pad_groupi_n_1072, csa_tree_add_83_21_pad_groupi_n_1073, csa_tree_add_83_21_pad_groupi_n_1074, csa_tree_add_83_21_pad_groupi_n_1075;
  wire csa_tree_add_83_21_pad_groupi_n_1076, csa_tree_add_83_21_pad_groupi_n_1077, csa_tree_add_83_21_pad_groupi_n_1078, csa_tree_add_83_21_pad_groupi_n_1079, csa_tree_add_83_21_pad_groupi_n_1080, csa_tree_add_83_21_pad_groupi_n_1081, csa_tree_add_83_21_pad_groupi_n_1082, csa_tree_add_83_21_pad_groupi_n_1083;
  wire csa_tree_add_83_21_pad_groupi_n_1084, csa_tree_add_83_21_pad_groupi_n_1085, csa_tree_add_83_21_pad_groupi_n_1086, csa_tree_add_83_21_pad_groupi_n_1087, csa_tree_add_83_21_pad_groupi_n_1088, csa_tree_add_83_21_pad_groupi_n_1089, csa_tree_add_83_21_pad_groupi_n_1090, csa_tree_add_83_21_pad_groupi_n_1091;
  wire csa_tree_add_83_21_pad_groupi_n_1092, csa_tree_add_83_21_pad_groupi_n_1093, csa_tree_add_83_21_pad_groupi_n_1094, csa_tree_add_83_21_pad_groupi_n_1095, csa_tree_add_83_21_pad_groupi_n_1096, csa_tree_add_83_21_pad_groupi_n_1097, csa_tree_add_83_21_pad_groupi_n_1098, csa_tree_add_83_21_pad_groupi_n_1099;
  wire csa_tree_add_83_21_pad_groupi_n_1100, csa_tree_add_83_21_pad_groupi_n_1101, csa_tree_add_83_21_pad_groupi_n_1102, csa_tree_add_83_21_pad_groupi_n_1103, csa_tree_add_83_21_pad_groupi_n_1104, csa_tree_add_83_21_pad_groupi_n_1105, csa_tree_add_83_21_pad_groupi_n_1106, csa_tree_add_83_21_pad_groupi_n_1107;
  wire csa_tree_add_83_21_pad_groupi_n_1108, csa_tree_add_83_21_pad_groupi_n_1109, csa_tree_add_83_21_pad_groupi_n_1110, csa_tree_add_83_21_pad_groupi_n_1111, csa_tree_add_83_21_pad_groupi_n_1112, csa_tree_add_83_21_pad_groupi_n_1113, csa_tree_add_83_21_pad_groupi_n_1114, csa_tree_add_83_21_pad_groupi_n_1115;
  wire csa_tree_add_83_21_pad_groupi_n_1116, csa_tree_add_83_21_pad_groupi_n_1117, csa_tree_add_83_21_pad_groupi_n_1118, csa_tree_add_83_21_pad_groupi_n_1119, csa_tree_add_83_21_pad_groupi_n_1120, csa_tree_add_83_21_pad_groupi_n_1121, csa_tree_add_83_21_pad_groupi_n_1122, csa_tree_add_83_21_pad_groupi_n_1123;
  wire csa_tree_add_83_21_pad_groupi_n_1124, csa_tree_add_83_21_pad_groupi_n_1125, csa_tree_add_83_21_pad_groupi_n_1126, csa_tree_add_83_21_pad_groupi_n_1127, csa_tree_add_83_21_pad_groupi_n_1128, csa_tree_add_83_21_pad_groupi_n_1129, csa_tree_add_83_21_pad_groupi_n_1130, csa_tree_add_83_21_pad_groupi_n_1131;
  wire csa_tree_add_83_21_pad_groupi_n_1132, csa_tree_add_83_21_pad_groupi_n_1133, csa_tree_add_83_21_pad_groupi_n_1134, csa_tree_add_83_21_pad_groupi_n_1135, csa_tree_add_83_21_pad_groupi_n_1136, csa_tree_add_83_21_pad_groupi_n_1137, csa_tree_add_83_21_pad_groupi_n_1138, csa_tree_add_83_21_pad_groupi_n_1139;
  wire csa_tree_add_83_21_pad_groupi_n_1140, csa_tree_add_83_21_pad_groupi_n_1141, csa_tree_add_83_21_pad_groupi_n_1142, csa_tree_add_83_21_pad_groupi_n_1143, csa_tree_add_83_21_pad_groupi_n_1144, csa_tree_add_83_21_pad_groupi_n_1145, csa_tree_add_83_21_pad_groupi_n_1146, csa_tree_add_83_21_pad_groupi_n_1147;
  wire csa_tree_add_83_21_pad_groupi_n_1148, csa_tree_add_83_21_pad_groupi_n_1149, csa_tree_add_83_21_pad_groupi_n_1150, csa_tree_add_83_21_pad_groupi_n_1151, csa_tree_add_83_21_pad_groupi_n_1152, csa_tree_add_83_21_pad_groupi_n_1153, csa_tree_add_83_21_pad_groupi_n_1154, csa_tree_add_83_21_pad_groupi_n_1155;
  wire csa_tree_add_83_21_pad_groupi_n_1156, csa_tree_add_83_21_pad_groupi_n_1157, csa_tree_add_83_21_pad_groupi_n_1158, csa_tree_add_83_21_pad_groupi_n_1159, csa_tree_add_83_21_pad_groupi_n_1160, csa_tree_add_83_21_pad_groupi_n_1161, csa_tree_add_83_21_pad_groupi_n_1162, csa_tree_add_83_21_pad_groupi_n_1163;
  wire csa_tree_add_83_21_pad_groupi_n_1164, csa_tree_add_83_21_pad_groupi_n_1165, csa_tree_add_83_21_pad_groupi_n_1166, csa_tree_add_83_21_pad_groupi_n_1167, csa_tree_add_83_21_pad_groupi_n_1168, csa_tree_add_83_21_pad_groupi_n_1169, csa_tree_add_83_21_pad_groupi_n_1170, csa_tree_add_83_21_pad_groupi_n_1171;
  wire csa_tree_add_83_21_pad_groupi_n_1172, csa_tree_add_83_21_pad_groupi_n_1173, csa_tree_add_83_21_pad_groupi_n_1174, csa_tree_add_83_21_pad_groupi_n_1175, csa_tree_add_83_21_pad_groupi_n_1176, csa_tree_add_83_21_pad_groupi_n_1177, csa_tree_add_83_21_pad_groupi_n_1178, csa_tree_add_83_21_pad_groupi_n_1179;
  wire csa_tree_add_83_21_pad_groupi_n_1180, csa_tree_add_83_21_pad_groupi_n_1181, csa_tree_add_83_21_pad_groupi_n_1182, csa_tree_add_83_21_pad_groupi_n_1183, csa_tree_add_83_21_pad_groupi_n_1184, csa_tree_add_83_21_pad_groupi_n_1185, csa_tree_add_83_21_pad_groupi_n_1186, csa_tree_add_83_21_pad_groupi_n_1187;
  wire csa_tree_add_83_21_pad_groupi_n_1188, csa_tree_add_83_21_pad_groupi_n_1189, csa_tree_add_83_21_pad_groupi_n_1190, csa_tree_add_83_21_pad_groupi_n_1191, csa_tree_add_83_21_pad_groupi_n_1192, csa_tree_add_83_21_pad_groupi_n_1193, csa_tree_add_83_21_pad_groupi_n_1194, csa_tree_add_83_21_pad_groupi_n_1195;
  wire csa_tree_add_83_21_pad_groupi_n_1196, csa_tree_add_83_21_pad_groupi_n_1197, csa_tree_add_83_21_pad_groupi_n_1198, csa_tree_add_83_21_pad_groupi_n_1199, csa_tree_add_83_21_pad_groupi_n_1200, csa_tree_add_83_21_pad_groupi_n_1201, csa_tree_add_83_21_pad_groupi_n_1202, csa_tree_add_83_21_pad_groupi_n_1203;
  wire csa_tree_add_83_21_pad_groupi_n_1204, csa_tree_add_83_21_pad_groupi_n_1205, csa_tree_add_83_21_pad_groupi_n_1206, csa_tree_add_83_21_pad_groupi_n_1207, csa_tree_add_83_21_pad_groupi_n_1208, csa_tree_add_83_21_pad_groupi_n_1209, csa_tree_add_83_21_pad_groupi_n_1210, csa_tree_add_83_21_pad_groupi_n_1211;
  wire csa_tree_add_83_21_pad_groupi_n_1212, csa_tree_add_83_21_pad_groupi_n_1213, csa_tree_add_83_21_pad_groupi_n_1214, csa_tree_add_83_21_pad_groupi_n_1215, csa_tree_add_83_21_pad_groupi_n_1216, csa_tree_add_83_21_pad_groupi_n_1217, csa_tree_add_83_21_pad_groupi_n_1218, csa_tree_add_83_21_pad_groupi_n_1219;
  wire csa_tree_add_83_21_pad_groupi_n_1220, csa_tree_add_83_21_pad_groupi_n_1221, csa_tree_add_83_21_pad_groupi_n_1222, csa_tree_add_83_21_pad_groupi_n_1223, csa_tree_add_83_21_pad_groupi_n_1224, csa_tree_add_83_21_pad_groupi_n_1225, csa_tree_add_83_21_pad_groupi_n_1226, csa_tree_add_83_21_pad_groupi_n_1227;
  wire csa_tree_add_83_21_pad_groupi_n_1228, csa_tree_add_83_21_pad_groupi_n_1229, csa_tree_add_83_21_pad_groupi_n_1230, csa_tree_add_83_21_pad_groupi_n_1231, csa_tree_add_83_21_pad_groupi_n_1232, csa_tree_add_83_21_pad_groupi_n_1233, csa_tree_add_83_21_pad_groupi_n_1234, csa_tree_add_83_21_pad_groupi_n_1235;
  wire csa_tree_add_83_21_pad_groupi_n_1236, csa_tree_add_83_21_pad_groupi_n_1237, csa_tree_add_83_21_pad_groupi_n_1238, csa_tree_add_83_21_pad_groupi_n_1239, csa_tree_add_83_21_pad_groupi_n_1240, csa_tree_add_83_21_pad_groupi_n_1241, csa_tree_add_83_21_pad_groupi_n_1242, csa_tree_add_83_21_pad_groupi_n_1243;
  wire csa_tree_add_83_21_pad_groupi_n_1244, csa_tree_add_83_21_pad_groupi_n_1245, csa_tree_add_83_21_pad_groupi_n_1246, csa_tree_add_83_21_pad_groupi_n_1247, csa_tree_add_83_21_pad_groupi_n_1248, csa_tree_add_83_21_pad_groupi_n_1249, csa_tree_add_83_21_pad_groupi_n_1250, csa_tree_add_83_21_pad_groupi_n_1251;
  wire csa_tree_add_83_21_pad_groupi_n_1252, csa_tree_add_83_21_pad_groupi_n_1253, csa_tree_add_83_21_pad_groupi_n_1254, csa_tree_add_83_21_pad_groupi_n_1255, csa_tree_add_83_21_pad_groupi_n_1256, csa_tree_add_83_21_pad_groupi_n_1257, csa_tree_add_83_21_pad_groupi_n_1258, csa_tree_add_83_21_pad_groupi_n_1259;
  wire csa_tree_add_83_21_pad_groupi_n_1260, csa_tree_add_83_21_pad_groupi_n_1261, csa_tree_add_83_21_pad_groupi_n_1262, csa_tree_add_83_21_pad_groupi_n_1263, csa_tree_add_83_21_pad_groupi_n_1264, csa_tree_add_83_21_pad_groupi_n_1265, csa_tree_add_83_21_pad_groupi_n_1266, csa_tree_add_83_21_pad_groupi_n_1267;
  wire csa_tree_add_83_21_pad_groupi_n_1268, csa_tree_add_83_21_pad_groupi_n_1269, csa_tree_add_83_21_pad_groupi_n_1270, csa_tree_add_83_21_pad_groupi_n_1271, csa_tree_add_83_21_pad_groupi_n_1272, csa_tree_add_83_21_pad_groupi_n_1273, csa_tree_add_83_21_pad_groupi_n_1274, csa_tree_add_83_21_pad_groupi_n_1275;
  wire csa_tree_add_83_21_pad_groupi_n_1276, csa_tree_add_83_21_pad_groupi_n_1277, csa_tree_add_83_21_pad_groupi_n_1278, csa_tree_add_83_21_pad_groupi_n_1279, csa_tree_add_83_21_pad_groupi_n_1280, csa_tree_add_83_21_pad_groupi_n_1281, csa_tree_add_83_21_pad_groupi_n_1282, csa_tree_add_83_21_pad_groupi_n_1283;
  wire csa_tree_add_83_21_pad_groupi_n_1284, csa_tree_add_83_21_pad_groupi_n_1285, csa_tree_add_83_21_pad_groupi_n_1286, csa_tree_add_83_21_pad_groupi_n_1287, csa_tree_add_83_21_pad_groupi_n_1288, csa_tree_add_83_21_pad_groupi_n_1289, csa_tree_add_83_21_pad_groupi_n_1290, csa_tree_add_83_21_pad_groupi_n_1291;
  wire csa_tree_add_83_21_pad_groupi_n_1292, csa_tree_add_83_21_pad_groupi_n_1293, csa_tree_add_83_21_pad_groupi_n_1294, csa_tree_add_83_21_pad_groupi_n_1295, csa_tree_add_83_21_pad_groupi_n_1296, csa_tree_add_83_21_pad_groupi_n_1297, csa_tree_add_83_21_pad_groupi_n_1298, csa_tree_add_83_21_pad_groupi_n_1299;
  wire csa_tree_add_83_21_pad_groupi_n_1300, csa_tree_add_83_21_pad_groupi_n_1301, csa_tree_add_83_21_pad_groupi_n_1302, csa_tree_add_83_21_pad_groupi_n_1303, csa_tree_add_83_21_pad_groupi_n_1304, csa_tree_add_83_21_pad_groupi_n_1305, csa_tree_add_83_21_pad_groupi_n_1306, csa_tree_add_83_21_pad_groupi_n_1307;
  wire csa_tree_add_83_21_pad_groupi_n_1308, csa_tree_add_83_21_pad_groupi_n_1309, csa_tree_add_83_21_pad_groupi_n_1310, csa_tree_add_83_21_pad_groupi_n_1311, csa_tree_add_83_21_pad_groupi_n_1312, csa_tree_add_83_21_pad_groupi_n_1313, csa_tree_add_83_21_pad_groupi_n_1314, csa_tree_add_83_21_pad_groupi_n_1315;
  wire csa_tree_add_83_21_pad_groupi_n_1316, csa_tree_add_83_21_pad_groupi_n_1317, csa_tree_add_83_21_pad_groupi_n_1318, csa_tree_add_83_21_pad_groupi_n_1319, csa_tree_add_83_21_pad_groupi_n_1320, csa_tree_add_83_21_pad_groupi_n_1321, csa_tree_add_83_21_pad_groupi_n_1322, csa_tree_add_83_21_pad_groupi_n_1323;
  wire csa_tree_add_83_21_pad_groupi_n_1324, csa_tree_add_83_21_pad_groupi_n_1325, csa_tree_add_83_21_pad_groupi_n_1326, csa_tree_add_83_21_pad_groupi_n_1327, csa_tree_add_83_21_pad_groupi_n_1328, csa_tree_add_83_21_pad_groupi_n_1329, csa_tree_add_83_21_pad_groupi_n_1330, csa_tree_add_83_21_pad_groupi_n_1331;
  wire csa_tree_add_83_21_pad_groupi_n_1332, csa_tree_add_83_21_pad_groupi_n_1333, csa_tree_add_83_21_pad_groupi_n_1334, csa_tree_add_83_21_pad_groupi_n_1335, csa_tree_add_83_21_pad_groupi_n_1336, csa_tree_add_83_21_pad_groupi_n_1337, csa_tree_add_83_21_pad_groupi_n_1338, csa_tree_add_83_21_pad_groupi_n_1339;
  wire csa_tree_add_83_21_pad_groupi_n_1340, csa_tree_add_83_21_pad_groupi_n_1341, csa_tree_add_83_21_pad_groupi_n_1342, csa_tree_add_83_21_pad_groupi_n_1343, csa_tree_add_83_21_pad_groupi_n_1344, csa_tree_add_83_21_pad_groupi_n_1345, csa_tree_add_83_21_pad_groupi_n_1346, csa_tree_add_83_21_pad_groupi_n_1347;
  wire csa_tree_add_83_21_pad_groupi_n_1348, csa_tree_add_83_21_pad_groupi_n_1349, csa_tree_add_83_21_pad_groupi_n_1350, csa_tree_add_83_21_pad_groupi_n_1351, csa_tree_add_83_21_pad_groupi_n_1352, csa_tree_add_83_21_pad_groupi_n_1353, csa_tree_add_83_21_pad_groupi_n_1354, csa_tree_add_83_21_pad_groupi_n_1355;
  wire csa_tree_add_83_21_pad_groupi_n_1356, csa_tree_add_83_21_pad_groupi_n_1357, csa_tree_add_83_21_pad_groupi_n_1358, csa_tree_add_83_21_pad_groupi_n_1359, csa_tree_add_83_21_pad_groupi_n_1360, csa_tree_add_83_21_pad_groupi_n_1361, csa_tree_add_83_21_pad_groupi_n_1362, csa_tree_add_83_21_pad_groupi_n_1363;
  wire csa_tree_add_83_21_pad_groupi_n_1364, csa_tree_add_83_21_pad_groupi_n_1365, csa_tree_add_83_21_pad_groupi_n_1366, csa_tree_add_83_21_pad_groupi_n_1367, csa_tree_add_83_21_pad_groupi_n_1368, csa_tree_add_83_21_pad_groupi_n_1369, csa_tree_add_83_21_pad_groupi_n_1370, csa_tree_add_83_21_pad_groupi_n_1371;
  wire csa_tree_add_83_21_pad_groupi_n_1372, csa_tree_add_83_21_pad_groupi_n_1373, csa_tree_add_83_21_pad_groupi_n_1374, csa_tree_add_83_21_pad_groupi_n_1375, csa_tree_add_83_21_pad_groupi_n_1376, csa_tree_add_83_21_pad_groupi_n_1377, csa_tree_add_83_21_pad_groupi_n_1378, csa_tree_add_83_21_pad_groupi_n_1379;
  wire csa_tree_add_83_21_pad_groupi_n_1380, csa_tree_add_83_21_pad_groupi_n_1381, csa_tree_add_83_21_pad_groupi_n_1382, csa_tree_add_83_21_pad_groupi_n_1383, csa_tree_add_83_21_pad_groupi_n_1384, csa_tree_add_83_21_pad_groupi_n_1385, csa_tree_add_83_21_pad_groupi_n_1386, csa_tree_add_83_21_pad_groupi_n_1387;
  wire csa_tree_add_83_21_pad_groupi_n_1388, csa_tree_add_83_21_pad_groupi_n_1389, csa_tree_add_83_21_pad_groupi_n_1390, csa_tree_add_83_21_pad_groupi_n_1391, csa_tree_add_83_21_pad_groupi_n_1392, csa_tree_add_83_21_pad_groupi_n_1393, csa_tree_add_83_21_pad_groupi_n_1394, csa_tree_add_83_21_pad_groupi_n_1395;
  wire csa_tree_add_83_21_pad_groupi_n_1396, csa_tree_add_83_21_pad_groupi_n_1397, csa_tree_add_83_21_pad_groupi_n_1398, csa_tree_add_83_21_pad_groupi_n_1399, csa_tree_add_83_21_pad_groupi_n_1400, csa_tree_add_83_21_pad_groupi_n_1401, csa_tree_add_83_21_pad_groupi_n_1402, csa_tree_add_83_21_pad_groupi_n_1403;
  wire csa_tree_add_83_21_pad_groupi_n_1404, csa_tree_add_83_21_pad_groupi_n_1405, csa_tree_add_83_21_pad_groupi_n_1406, csa_tree_add_83_21_pad_groupi_n_1407, csa_tree_add_83_21_pad_groupi_n_1408, csa_tree_add_83_21_pad_groupi_n_1409, csa_tree_add_83_21_pad_groupi_n_1410, csa_tree_add_83_21_pad_groupi_n_1411;
  wire csa_tree_add_83_21_pad_groupi_n_1412, csa_tree_add_83_21_pad_groupi_n_1413, csa_tree_add_83_21_pad_groupi_n_1414, csa_tree_add_83_21_pad_groupi_n_1415, csa_tree_add_83_21_pad_groupi_n_1416, csa_tree_add_83_21_pad_groupi_n_1417, csa_tree_add_83_21_pad_groupi_n_1418, csa_tree_add_83_21_pad_groupi_n_1419;
  wire csa_tree_add_83_21_pad_groupi_n_1420, csa_tree_add_83_21_pad_groupi_n_1421, csa_tree_add_83_21_pad_groupi_n_1422, csa_tree_add_83_21_pad_groupi_n_1423, csa_tree_add_83_21_pad_groupi_n_1424, csa_tree_add_83_21_pad_groupi_n_1425, csa_tree_add_83_21_pad_groupi_n_1426, csa_tree_add_83_21_pad_groupi_n_1427;
  wire csa_tree_add_83_21_pad_groupi_n_1428, csa_tree_add_83_21_pad_groupi_n_1429, csa_tree_add_83_21_pad_groupi_n_1430, csa_tree_add_83_21_pad_groupi_n_1431, csa_tree_add_83_21_pad_groupi_n_1432, csa_tree_add_83_21_pad_groupi_n_1433, csa_tree_add_83_21_pad_groupi_n_1434, csa_tree_add_83_21_pad_groupi_n_1435;
  wire csa_tree_add_83_21_pad_groupi_n_1436, csa_tree_add_83_21_pad_groupi_n_1437, csa_tree_add_83_21_pad_groupi_n_1438, csa_tree_add_83_21_pad_groupi_n_1439, csa_tree_add_83_21_pad_groupi_n_1440, csa_tree_add_83_21_pad_groupi_n_1441, csa_tree_add_83_21_pad_groupi_n_1442, csa_tree_add_83_21_pad_groupi_n_1443;
  wire csa_tree_add_83_21_pad_groupi_n_1444, csa_tree_add_83_21_pad_groupi_n_1445, csa_tree_add_83_21_pad_groupi_n_1446, csa_tree_add_83_21_pad_groupi_n_1447, csa_tree_add_83_21_pad_groupi_n_1448, csa_tree_add_83_21_pad_groupi_n_1449, csa_tree_add_83_21_pad_groupi_n_1450, csa_tree_add_83_21_pad_groupi_n_1451;
  wire csa_tree_add_83_21_pad_groupi_n_1452, csa_tree_add_83_21_pad_groupi_n_1453, csa_tree_add_83_21_pad_groupi_n_1454, csa_tree_add_83_21_pad_groupi_n_1455, csa_tree_add_83_21_pad_groupi_n_1456, csa_tree_add_83_21_pad_groupi_n_1457, csa_tree_add_83_21_pad_groupi_n_1458, csa_tree_add_83_21_pad_groupi_n_1459;
  wire csa_tree_add_83_21_pad_groupi_n_1460, csa_tree_add_83_21_pad_groupi_n_1461, csa_tree_add_83_21_pad_groupi_n_1462, csa_tree_add_83_21_pad_groupi_n_1463, csa_tree_add_83_21_pad_groupi_n_1464, csa_tree_add_83_21_pad_groupi_n_1465, csa_tree_add_83_21_pad_groupi_n_1466, csa_tree_add_83_21_pad_groupi_n_1467;
  wire csa_tree_add_83_21_pad_groupi_n_1468, csa_tree_add_83_21_pad_groupi_n_1469, csa_tree_add_83_21_pad_groupi_n_1470, csa_tree_add_83_21_pad_groupi_n_1471, csa_tree_add_83_21_pad_groupi_n_1472, csa_tree_add_83_21_pad_groupi_n_1473, csa_tree_add_83_21_pad_groupi_n_1474, csa_tree_add_83_21_pad_groupi_n_1475;
  wire csa_tree_add_83_21_pad_groupi_n_1476, csa_tree_add_83_21_pad_groupi_n_1477, csa_tree_add_83_21_pad_groupi_n_1478, csa_tree_add_83_21_pad_groupi_n_1479, csa_tree_add_83_21_pad_groupi_n_1480, csa_tree_add_83_21_pad_groupi_n_1481, csa_tree_add_83_21_pad_groupi_n_1482, csa_tree_add_83_21_pad_groupi_n_1483;
  wire csa_tree_add_83_21_pad_groupi_n_1484, csa_tree_add_83_21_pad_groupi_n_1485, csa_tree_add_83_21_pad_groupi_n_1486, csa_tree_add_83_21_pad_groupi_n_1487, csa_tree_add_83_21_pad_groupi_n_1488, csa_tree_add_83_21_pad_groupi_n_1489, csa_tree_add_83_21_pad_groupi_n_1490, csa_tree_add_83_21_pad_groupi_n_1491;
  wire csa_tree_add_83_21_pad_groupi_n_1492, csa_tree_add_83_21_pad_groupi_n_1493, csa_tree_add_83_21_pad_groupi_n_1494, csa_tree_add_83_21_pad_groupi_n_1495, csa_tree_add_83_21_pad_groupi_n_1496, csa_tree_add_83_21_pad_groupi_n_1497, csa_tree_add_83_21_pad_groupi_n_1498, csa_tree_add_83_21_pad_groupi_n_1499;
  wire csa_tree_add_83_21_pad_groupi_n_1500, csa_tree_add_83_21_pad_groupi_n_1501, csa_tree_add_83_21_pad_groupi_n_1502, csa_tree_add_83_21_pad_groupi_n_1503, csa_tree_add_83_21_pad_groupi_n_1505, csa_tree_add_83_21_pad_groupi_n_1506, csa_tree_add_83_21_pad_groupi_n_1507, csa_tree_add_83_21_pad_groupi_n_1508;
  wire csa_tree_add_83_21_pad_groupi_n_1509, csa_tree_add_83_21_pad_groupi_n_1510, csa_tree_add_83_21_pad_groupi_n_1511, csa_tree_add_83_21_pad_groupi_n_1512, csa_tree_add_83_21_pad_groupi_n_1513, csa_tree_add_83_21_pad_groupi_n_1514, csa_tree_add_83_21_pad_groupi_n_1515, csa_tree_add_83_21_pad_groupi_n_1516;
  wire csa_tree_add_83_21_pad_groupi_n_1517, csa_tree_add_83_21_pad_groupi_n_1518, csa_tree_add_83_21_pad_groupi_n_1519, csa_tree_add_83_21_pad_groupi_n_1520, csa_tree_add_83_21_pad_groupi_n_1521, csa_tree_add_83_21_pad_groupi_n_1522, csa_tree_add_83_21_pad_groupi_n_1523, csa_tree_add_83_21_pad_groupi_n_1524;
  wire csa_tree_add_83_21_pad_groupi_n_1525, csa_tree_add_83_21_pad_groupi_n_1526, csa_tree_add_83_21_pad_groupi_n_1527, csa_tree_add_83_21_pad_groupi_n_1529, csa_tree_add_83_21_pad_groupi_n_1530, csa_tree_add_83_21_pad_groupi_n_1532, csa_tree_add_83_21_pad_groupi_n_1533, csa_tree_add_83_21_pad_groupi_n_1534;
  wire csa_tree_add_83_21_pad_groupi_n_1535, csa_tree_add_83_21_pad_groupi_n_1537, csa_tree_add_83_21_pad_groupi_n_1538, csa_tree_add_83_21_pad_groupi_n_1539, csa_tree_add_83_21_pad_groupi_n_1540, csa_tree_add_83_21_pad_groupi_n_1542, csa_tree_add_83_21_pad_groupi_n_1543, csa_tree_add_83_21_pad_groupi_n_1544;
  wire csa_tree_add_83_21_pad_groupi_n_1546, csa_tree_add_83_21_pad_groupi_n_1547, csa_tree_add_83_21_pad_groupi_n_1549, csa_tree_add_83_21_pad_groupi_n_1550, csa_tree_add_83_21_pad_groupi_n_1552, csa_tree_add_83_21_pad_groupi_n_1553, csa_tree_add_83_21_pad_groupi_n_1555, csa_tree_add_83_21_pad_groupi_n_1556;
  wire csa_tree_add_83_21_pad_groupi_n_1558, csa_tree_add_89_22_pad_groupi_n_0, csa_tree_add_89_22_pad_groupi_n_1, csa_tree_add_89_22_pad_groupi_n_2, csa_tree_add_89_22_pad_groupi_n_3, csa_tree_add_89_22_pad_groupi_n_4, csa_tree_add_89_22_pad_groupi_n_5, csa_tree_add_89_22_pad_groupi_n_6;
  wire csa_tree_add_89_22_pad_groupi_n_12, csa_tree_add_89_22_pad_groupi_n_13, csa_tree_add_89_22_pad_groupi_n_14, csa_tree_add_89_22_pad_groupi_n_15, csa_tree_add_89_22_pad_groupi_n_16, csa_tree_add_89_22_pad_groupi_n_17, csa_tree_add_89_22_pad_groupi_n_18, csa_tree_add_89_22_pad_groupi_n_19;
  wire csa_tree_add_89_22_pad_groupi_n_20, csa_tree_add_89_22_pad_groupi_n_21, csa_tree_add_89_22_pad_groupi_n_22, csa_tree_add_89_22_pad_groupi_n_23, csa_tree_add_89_22_pad_groupi_n_24, csa_tree_add_89_22_pad_groupi_n_25, csa_tree_add_89_22_pad_groupi_n_26, csa_tree_add_89_22_pad_groupi_n_27;
  wire csa_tree_add_89_22_pad_groupi_n_28, csa_tree_add_89_22_pad_groupi_n_29, csa_tree_add_89_22_pad_groupi_n_30, csa_tree_add_89_22_pad_groupi_n_31, csa_tree_add_89_22_pad_groupi_n_32, csa_tree_add_89_22_pad_groupi_n_33, csa_tree_add_89_22_pad_groupi_n_34, csa_tree_add_89_22_pad_groupi_n_35;
  wire csa_tree_add_89_22_pad_groupi_n_36, csa_tree_add_89_22_pad_groupi_n_37, csa_tree_add_89_22_pad_groupi_n_38, csa_tree_add_89_22_pad_groupi_n_39, csa_tree_add_89_22_pad_groupi_n_40, csa_tree_add_89_22_pad_groupi_n_41, csa_tree_add_89_22_pad_groupi_n_42, csa_tree_add_89_22_pad_groupi_n_43;
  wire csa_tree_add_89_22_pad_groupi_n_45, csa_tree_add_89_22_pad_groupi_n_46, csa_tree_add_89_22_pad_groupi_n_47, csa_tree_add_89_22_pad_groupi_n_48, csa_tree_add_89_22_pad_groupi_n_50, csa_tree_add_89_22_pad_groupi_n_51, csa_tree_add_89_22_pad_groupi_n_52, csa_tree_add_89_22_pad_groupi_n_53;
  wire csa_tree_add_89_22_pad_groupi_n_54, csa_tree_add_89_22_pad_groupi_n_55, csa_tree_add_89_22_pad_groupi_n_56, csa_tree_add_89_22_pad_groupi_n_57, csa_tree_add_89_22_pad_groupi_n_58, csa_tree_add_89_22_pad_groupi_n_59, csa_tree_add_89_22_pad_groupi_n_60, csa_tree_add_89_22_pad_groupi_n_61;
  wire csa_tree_add_89_22_pad_groupi_n_62, csa_tree_add_89_22_pad_groupi_n_64, csa_tree_add_89_22_pad_groupi_n_65, csa_tree_add_89_22_pad_groupi_n_66, csa_tree_add_89_22_pad_groupi_n_67, csa_tree_add_89_22_pad_groupi_n_68, csa_tree_add_89_22_pad_groupi_n_69, csa_tree_add_89_22_pad_groupi_n_70;
  wire csa_tree_add_89_22_pad_groupi_n_71, csa_tree_add_89_22_pad_groupi_n_72, csa_tree_add_89_22_pad_groupi_n_73, csa_tree_add_89_22_pad_groupi_n_74, csa_tree_add_89_22_pad_groupi_n_75, csa_tree_add_89_22_pad_groupi_n_76, csa_tree_add_89_22_pad_groupi_n_77, csa_tree_add_89_22_pad_groupi_n_78;
  wire csa_tree_add_89_22_pad_groupi_n_79, csa_tree_add_89_22_pad_groupi_n_80, csa_tree_add_89_22_pad_groupi_n_82, csa_tree_add_89_22_pad_groupi_n_83, csa_tree_add_89_22_pad_groupi_n_84, csa_tree_add_89_22_pad_groupi_n_85, csa_tree_add_89_22_pad_groupi_n_86, csa_tree_add_89_22_pad_groupi_n_87;
  wire csa_tree_add_89_22_pad_groupi_n_88, csa_tree_add_89_22_pad_groupi_n_89, csa_tree_add_89_22_pad_groupi_n_90, csa_tree_add_89_22_pad_groupi_n_91, csa_tree_add_89_22_pad_groupi_n_92, csa_tree_add_89_22_pad_groupi_n_93, csa_tree_add_89_22_pad_groupi_n_94, csa_tree_add_89_22_pad_groupi_n_95;
  wire csa_tree_add_89_22_pad_groupi_n_96, csa_tree_add_89_22_pad_groupi_n_97, csa_tree_add_89_22_pad_groupi_n_98, csa_tree_add_89_22_pad_groupi_n_99, csa_tree_add_89_22_pad_groupi_n_100, csa_tree_add_89_22_pad_groupi_n_101, csa_tree_add_89_22_pad_groupi_n_102, csa_tree_add_89_22_pad_groupi_n_103;
  wire csa_tree_add_89_22_pad_groupi_n_104, csa_tree_add_89_22_pad_groupi_n_105, csa_tree_add_89_22_pad_groupi_n_106, csa_tree_add_89_22_pad_groupi_n_107, csa_tree_add_89_22_pad_groupi_n_108, csa_tree_add_89_22_pad_groupi_n_109, csa_tree_add_89_22_pad_groupi_n_110, csa_tree_add_89_22_pad_groupi_n_111;
  wire csa_tree_add_89_22_pad_groupi_n_112, csa_tree_add_89_22_pad_groupi_n_113, csa_tree_add_89_22_pad_groupi_n_114, csa_tree_add_89_22_pad_groupi_n_115, csa_tree_add_89_22_pad_groupi_n_116, csa_tree_add_89_22_pad_groupi_n_117, csa_tree_add_89_22_pad_groupi_n_118, csa_tree_add_89_22_pad_groupi_n_119;
  wire csa_tree_add_89_22_pad_groupi_n_120, csa_tree_add_89_22_pad_groupi_n_121, csa_tree_add_89_22_pad_groupi_n_122, csa_tree_add_89_22_pad_groupi_n_123, csa_tree_add_89_22_pad_groupi_n_124, csa_tree_add_89_22_pad_groupi_n_125, csa_tree_add_89_22_pad_groupi_n_126, csa_tree_add_89_22_pad_groupi_n_127;
  wire csa_tree_add_89_22_pad_groupi_n_128, csa_tree_add_89_22_pad_groupi_n_129, csa_tree_add_89_22_pad_groupi_n_130, csa_tree_add_89_22_pad_groupi_n_131, csa_tree_add_89_22_pad_groupi_n_132, csa_tree_add_89_22_pad_groupi_n_133, csa_tree_add_89_22_pad_groupi_n_134, csa_tree_add_89_22_pad_groupi_n_135;
  wire csa_tree_add_89_22_pad_groupi_n_136, csa_tree_add_89_22_pad_groupi_n_137, csa_tree_add_89_22_pad_groupi_n_138, csa_tree_add_89_22_pad_groupi_n_139, csa_tree_add_89_22_pad_groupi_n_140, csa_tree_add_89_22_pad_groupi_n_141, csa_tree_add_89_22_pad_groupi_n_142, csa_tree_add_89_22_pad_groupi_n_143;
  wire csa_tree_add_89_22_pad_groupi_n_144, csa_tree_add_89_22_pad_groupi_n_145, csa_tree_add_89_22_pad_groupi_n_146, csa_tree_add_89_22_pad_groupi_n_147, csa_tree_add_89_22_pad_groupi_n_148, csa_tree_add_89_22_pad_groupi_n_149, csa_tree_add_89_22_pad_groupi_n_150, csa_tree_add_89_22_pad_groupi_n_151;
  wire csa_tree_add_89_22_pad_groupi_n_152, csa_tree_add_89_22_pad_groupi_n_153, csa_tree_add_89_22_pad_groupi_n_154, csa_tree_add_89_22_pad_groupi_n_155, csa_tree_add_89_22_pad_groupi_n_156, csa_tree_add_89_22_pad_groupi_n_158, csa_tree_add_89_22_pad_groupi_n_159, csa_tree_add_89_22_pad_groupi_n_160;
  wire csa_tree_add_89_22_pad_groupi_n_161, csa_tree_add_89_22_pad_groupi_n_162, csa_tree_add_89_22_pad_groupi_n_163, csa_tree_add_89_22_pad_groupi_n_164, csa_tree_add_89_22_pad_groupi_n_165, csa_tree_add_89_22_pad_groupi_n_166, csa_tree_add_89_22_pad_groupi_n_167, csa_tree_add_89_22_pad_groupi_n_168;
  wire csa_tree_add_89_22_pad_groupi_n_169, csa_tree_add_89_22_pad_groupi_n_170, csa_tree_add_89_22_pad_groupi_n_171, csa_tree_add_89_22_pad_groupi_n_172, csa_tree_add_89_22_pad_groupi_n_173, csa_tree_add_89_22_pad_groupi_n_174, csa_tree_add_89_22_pad_groupi_n_175, csa_tree_add_89_22_pad_groupi_n_176;
  wire csa_tree_add_89_22_pad_groupi_n_177, csa_tree_add_89_22_pad_groupi_n_178, csa_tree_add_89_22_pad_groupi_n_179, csa_tree_add_89_22_pad_groupi_n_180, csa_tree_add_89_22_pad_groupi_n_181, csa_tree_add_89_22_pad_groupi_n_182, csa_tree_add_89_22_pad_groupi_n_183, csa_tree_add_89_22_pad_groupi_n_184;
  wire csa_tree_add_89_22_pad_groupi_n_185, csa_tree_add_89_22_pad_groupi_n_186, csa_tree_add_89_22_pad_groupi_n_187, csa_tree_add_89_22_pad_groupi_n_188, csa_tree_add_89_22_pad_groupi_n_189, csa_tree_add_89_22_pad_groupi_n_190, csa_tree_add_89_22_pad_groupi_n_191, csa_tree_add_89_22_pad_groupi_n_192;
  wire csa_tree_add_89_22_pad_groupi_n_193, csa_tree_add_89_22_pad_groupi_n_194, csa_tree_add_89_22_pad_groupi_n_195, csa_tree_add_89_22_pad_groupi_n_196, csa_tree_add_89_22_pad_groupi_n_197, csa_tree_add_89_22_pad_groupi_n_198, csa_tree_add_89_22_pad_groupi_n_200, csa_tree_add_89_22_pad_groupi_n_201;
  wire csa_tree_add_89_22_pad_groupi_n_202, csa_tree_add_89_22_pad_groupi_n_203, csa_tree_add_89_22_pad_groupi_n_204, csa_tree_add_89_22_pad_groupi_n_205, csa_tree_add_89_22_pad_groupi_n_206, csa_tree_add_89_22_pad_groupi_n_207, csa_tree_add_89_22_pad_groupi_n_208, csa_tree_add_89_22_pad_groupi_n_209;
  wire csa_tree_add_89_22_pad_groupi_n_210, csa_tree_add_89_22_pad_groupi_n_211, csa_tree_add_89_22_pad_groupi_n_212, csa_tree_add_89_22_pad_groupi_n_213, csa_tree_add_89_22_pad_groupi_n_214, csa_tree_add_89_22_pad_groupi_n_215, csa_tree_add_89_22_pad_groupi_n_216, csa_tree_add_89_22_pad_groupi_n_217;
  wire csa_tree_add_89_22_pad_groupi_n_218, csa_tree_add_89_22_pad_groupi_n_219, csa_tree_add_89_22_pad_groupi_n_220, csa_tree_add_89_22_pad_groupi_n_221, csa_tree_add_89_22_pad_groupi_n_222, csa_tree_add_89_22_pad_groupi_n_223, csa_tree_add_89_22_pad_groupi_n_224, csa_tree_add_89_22_pad_groupi_n_225;
  wire csa_tree_add_89_22_pad_groupi_n_226, csa_tree_add_89_22_pad_groupi_n_227, csa_tree_add_89_22_pad_groupi_n_228, csa_tree_add_89_22_pad_groupi_n_229, csa_tree_add_89_22_pad_groupi_n_230, csa_tree_add_89_22_pad_groupi_n_231, csa_tree_add_89_22_pad_groupi_n_232, csa_tree_add_89_22_pad_groupi_n_233;
  wire csa_tree_add_89_22_pad_groupi_n_234, csa_tree_add_89_22_pad_groupi_n_235, csa_tree_add_89_22_pad_groupi_n_236, csa_tree_add_89_22_pad_groupi_n_237, csa_tree_add_89_22_pad_groupi_n_238, csa_tree_add_89_22_pad_groupi_n_239, csa_tree_add_89_22_pad_groupi_n_240, csa_tree_add_89_22_pad_groupi_n_241;
  wire csa_tree_add_89_22_pad_groupi_n_242, csa_tree_add_89_22_pad_groupi_n_243, csa_tree_add_89_22_pad_groupi_n_244, csa_tree_add_89_22_pad_groupi_n_245, csa_tree_add_89_22_pad_groupi_n_246, csa_tree_add_89_22_pad_groupi_n_247, csa_tree_add_89_22_pad_groupi_n_248, csa_tree_add_89_22_pad_groupi_n_249;
  wire csa_tree_add_89_22_pad_groupi_n_250, csa_tree_add_89_22_pad_groupi_n_251, csa_tree_add_89_22_pad_groupi_n_252, csa_tree_add_89_22_pad_groupi_n_253, csa_tree_add_89_22_pad_groupi_n_254, csa_tree_add_89_22_pad_groupi_n_255, csa_tree_add_89_22_pad_groupi_n_256, csa_tree_add_89_22_pad_groupi_n_257;
  wire csa_tree_add_89_22_pad_groupi_n_258, csa_tree_add_89_22_pad_groupi_n_259, csa_tree_add_89_22_pad_groupi_n_260, csa_tree_add_89_22_pad_groupi_n_261, csa_tree_add_89_22_pad_groupi_n_262, csa_tree_add_89_22_pad_groupi_n_263, csa_tree_add_89_22_pad_groupi_n_264, csa_tree_add_89_22_pad_groupi_n_265;
  wire csa_tree_add_89_22_pad_groupi_n_266, csa_tree_add_89_22_pad_groupi_n_267, csa_tree_add_89_22_pad_groupi_n_268, csa_tree_add_89_22_pad_groupi_n_269, csa_tree_add_89_22_pad_groupi_n_270, csa_tree_add_89_22_pad_groupi_n_271, csa_tree_add_89_22_pad_groupi_n_272, csa_tree_add_89_22_pad_groupi_n_273;
  wire csa_tree_add_89_22_pad_groupi_n_274, csa_tree_add_89_22_pad_groupi_n_275, csa_tree_add_89_22_pad_groupi_n_276, csa_tree_add_89_22_pad_groupi_n_277, csa_tree_add_89_22_pad_groupi_n_278, csa_tree_add_89_22_pad_groupi_n_279, csa_tree_add_89_22_pad_groupi_n_280, csa_tree_add_89_22_pad_groupi_n_281;
  wire csa_tree_add_89_22_pad_groupi_n_282, csa_tree_add_89_22_pad_groupi_n_283, csa_tree_add_89_22_pad_groupi_n_284, csa_tree_add_89_22_pad_groupi_n_285, csa_tree_add_89_22_pad_groupi_n_286, csa_tree_add_89_22_pad_groupi_n_287, csa_tree_add_89_22_pad_groupi_n_288, csa_tree_add_89_22_pad_groupi_n_289;
  wire csa_tree_add_89_22_pad_groupi_n_290, csa_tree_add_89_22_pad_groupi_n_291, csa_tree_add_89_22_pad_groupi_n_292, csa_tree_add_89_22_pad_groupi_n_293, csa_tree_add_89_22_pad_groupi_n_294, csa_tree_add_89_22_pad_groupi_n_295, csa_tree_add_89_22_pad_groupi_n_296, csa_tree_add_89_22_pad_groupi_n_297;
  wire csa_tree_add_89_22_pad_groupi_n_298, csa_tree_add_89_22_pad_groupi_n_299, csa_tree_add_89_22_pad_groupi_n_300, csa_tree_add_89_22_pad_groupi_n_301, csa_tree_add_89_22_pad_groupi_n_302, csa_tree_add_89_22_pad_groupi_n_303, csa_tree_add_89_22_pad_groupi_n_304, csa_tree_add_89_22_pad_groupi_n_305;
  wire csa_tree_add_89_22_pad_groupi_n_306, csa_tree_add_89_22_pad_groupi_n_307, csa_tree_add_89_22_pad_groupi_n_308, csa_tree_add_89_22_pad_groupi_n_309, csa_tree_add_89_22_pad_groupi_n_310, csa_tree_add_89_22_pad_groupi_n_311, csa_tree_add_89_22_pad_groupi_n_312, csa_tree_add_89_22_pad_groupi_n_313;
  wire csa_tree_add_89_22_pad_groupi_n_314, csa_tree_add_89_22_pad_groupi_n_315, csa_tree_add_89_22_pad_groupi_n_316, csa_tree_add_89_22_pad_groupi_n_317, csa_tree_add_89_22_pad_groupi_n_318, csa_tree_add_89_22_pad_groupi_n_319, csa_tree_add_89_22_pad_groupi_n_320, csa_tree_add_89_22_pad_groupi_n_321;
  wire csa_tree_add_89_22_pad_groupi_n_322, csa_tree_add_89_22_pad_groupi_n_323, csa_tree_add_89_22_pad_groupi_n_324, csa_tree_add_89_22_pad_groupi_n_325, csa_tree_add_89_22_pad_groupi_n_326, csa_tree_add_89_22_pad_groupi_n_327, csa_tree_add_89_22_pad_groupi_n_328, csa_tree_add_89_22_pad_groupi_n_329;
  wire csa_tree_add_89_22_pad_groupi_n_330, csa_tree_add_89_22_pad_groupi_n_331, csa_tree_add_89_22_pad_groupi_n_332, csa_tree_add_89_22_pad_groupi_n_333, csa_tree_add_89_22_pad_groupi_n_334, csa_tree_add_89_22_pad_groupi_n_335, csa_tree_add_89_22_pad_groupi_n_336, csa_tree_add_89_22_pad_groupi_n_337;
  wire csa_tree_add_89_22_pad_groupi_n_338, csa_tree_add_89_22_pad_groupi_n_339, csa_tree_add_89_22_pad_groupi_n_340, csa_tree_add_89_22_pad_groupi_n_341, csa_tree_add_89_22_pad_groupi_n_342, csa_tree_add_89_22_pad_groupi_n_343, csa_tree_add_89_22_pad_groupi_n_344, csa_tree_add_89_22_pad_groupi_n_345;
  wire csa_tree_add_89_22_pad_groupi_n_346, csa_tree_add_89_22_pad_groupi_n_347, csa_tree_add_89_22_pad_groupi_n_348, csa_tree_add_89_22_pad_groupi_n_349, csa_tree_add_89_22_pad_groupi_n_350, csa_tree_add_89_22_pad_groupi_n_351, csa_tree_add_89_22_pad_groupi_n_352, csa_tree_add_89_22_pad_groupi_n_353;
  wire csa_tree_add_89_22_pad_groupi_n_354, csa_tree_add_89_22_pad_groupi_n_355, csa_tree_add_89_22_pad_groupi_n_356, csa_tree_add_89_22_pad_groupi_n_357, csa_tree_add_89_22_pad_groupi_n_358, csa_tree_add_89_22_pad_groupi_n_359, csa_tree_add_89_22_pad_groupi_n_361, csa_tree_add_89_22_pad_groupi_n_362;
  wire csa_tree_add_89_22_pad_groupi_n_363, csa_tree_add_89_22_pad_groupi_n_364, csa_tree_add_89_22_pad_groupi_n_365, csa_tree_add_89_22_pad_groupi_n_366, csa_tree_add_89_22_pad_groupi_n_367, csa_tree_add_89_22_pad_groupi_n_368, csa_tree_add_89_22_pad_groupi_n_369, csa_tree_add_89_22_pad_groupi_n_370;
  wire csa_tree_add_89_22_pad_groupi_n_371, csa_tree_add_89_22_pad_groupi_n_372, csa_tree_add_89_22_pad_groupi_n_373, csa_tree_add_89_22_pad_groupi_n_374, csa_tree_add_89_22_pad_groupi_n_375, csa_tree_add_89_22_pad_groupi_n_376, csa_tree_add_89_22_pad_groupi_n_377, csa_tree_add_89_22_pad_groupi_n_378;
  wire csa_tree_add_89_22_pad_groupi_n_379, csa_tree_add_89_22_pad_groupi_n_380, csa_tree_add_89_22_pad_groupi_n_381, csa_tree_add_89_22_pad_groupi_n_382, csa_tree_add_89_22_pad_groupi_n_383, csa_tree_add_89_22_pad_groupi_n_384, csa_tree_add_89_22_pad_groupi_n_385, csa_tree_add_89_22_pad_groupi_n_386;
  wire csa_tree_add_89_22_pad_groupi_n_387, csa_tree_add_89_22_pad_groupi_n_388, csa_tree_add_89_22_pad_groupi_n_389, csa_tree_add_89_22_pad_groupi_n_390, csa_tree_add_89_22_pad_groupi_n_391, csa_tree_add_89_22_pad_groupi_n_392, csa_tree_add_89_22_pad_groupi_n_393, csa_tree_add_89_22_pad_groupi_n_394;
  wire csa_tree_add_89_22_pad_groupi_n_395, csa_tree_add_89_22_pad_groupi_n_396, csa_tree_add_89_22_pad_groupi_n_397, csa_tree_add_89_22_pad_groupi_n_398, csa_tree_add_89_22_pad_groupi_n_399, csa_tree_add_89_22_pad_groupi_n_401, csa_tree_add_89_22_pad_groupi_n_402, csa_tree_add_89_22_pad_groupi_n_403;
  wire csa_tree_add_89_22_pad_groupi_n_404, csa_tree_add_89_22_pad_groupi_n_406, csa_tree_add_89_22_pad_groupi_n_409, csa_tree_add_89_22_pad_groupi_n_410, csa_tree_add_89_22_pad_groupi_n_411, csa_tree_add_89_22_pad_groupi_n_412, csa_tree_add_89_22_pad_groupi_n_413, csa_tree_add_89_22_pad_groupi_n_414;
  wire csa_tree_add_89_22_pad_groupi_n_415, csa_tree_add_89_22_pad_groupi_n_416, csa_tree_add_89_22_pad_groupi_n_417, csa_tree_add_89_22_pad_groupi_n_418, csa_tree_add_89_22_pad_groupi_n_419, csa_tree_add_89_22_pad_groupi_n_420, csa_tree_add_89_22_pad_groupi_n_421, csa_tree_add_89_22_pad_groupi_n_422;
  wire csa_tree_add_89_22_pad_groupi_n_423, csa_tree_add_89_22_pad_groupi_n_424, csa_tree_add_89_22_pad_groupi_n_425, csa_tree_add_89_22_pad_groupi_n_426, csa_tree_add_89_22_pad_groupi_n_427, csa_tree_add_89_22_pad_groupi_n_428, csa_tree_add_89_22_pad_groupi_n_429, csa_tree_add_89_22_pad_groupi_n_430;
  wire csa_tree_add_89_22_pad_groupi_n_431, csa_tree_add_89_22_pad_groupi_n_432, csa_tree_add_89_22_pad_groupi_n_433, csa_tree_add_89_22_pad_groupi_n_434, csa_tree_add_89_22_pad_groupi_n_435, csa_tree_add_89_22_pad_groupi_n_438, csa_tree_add_89_22_pad_groupi_n_439, csa_tree_add_89_22_pad_groupi_n_445;
  wire csa_tree_add_89_22_pad_groupi_n_455, csa_tree_add_89_22_pad_groupi_n_456, csa_tree_add_89_22_pad_groupi_n_457, csa_tree_add_89_22_pad_groupi_n_458, csa_tree_add_89_22_pad_groupi_n_459, csa_tree_add_89_22_pad_groupi_n_460, csa_tree_add_89_22_pad_groupi_n_461, csa_tree_add_89_22_pad_groupi_n_462;
  wire csa_tree_add_89_22_pad_groupi_n_463, csa_tree_add_89_22_pad_groupi_n_464, csa_tree_add_89_22_pad_groupi_n_465, csa_tree_add_89_22_pad_groupi_n_466, csa_tree_add_89_22_pad_groupi_n_467, csa_tree_add_89_22_pad_groupi_n_468, csa_tree_add_89_22_pad_groupi_n_469, csa_tree_add_89_22_pad_groupi_n_470;
  wire csa_tree_add_89_22_pad_groupi_n_471, csa_tree_add_89_22_pad_groupi_n_472, csa_tree_add_89_22_pad_groupi_n_473, csa_tree_add_89_22_pad_groupi_n_474, csa_tree_add_89_22_pad_groupi_n_475, csa_tree_add_89_22_pad_groupi_n_476, csa_tree_add_89_22_pad_groupi_n_477, csa_tree_add_89_22_pad_groupi_n_478;
  wire csa_tree_add_89_22_pad_groupi_n_479, csa_tree_add_89_22_pad_groupi_n_480, csa_tree_add_89_22_pad_groupi_n_481, csa_tree_add_89_22_pad_groupi_n_482, csa_tree_add_89_22_pad_groupi_n_483, csa_tree_add_89_22_pad_groupi_n_484, csa_tree_add_89_22_pad_groupi_n_485, csa_tree_add_89_22_pad_groupi_n_486;
  wire csa_tree_add_89_22_pad_groupi_n_487, csa_tree_add_89_22_pad_groupi_n_488, csa_tree_add_89_22_pad_groupi_n_489, csa_tree_add_89_22_pad_groupi_n_490, csa_tree_add_89_22_pad_groupi_n_491, csa_tree_add_89_22_pad_groupi_n_492, csa_tree_add_89_22_pad_groupi_n_493, csa_tree_add_89_22_pad_groupi_n_494;
  wire csa_tree_add_89_22_pad_groupi_n_495, csa_tree_add_89_22_pad_groupi_n_496, csa_tree_add_89_22_pad_groupi_n_497, csa_tree_add_89_22_pad_groupi_n_498, csa_tree_add_89_22_pad_groupi_n_499, csa_tree_add_89_22_pad_groupi_n_500, csa_tree_add_89_22_pad_groupi_n_501, csa_tree_add_89_22_pad_groupi_n_502;
  wire csa_tree_add_89_22_pad_groupi_n_503, csa_tree_add_89_22_pad_groupi_n_504, csa_tree_add_89_22_pad_groupi_n_505, csa_tree_add_89_22_pad_groupi_n_506, csa_tree_add_89_22_pad_groupi_n_507, csa_tree_add_89_22_pad_groupi_n_508, csa_tree_add_89_22_pad_groupi_n_509, csa_tree_add_89_22_pad_groupi_n_510;
  wire csa_tree_add_89_22_pad_groupi_n_511, csa_tree_add_89_22_pad_groupi_n_512, csa_tree_add_89_22_pad_groupi_n_513, csa_tree_add_89_22_pad_groupi_n_514, csa_tree_add_89_22_pad_groupi_n_515, csa_tree_add_89_22_pad_groupi_n_516, csa_tree_add_89_22_pad_groupi_n_517, csa_tree_add_89_22_pad_groupi_n_518;
  wire csa_tree_add_89_22_pad_groupi_n_519, csa_tree_add_89_22_pad_groupi_n_520, csa_tree_add_89_22_pad_groupi_n_521, csa_tree_add_89_22_pad_groupi_n_522, csa_tree_add_89_22_pad_groupi_n_523, csa_tree_add_89_22_pad_groupi_n_524, csa_tree_add_89_22_pad_groupi_n_525, csa_tree_add_89_22_pad_groupi_n_526;
  wire csa_tree_add_89_22_pad_groupi_n_527, csa_tree_add_89_22_pad_groupi_n_528, csa_tree_add_89_22_pad_groupi_n_529, csa_tree_add_89_22_pad_groupi_n_530, csa_tree_add_89_22_pad_groupi_n_531, csa_tree_add_89_22_pad_groupi_n_532, csa_tree_add_89_22_pad_groupi_n_533, csa_tree_add_89_22_pad_groupi_n_534;
  wire csa_tree_add_89_22_pad_groupi_n_535, csa_tree_add_89_22_pad_groupi_n_536, csa_tree_add_89_22_pad_groupi_n_537, csa_tree_add_89_22_pad_groupi_n_538, csa_tree_add_89_22_pad_groupi_n_539, csa_tree_add_89_22_pad_groupi_n_540, csa_tree_add_89_22_pad_groupi_n_541, csa_tree_add_89_22_pad_groupi_n_542;
  wire csa_tree_add_89_22_pad_groupi_n_543, csa_tree_add_89_22_pad_groupi_n_544, csa_tree_add_89_22_pad_groupi_n_545, csa_tree_add_89_22_pad_groupi_n_546, csa_tree_add_89_22_pad_groupi_n_547, csa_tree_add_89_22_pad_groupi_n_548, csa_tree_add_89_22_pad_groupi_n_549, csa_tree_add_89_22_pad_groupi_n_550;
  wire csa_tree_add_89_22_pad_groupi_n_551, csa_tree_add_89_22_pad_groupi_n_552, csa_tree_add_89_22_pad_groupi_n_553, csa_tree_add_89_22_pad_groupi_n_554, csa_tree_add_89_22_pad_groupi_n_555, csa_tree_add_89_22_pad_groupi_n_556, csa_tree_add_89_22_pad_groupi_n_557, csa_tree_add_89_22_pad_groupi_n_559;
  wire csa_tree_add_89_22_pad_groupi_n_561, csa_tree_add_89_22_pad_groupi_n_562, csa_tree_add_89_22_pad_groupi_n_563, csa_tree_add_89_22_pad_groupi_n_564, csa_tree_add_89_22_pad_groupi_n_565, csa_tree_add_89_22_pad_groupi_n_566, csa_tree_add_89_22_pad_groupi_n_567, csa_tree_add_89_22_pad_groupi_n_568;
  wire csa_tree_add_89_22_pad_groupi_n_569, csa_tree_add_89_22_pad_groupi_n_570, csa_tree_add_89_22_pad_groupi_n_572, csa_tree_add_89_22_pad_groupi_n_573, csa_tree_add_89_22_pad_groupi_n_574, csa_tree_add_89_22_pad_groupi_n_575, csa_tree_add_89_22_pad_groupi_n_576, csa_tree_add_89_22_pad_groupi_n_577;
  wire csa_tree_add_89_22_pad_groupi_n_578, csa_tree_add_89_22_pad_groupi_n_579, csa_tree_add_89_22_pad_groupi_n_580, csa_tree_add_89_22_pad_groupi_n_581, csa_tree_add_89_22_pad_groupi_n_582, csa_tree_add_89_22_pad_groupi_n_583, csa_tree_add_89_22_pad_groupi_n_584, csa_tree_add_89_22_pad_groupi_n_586;
  wire csa_tree_add_89_22_pad_groupi_n_587, csa_tree_add_89_22_pad_groupi_n_588, csa_tree_add_89_22_pad_groupi_n_589, csa_tree_add_89_22_pad_groupi_n_590, csa_tree_add_89_22_pad_groupi_n_591, csa_tree_add_89_22_pad_groupi_n_592, csa_tree_add_89_22_pad_groupi_n_593, csa_tree_add_89_22_pad_groupi_n_594;
  wire csa_tree_add_89_22_pad_groupi_n_595, csa_tree_add_89_22_pad_groupi_n_598, csa_tree_add_89_22_pad_groupi_n_599, csa_tree_add_89_22_pad_groupi_n_600, csa_tree_add_89_22_pad_groupi_n_601, csa_tree_add_89_22_pad_groupi_n_602, csa_tree_add_89_22_pad_groupi_n_603, csa_tree_add_89_22_pad_groupi_n_604;
  wire csa_tree_add_89_22_pad_groupi_n_605, csa_tree_add_89_22_pad_groupi_n_606, csa_tree_add_89_22_pad_groupi_n_607, csa_tree_add_89_22_pad_groupi_n_608, csa_tree_add_89_22_pad_groupi_n_609, csa_tree_add_89_22_pad_groupi_n_610, csa_tree_add_89_22_pad_groupi_n_611, csa_tree_add_89_22_pad_groupi_n_612;
  wire csa_tree_add_89_22_pad_groupi_n_613, csa_tree_add_89_22_pad_groupi_n_614, csa_tree_add_89_22_pad_groupi_n_615, csa_tree_add_89_22_pad_groupi_n_616, csa_tree_add_89_22_pad_groupi_n_617, csa_tree_add_89_22_pad_groupi_n_618, csa_tree_add_89_22_pad_groupi_n_619, csa_tree_add_89_22_pad_groupi_n_620;
  wire csa_tree_add_89_22_pad_groupi_n_621, csa_tree_add_89_22_pad_groupi_n_622, csa_tree_add_89_22_pad_groupi_n_623, csa_tree_add_89_22_pad_groupi_n_624, csa_tree_add_89_22_pad_groupi_n_625, csa_tree_add_89_22_pad_groupi_n_626, csa_tree_add_89_22_pad_groupi_n_627, csa_tree_add_89_22_pad_groupi_n_628;
  wire csa_tree_add_89_22_pad_groupi_n_629, csa_tree_add_89_22_pad_groupi_n_630, csa_tree_add_89_22_pad_groupi_n_631, csa_tree_add_89_22_pad_groupi_n_633, csa_tree_add_89_22_pad_groupi_n_634, csa_tree_add_89_22_pad_groupi_n_635, csa_tree_add_89_22_pad_groupi_n_637, csa_tree_add_89_22_pad_groupi_n_638;
  wire csa_tree_add_89_22_pad_groupi_n_639, csa_tree_add_89_22_pad_groupi_n_640, csa_tree_add_89_22_pad_groupi_n_641, csa_tree_add_89_22_pad_groupi_n_642, csa_tree_add_89_22_pad_groupi_n_643, csa_tree_add_89_22_pad_groupi_n_644, csa_tree_add_89_22_pad_groupi_n_645, csa_tree_add_89_22_pad_groupi_n_646;
  wire csa_tree_add_89_22_pad_groupi_n_647, csa_tree_add_89_22_pad_groupi_n_648, csa_tree_add_89_22_pad_groupi_n_649, csa_tree_add_89_22_pad_groupi_n_650, csa_tree_add_89_22_pad_groupi_n_651, csa_tree_add_89_22_pad_groupi_n_652, csa_tree_add_89_22_pad_groupi_n_653, csa_tree_add_89_22_pad_groupi_n_654;
  wire csa_tree_add_89_22_pad_groupi_n_655, csa_tree_add_89_22_pad_groupi_n_656, csa_tree_add_89_22_pad_groupi_n_657, csa_tree_add_89_22_pad_groupi_n_658, csa_tree_add_89_22_pad_groupi_n_659, csa_tree_add_89_22_pad_groupi_n_660, csa_tree_add_89_22_pad_groupi_n_661, csa_tree_add_89_22_pad_groupi_n_662;
  wire csa_tree_add_89_22_pad_groupi_n_663, csa_tree_add_89_22_pad_groupi_n_664, csa_tree_add_89_22_pad_groupi_n_665, csa_tree_add_89_22_pad_groupi_n_666, csa_tree_add_89_22_pad_groupi_n_667, csa_tree_add_89_22_pad_groupi_n_668, csa_tree_add_89_22_pad_groupi_n_669, csa_tree_add_89_22_pad_groupi_n_670;
  wire csa_tree_add_89_22_pad_groupi_n_671, csa_tree_add_89_22_pad_groupi_n_672, csa_tree_add_89_22_pad_groupi_n_673, csa_tree_add_89_22_pad_groupi_n_674, csa_tree_add_89_22_pad_groupi_n_675, csa_tree_add_89_22_pad_groupi_n_676, csa_tree_add_89_22_pad_groupi_n_677, csa_tree_add_89_22_pad_groupi_n_678;
  wire csa_tree_add_89_22_pad_groupi_n_679, csa_tree_add_89_22_pad_groupi_n_680, csa_tree_add_89_22_pad_groupi_n_681, csa_tree_add_89_22_pad_groupi_n_682, csa_tree_add_89_22_pad_groupi_n_683, csa_tree_add_89_22_pad_groupi_n_684, csa_tree_add_89_22_pad_groupi_n_685, csa_tree_add_89_22_pad_groupi_n_686;
  wire csa_tree_add_89_22_pad_groupi_n_688, csa_tree_add_89_22_pad_groupi_n_689, csa_tree_add_89_22_pad_groupi_n_690, csa_tree_add_89_22_pad_groupi_n_691, csa_tree_add_89_22_pad_groupi_n_692, csa_tree_add_89_22_pad_groupi_n_693, csa_tree_add_89_22_pad_groupi_n_694, csa_tree_add_89_22_pad_groupi_n_695;
  wire csa_tree_add_89_22_pad_groupi_n_696, csa_tree_add_89_22_pad_groupi_n_697, csa_tree_add_89_22_pad_groupi_n_698, csa_tree_add_89_22_pad_groupi_n_699, csa_tree_add_89_22_pad_groupi_n_700, csa_tree_add_89_22_pad_groupi_n_702, csa_tree_add_89_22_pad_groupi_n_703, csa_tree_add_89_22_pad_groupi_n_704;
  wire csa_tree_add_89_22_pad_groupi_n_705, csa_tree_add_89_22_pad_groupi_n_706, csa_tree_add_89_22_pad_groupi_n_707, csa_tree_add_89_22_pad_groupi_n_708, csa_tree_add_89_22_pad_groupi_n_709, csa_tree_add_89_22_pad_groupi_n_710, csa_tree_add_89_22_pad_groupi_n_711, csa_tree_add_89_22_pad_groupi_n_712;
  wire csa_tree_add_89_22_pad_groupi_n_713, csa_tree_add_89_22_pad_groupi_n_714, csa_tree_add_89_22_pad_groupi_n_715, csa_tree_add_89_22_pad_groupi_n_716, csa_tree_add_89_22_pad_groupi_n_717, csa_tree_add_89_22_pad_groupi_n_718, csa_tree_add_89_22_pad_groupi_n_719, csa_tree_add_89_22_pad_groupi_n_720;
  wire csa_tree_add_89_22_pad_groupi_n_721, csa_tree_add_89_22_pad_groupi_n_722, csa_tree_add_89_22_pad_groupi_n_723, csa_tree_add_89_22_pad_groupi_n_724, csa_tree_add_89_22_pad_groupi_n_725, csa_tree_add_89_22_pad_groupi_n_726, csa_tree_add_89_22_pad_groupi_n_727, csa_tree_add_89_22_pad_groupi_n_728;
  wire csa_tree_add_89_22_pad_groupi_n_729, csa_tree_add_89_22_pad_groupi_n_730, csa_tree_add_89_22_pad_groupi_n_731, csa_tree_add_89_22_pad_groupi_n_732, csa_tree_add_89_22_pad_groupi_n_733, csa_tree_add_89_22_pad_groupi_n_734, csa_tree_add_89_22_pad_groupi_n_735, csa_tree_add_89_22_pad_groupi_n_736;
  wire csa_tree_add_89_22_pad_groupi_n_737, csa_tree_add_89_22_pad_groupi_n_738, csa_tree_add_89_22_pad_groupi_n_739, csa_tree_add_89_22_pad_groupi_n_740, csa_tree_add_89_22_pad_groupi_n_741, csa_tree_add_89_22_pad_groupi_n_742, csa_tree_add_89_22_pad_groupi_n_743, csa_tree_add_89_22_pad_groupi_n_744;
  wire csa_tree_add_89_22_pad_groupi_n_745, csa_tree_add_89_22_pad_groupi_n_746, csa_tree_add_89_22_pad_groupi_n_747, csa_tree_add_89_22_pad_groupi_n_748, csa_tree_add_89_22_pad_groupi_n_749, csa_tree_add_89_22_pad_groupi_n_750, csa_tree_add_89_22_pad_groupi_n_751, csa_tree_add_89_22_pad_groupi_n_752;
  wire csa_tree_add_89_22_pad_groupi_n_753, csa_tree_add_89_22_pad_groupi_n_754, csa_tree_add_89_22_pad_groupi_n_755, csa_tree_add_89_22_pad_groupi_n_756, csa_tree_add_89_22_pad_groupi_n_757, csa_tree_add_89_22_pad_groupi_n_758, csa_tree_add_89_22_pad_groupi_n_759, csa_tree_add_89_22_pad_groupi_n_760;
  wire csa_tree_add_89_22_pad_groupi_n_761, csa_tree_add_89_22_pad_groupi_n_762, csa_tree_add_89_22_pad_groupi_n_763, csa_tree_add_89_22_pad_groupi_n_764, csa_tree_add_89_22_pad_groupi_n_765, csa_tree_add_89_22_pad_groupi_n_766, csa_tree_add_89_22_pad_groupi_n_767, csa_tree_add_89_22_pad_groupi_n_768;
  wire csa_tree_add_89_22_pad_groupi_n_769, csa_tree_add_89_22_pad_groupi_n_770, csa_tree_add_89_22_pad_groupi_n_771, csa_tree_add_89_22_pad_groupi_n_772, csa_tree_add_89_22_pad_groupi_n_773, csa_tree_add_89_22_pad_groupi_n_774, csa_tree_add_89_22_pad_groupi_n_775, csa_tree_add_89_22_pad_groupi_n_776;
  wire csa_tree_add_89_22_pad_groupi_n_777, csa_tree_add_89_22_pad_groupi_n_778, csa_tree_add_89_22_pad_groupi_n_779, csa_tree_add_89_22_pad_groupi_n_780, csa_tree_add_89_22_pad_groupi_n_781, csa_tree_add_89_22_pad_groupi_n_782, csa_tree_add_89_22_pad_groupi_n_783, csa_tree_add_89_22_pad_groupi_n_784;
  wire csa_tree_add_89_22_pad_groupi_n_785, csa_tree_add_89_22_pad_groupi_n_786, csa_tree_add_89_22_pad_groupi_n_787, csa_tree_add_89_22_pad_groupi_n_788, csa_tree_add_89_22_pad_groupi_n_789, csa_tree_add_89_22_pad_groupi_n_790, csa_tree_add_89_22_pad_groupi_n_791, csa_tree_add_89_22_pad_groupi_n_792;
  wire csa_tree_add_89_22_pad_groupi_n_793, csa_tree_add_89_22_pad_groupi_n_794, csa_tree_add_89_22_pad_groupi_n_795, csa_tree_add_89_22_pad_groupi_n_796, csa_tree_add_89_22_pad_groupi_n_797, csa_tree_add_89_22_pad_groupi_n_798, csa_tree_add_89_22_pad_groupi_n_799, csa_tree_add_89_22_pad_groupi_n_800;
  wire csa_tree_add_89_22_pad_groupi_n_801, csa_tree_add_89_22_pad_groupi_n_802, csa_tree_add_89_22_pad_groupi_n_803, csa_tree_add_89_22_pad_groupi_n_804, csa_tree_add_89_22_pad_groupi_n_805, csa_tree_add_89_22_pad_groupi_n_806, csa_tree_add_89_22_pad_groupi_n_807, csa_tree_add_89_22_pad_groupi_n_808;
  wire csa_tree_add_89_22_pad_groupi_n_809, csa_tree_add_89_22_pad_groupi_n_810, csa_tree_add_89_22_pad_groupi_n_811, csa_tree_add_89_22_pad_groupi_n_812, csa_tree_add_89_22_pad_groupi_n_813, csa_tree_add_89_22_pad_groupi_n_814, csa_tree_add_89_22_pad_groupi_n_815, csa_tree_add_89_22_pad_groupi_n_816;
  wire csa_tree_add_89_22_pad_groupi_n_817, csa_tree_add_89_22_pad_groupi_n_818, csa_tree_add_89_22_pad_groupi_n_819, csa_tree_add_89_22_pad_groupi_n_820, csa_tree_add_89_22_pad_groupi_n_821, csa_tree_add_89_22_pad_groupi_n_822, csa_tree_add_89_22_pad_groupi_n_823, csa_tree_add_89_22_pad_groupi_n_824;
  wire csa_tree_add_89_22_pad_groupi_n_825, csa_tree_add_89_22_pad_groupi_n_826, csa_tree_add_89_22_pad_groupi_n_827, csa_tree_add_89_22_pad_groupi_n_828, csa_tree_add_89_22_pad_groupi_n_829, csa_tree_add_89_22_pad_groupi_n_830, csa_tree_add_89_22_pad_groupi_n_831, csa_tree_add_89_22_pad_groupi_n_832;
  wire csa_tree_add_89_22_pad_groupi_n_833, csa_tree_add_89_22_pad_groupi_n_834, csa_tree_add_89_22_pad_groupi_n_835, csa_tree_add_89_22_pad_groupi_n_836, csa_tree_add_89_22_pad_groupi_n_837, csa_tree_add_89_22_pad_groupi_n_838, csa_tree_add_89_22_pad_groupi_n_839, csa_tree_add_89_22_pad_groupi_n_840;
  wire csa_tree_add_89_22_pad_groupi_n_841, csa_tree_add_89_22_pad_groupi_n_842, csa_tree_add_89_22_pad_groupi_n_843, csa_tree_add_89_22_pad_groupi_n_844, csa_tree_add_89_22_pad_groupi_n_845, csa_tree_add_89_22_pad_groupi_n_846, csa_tree_add_89_22_pad_groupi_n_847, csa_tree_add_89_22_pad_groupi_n_848;
  wire csa_tree_add_89_22_pad_groupi_n_849, csa_tree_add_89_22_pad_groupi_n_851, csa_tree_add_89_22_pad_groupi_n_852, csa_tree_add_89_22_pad_groupi_n_853, csa_tree_add_89_22_pad_groupi_n_854, csa_tree_add_89_22_pad_groupi_n_855, csa_tree_add_89_22_pad_groupi_n_856, csa_tree_add_89_22_pad_groupi_n_857;
  wire csa_tree_add_89_22_pad_groupi_n_858, csa_tree_add_89_22_pad_groupi_n_859, csa_tree_add_89_22_pad_groupi_n_860, csa_tree_add_89_22_pad_groupi_n_861, csa_tree_add_89_22_pad_groupi_n_862, csa_tree_add_89_22_pad_groupi_n_863, csa_tree_add_89_22_pad_groupi_n_864, csa_tree_add_89_22_pad_groupi_n_865;
  wire csa_tree_add_89_22_pad_groupi_n_866, csa_tree_add_89_22_pad_groupi_n_867, csa_tree_add_89_22_pad_groupi_n_868, csa_tree_add_89_22_pad_groupi_n_869, csa_tree_add_89_22_pad_groupi_n_870, csa_tree_add_89_22_pad_groupi_n_871, csa_tree_add_89_22_pad_groupi_n_872, csa_tree_add_89_22_pad_groupi_n_873;
  wire csa_tree_add_89_22_pad_groupi_n_874, csa_tree_add_89_22_pad_groupi_n_875, csa_tree_add_89_22_pad_groupi_n_876, csa_tree_add_89_22_pad_groupi_n_877, csa_tree_add_89_22_pad_groupi_n_878, csa_tree_add_89_22_pad_groupi_n_879, csa_tree_add_89_22_pad_groupi_n_880, csa_tree_add_89_22_pad_groupi_n_881;
  wire csa_tree_add_89_22_pad_groupi_n_882, csa_tree_add_89_22_pad_groupi_n_883, csa_tree_add_89_22_pad_groupi_n_884, csa_tree_add_89_22_pad_groupi_n_885, csa_tree_add_89_22_pad_groupi_n_886, csa_tree_add_89_22_pad_groupi_n_887, csa_tree_add_89_22_pad_groupi_n_888, csa_tree_add_89_22_pad_groupi_n_889;
  wire csa_tree_add_89_22_pad_groupi_n_890, csa_tree_add_89_22_pad_groupi_n_891, csa_tree_add_89_22_pad_groupi_n_892, csa_tree_add_89_22_pad_groupi_n_893, csa_tree_add_89_22_pad_groupi_n_894, csa_tree_add_89_22_pad_groupi_n_895, csa_tree_add_89_22_pad_groupi_n_896, csa_tree_add_89_22_pad_groupi_n_897;
  wire csa_tree_add_89_22_pad_groupi_n_898, csa_tree_add_89_22_pad_groupi_n_899, csa_tree_add_89_22_pad_groupi_n_900, csa_tree_add_89_22_pad_groupi_n_901, csa_tree_add_89_22_pad_groupi_n_902, csa_tree_add_89_22_pad_groupi_n_903, csa_tree_add_89_22_pad_groupi_n_904, csa_tree_add_89_22_pad_groupi_n_905;
  wire csa_tree_add_89_22_pad_groupi_n_906, csa_tree_add_89_22_pad_groupi_n_907, csa_tree_add_89_22_pad_groupi_n_908, csa_tree_add_89_22_pad_groupi_n_909, csa_tree_add_89_22_pad_groupi_n_910, csa_tree_add_89_22_pad_groupi_n_911, csa_tree_add_89_22_pad_groupi_n_912, csa_tree_add_89_22_pad_groupi_n_913;
  wire csa_tree_add_89_22_pad_groupi_n_914, csa_tree_add_89_22_pad_groupi_n_915, csa_tree_add_89_22_pad_groupi_n_916, csa_tree_add_89_22_pad_groupi_n_917, csa_tree_add_89_22_pad_groupi_n_918, csa_tree_add_89_22_pad_groupi_n_919, csa_tree_add_89_22_pad_groupi_n_920, csa_tree_add_89_22_pad_groupi_n_921;
  wire csa_tree_add_89_22_pad_groupi_n_922, csa_tree_add_89_22_pad_groupi_n_923, csa_tree_add_89_22_pad_groupi_n_924, csa_tree_add_89_22_pad_groupi_n_925, csa_tree_add_89_22_pad_groupi_n_926, csa_tree_add_89_22_pad_groupi_n_927, csa_tree_add_89_22_pad_groupi_n_928, csa_tree_add_89_22_pad_groupi_n_929;
  wire csa_tree_add_89_22_pad_groupi_n_930, csa_tree_add_89_22_pad_groupi_n_931, csa_tree_add_89_22_pad_groupi_n_932, csa_tree_add_89_22_pad_groupi_n_933, csa_tree_add_89_22_pad_groupi_n_934, csa_tree_add_89_22_pad_groupi_n_935, csa_tree_add_89_22_pad_groupi_n_936, csa_tree_add_89_22_pad_groupi_n_937;
  wire csa_tree_add_89_22_pad_groupi_n_938, csa_tree_add_89_22_pad_groupi_n_939, csa_tree_add_89_22_pad_groupi_n_940, csa_tree_add_89_22_pad_groupi_n_941, csa_tree_add_89_22_pad_groupi_n_942, csa_tree_add_89_22_pad_groupi_n_943, csa_tree_add_89_22_pad_groupi_n_944, csa_tree_add_89_22_pad_groupi_n_945;
  wire csa_tree_add_89_22_pad_groupi_n_946, csa_tree_add_89_22_pad_groupi_n_947, csa_tree_add_89_22_pad_groupi_n_948, csa_tree_add_89_22_pad_groupi_n_949, csa_tree_add_89_22_pad_groupi_n_950, csa_tree_add_89_22_pad_groupi_n_951, csa_tree_add_89_22_pad_groupi_n_952, csa_tree_add_89_22_pad_groupi_n_953;
  wire csa_tree_add_89_22_pad_groupi_n_954, csa_tree_add_89_22_pad_groupi_n_955, csa_tree_add_89_22_pad_groupi_n_956, csa_tree_add_89_22_pad_groupi_n_957, csa_tree_add_89_22_pad_groupi_n_958, csa_tree_add_89_22_pad_groupi_n_959, csa_tree_add_89_22_pad_groupi_n_960, csa_tree_add_89_22_pad_groupi_n_961;
  wire csa_tree_add_89_22_pad_groupi_n_962, csa_tree_add_89_22_pad_groupi_n_963, csa_tree_add_89_22_pad_groupi_n_964, csa_tree_add_89_22_pad_groupi_n_965, csa_tree_add_89_22_pad_groupi_n_966, csa_tree_add_89_22_pad_groupi_n_967, csa_tree_add_89_22_pad_groupi_n_968, csa_tree_add_89_22_pad_groupi_n_969;
  wire csa_tree_add_89_22_pad_groupi_n_970, csa_tree_add_89_22_pad_groupi_n_971, csa_tree_add_89_22_pad_groupi_n_972, csa_tree_add_89_22_pad_groupi_n_973, csa_tree_add_89_22_pad_groupi_n_974, csa_tree_add_89_22_pad_groupi_n_975, csa_tree_add_89_22_pad_groupi_n_976, csa_tree_add_89_22_pad_groupi_n_977;
  wire csa_tree_add_89_22_pad_groupi_n_978, csa_tree_add_89_22_pad_groupi_n_979, csa_tree_add_89_22_pad_groupi_n_980, csa_tree_add_89_22_pad_groupi_n_981, csa_tree_add_89_22_pad_groupi_n_982, csa_tree_add_89_22_pad_groupi_n_983, csa_tree_add_89_22_pad_groupi_n_984, csa_tree_add_89_22_pad_groupi_n_985;
  wire csa_tree_add_89_22_pad_groupi_n_986, csa_tree_add_89_22_pad_groupi_n_987, csa_tree_add_89_22_pad_groupi_n_988, csa_tree_add_89_22_pad_groupi_n_989, csa_tree_add_89_22_pad_groupi_n_990, csa_tree_add_89_22_pad_groupi_n_991, csa_tree_add_89_22_pad_groupi_n_992, csa_tree_add_89_22_pad_groupi_n_993;
  wire csa_tree_add_89_22_pad_groupi_n_994, csa_tree_add_89_22_pad_groupi_n_995, csa_tree_add_89_22_pad_groupi_n_996, csa_tree_add_89_22_pad_groupi_n_997, csa_tree_add_89_22_pad_groupi_n_998, csa_tree_add_89_22_pad_groupi_n_999, csa_tree_add_89_22_pad_groupi_n_1000, csa_tree_add_89_22_pad_groupi_n_1001;
  wire csa_tree_add_89_22_pad_groupi_n_1002, csa_tree_add_89_22_pad_groupi_n_1003, csa_tree_add_89_22_pad_groupi_n_1004, csa_tree_add_89_22_pad_groupi_n_1005, csa_tree_add_89_22_pad_groupi_n_1006, csa_tree_add_89_22_pad_groupi_n_1007, csa_tree_add_89_22_pad_groupi_n_1008, csa_tree_add_89_22_pad_groupi_n_1009;
  wire csa_tree_add_89_22_pad_groupi_n_1010, csa_tree_add_89_22_pad_groupi_n_1011, csa_tree_add_89_22_pad_groupi_n_1012, csa_tree_add_89_22_pad_groupi_n_1013, csa_tree_add_89_22_pad_groupi_n_1014, csa_tree_add_89_22_pad_groupi_n_1015, csa_tree_add_89_22_pad_groupi_n_1016, csa_tree_add_89_22_pad_groupi_n_1017;
  wire csa_tree_add_89_22_pad_groupi_n_1018, csa_tree_add_89_22_pad_groupi_n_1019, csa_tree_add_89_22_pad_groupi_n_1020, csa_tree_add_89_22_pad_groupi_n_1021, csa_tree_add_89_22_pad_groupi_n_1022, csa_tree_add_89_22_pad_groupi_n_1023, csa_tree_add_89_22_pad_groupi_n_1024, csa_tree_add_89_22_pad_groupi_n_1025;
  wire csa_tree_add_89_22_pad_groupi_n_1026, csa_tree_add_89_22_pad_groupi_n_1027, csa_tree_add_89_22_pad_groupi_n_1028, csa_tree_add_89_22_pad_groupi_n_1029, csa_tree_add_89_22_pad_groupi_n_1030, csa_tree_add_89_22_pad_groupi_n_1031, csa_tree_add_89_22_pad_groupi_n_1032, csa_tree_add_89_22_pad_groupi_n_1033;
  wire csa_tree_add_89_22_pad_groupi_n_1034, csa_tree_add_89_22_pad_groupi_n_1035, csa_tree_add_89_22_pad_groupi_n_1036, csa_tree_add_89_22_pad_groupi_n_1037, csa_tree_add_89_22_pad_groupi_n_1038, csa_tree_add_89_22_pad_groupi_n_1039, csa_tree_add_89_22_pad_groupi_n_1040, csa_tree_add_89_22_pad_groupi_n_1041;
  wire csa_tree_add_89_22_pad_groupi_n_1042, csa_tree_add_89_22_pad_groupi_n_1043, csa_tree_add_89_22_pad_groupi_n_1044, csa_tree_add_89_22_pad_groupi_n_1045, csa_tree_add_89_22_pad_groupi_n_1046, csa_tree_add_89_22_pad_groupi_n_1047, csa_tree_add_89_22_pad_groupi_n_1048, csa_tree_add_89_22_pad_groupi_n_1049;
  wire csa_tree_add_89_22_pad_groupi_n_1050, csa_tree_add_89_22_pad_groupi_n_1051, csa_tree_add_89_22_pad_groupi_n_1052, csa_tree_add_89_22_pad_groupi_n_1053, csa_tree_add_89_22_pad_groupi_n_1054, csa_tree_add_89_22_pad_groupi_n_1055, csa_tree_add_89_22_pad_groupi_n_1056, csa_tree_add_89_22_pad_groupi_n_1057;
  wire csa_tree_add_89_22_pad_groupi_n_1058, csa_tree_add_89_22_pad_groupi_n_1059, csa_tree_add_89_22_pad_groupi_n_1060, csa_tree_add_89_22_pad_groupi_n_1061, csa_tree_add_89_22_pad_groupi_n_1062, csa_tree_add_89_22_pad_groupi_n_1063, csa_tree_add_89_22_pad_groupi_n_1064, csa_tree_add_89_22_pad_groupi_n_1065;
  wire csa_tree_add_89_22_pad_groupi_n_1066, csa_tree_add_89_22_pad_groupi_n_1067, csa_tree_add_89_22_pad_groupi_n_1068, csa_tree_add_89_22_pad_groupi_n_1069, csa_tree_add_89_22_pad_groupi_n_1070, csa_tree_add_89_22_pad_groupi_n_1071, csa_tree_add_89_22_pad_groupi_n_1072, csa_tree_add_89_22_pad_groupi_n_1073;
  wire csa_tree_add_89_22_pad_groupi_n_1074, csa_tree_add_89_22_pad_groupi_n_1075, csa_tree_add_89_22_pad_groupi_n_1076, csa_tree_add_89_22_pad_groupi_n_1077, csa_tree_add_89_22_pad_groupi_n_1078, csa_tree_add_89_22_pad_groupi_n_1079, csa_tree_add_89_22_pad_groupi_n_1080, csa_tree_add_89_22_pad_groupi_n_1081;
  wire csa_tree_add_89_22_pad_groupi_n_1082, csa_tree_add_89_22_pad_groupi_n_1083, csa_tree_add_89_22_pad_groupi_n_1084, csa_tree_add_89_22_pad_groupi_n_1085, csa_tree_add_89_22_pad_groupi_n_1086, csa_tree_add_89_22_pad_groupi_n_1087, csa_tree_add_89_22_pad_groupi_n_1088, csa_tree_add_89_22_pad_groupi_n_1089;
  wire csa_tree_add_89_22_pad_groupi_n_1090, csa_tree_add_89_22_pad_groupi_n_1091, csa_tree_add_89_22_pad_groupi_n_1092, csa_tree_add_89_22_pad_groupi_n_1093, csa_tree_add_89_22_pad_groupi_n_1094, csa_tree_add_89_22_pad_groupi_n_1095, csa_tree_add_89_22_pad_groupi_n_1096, csa_tree_add_89_22_pad_groupi_n_1097;
  wire csa_tree_add_89_22_pad_groupi_n_1098, csa_tree_add_89_22_pad_groupi_n_1099, csa_tree_add_89_22_pad_groupi_n_1100, csa_tree_add_89_22_pad_groupi_n_1101, csa_tree_add_89_22_pad_groupi_n_1102, csa_tree_add_89_22_pad_groupi_n_1103, csa_tree_add_89_22_pad_groupi_n_1104, csa_tree_add_89_22_pad_groupi_n_1105;
  wire csa_tree_add_89_22_pad_groupi_n_1106, csa_tree_add_89_22_pad_groupi_n_1107, csa_tree_add_89_22_pad_groupi_n_1108, csa_tree_add_89_22_pad_groupi_n_1109, csa_tree_add_89_22_pad_groupi_n_1110, csa_tree_add_89_22_pad_groupi_n_1111, csa_tree_add_89_22_pad_groupi_n_1112, csa_tree_add_89_22_pad_groupi_n_1113;
  wire csa_tree_add_89_22_pad_groupi_n_1114, csa_tree_add_89_22_pad_groupi_n_1115, csa_tree_add_89_22_pad_groupi_n_1116, csa_tree_add_89_22_pad_groupi_n_1117, csa_tree_add_89_22_pad_groupi_n_1118, csa_tree_add_89_22_pad_groupi_n_1119, csa_tree_add_89_22_pad_groupi_n_1120, csa_tree_add_89_22_pad_groupi_n_1121;
  wire csa_tree_add_89_22_pad_groupi_n_1122, csa_tree_add_89_22_pad_groupi_n_1123, csa_tree_add_89_22_pad_groupi_n_1124, csa_tree_add_89_22_pad_groupi_n_1125, csa_tree_add_89_22_pad_groupi_n_1126, csa_tree_add_89_22_pad_groupi_n_1127, csa_tree_add_89_22_pad_groupi_n_1128, csa_tree_add_89_22_pad_groupi_n_1129;
  wire csa_tree_add_89_22_pad_groupi_n_1130, csa_tree_add_89_22_pad_groupi_n_1131, csa_tree_add_89_22_pad_groupi_n_1132, csa_tree_add_89_22_pad_groupi_n_1133, csa_tree_add_89_22_pad_groupi_n_1134, csa_tree_add_89_22_pad_groupi_n_1135, csa_tree_add_89_22_pad_groupi_n_1136, csa_tree_add_89_22_pad_groupi_n_1137;
  wire csa_tree_add_89_22_pad_groupi_n_1138, csa_tree_add_89_22_pad_groupi_n_1139, csa_tree_add_89_22_pad_groupi_n_1140, csa_tree_add_89_22_pad_groupi_n_1141, csa_tree_add_89_22_pad_groupi_n_1142, csa_tree_add_89_22_pad_groupi_n_1143, csa_tree_add_89_22_pad_groupi_n_1144, csa_tree_add_89_22_pad_groupi_n_1145;
  wire csa_tree_add_89_22_pad_groupi_n_1146, csa_tree_add_89_22_pad_groupi_n_1147, csa_tree_add_89_22_pad_groupi_n_1148, csa_tree_add_89_22_pad_groupi_n_1149, csa_tree_add_89_22_pad_groupi_n_1150, csa_tree_add_89_22_pad_groupi_n_1151, csa_tree_add_89_22_pad_groupi_n_1152, csa_tree_add_89_22_pad_groupi_n_1153;
  wire csa_tree_add_89_22_pad_groupi_n_1154, csa_tree_add_89_22_pad_groupi_n_1155, csa_tree_add_89_22_pad_groupi_n_1156, csa_tree_add_89_22_pad_groupi_n_1157, csa_tree_add_89_22_pad_groupi_n_1158, csa_tree_add_89_22_pad_groupi_n_1159, csa_tree_add_89_22_pad_groupi_n_1160, csa_tree_add_89_22_pad_groupi_n_1161;
  wire csa_tree_add_89_22_pad_groupi_n_1162, csa_tree_add_89_22_pad_groupi_n_1163, csa_tree_add_89_22_pad_groupi_n_1164, csa_tree_add_89_22_pad_groupi_n_1165, csa_tree_add_89_22_pad_groupi_n_1166, csa_tree_add_89_22_pad_groupi_n_1167, csa_tree_add_89_22_pad_groupi_n_1168, csa_tree_add_89_22_pad_groupi_n_1169;
  wire csa_tree_add_89_22_pad_groupi_n_1170, csa_tree_add_89_22_pad_groupi_n_1171, csa_tree_add_89_22_pad_groupi_n_1172, csa_tree_add_89_22_pad_groupi_n_1173, csa_tree_add_89_22_pad_groupi_n_1174, csa_tree_add_89_22_pad_groupi_n_1175, csa_tree_add_89_22_pad_groupi_n_1176, csa_tree_add_89_22_pad_groupi_n_1177;
  wire csa_tree_add_89_22_pad_groupi_n_1178, csa_tree_add_89_22_pad_groupi_n_1179, csa_tree_add_89_22_pad_groupi_n_1180, csa_tree_add_89_22_pad_groupi_n_1181, csa_tree_add_89_22_pad_groupi_n_1182, csa_tree_add_89_22_pad_groupi_n_1183, csa_tree_add_89_22_pad_groupi_n_1184, csa_tree_add_89_22_pad_groupi_n_1185;
  wire csa_tree_add_89_22_pad_groupi_n_1186, csa_tree_add_89_22_pad_groupi_n_1187, csa_tree_add_89_22_pad_groupi_n_1188, csa_tree_add_89_22_pad_groupi_n_1189, csa_tree_add_89_22_pad_groupi_n_1190, csa_tree_add_89_22_pad_groupi_n_1191, csa_tree_add_89_22_pad_groupi_n_1192, csa_tree_add_89_22_pad_groupi_n_1193;
  wire csa_tree_add_89_22_pad_groupi_n_1194, csa_tree_add_89_22_pad_groupi_n_1195, csa_tree_add_89_22_pad_groupi_n_1196, csa_tree_add_89_22_pad_groupi_n_1197, csa_tree_add_89_22_pad_groupi_n_1198, csa_tree_add_89_22_pad_groupi_n_1199, csa_tree_add_89_22_pad_groupi_n_1200, csa_tree_add_89_22_pad_groupi_n_1201;
  wire csa_tree_add_89_22_pad_groupi_n_1202, csa_tree_add_89_22_pad_groupi_n_1203, csa_tree_add_89_22_pad_groupi_n_1204, csa_tree_add_89_22_pad_groupi_n_1205, csa_tree_add_89_22_pad_groupi_n_1206, csa_tree_add_89_22_pad_groupi_n_1207, csa_tree_add_89_22_pad_groupi_n_1208, csa_tree_add_89_22_pad_groupi_n_1209;
  wire csa_tree_add_89_22_pad_groupi_n_1210, csa_tree_add_89_22_pad_groupi_n_1211, csa_tree_add_89_22_pad_groupi_n_1212, csa_tree_add_89_22_pad_groupi_n_1213, csa_tree_add_89_22_pad_groupi_n_1214, csa_tree_add_89_22_pad_groupi_n_1215, csa_tree_add_89_22_pad_groupi_n_1216, csa_tree_add_89_22_pad_groupi_n_1217;
  wire csa_tree_add_89_22_pad_groupi_n_1218, csa_tree_add_89_22_pad_groupi_n_1219, csa_tree_add_89_22_pad_groupi_n_1220, csa_tree_add_89_22_pad_groupi_n_1221, csa_tree_add_89_22_pad_groupi_n_1222, csa_tree_add_89_22_pad_groupi_n_1223, csa_tree_add_89_22_pad_groupi_n_1224, csa_tree_add_89_22_pad_groupi_n_1225;
  wire csa_tree_add_89_22_pad_groupi_n_1226, csa_tree_add_89_22_pad_groupi_n_1227, csa_tree_add_89_22_pad_groupi_n_1228, csa_tree_add_89_22_pad_groupi_n_1229, csa_tree_add_89_22_pad_groupi_n_1230, csa_tree_add_89_22_pad_groupi_n_1231, csa_tree_add_89_22_pad_groupi_n_1232, csa_tree_add_89_22_pad_groupi_n_1233;
  wire csa_tree_add_89_22_pad_groupi_n_1234, csa_tree_add_89_22_pad_groupi_n_1235, csa_tree_add_89_22_pad_groupi_n_1236, csa_tree_add_89_22_pad_groupi_n_1237, csa_tree_add_89_22_pad_groupi_n_1238, csa_tree_add_89_22_pad_groupi_n_1239, csa_tree_add_89_22_pad_groupi_n_1240, csa_tree_add_89_22_pad_groupi_n_1241;
  wire csa_tree_add_89_22_pad_groupi_n_1242, csa_tree_add_89_22_pad_groupi_n_1243, csa_tree_add_89_22_pad_groupi_n_1244, csa_tree_add_89_22_pad_groupi_n_1245, csa_tree_add_89_22_pad_groupi_n_1246, csa_tree_add_89_22_pad_groupi_n_1247, csa_tree_add_89_22_pad_groupi_n_1248, csa_tree_add_89_22_pad_groupi_n_1249;
  wire csa_tree_add_89_22_pad_groupi_n_1250, csa_tree_add_89_22_pad_groupi_n_1251, csa_tree_add_89_22_pad_groupi_n_1252, csa_tree_add_89_22_pad_groupi_n_1253, csa_tree_add_89_22_pad_groupi_n_1254, csa_tree_add_89_22_pad_groupi_n_1255, csa_tree_add_89_22_pad_groupi_n_1256, csa_tree_add_89_22_pad_groupi_n_1257;
  wire csa_tree_add_89_22_pad_groupi_n_1258, csa_tree_add_89_22_pad_groupi_n_1259, csa_tree_add_89_22_pad_groupi_n_1260, csa_tree_add_89_22_pad_groupi_n_1261, csa_tree_add_89_22_pad_groupi_n_1262, csa_tree_add_89_22_pad_groupi_n_1263, csa_tree_add_89_22_pad_groupi_n_1264, csa_tree_add_89_22_pad_groupi_n_1265;
  wire csa_tree_add_89_22_pad_groupi_n_1266, csa_tree_add_89_22_pad_groupi_n_1267, csa_tree_add_89_22_pad_groupi_n_1268, csa_tree_add_89_22_pad_groupi_n_1269, csa_tree_add_89_22_pad_groupi_n_1270, csa_tree_add_89_22_pad_groupi_n_1271, csa_tree_add_89_22_pad_groupi_n_1272, csa_tree_add_89_22_pad_groupi_n_1273;
  wire csa_tree_add_89_22_pad_groupi_n_1274, csa_tree_add_89_22_pad_groupi_n_1275, csa_tree_add_89_22_pad_groupi_n_1276, csa_tree_add_89_22_pad_groupi_n_1277, csa_tree_add_89_22_pad_groupi_n_1278, csa_tree_add_89_22_pad_groupi_n_1279, csa_tree_add_89_22_pad_groupi_n_1280, csa_tree_add_89_22_pad_groupi_n_1281;
  wire csa_tree_add_89_22_pad_groupi_n_1282, csa_tree_add_89_22_pad_groupi_n_1283, csa_tree_add_89_22_pad_groupi_n_1284, csa_tree_add_89_22_pad_groupi_n_1285, csa_tree_add_89_22_pad_groupi_n_1286, csa_tree_add_89_22_pad_groupi_n_1287, csa_tree_add_89_22_pad_groupi_n_1288, csa_tree_add_89_22_pad_groupi_n_1289;
  wire csa_tree_add_89_22_pad_groupi_n_1290, csa_tree_add_89_22_pad_groupi_n_1291, csa_tree_add_89_22_pad_groupi_n_1292, csa_tree_add_89_22_pad_groupi_n_1293, csa_tree_add_89_22_pad_groupi_n_1294, csa_tree_add_89_22_pad_groupi_n_1295, csa_tree_add_89_22_pad_groupi_n_1296, csa_tree_add_89_22_pad_groupi_n_1297;
  wire csa_tree_add_89_22_pad_groupi_n_1298, csa_tree_add_89_22_pad_groupi_n_1299, csa_tree_add_89_22_pad_groupi_n_1300, csa_tree_add_89_22_pad_groupi_n_1301, csa_tree_add_89_22_pad_groupi_n_1302, csa_tree_add_89_22_pad_groupi_n_1303, csa_tree_add_89_22_pad_groupi_n_1304, csa_tree_add_89_22_pad_groupi_n_1305;
  wire csa_tree_add_89_22_pad_groupi_n_1306, csa_tree_add_89_22_pad_groupi_n_1307, csa_tree_add_89_22_pad_groupi_n_1308, csa_tree_add_89_22_pad_groupi_n_1309, csa_tree_add_89_22_pad_groupi_n_1310, csa_tree_add_89_22_pad_groupi_n_1311, csa_tree_add_89_22_pad_groupi_n_1312, csa_tree_add_89_22_pad_groupi_n_1313;
  wire csa_tree_add_89_22_pad_groupi_n_1314, csa_tree_add_89_22_pad_groupi_n_1315, csa_tree_add_89_22_pad_groupi_n_1316, csa_tree_add_89_22_pad_groupi_n_1317, csa_tree_add_89_22_pad_groupi_n_1318, csa_tree_add_89_22_pad_groupi_n_1319, csa_tree_add_89_22_pad_groupi_n_1320, csa_tree_add_89_22_pad_groupi_n_1321;
  wire csa_tree_add_89_22_pad_groupi_n_1322, csa_tree_add_89_22_pad_groupi_n_1323, csa_tree_add_89_22_pad_groupi_n_1324, csa_tree_add_89_22_pad_groupi_n_1325, csa_tree_add_89_22_pad_groupi_n_1326, csa_tree_add_89_22_pad_groupi_n_1327, csa_tree_add_89_22_pad_groupi_n_1328, csa_tree_add_89_22_pad_groupi_n_1329;
  wire csa_tree_add_89_22_pad_groupi_n_1330, csa_tree_add_89_22_pad_groupi_n_1331, csa_tree_add_89_22_pad_groupi_n_1332, csa_tree_add_89_22_pad_groupi_n_1333, csa_tree_add_89_22_pad_groupi_n_1334, csa_tree_add_89_22_pad_groupi_n_1335, csa_tree_add_89_22_pad_groupi_n_1336, csa_tree_add_89_22_pad_groupi_n_1337;
  wire csa_tree_add_89_22_pad_groupi_n_1338, csa_tree_add_89_22_pad_groupi_n_1339, csa_tree_add_89_22_pad_groupi_n_1340, csa_tree_add_89_22_pad_groupi_n_1341, csa_tree_add_89_22_pad_groupi_n_1342, csa_tree_add_89_22_pad_groupi_n_1343, csa_tree_add_89_22_pad_groupi_n_1344, csa_tree_add_89_22_pad_groupi_n_1345;
  wire csa_tree_add_89_22_pad_groupi_n_1346, csa_tree_add_89_22_pad_groupi_n_1347, csa_tree_add_89_22_pad_groupi_n_1348, csa_tree_add_89_22_pad_groupi_n_1349, csa_tree_add_89_22_pad_groupi_n_1350, csa_tree_add_89_22_pad_groupi_n_1351, csa_tree_add_89_22_pad_groupi_n_1352, csa_tree_add_89_22_pad_groupi_n_1353;
  wire csa_tree_add_89_22_pad_groupi_n_1354, csa_tree_add_89_22_pad_groupi_n_1355, csa_tree_add_89_22_pad_groupi_n_1356, csa_tree_add_89_22_pad_groupi_n_1357, csa_tree_add_89_22_pad_groupi_n_1358, csa_tree_add_89_22_pad_groupi_n_1359, csa_tree_add_89_22_pad_groupi_n_1360, csa_tree_add_89_22_pad_groupi_n_1361;
  wire csa_tree_add_89_22_pad_groupi_n_1362, csa_tree_add_89_22_pad_groupi_n_1363, csa_tree_add_89_22_pad_groupi_n_1364, csa_tree_add_89_22_pad_groupi_n_1365, csa_tree_add_89_22_pad_groupi_n_1366, csa_tree_add_89_22_pad_groupi_n_1367, csa_tree_add_89_22_pad_groupi_n_1368, csa_tree_add_89_22_pad_groupi_n_1369;
  wire csa_tree_add_89_22_pad_groupi_n_1370, csa_tree_add_89_22_pad_groupi_n_1371, csa_tree_add_89_22_pad_groupi_n_1372, csa_tree_add_89_22_pad_groupi_n_1373, csa_tree_add_89_22_pad_groupi_n_1374, csa_tree_add_89_22_pad_groupi_n_1375, csa_tree_add_89_22_pad_groupi_n_1376, csa_tree_add_89_22_pad_groupi_n_1377;
  wire csa_tree_add_89_22_pad_groupi_n_1378, csa_tree_add_89_22_pad_groupi_n_1379, csa_tree_add_89_22_pad_groupi_n_1380, csa_tree_add_89_22_pad_groupi_n_1381, csa_tree_add_89_22_pad_groupi_n_1382, csa_tree_add_89_22_pad_groupi_n_1383, csa_tree_add_89_22_pad_groupi_n_1384, csa_tree_add_89_22_pad_groupi_n_1385;
  wire csa_tree_add_89_22_pad_groupi_n_1386, csa_tree_add_89_22_pad_groupi_n_1387, csa_tree_add_89_22_pad_groupi_n_1388, csa_tree_add_89_22_pad_groupi_n_1389, csa_tree_add_89_22_pad_groupi_n_1390, csa_tree_add_89_22_pad_groupi_n_1391, csa_tree_add_89_22_pad_groupi_n_1392, csa_tree_add_89_22_pad_groupi_n_1393;
  wire csa_tree_add_89_22_pad_groupi_n_1394, csa_tree_add_89_22_pad_groupi_n_1395, csa_tree_add_89_22_pad_groupi_n_1396, csa_tree_add_89_22_pad_groupi_n_1397, csa_tree_add_89_22_pad_groupi_n_1398, csa_tree_add_89_22_pad_groupi_n_1399, csa_tree_add_89_22_pad_groupi_n_1400, csa_tree_add_89_22_pad_groupi_n_1401;
  wire csa_tree_add_89_22_pad_groupi_n_1402, csa_tree_add_89_22_pad_groupi_n_1403, csa_tree_add_89_22_pad_groupi_n_1404, csa_tree_add_89_22_pad_groupi_n_1405, csa_tree_add_89_22_pad_groupi_n_1406, csa_tree_add_89_22_pad_groupi_n_1407, csa_tree_add_89_22_pad_groupi_n_1408, csa_tree_add_89_22_pad_groupi_n_1409;
  wire csa_tree_add_89_22_pad_groupi_n_1410, csa_tree_add_89_22_pad_groupi_n_1411, csa_tree_add_89_22_pad_groupi_n_1412, csa_tree_add_89_22_pad_groupi_n_1413, csa_tree_add_89_22_pad_groupi_n_1414, csa_tree_add_89_22_pad_groupi_n_1415, csa_tree_add_89_22_pad_groupi_n_1416, csa_tree_add_89_22_pad_groupi_n_1417;
  wire csa_tree_add_89_22_pad_groupi_n_1418, csa_tree_add_89_22_pad_groupi_n_1419, csa_tree_add_89_22_pad_groupi_n_1420, csa_tree_add_89_22_pad_groupi_n_1421, csa_tree_add_89_22_pad_groupi_n_1422, csa_tree_add_89_22_pad_groupi_n_1423, csa_tree_add_89_22_pad_groupi_n_1424, csa_tree_add_89_22_pad_groupi_n_1425;
  wire csa_tree_add_89_22_pad_groupi_n_1426, csa_tree_add_89_22_pad_groupi_n_1427, csa_tree_add_89_22_pad_groupi_n_1428, csa_tree_add_89_22_pad_groupi_n_1429, csa_tree_add_89_22_pad_groupi_n_1430, csa_tree_add_89_22_pad_groupi_n_1431, csa_tree_add_89_22_pad_groupi_n_1432, csa_tree_add_89_22_pad_groupi_n_1433;
  wire csa_tree_add_89_22_pad_groupi_n_1434, csa_tree_add_89_22_pad_groupi_n_1435, csa_tree_add_89_22_pad_groupi_n_1436, csa_tree_add_89_22_pad_groupi_n_1437, csa_tree_add_89_22_pad_groupi_n_1438, csa_tree_add_89_22_pad_groupi_n_1439, csa_tree_add_89_22_pad_groupi_n_1440, csa_tree_add_89_22_pad_groupi_n_1441;
  wire csa_tree_add_89_22_pad_groupi_n_1442, csa_tree_add_89_22_pad_groupi_n_1443, csa_tree_add_89_22_pad_groupi_n_1444, csa_tree_add_89_22_pad_groupi_n_1445, csa_tree_add_89_22_pad_groupi_n_1446, csa_tree_add_89_22_pad_groupi_n_1447, csa_tree_add_89_22_pad_groupi_n_1448, csa_tree_add_89_22_pad_groupi_n_1449;
  wire csa_tree_add_89_22_pad_groupi_n_1450, csa_tree_add_89_22_pad_groupi_n_1451, csa_tree_add_89_22_pad_groupi_n_1452, csa_tree_add_89_22_pad_groupi_n_1453, csa_tree_add_89_22_pad_groupi_n_1454, csa_tree_add_89_22_pad_groupi_n_1455, csa_tree_add_89_22_pad_groupi_n_1456, csa_tree_add_89_22_pad_groupi_n_1457;
  wire csa_tree_add_89_22_pad_groupi_n_1458, csa_tree_add_89_22_pad_groupi_n_1459, csa_tree_add_89_22_pad_groupi_n_1460, csa_tree_add_89_22_pad_groupi_n_1461, csa_tree_add_89_22_pad_groupi_n_1462, csa_tree_add_89_22_pad_groupi_n_1463, csa_tree_add_89_22_pad_groupi_n_1464, csa_tree_add_89_22_pad_groupi_n_1465;
  wire csa_tree_add_89_22_pad_groupi_n_1466, csa_tree_add_89_22_pad_groupi_n_1467, csa_tree_add_89_22_pad_groupi_n_1468, csa_tree_add_89_22_pad_groupi_n_1469, csa_tree_add_89_22_pad_groupi_n_1470, csa_tree_add_89_22_pad_groupi_n_1471, csa_tree_add_89_22_pad_groupi_n_1472, csa_tree_add_89_22_pad_groupi_n_1473;
  wire csa_tree_add_89_22_pad_groupi_n_1474, csa_tree_add_89_22_pad_groupi_n_1475, csa_tree_add_89_22_pad_groupi_n_1476, csa_tree_add_89_22_pad_groupi_n_1477, csa_tree_add_89_22_pad_groupi_n_1478, csa_tree_add_89_22_pad_groupi_n_1479, csa_tree_add_89_22_pad_groupi_n_1480, csa_tree_add_89_22_pad_groupi_n_1481;
  wire csa_tree_add_89_22_pad_groupi_n_1482, csa_tree_add_89_22_pad_groupi_n_1483, csa_tree_add_89_22_pad_groupi_n_1484, csa_tree_add_89_22_pad_groupi_n_1485, csa_tree_add_89_22_pad_groupi_n_1486, csa_tree_add_89_22_pad_groupi_n_1487, csa_tree_add_89_22_pad_groupi_n_1488, csa_tree_add_89_22_pad_groupi_n_1489;
  wire csa_tree_add_89_22_pad_groupi_n_1490, csa_tree_add_89_22_pad_groupi_n_1491, csa_tree_add_89_22_pad_groupi_n_1492, csa_tree_add_89_22_pad_groupi_n_1493, csa_tree_add_89_22_pad_groupi_n_1494, csa_tree_add_89_22_pad_groupi_n_1495, csa_tree_add_89_22_pad_groupi_n_1496, csa_tree_add_89_22_pad_groupi_n_1497;
  wire csa_tree_add_89_22_pad_groupi_n_1498, csa_tree_add_89_22_pad_groupi_n_1499, csa_tree_add_89_22_pad_groupi_n_1500, csa_tree_add_89_22_pad_groupi_n_1501, csa_tree_add_89_22_pad_groupi_n_1502, csa_tree_add_89_22_pad_groupi_n_1503, csa_tree_add_89_22_pad_groupi_n_1505, csa_tree_add_89_22_pad_groupi_n_1506;
  wire csa_tree_add_89_22_pad_groupi_n_1507, csa_tree_add_89_22_pad_groupi_n_1508, csa_tree_add_89_22_pad_groupi_n_1509, csa_tree_add_89_22_pad_groupi_n_1510, csa_tree_add_89_22_pad_groupi_n_1511, csa_tree_add_89_22_pad_groupi_n_1512, csa_tree_add_89_22_pad_groupi_n_1513, csa_tree_add_89_22_pad_groupi_n_1514;
  wire csa_tree_add_89_22_pad_groupi_n_1515, csa_tree_add_89_22_pad_groupi_n_1516, csa_tree_add_89_22_pad_groupi_n_1517, csa_tree_add_89_22_pad_groupi_n_1518, csa_tree_add_89_22_pad_groupi_n_1519, csa_tree_add_89_22_pad_groupi_n_1520, csa_tree_add_89_22_pad_groupi_n_1521, csa_tree_add_89_22_pad_groupi_n_1522;
  wire csa_tree_add_89_22_pad_groupi_n_1523, csa_tree_add_89_22_pad_groupi_n_1524, csa_tree_add_89_22_pad_groupi_n_1525, csa_tree_add_89_22_pad_groupi_n_1526, csa_tree_add_89_22_pad_groupi_n_1527, csa_tree_add_89_22_pad_groupi_n_1529, csa_tree_add_89_22_pad_groupi_n_1530, csa_tree_add_89_22_pad_groupi_n_1532;
  wire csa_tree_add_89_22_pad_groupi_n_1533, csa_tree_add_89_22_pad_groupi_n_1534, csa_tree_add_89_22_pad_groupi_n_1535, csa_tree_add_89_22_pad_groupi_n_1537, csa_tree_add_89_22_pad_groupi_n_1538, csa_tree_add_89_22_pad_groupi_n_1539, csa_tree_add_89_22_pad_groupi_n_1540, csa_tree_add_89_22_pad_groupi_n_1542;
  wire csa_tree_add_89_22_pad_groupi_n_1543, csa_tree_add_89_22_pad_groupi_n_1544, csa_tree_add_89_22_pad_groupi_n_1546, csa_tree_add_89_22_pad_groupi_n_1547, csa_tree_add_89_22_pad_groupi_n_1549, csa_tree_add_89_22_pad_groupi_n_1550, csa_tree_add_89_22_pad_groupi_n_1552, csa_tree_add_89_22_pad_groupi_n_1553;
  wire csa_tree_add_89_22_pad_groupi_n_1555, csa_tree_add_89_22_pad_groupi_n_1556, csa_tree_add_89_22_pad_groupi_n_1558, csa_tree_add_95_22_pad_groupi_n_0, csa_tree_add_95_22_pad_groupi_n_1, csa_tree_add_95_22_pad_groupi_n_3, csa_tree_add_95_22_pad_groupi_n_4, csa_tree_add_95_22_pad_groupi_n_5;
  wire csa_tree_add_95_22_pad_groupi_n_6, csa_tree_add_95_22_pad_groupi_n_12, csa_tree_add_95_22_pad_groupi_n_13, csa_tree_add_95_22_pad_groupi_n_14, csa_tree_add_95_22_pad_groupi_n_15, csa_tree_add_95_22_pad_groupi_n_16, csa_tree_add_95_22_pad_groupi_n_17, csa_tree_add_95_22_pad_groupi_n_18;
  wire csa_tree_add_95_22_pad_groupi_n_19, csa_tree_add_95_22_pad_groupi_n_20, csa_tree_add_95_22_pad_groupi_n_21, csa_tree_add_95_22_pad_groupi_n_22, csa_tree_add_95_22_pad_groupi_n_23, csa_tree_add_95_22_pad_groupi_n_24, csa_tree_add_95_22_pad_groupi_n_25, csa_tree_add_95_22_pad_groupi_n_26;
  wire csa_tree_add_95_22_pad_groupi_n_27, csa_tree_add_95_22_pad_groupi_n_28, csa_tree_add_95_22_pad_groupi_n_29, csa_tree_add_95_22_pad_groupi_n_30, csa_tree_add_95_22_pad_groupi_n_31, csa_tree_add_95_22_pad_groupi_n_32, csa_tree_add_95_22_pad_groupi_n_33, csa_tree_add_95_22_pad_groupi_n_34;
  wire csa_tree_add_95_22_pad_groupi_n_35, csa_tree_add_95_22_pad_groupi_n_36, csa_tree_add_95_22_pad_groupi_n_37, csa_tree_add_95_22_pad_groupi_n_38, csa_tree_add_95_22_pad_groupi_n_39, csa_tree_add_95_22_pad_groupi_n_40, csa_tree_add_95_22_pad_groupi_n_41, csa_tree_add_95_22_pad_groupi_n_42;
  wire csa_tree_add_95_22_pad_groupi_n_43, csa_tree_add_95_22_pad_groupi_n_45, csa_tree_add_95_22_pad_groupi_n_46, csa_tree_add_95_22_pad_groupi_n_47, csa_tree_add_95_22_pad_groupi_n_48, csa_tree_add_95_22_pad_groupi_n_50, csa_tree_add_95_22_pad_groupi_n_51, csa_tree_add_95_22_pad_groupi_n_52;
  wire csa_tree_add_95_22_pad_groupi_n_53, csa_tree_add_95_22_pad_groupi_n_54, csa_tree_add_95_22_pad_groupi_n_55, csa_tree_add_95_22_pad_groupi_n_56, csa_tree_add_95_22_pad_groupi_n_57, csa_tree_add_95_22_pad_groupi_n_58, csa_tree_add_95_22_pad_groupi_n_59, csa_tree_add_95_22_pad_groupi_n_60;
  wire csa_tree_add_95_22_pad_groupi_n_61, csa_tree_add_95_22_pad_groupi_n_62, csa_tree_add_95_22_pad_groupi_n_64, csa_tree_add_95_22_pad_groupi_n_65, csa_tree_add_95_22_pad_groupi_n_66, csa_tree_add_95_22_pad_groupi_n_67, csa_tree_add_95_22_pad_groupi_n_68, csa_tree_add_95_22_pad_groupi_n_69;
  wire csa_tree_add_95_22_pad_groupi_n_70, csa_tree_add_95_22_pad_groupi_n_71, csa_tree_add_95_22_pad_groupi_n_72, csa_tree_add_95_22_pad_groupi_n_73, csa_tree_add_95_22_pad_groupi_n_74, csa_tree_add_95_22_pad_groupi_n_75, csa_tree_add_95_22_pad_groupi_n_76, csa_tree_add_95_22_pad_groupi_n_77;
  wire csa_tree_add_95_22_pad_groupi_n_78, csa_tree_add_95_22_pad_groupi_n_79, csa_tree_add_95_22_pad_groupi_n_80, csa_tree_add_95_22_pad_groupi_n_82, csa_tree_add_95_22_pad_groupi_n_83, csa_tree_add_95_22_pad_groupi_n_84, csa_tree_add_95_22_pad_groupi_n_85, csa_tree_add_95_22_pad_groupi_n_86;
  wire csa_tree_add_95_22_pad_groupi_n_87, csa_tree_add_95_22_pad_groupi_n_88, csa_tree_add_95_22_pad_groupi_n_89, csa_tree_add_95_22_pad_groupi_n_90, csa_tree_add_95_22_pad_groupi_n_91, csa_tree_add_95_22_pad_groupi_n_92, csa_tree_add_95_22_pad_groupi_n_93, csa_tree_add_95_22_pad_groupi_n_94;
  wire csa_tree_add_95_22_pad_groupi_n_95, csa_tree_add_95_22_pad_groupi_n_96, csa_tree_add_95_22_pad_groupi_n_97, csa_tree_add_95_22_pad_groupi_n_98, csa_tree_add_95_22_pad_groupi_n_99, csa_tree_add_95_22_pad_groupi_n_100, csa_tree_add_95_22_pad_groupi_n_101, csa_tree_add_95_22_pad_groupi_n_102;
  wire csa_tree_add_95_22_pad_groupi_n_103, csa_tree_add_95_22_pad_groupi_n_104, csa_tree_add_95_22_pad_groupi_n_105, csa_tree_add_95_22_pad_groupi_n_106, csa_tree_add_95_22_pad_groupi_n_107, csa_tree_add_95_22_pad_groupi_n_108, csa_tree_add_95_22_pad_groupi_n_109, csa_tree_add_95_22_pad_groupi_n_110;
  wire csa_tree_add_95_22_pad_groupi_n_111, csa_tree_add_95_22_pad_groupi_n_112, csa_tree_add_95_22_pad_groupi_n_113, csa_tree_add_95_22_pad_groupi_n_114, csa_tree_add_95_22_pad_groupi_n_115, csa_tree_add_95_22_pad_groupi_n_116, csa_tree_add_95_22_pad_groupi_n_117, csa_tree_add_95_22_pad_groupi_n_118;
  wire csa_tree_add_95_22_pad_groupi_n_119, csa_tree_add_95_22_pad_groupi_n_120, csa_tree_add_95_22_pad_groupi_n_121, csa_tree_add_95_22_pad_groupi_n_122, csa_tree_add_95_22_pad_groupi_n_123, csa_tree_add_95_22_pad_groupi_n_124, csa_tree_add_95_22_pad_groupi_n_125, csa_tree_add_95_22_pad_groupi_n_126;
  wire csa_tree_add_95_22_pad_groupi_n_127, csa_tree_add_95_22_pad_groupi_n_128, csa_tree_add_95_22_pad_groupi_n_129, csa_tree_add_95_22_pad_groupi_n_130, csa_tree_add_95_22_pad_groupi_n_131, csa_tree_add_95_22_pad_groupi_n_132, csa_tree_add_95_22_pad_groupi_n_133, csa_tree_add_95_22_pad_groupi_n_134;
  wire csa_tree_add_95_22_pad_groupi_n_135, csa_tree_add_95_22_pad_groupi_n_136, csa_tree_add_95_22_pad_groupi_n_137, csa_tree_add_95_22_pad_groupi_n_138, csa_tree_add_95_22_pad_groupi_n_139, csa_tree_add_95_22_pad_groupi_n_140, csa_tree_add_95_22_pad_groupi_n_141, csa_tree_add_95_22_pad_groupi_n_142;
  wire csa_tree_add_95_22_pad_groupi_n_143, csa_tree_add_95_22_pad_groupi_n_144, csa_tree_add_95_22_pad_groupi_n_145, csa_tree_add_95_22_pad_groupi_n_146, csa_tree_add_95_22_pad_groupi_n_147, csa_tree_add_95_22_pad_groupi_n_148, csa_tree_add_95_22_pad_groupi_n_149, csa_tree_add_95_22_pad_groupi_n_150;
  wire csa_tree_add_95_22_pad_groupi_n_151, csa_tree_add_95_22_pad_groupi_n_152, csa_tree_add_95_22_pad_groupi_n_153, csa_tree_add_95_22_pad_groupi_n_154, csa_tree_add_95_22_pad_groupi_n_155, csa_tree_add_95_22_pad_groupi_n_158, csa_tree_add_95_22_pad_groupi_n_159, csa_tree_add_95_22_pad_groupi_n_160;
  wire csa_tree_add_95_22_pad_groupi_n_161, csa_tree_add_95_22_pad_groupi_n_162, csa_tree_add_95_22_pad_groupi_n_163, csa_tree_add_95_22_pad_groupi_n_164, csa_tree_add_95_22_pad_groupi_n_165, csa_tree_add_95_22_pad_groupi_n_166, csa_tree_add_95_22_pad_groupi_n_167, csa_tree_add_95_22_pad_groupi_n_168;
  wire csa_tree_add_95_22_pad_groupi_n_169, csa_tree_add_95_22_pad_groupi_n_170, csa_tree_add_95_22_pad_groupi_n_171, csa_tree_add_95_22_pad_groupi_n_172, csa_tree_add_95_22_pad_groupi_n_173, csa_tree_add_95_22_pad_groupi_n_174, csa_tree_add_95_22_pad_groupi_n_175, csa_tree_add_95_22_pad_groupi_n_176;
  wire csa_tree_add_95_22_pad_groupi_n_177, csa_tree_add_95_22_pad_groupi_n_178, csa_tree_add_95_22_pad_groupi_n_179, csa_tree_add_95_22_pad_groupi_n_180, csa_tree_add_95_22_pad_groupi_n_181, csa_tree_add_95_22_pad_groupi_n_182, csa_tree_add_95_22_pad_groupi_n_183, csa_tree_add_95_22_pad_groupi_n_184;
  wire csa_tree_add_95_22_pad_groupi_n_185, csa_tree_add_95_22_pad_groupi_n_186, csa_tree_add_95_22_pad_groupi_n_187, csa_tree_add_95_22_pad_groupi_n_188, csa_tree_add_95_22_pad_groupi_n_189, csa_tree_add_95_22_pad_groupi_n_190, csa_tree_add_95_22_pad_groupi_n_191, csa_tree_add_95_22_pad_groupi_n_192;
  wire csa_tree_add_95_22_pad_groupi_n_193, csa_tree_add_95_22_pad_groupi_n_194, csa_tree_add_95_22_pad_groupi_n_195, csa_tree_add_95_22_pad_groupi_n_196, csa_tree_add_95_22_pad_groupi_n_197, csa_tree_add_95_22_pad_groupi_n_198, csa_tree_add_95_22_pad_groupi_n_200, csa_tree_add_95_22_pad_groupi_n_201;
  wire csa_tree_add_95_22_pad_groupi_n_202, csa_tree_add_95_22_pad_groupi_n_203, csa_tree_add_95_22_pad_groupi_n_204, csa_tree_add_95_22_pad_groupi_n_205, csa_tree_add_95_22_pad_groupi_n_206, csa_tree_add_95_22_pad_groupi_n_207, csa_tree_add_95_22_pad_groupi_n_208, csa_tree_add_95_22_pad_groupi_n_209;
  wire csa_tree_add_95_22_pad_groupi_n_210, csa_tree_add_95_22_pad_groupi_n_211, csa_tree_add_95_22_pad_groupi_n_212, csa_tree_add_95_22_pad_groupi_n_213, csa_tree_add_95_22_pad_groupi_n_214, csa_tree_add_95_22_pad_groupi_n_215, csa_tree_add_95_22_pad_groupi_n_216, csa_tree_add_95_22_pad_groupi_n_217;
  wire csa_tree_add_95_22_pad_groupi_n_218, csa_tree_add_95_22_pad_groupi_n_219, csa_tree_add_95_22_pad_groupi_n_220, csa_tree_add_95_22_pad_groupi_n_221, csa_tree_add_95_22_pad_groupi_n_222, csa_tree_add_95_22_pad_groupi_n_223, csa_tree_add_95_22_pad_groupi_n_224, csa_tree_add_95_22_pad_groupi_n_225;
  wire csa_tree_add_95_22_pad_groupi_n_226, csa_tree_add_95_22_pad_groupi_n_227, csa_tree_add_95_22_pad_groupi_n_228, csa_tree_add_95_22_pad_groupi_n_229, csa_tree_add_95_22_pad_groupi_n_230, csa_tree_add_95_22_pad_groupi_n_231, csa_tree_add_95_22_pad_groupi_n_232, csa_tree_add_95_22_pad_groupi_n_233;
  wire csa_tree_add_95_22_pad_groupi_n_234, csa_tree_add_95_22_pad_groupi_n_235, csa_tree_add_95_22_pad_groupi_n_236, csa_tree_add_95_22_pad_groupi_n_237, csa_tree_add_95_22_pad_groupi_n_238, csa_tree_add_95_22_pad_groupi_n_239, csa_tree_add_95_22_pad_groupi_n_240, csa_tree_add_95_22_pad_groupi_n_241;
  wire csa_tree_add_95_22_pad_groupi_n_242, csa_tree_add_95_22_pad_groupi_n_243, csa_tree_add_95_22_pad_groupi_n_244, csa_tree_add_95_22_pad_groupi_n_245, csa_tree_add_95_22_pad_groupi_n_246, csa_tree_add_95_22_pad_groupi_n_247, csa_tree_add_95_22_pad_groupi_n_248, csa_tree_add_95_22_pad_groupi_n_249;
  wire csa_tree_add_95_22_pad_groupi_n_250, csa_tree_add_95_22_pad_groupi_n_251, csa_tree_add_95_22_pad_groupi_n_252, csa_tree_add_95_22_pad_groupi_n_253, csa_tree_add_95_22_pad_groupi_n_254, csa_tree_add_95_22_pad_groupi_n_255, csa_tree_add_95_22_pad_groupi_n_256, csa_tree_add_95_22_pad_groupi_n_257;
  wire csa_tree_add_95_22_pad_groupi_n_258, csa_tree_add_95_22_pad_groupi_n_259, csa_tree_add_95_22_pad_groupi_n_260, csa_tree_add_95_22_pad_groupi_n_261, csa_tree_add_95_22_pad_groupi_n_262, csa_tree_add_95_22_pad_groupi_n_263, csa_tree_add_95_22_pad_groupi_n_264, csa_tree_add_95_22_pad_groupi_n_265;
  wire csa_tree_add_95_22_pad_groupi_n_266, csa_tree_add_95_22_pad_groupi_n_267, csa_tree_add_95_22_pad_groupi_n_268, csa_tree_add_95_22_pad_groupi_n_269, csa_tree_add_95_22_pad_groupi_n_270, csa_tree_add_95_22_pad_groupi_n_271, csa_tree_add_95_22_pad_groupi_n_272, csa_tree_add_95_22_pad_groupi_n_273;
  wire csa_tree_add_95_22_pad_groupi_n_274, csa_tree_add_95_22_pad_groupi_n_275, csa_tree_add_95_22_pad_groupi_n_276, csa_tree_add_95_22_pad_groupi_n_277, csa_tree_add_95_22_pad_groupi_n_278, csa_tree_add_95_22_pad_groupi_n_279, csa_tree_add_95_22_pad_groupi_n_280, csa_tree_add_95_22_pad_groupi_n_281;
  wire csa_tree_add_95_22_pad_groupi_n_282, csa_tree_add_95_22_pad_groupi_n_283, csa_tree_add_95_22_pad_groupi_n_284, csa_tree_add_95_22_pad_groupi_n_285, csa_tree_add_95_22_pad_groupi_n_286, csa_tree_add_95_22_pad_groupi_n_287, csa_tree_add_95_22_pad_groupi_n_288, csa_tree_add_95_22_pad_groupi_n_289;
  wire csa_tree_add_95_22_pad_groupi_n_290, csa_tree_add_95_22_pad_groupi_n_291, csa_tree_add_95_22_pad_groupi_n_292, csa_tree_add_95_22_pad_groupi_n_293, csa_tree_add_95_22_pad_groupi_n_294, csa_tree_add_95_22_pad_groupi_n_295, csa_tree_add_95_22_pad_groupi_n_296, csa_tree_add_95_22_pad_groupi_n_297;
  wire csa_tree_add_95_22_pad_groupi_n_298, csa_tree_add_95_22_pad_groupi_n_299, csa_tree_add_95_22_pad_groupi_n_300, csa_tree_add_95_22_pad_groupi_n_301, csa_tree_add_95_22_pad_groupi_n_302, csa_tree_add_95_22_pad_groupi_n_303, csa_tree_add_95_22_pad_groupi_n_304, csa_tree_add_95_22_pad_groupi_n_305;
  wire csa_tree_add_95_22_pad_groupi_n_306, csa_tree_add_95_22_pad_groupi_n_307, csa_tree_add_95_22_pad_groupi_n_308, csa_tree_add_95_22_pad_groupi_n_309, csa_tree_add_95_22_pad_groupi_n_310, csa_tree_add_95_22_pad_groupi_n_311, csa_tree_add_95_22_pad_groupi_n_312, csa_tree_add_95_22_pad_groupi_n_313;
  wire csa_tree_add_95_22_pad_groupi_n_314, csa_tree_add_95_22_pad_groupi_n_315, csa_tree_add_95_22_pad_groupi_n_316, csa_tree_add_95_22_pad_groupi_n_317, csa_tree_add_95_22_pad_groupi_n_318, csa_tree_add_95_22_pad_groupi_n_319, csa_tree_add_95_22_pad_groupi_n_320, csa_tree_add_95_22_pad_groupi_n_321;
  wire csa_tree_add_95_22_pad_groupi_n_322, csa_tree_add_95_22_pad_groupi_n_323, csa_tree_add_95_22_pad_groupi_n_324, csa_tree_add_95_22_pad_groupi_n_325, csa_tree_add_95_22_pad_groupi_n_326, csa_tree_add_95_22_pad_groupi_n_327, csa_tree_add_95_22_pad_groupi_n_328, csa_tree_add_95_22_pad_groupi_n_329;
  wire csa_tree_add_95_22_pad_groupi_n_330, csa_tree_add_95_22_pad_groupi_n_331, csa_tree_add_95_22_pad_groupi_n_332, csa_tree_add_95_22_pad_groupi_n_333, csa_tree_add_95_22_pad_groupi_n_334, csa_tree_add_95_22_pad_groupi_n_335, csa_tree_add_95_22_pad_groupi_n_336, csa_tree_add_95_22_pad_groupi_n_337;
  wire csa_tree_add_95_22_pad_groupi_n_338, csa_tree_add_95_22_pad_groupi_n_339, csa_tree_add_95_22_pad_groupi_n_340, csa_tree_add_95_22_pad_groupi_n_341, csa_tree_add_95_22_pad_groupi_n_342, csa_tree_add_95_22_pad_groupi_n_343, csa_tree_add_95_22_pad_groupi_n_344, csa_tree_add_95_22_pad_groupi_n_345;
  wire csa_tree_add_95_22_pad_groupi_n_346, csa_tree_add_95_22_pad_groupi_n_347, csa_tree_add_95_22_pad_groupi_n_348, csa_tree_add_95_22_pad_groupi_n_349, csa_tree_add_95_22_pad_groupi_n_350, csa_tree_add_95_22_pad_groupi_n_351, csa_tree_add_95_22_pad_groupi_n_352, csa_tree_add_95_22_pad_groupi_n_353;
  wire csa_tree_add_95_22_pad_groupi_n_354, csa_tree_add_95_22_pad_groupi_n_355, csa_tree_add_95_22_pad_groupi_n_356, csa_tree_add_95_22_pad_groupi_n_357, csa_tree_add_95_22_pad_groupi_n_358, csa_tree_add_95_22_pad_groupi_n_359, csa_tree_add_95_22_pad_groupi_n_361, csa_tree_add_95_22_pad_groupi_n_362;
  wire csa_tree_add_95_22_pad_groupi_n_363, csa_tree_add_95_22_pad_groupi_n_364, csa_tree_add_95_22_pad_groupi_n_365, csa_tree_add_95_22_pad_groupi_n_366, csa_tree_add_95_22_pad_groupi_n_367, csa_tree_add_95_22_pad_groupi_n_368, csa_tree_add_95_22_pad_groupi_n_369, csa_tree_add_95_22_pad_groupi_n_370;
  wire csa_tree_add_95_22_pad_groupi_n_371, csa_tree_add_95_22_pad_groupi_n_372, csa_tree_add_95_22_pad_groupi_n_373, csa_tree_add_95_22_pad_groupi_n_374, csa_tree_add_95_22_pad_groupi_n_375, csa_tree_add_95_22_pad_groupi_n_376, csa_tree_add_95_22_pad_groupi_n_377, csa_tree_add_95_22_pad_groupi_n_378;
  wire csa_tree_add_95_22_pad_groupi_n_379, csa_tree_add_95_22_pad_groupi_n_380, csa_tree_add_95_22_pad_groupi_n_381, csa_tree_add_95_22_pad_groupi_n_382, csa_tree_add_95_22_pad_groupi_n_383, csa_tree_add_95_22_pad_groupi_n_384, csa_tree_add_95_22_pad_groupi_n_385, csa_tree_add_95_22_pad_groupi_n_386;
  wire csa_tree_add_95_22_pad_groupi_n_387, csa_tree_add_95_22_pad_groupi_n_388, csa_tree_add_95_22_pad_groupi_n_389, csa_tree_add_95_22_pad_groupi_n_390, csa_tree_add_95_22_pad_groupi_n_391, csa_tree_add_95_22_pad_groupi_n_392, csa_tree_add_95_22_pad_groupi_n_393, csa_tree_add_95_22_pad_groupi_n_394;
  wire csa_tree_add_95_22_pad_groupi_n_395, csa_tree_add_95_22_pad_groupi_n_396, csa_tree_add_95_22_pad_groupi_n_397, csa_tree_add_95_22_pad_groupi_n_398, csa_tree_add_95_22_pad_groupi_n_399, csa_tree_add_95_22_pad_groupi_n_401, csa_tree_add_95_22_pad_groupi_n_402, csa_tree_add_95_22_pad_groupi_n_403;
  wire csa_tree_add_95_22_pad_groupi_n_404, csa_tree_add_95_22_pad_groupi_n_406, csa_tree_add_95_22_pad_groupi_n_409, csa_tree_add_95_22_pad_groupi_n_410, csa_tree_add_95_22_pad_groupi_n_411, csa_tree_add_95_22_pad_groupi_n_412, csa_tree_add_95_22_pad_groupi_n_413, csa_tree_add_95_22_pad_groupi_n_414;
  wire csa_tree_add_95_22_pad_groupi_n_415, csa_tree_add_95_22_pad_groupi_n_416, csa_tree_add_95_22_pad_groupi_n_417, csa_tree_add_95_22_pad_groupi_n_418, csa_tree_add_95_22_pad_groupi_n_419, csa_tree_add_95_22_pad_groupi_n_420, csa_tree_add_95_22_pad_groupi_n_421, csa_tree_add_95_22_pad_groupi_n_422;
  wire csa_tree_add_95_22_pad_groupi_n_423, csa_tree_add_95_22_pad_groupi_n_424, csa_tree_add_95_22_pad_groupi_n_425, csa_tree_add_95_22_pad_groupi_n_426, csa_tree_add_95_22_pad_groupi_n_427, csa_tree_add_95_22_pad_groupi_n_428, csa_tree_add_95_22_pad_groupi_n_429, csa_tree_add_95_22_pad_groupi_n_430;
  wire csa_tree_add_95_22_pad_groupi_n_431, csa_tree_add_95_22_pad_groupi_n_432, csa_tree_add_95_22_pad_groupi_n_433, csa_tree_add_95_22_pad_groupi_n_434, csa_tree_add_95_22_pad_groupi_n_435, csa_tree_add_95_22_pad_groupi_n_438, csa_tree_add_95_22_pad_groupi_n_439, csa_tree_add_95_22_pad_groupi_n_445;
  wire csa_tree_add_95_22_pad_groupi_n_455, csa_tree_add_95_22_pad_groupi_n_456, csa_tree_add_95_22_pad_groupi_n_457, csa_tree_add_95_22_pad_groupi_n_458, csa_tree_add_95_22_pad_groupi_n_459, csa_tree_add_95_22_pad_groupi_n_460, csa_tree_add_95_22_pad_groupi_n_461, csa_tree_add_95_22_pad_groupi_n_462;
  wire csa_tree_add_95_22_pad_groupi_n_463, csa_tree_add_95_22_pad_groupi_n_464, csa_tree_add_95_22_pad_groupi_n_465, csa_tree_add_95_22_pad_groupi_n_466, csa_tree_add_95_22_pad_groupi_n_467, csa_tree_add_95_22_pad_groupi_n_468, csa_tree_add_95_22_pad_groupi_n_469, csa_tree_add_95_22_pad_groupi_n_470;
  wire csa_tree_add_95_22_pad_groupi_n_471, csa_tree_add_95_22_pad_groupi_n_472, csa_tree_add_95_22_pad_groupi_n_473, csa_tree_add_95_22_pad_groupi_n_474, csa_tree_add_95_22_pad_groupi_n_475, csa_tree_add_95_22_pad_groupi_n_476, csa_tree_add_95_22_pad_groupi_n_477, csa_tree_add_95_22_pad_groupi_n_478;
  wire csa_tree_add_95_22_pad_groupi_n_479, csa_tree_add_95_22_pad_groupi_n_480, csa_tree_add_95_22_pad_groupi_n_481, csa_tree_add_95_22_pad_groupi_n_482, csa_tree_add_95_22_pad_groupi_n_483, csa_tree_add_95_22_pad_groupi_n_484, csa_tree_add_95_22_pad_groupi_n_485, csa_tree_add_95_22_pad_groupi_n_486;
  wire csa_tree_add_95_22_pad_groupi_n_487, csa_tree_add_95_22_pad_groupi_n_488, csa_tree_add_95_22_pad_groupi_n_489, csa_tree_add_95_22_pad_groupi_n_490, csa_tree_add_95_22_pad_groupi_n_491, csa_tree_add_95_22_pad_groupi_n_492, csa_tree_add_95_22_pad_groupi_n_493, csa_tree_add_95_22_pad_groupi_n_494;
  wire csa_tree_add_95_22_pad_groupi_n_495, csa_tree_add_95_22_pad_groupi_n_496, csa_tree_add_95_22_pad_groupi_n_497, csa_tree_add_95_22_pad_groupi_n_498, csa_tree_add_95_22_pad_groupi_n_499, csa_tree_add_95_22_pad_groupi_n_500, csa_tree_add_95_22_pad_groupi_n_501, csa_tree_add_95_22_pad_groupi_n_502;
  wire csa_tree_add_95_22_pad_groupi_n_503, csa_tree_add_95_22_pad_groupi_n_504, csa_tree_add_95_22_pad_groupi_n_505, csa_tree_add_95_22_pad_groupi_n_506, csa_tree_add_95_22_pad_groupi_n_507, csa_tree_add_95_22_pad_groupi_n_508, csa_tree_add_95_22_pad_groupi_n_509, csa_tree_add_95_22_pad_groupi_n_510;
  wire csa_tree_add_95_22_pad_groupi_n_511, csa_tree_add_95_22_pad_groupi_n_512, csa_tree_add_95_22_pad_groupi_n_513, csa_tree_add_95_22_pad_groupi_n_514, csa_tree_add_95_22_pad_groupi_n_515, csa_tree_add_95_22_pad_groupi_n_516, csa_tree_add_95_22_pad_groupi_n_517, csa_tree_add_95_22_pad_groupi_n_518;
  wire csa_tree_add_95_22_pad_groupi_n_519, csa_tree_add_95_22_pad_groupi_n_520, csa_tree_add_95_22_pad_groupi_n_521, csa_tree_add_95_22_pad_groupi_n_522, csa_tree_add_95_22_pad_groupi_n_523, csa_tree_add_95_22_pad_groupi_n_524, csa_tree_add_95_22_pad_groupi_n_525, csa_tree_add_95_22_pad_groupi_n_526;
  wire csa_tree_add_95_22_pad_groupi_n_527, csa_tree_add_95_22_pad_groupi_n_528, csa_tree_add_95_22_pad_groupi_n_529, csa_tree_add_95_22_pad_groupi_n_530, csa_tree_add_95_22_pad_groupi_n_531, csa_tree_add_95_22_pad_groupi_n_532, csa_tree_add_95_22_pad_groupi_n_533, csa_tree_add_95_22_pad_groupi_n_534;
  wire csa_tree_add_95_22_pad_groupi_n_535, csa_tree_add_95_22_pad_groupi_n_536, csa_tree_add_95_22_pad_groupi_n_537, csa_tree_add_95_22_pad_groupi_n_538, csa_tree_add_95_22_pad_groupi_n_539, csa_tree_add_95_22_pad_groupi_n_540, csa_tree_add_95_22_pad_groupi_n_541, csa_tree_add_95_22_pad_groupi_n_542;
  wire csa_tree_add_95_22_pad_groupi_n_543, csa_tree_add_95_22_pad_groupi_n_544, csa_tree_add_95_22_pad_groupi_n_545, csa_tree_add_95_22_pad_groupi_n_546, csa_tree_add_95_22_pad_groupi_n_547, csa_tree_add_95_22_pad_groupi_n_548, csa_tree_add_95_22_pad_groupi_n_549, csa_tree_add_95_22_pad_groupi_n_550;
  wire csa_tree_add_95_22_pad_groupi_n_551, csa_tree_add_95_22_pad_groupi_n_552, csa_tree_add_95_22_pad_groupi_n_553, csa_tree_add_95_22_pad_groupi_n_554, csa_tree_add_95_22_pad_groupi_n_555, csa_tree_add_95_22_pad_groupi_n_556, csa_tree_add_95_22_pad_groupi_n_557, csa_tree_add_95_22_pad_groupi_n_559;
  wire csa_tree_add_95_22_pad_groupi_n_561, csa_tree_add_95_22_pad_groupi_n_562, csa_tree_add_95_22_pad_groupi_n_563, csa_tree_add_95_22_pad_groupi_n_564, csa_tree_add_95_22_pad_groupi_n_565, csa_tree_add_95_22_pad_groupi_n_566, csa_tree_add_95_22_pad_groupi_n_567, csa_tree_add_95_22_pad_groupi_n_568;
  wire csa_tree_add_95_22_pad_groupi_n_569, csa_tree_add_95_22_pad_groupi_n_570, csa_tree_add_95_22_pad_groupi_n_572, csa_tree_add_95_22_pad_groupi_n_573, csa_tree_add_95_22_pad_groupi_n_574, csa_tree_add_95_22_pad_groupi_n_575, csa_tree_add_95_22_pad_groupi_n_576, csa_tree_add_95_22_pad_groupi_n_577;
  wire csa_tree_add_95_22_pad_groupi_n_578, csa_tree_add_95_22_pad_groupi_n_579, csa_tree_add_95_22_pad_groupi_n_580, csa_tree_add_95_22_pad_groupi_n_581, csa_tree_add_95_22_pad_groupi_n_582, csa_tree_add_95_22_pad_groupi_n_583, csa_tree_add_95_22_pad_groupi_n_584, csa_tree_add_95_22_pad_groupi_n_586;
  wire csa_tree_add_95_22_pad_groupi_n_587, csa_tree_add_95_22_pad_groupi_n_588, csa_tree_add_95_22_pad_groupi_n_589, csa_tree_add_95_22_pad_groupi_n_590, csa_tree_add_95_22_pad_groupi_n_591, csa_tree_add_95_22_pad_groupi_n_592, csa_tree_add_95_22_pad_groupi_n_593, csa_tree_add_95_22_pad_groupi_n_594;
  wire csa_tree_add_95_22_pad_groupi_n_595, csa_tree_add_95_22_pad_groupi_n_598, csa_tree_add_95_22_pad_groupi_n_599, csa_tree_add_95_22_pad_groupi_n_600, csa_tree_add_95_22_pad_groupi_n_601, csa_tree_add_95_22_pad_groupi_n_602, csa_tree_add_95_22_pad_groupi_n_603, csa_tree_add_95_22_pad_groupi_n_604;
  wire csa_tree_add_95_22_pad_groupi_n_605, csa_tree_add_95_22_pad_groupi_n_606, csa_tree_add_95_22_pad_groupi_n_607, csa_tree_add_95_22_pad_groupi_n_608, csa_tree_add_95_22_pad_groupi_n_609, csa_tree_add_95_22_pad_groupi_n_610, csa_tree_add_95_22_pad_groupi_n_611, csa_tree_add_95_22_pad_groupi_n_612;
  wire csa_tree_add_95_22_pad_groupi_n_613, csa_tree_add_95_22_pad_groupi_n_614, csa_tree_add_95_22_pad_groupi_n_615, csa_tree_add_95_22_pad_groupi_n_616, csa_tree_add_95_22_pad_groupi_n_617, csa_tree_add_95_22_pad_groupi_n_618, csa_tree_add_95_22_pad_groupi_n_619, csa_tree_add_95_22_pad_groupi_n_620;
  wire csa_tree_add_95_22_pad_groupi_n_621, csa_tree_add_95_22_pad_groupi_n_622, csa_tree_add_95_22_pad_groupi_n_623, csa_tree_add_95_22_pad_groupi_n_624, csa_tree_add_95_22_pad_groupi_n_625, csa_tree_add_95_22_pad_groupi_n_626, csa_tree_add_95_22_pad_groupi_n_627, csa_tree_add_95_22_pad_groupi_n_628;
  wire csa_tree_add_95_22_pad_groupi_n_629, csa_tree_add_95_22_pad_groupi_n_630, csa_tree_add_95_22_pad_groupi_n_631, csa_tree_add_95_22_pad_groupi_n_633, csa_tree_add_95_22_pad_groupi_n_634, csa_tree_add_95_22_pad_groupi_n_635, csa_tree_add_95_22_pad_groupi_n_637, csa_tree_add_95_22_pad_groupi_n_638;
  wire csa_tree_add_95_22_pad_groupi_n_639, csa_tree_add_95_22_pad_groupi_n_640, csa_tree_add_95_22_pad_groupi_n_641, csa_tree_add_95_22_pad_groupi_n_642, csa_tree_add_95_22_pad_groupi_n_643, csa_tree_add_95_22_pad_groupi_n_644, csa_tree_add_95_22_pad_groupi_n_645, csa_tree_add_95_22_pad_groupi_n_646;
  wire csa_tree_add_95_22_pad_groupi_n_647, csa_tree_add_95_22_pad_groupi_n_648, csa_tree_add_95_22_pad_groupi_n_649, csa_tree_add_95_22_pad_groupi_n_650, csa_tree_add_95_22_pad_groupi_n_651, csa_tree_add_95_22_pad_groupi_n_652, csa_tree_add_95_22_pad_groupi_n_653, csa_tree_add_95_22_pad_groupi_n_654;
  wire csa_tree_add_95_22_pad_groupi_n_655, csa_tree_add_95_22_pad_groupi_n_656, csa_tree_add_95_22_pad_groupi_n_657, csa_tree_add_95_22_pad_groupi_n_658, csa_tree_add_95_22_pad_groupi_n_659, csa_tree_add_95_22_pad_groupi_n_660, csa_tree_add_95_22_pad_groupi_n_661, csa_tree_add_95_22_pad_groupi_n_662;
  wire csa_tree_add_95_22_pad_groupi_n_663, csa_tree_add_95_22_pad_groupi_n_664, csa_tree_add_95_22_pad_groupi_n_665, csa_tree_add_95_22_pad_groupi_n_666, csa_tree_add_95_22_pad_groupi_n_667, csa_tree_add_95_22_pad_groupi_n_668, csa_tree_add_95_22_pad_groupi_n_669, csa_tree_add_95_22_pad_groupi_n_670;
  wire csa_tree_add_95_22_pad_groupi_n_671, csa_tree_add_95_22_pad_groupi_n_672, csa_tree_add_95_22_pad_groupi_n_673, csa_tree_add_95_22_pad_groupi_n_674, csa_tree_add_95_22_pad_groupi_n_675, csa_tree_add_95_22_pad_groupi_n_676, csa_tree_add_95_22_pad_groupi_n_677, csa_tree_add_95_22_pad_groupi_n_678;
  wire csa_tree_add_95_22_pad_groupi_n_679, csa_tree_add_95_22_pad_groupi_n_680, csa_tree_add_95_22_pad_groupi_n_681, csa_tree_add_95_22_pad_groupi_n_682, csa_tree_add_95_22_pad_groupi_n_683, csa_tree_add_95_22_pad_groupi_n_684, csa_tree_add_95_22_pad_groupi_n_685, csa_tree_add_95_22_pad_groupi_n_686;
  wire csa_tree_add_95_22_pad_groupi_n_688, csa_tree_add_95_22_pad_groupi_n_689, csa_tree_add_95_22_pad_groupi_n_690, csa_tree_add_95_22_pad_groupi_n_691, csa_tree_add_95_22_pad_groupi_n_692, csa_tree_add_95_22_pad_groupi_n_693, csa_tree_add_95_22_pad_groupi_n_694, csa_tree_add_95_22_pad_groupi_n_695;
  wire csa_tree_add_95_22_pad_groupi_n_696, csa_tree_add_95_22_pad_groupi_n_697, csa_tree_add_95_22_pad_groupi_n_698, csa_tree_add_95_22_pad_groupi_n_699, csa_tree_add_95_22_pad_groupi_n_700, csa_tree_add_95_22_pad_groupi_n_702, csa_tree_add_95_22_pad_groupi_n_703, csa_tree_add_95_22_pad_groupi_n_704;
  wire csa_tree_add_95_22_pad_groupi_n_705, csa_tree_add_95_22_pad_groupi_n_706, csa_tree_add_95_22_pad_groupi_n_707, csa_tree_add_95_22_pad_groupi_n_708, csa_tree_add_95_22_pad_groupi_n_709, csa_tree_add_95_22_pad_groupi_n_710, csa_tree_add_95_22_pad_groupi_n_711, csa_tree_add_95_22_pad_groupi_n_712;
  wire csa_tree_add_95_22_pad_groupi_n_713, csa_tree_add_95_22_pad_groupi_n_714, csa_tree_add_95_22_pad_groupi_n_715, csa_tree_add_95_22_pad_groupi_n_716, csa_tree_add_95_22_pad_groupi_n_717, csa_tree_add_95_22_pad_groupi_n_718, csa_tree_add_95_22_pad_groupi_n_719, csa_tree_add_95_22_pad_groupi_n_720;
  wire csa_tree_add_95_22_pad_groupi_n_721, csa_tree_add_95_22_pad_groupi_n_722, csa_tree_add_95_22_pad_groupi_n_723, csa_tree_add_95_22_pad_groupi_n_724, csa_tree_add_95_22_pad_groupi_n_725, csa_tree_add_95_22_pad_groupi_n_726, csa_tree_add_95_22_pad_groupi_n_727, csa_tree_add_95_22_pad_groupi_n_728;
  wire csa_tree_add_95_22_pad_groupi_n_729, csa_tree_add_95_22_pad_groupi_n_730, csa_tree_add_95_22_pad_groupi_n_731, csa_tree_add_95_22_pad_groupi_n_732, csa_tree_add_95_22_pad_groupi_n_733, csa_tree_add_95_22_pad_groupi_n_734, csa_tree_add_95_22_pad_groupi_n_735, csa_tree_add_95_22_pad_groupi_n_736;
  wire csa_tree_add_95_22_pad_groupi_n_737, csa_tree_add_95_22_pad_groupi_n_738, csa_tree_add_95_22_pad_groupi_n_739, csa_tree_add_95_22_pad_groupi_n_740, csa_tree_add_95_22_pad_groupi_n_741, csa_tree_add_95_22_pad_groupi_n_742, csa_tree_add_95_22_pad_groupi_n_743, csa_tree_add_95_22_pad_groupi_n_744;
  wire csa_tree_add_95_22_pad_groupi_n_745, csa_tree_add_95_22_pad_groupi_n_746, csa_tree_add_95_22_pad_groupi_n_747, csa_tree_add_95_22_pad_groupi_n_748, csa_tree_add_95_22_pad_groupi_n_749, csa_tree_add_95_22_pad_groupi_n_750, csa_tree_add_95_22_pad_groupi_n_751, csa_tree_add_95_22_pad_groupi_n_752;
  wire csa_tree_add_95_22_pad_groupi_n_753, csa_tree_add_95_22_pad_groupi_n_754, csa_tree_add_95_22_pad_groupi_n_755, csa_tree_add_95_22_pad_groupi_n_756, csa_tree_add_95_22_pad_groupi_n_757, csa_tree_add_95_22_pad_groupi_n_758, csa_tree_add_95_22_pad_groupi_n_759, csa_tree_add_95_22_pad_groupi_n_760;
  wire csa_tree_add_95_22_pad_groupi_n_761, csa_tree_add_95_22_pad_groupi_n_762, csa_tree_add_95_22_pad_groupi_n_763, csa_tree_add_95_22_pad_groupi_n_764, csa_tree_add_95_22_pad_groupi_n_765, csa_tree_add_95_22_pad_groupi_n_766, csa_tree_add_95_22_pad_groupi_n_767, csa_tree_add_95_22_pad_groupi_n_768;
  wire csa_tree_add_95_22_pad_groupi_n_769, csa_tree_add_95_22_pad_groupi_n_770, csa_tree_add_95_22_pad_groupi_n_771, csa_tree_add_95_22_pad_groupi_n_772, csa_tree_add_95_22_pad_groupi_n_773, csa_tree_add_95_22_pad_groupi_n_774, csa_tree_add_95_22_pad_groupi_n_775, csa_tree_add_95_22_pad_groupi_n_776;
  wire csa_tree_add_95_22_pad_groupi_n_777, csa_tree_add_95_22_pad_groupi_n_778, csa_tree_add_95_22_pad_groupi_n_779, csa_tree_add_95_22_pad_groupi_n_780, csa_tree_add_95_22_pad_groupi_n_781, csa_tree_add_95_22_pad_groupi_n_782, csa_tree_add_95_22_pad_groupi_n_783, csa_tree_add_95_22_pad_groupi_n_784;
  wire csa_tree_add_95_22_pad_groupi_n_785, csa_tree_add_95_22_pad_groupi_n_786, csa_tree_add_95_22_pad_groupi_n_787, csa_tree_add_95_22_pad_groupi_n_788, csa_tree_add_95_22_pad_groupi_n_789, csa_tree_add_95_22_pad_groupi_n_790, csa_tree_add_95_22_pad_groupi_n_791, csa_tree_add_95_22_pad_groupi_n_792;
  wire csa_tree_add_95_22_pad_groupi_n_793, csa_tree_add_95_22_pad_groupi_n_794, csa_tree_add_95_22_pad_groupi_n_795, csa_tree_add_95_22_pad_groupi_n_796, csa_tree_add_95_22_pad_groupi_n_797, csa_tree_add_95_22_pad_groupi_n_798, csa_tree_add_95_22_pad_groupi_n_799, csa_tree_add_95_22_pad_groupi_n_800;
  wire csa_tree_add_95_22_pad_groupi_n_801, csa_tree_add_95_22_pad_groupi_n_802, csa_tree_add_95_22_pad_groupi_n_803, csa_tree_add_95_22_pad_groupi_n_804, csa_tree_add_95_22_pad_groupi_n_805, csa_tree_add_95_22_pad_groupi_n_806, csa_tree_add_95_22_pad_groupi_n_807, csa_tree_add_95_22_pad_groupi_n_808;
  wire csa_tree_add_95_22_pad_groupi_n_809, csa_tree_add_95_22_pad_groupi_n_810, csa_tree_add_95_22_pad_groupi_n_811, csa_tree_add_95_22_pad_groupi_n_812, csa_tree_add_95_22_pad_groupi_n_813, csa_tree_add_95_22_pad_groupi_n_814, csa_tree_add_95_22_pad_groupi_n_815, csa_tree_add_95_22_pad_groupi_n_816;
  wire csa_tree_add_95_22_pad_groupi_n_817, csa_tree_add_95_22_pad_groupi_n_818, csa_tree_add_95_22_pad_groupi_n_819, csa_tree_add_95_22_pad_groupi_n_820, csa_tree_add_95_22_pad_groupi_n_821, csa_tree_add_95_22_pad_groupi_n_822, csa_tree_add_95_22_pad_groupi_n_823, csa_tree_add_95_22_pad_groupi_n_824;
  wire csa_tree_add_95_22_pad_groupi_n_825, csa_tree_add_95_22_pad_groupi_n_826, csa_tree_add_95_22_pad_groupi_n_827, csa_tree_add_95_22_pad_groupi_n_828, csa_tree_add_95_22_pad_groupi_n_829, csa_tree_add_95_22_pad_groupi_n_830, csa_tree_add_95_22_pad_groupi_n_831, csa_tree_add_95_22_pad_groupi_n_832;
  wire csa_tree_add_95_22_pad_groupi_n_833, csa_tree_add_95_22_pad_groupi_n_834, csa_tree_add_95_22_pad_groupi_n_835, csa_tree_add_95_22_pad_groupi_n_836, csa_tree_add_95_22_pad_groupi_n_837, csa_tree_add_95_22_pad_groupi_n_838, csa_tree_add_95_22_pad_groupi_n_839, csa_tree_add_95_22_pad_groupi_n_840;
  wire csa_tree_add_95_22_pad_groupi_n_841, csa_tree_add_95_22_pad_groupi_n_842, csa_tree_add_95_22_pad_groupi_n_843, csa_tree_add_95_22_pad_groupi_n_844, csa_tree_add_95_22_pad_groupi_n_845, csa_tree_add_95_22_pad_groupi_n_846, csa_tree_add_95_22_pad_groupi_n_847, csa_tree_add_95_22_pad_groupi_n_848;
  wire csa_tree_add_95_22_pad_groupi_n_849, csa_tree_add_95_22_pad_groupi_n_851, csa_tree_add_95_22_pad_groupi_n_852, csa_tree_add_95_22_pad_groupi_n_853, csa_tree_add_95_22_pad_groupi_n_854, csa_tree_add_95_22_pad_groupi_n_855, csa_tree_add_95_22_pad_groupi_n_856, csa_tree_add_95_22_pad_groupi_n_857;
  wire csa_tree_add_95_22_pad_groupi_n_858, csa_tree_add_95_22_pad_groupi_n_859, csa_tree_add_95_22_pad_groupi_n_860, csa_tree_add_95_22_pad_groupi_n_861, csa_tree_add_95_22_pad_groupi_n_862, csa_tree_add_95_22_pad_groupi_n_863, csa_tree_add_95_22_pad_groupi_n_864, csa_tree_add_95_22_pad_groupi_n_865;
  wire csa_tree_add_95_22_pad_groupi_n_866, csa_tree_add_95_22_pad_groupi_n_867, csa_tree_add_95_22_pad_groupi_n_868, csa_tree_add_95_22_pad_groupi_n_869, csa_tree_add_95_22_pad_groupi_n_870, csa_tree_add_95_22_pad_groupi_n_871, csa_tree_add_95_22_pad_groupi_n_872, csa_tree_add_95_22_pad_groupi_n_873;
  wire csa_tree_add_95_22_pad_groupi_n_874, csa_tree_add_95_22_pad_groupi_n_875, csa_tree_add_95_22_pad_groupi_n_876, csa_tree_add_95_22_pad_groupi_n_877, csa_tree_add_95_22_pad_groupi_n_878, csa_tree_add_95_22_pad_groupi_n_879, csa_tree_add_95_22_pad_groupi_n_880, csa_tree_add_95_22_pad_groupi_n_881;
  wire csa_tree_add_95_22_pad_groupi_n_882, csa_tree_add_95_22_pad_groupi_n_883, csa_tree_add_95_22_pad_groupi_n_884, csa_tree_add_95_22_pad_groupi_n_885, csa_tree_add_95_22_pad_groupi_n_886, csa_tree_add_95_22_pad_groupi_n_887, csa_tree_add_95_22_pad_groupi_n_888, csa_tree_add_95_22_pad_groupi_n_889;
  wire csa_tree_add_95_22_pad_groupi_n_890, csa_tree_add_95_22_pad_groupi_n_891, csa_tree_add_95_22_pad_groupi_n_892, csa_tree_add_95_22_pad_groupi_n_893, csa_tree_add_95_22_pad_groupi_n_894, csa_tree_add_95_22_pad_groupi_n_895, csa_tree_add_95_22_pad_groupi_n_896, csa_tree_add_95_22_pad_groupi_n_897;
  wire csa_tree_add_95_22_pad_groupi_n_898, csa_tree_add_95_22_pad_groupi_n_899, csa_tree_add_95_22_pad_groupi_n_900, csa_tree_add_95_22_pad_groupi_n_901, csa_tree_add_95_22_pad_groupi_n_902, csa_tree_add_95_22_pad_groupi_n_903, csa_tree_add_95_22_pad_groupi_n_904, csa_tree_add_95_22_pad_groupi_n_905;
  wire csa_tree_add_95_22_pad_groupi_n_906, csa_tree_add_95_22_pad_groupi_n_907, csa_tree_add_95_22_pad_groupi_n_908, csa_tree_add_95_22_pad_groupi_n_909, csa_tree_add_95_22_pad_groupi_n_910, csa_tree_add_95_22_pad_groupi_n_911, csa_tree_add_95_22_pad_groupi_n_912, csa_tree_add_95_22_pad_groupi_n_913;
  wire csa_tree_add_95_22_pad_groupi_n_914, csa_tree_add_95_22_pad_groupi_n_915, csa_tree_add_95_22_pad_groupi_n_916, csa_tree_add_95_22_pad_groupi_n_917, csa_tree_add_95_22_pad_groupi_n_918, csa_tree_add_95_22_pad_groupi_n_919, csa_tree_add_95_22_pad_groupi_n_920, csa_tree_add_95_22_pad_groupi_n_921;
  wire csa_tree_add_95_22_pad_groupi_n_922, csa_tree_add_95_22_pad_groupi_n_923, csa_tree_add_95_22_pad_groupi_n_924, csa_tree_add_95_22_pad_groupi_n_925, csa_tree_add_95_22_pad_groupi_n_926, csa_tree_add_95_22_pad_groupi_n_927, csa_tree_add_95_22_pad_groupi_n_928, csa_tree_add_95_22_pad_groupi_n_929;
  wire csa_tree_add_95_22_pad_groupi_n_930, csa_tree_add_95_22_pad_groupi_n_931, csa_tree_add_95_22_pad_groupi_n_932, csa_tree_add_95_22_pad_groupi_n_933, csa_tree_add_95_22_pad_groupi_n_934, csa_tree_add_95_22_pad_groupi_n_935, csa_tree_add_95_22_pad_groupi_n_936, csa_tree_add_95_22_pad_groupi_n_937;
  wire csa_tree_add_95_22_pad_groupi_n_938, csa_tree_add_95_22_pad_groupi_n_939, csa_tree_add_95_22_pad_groupi_n_940, csa_tree_add_95_22_pad_groupi_n_941, csa_tree_add_95_22_pad_groupi_n_942, csa_tree_add_95_22_pad_groupi_n_943, csa_tree_add_95_22_pad_groupi_n_944, csa_tree_add_95_22_pad_groupi_n_945;
  wire csa_tree_add_95_22_pad_groupi_n_946, csa_tree_add_95_22_pad_groupi_n_947, csa_tree_add_95_22_pad_groupi_n_948, csa_tree_add_95_22_pad_groupi_n_949, csa_tree_add_95_22_pad_groupi_n_950, csa_tree_add_95_22_pad_groupi_n_951, csa_tree_add_95_22_pad_groupi_n_952, csa_tree_add_95_22_pad_groupi_n_953;
  wire csa_tree_add_95_22_pad_groupi_n_954, csa_tree_add_95_22_pad_groupi_n_955, csa_tree_add_95_22_pad_groupi_n_956, csa_tree_add_95_22_pad_groupi_n_957, csa_tree_add_95_22_pad_groupi_n_958, csa_tree_add_95_22_pad_groupi_n_959, csa_tree_add_95_22_pad_groupi_n_960, csa_tree_add_95_22_pad_groupi_n_961;
  wire csa_tree_add_95_22_pad_groupi_n_962, csa_tree_add_95_22_pad_groupi_n_963, csa_tree_add_95_22_pad_groupi_n_964, csa_tree_add_95_22_pad_groupi_n_965, csa_tree_add_95_22_pad_groupi_n_966, csa_tree_add_95_22_pad_groupi_n_967, csa_tree_add_95_22_pad_groupi_n_968, csa_tree_add_95_22_pad_groupi_n_969;
  wire csa_tree_add_95_22_pad_groupi_n_970, csa_tree_add_95_22_pad_groupi_n_971, csa_tree_add_95_22_pad_groupi_n_972, csa_tree_add_95_22_pad_groupi_n_973, csa_tree_add_95_22_pad_groupi_n_974, csa_tree_add_95_22_pad_groupi_n_975, csa_tree_add_95_22_pad_groupi_n_976, csa_tree_add_95_22_pad_groupi_n_977;
  wire csa_tree_add_95_22_pad_groupi_n_978, csa_tree_add_95_22_pad_groupi_n_979, csa_tree_add_95_22_pad_groupi_n_980, csa_tree_add_95_22_pad_groupi_n_981, csa_tree_add_95_22_pad_groupi_n_982, csa_tree_add_95_22_pad_groupi_n_983, csa_tree_add_95_22_pad_groupi_n_984, csa_tree_add_95_22_pad_groupi_n_985;
  wire csa_tree_add_95_22_pad_groupi_n_986, csa_tree_add_95_22_pad_groupi_n_987, csa_tree_add_95_22_pad_groupi_n_988, csa_tree_add_95_22_pad_groupi_n_989, csa_tree_add_95_22_pad_groupi_n_990, csa_tree_add_95_22_pad_groupi_n_991, csa_tree_add_95_22_pad_groupi_n_992, csa_tree_add_95_22_pad_groupi_n_993;
  wire csa_tree_add_95_22_pad_groupi_n_994, csa_tree_add_95_22_pad_groupi_n_995, csa_tree_add_95_22_pad_groupi_n_996, csa_tree_add_95_22_pad_groupi_n_997, csa_tree_add_95_22_pad_groupi_n_998, csa_tree_add_95_22_pad_groupi_n_999, csa_tree_add_95_22_pad_groupi_n_1000, csa_tree_add_95_22_pad_groupi_n_1001;
  wire csa_tree_add_95_22_pad_groupi_n_1002, csa_tree_add_95_22_pad_groupi_n_1003, csa_tree_add_95_22_pad_groupi_n_1004, csa_tree_add_95_22_pad_groupi_n_1005, csa_tree_add_95_22_pad_groupi_n_1006, csa_tree_add_95_22_pad_groupi_n_1007, csa_tree_add_95_22_pad_groupi_n_1008, csa_tree_add_95_22_pad_groupi_n_1009;
  wire csa_tree_add_95_22_pad_groupi_n_1010, csa_tree_add_95_22_pad_groupi_n_1011, csa_tree_add_95_22_pad_groupi_n_1012, csa_tree_add_95_22_pad_groupi_n_1013, csa_tree_add_95_22_pad_groupi_n_1014, csa_tree_add_95_22_pad_groupi_n_1015, csa_tree_add_95_22_pad_groupi_n_1016, csa_tree_add_95_22_pad_groupi_n_1017;
  wire csa_tree_add_95_22_pad_groupi_n_1018, csa_tree_add_95_22_pad_groupi_n_1019, csa_tree_add_95_22_pad_groupi_n_1020, csa_tree_add_95_22_pad_groupi_n_1021, csa_tree_add_95_22_pad_groupi_n_1022, csa_tree_add_95_22_pad_groupi_n_1023, csa_tree_add_95_22_pad_groupi_n_1024, csa_tree_add_95_22_pad_groupi_n_1025;
  wire csa_tree_add_95_22_pad_groupi_n_1026, csa_tree_add_95_22_pad_groupi_n_1027, csa_tree_add_95_22_pad_groupi_n_1028, csa_tree_add_95_22_pad_groupi_n_1029, csa_tree_add_95_22_pad_groupi_n_1030, csa_tree_add_95_22_pad_groupi_n_1031, csa_tree_add_95_22_pad_groupi_n_1032, csa_tree_add_95_22_pad_groupi_n_1033;
  wire csa_tree_add_95_22_pad_groupi_n_1034, csa_tree_add_95_22_pad_groupi_n_1035, csa_tree_add_95_22_pad_groupi_n_1036, csa_tree_add_95_22_pad_groupi_n_1037, csa_tree_add_95_22_pad_groupi_n_1038, csa_tree_add_95_22_pad_groupi_n_1039, csa_tree_add_95_22_pad_groupi_n_1040, csa_tree_add_95_22_pad_groupi_n_1041;
  wire csa_tree_add_95_22_pad_groupi_n_1042, csa_tree_add_95_22_pad_groupi_n_1043, csa_tree_add_95_22_pad_groupi_n_1044, csa_tree_add_95_22_pad_groupi_n_1045, csa_tree_add_95_22_pad_groupi_n_1046, csa_tree_add_95_22_pad_groupi_n_1047, csa_tree_add_95_22_pad_groupi_n_1048, csa_tree_add_95_22_pad_groupi_n_1049;
  wire csa_tree_add_95_22_pad_groupi_n_1050, csa_tree_add_95_22_pad_groupi_n_1051, csa_tree_add_95_22_pad_groupi_n_1052, csa_tree_add_95_22_pad_groupi_n_1053, csa_tree_add_95_22_pad_groupi_n_1054, csa_tree_add_95_22_pad_groupi_n_1055, csa_tree_add_95_22_pad_groupi_n_1056, csa_tree_add_95_22_pad_groupi_n_1057;
  wire csa_tree_add_95_22_pad_groupi_n_1058, csa_tree_add_95_22_pad_groupi_n_1059, csa_tree_add_95_22_pad_groupi_n_1060, csa_tree_add_95_22_pad_groupi_n_1061, csa_tree_add_95_22_pad_groupi_n_1062, csa_tree_add_95_22_pad_groupi_n_1063, csa_tree_add_95_22_pad_groupi_n_1064, csa_tree_add_95_22_pad_groupi_n_1065;
  wire csa_tree_add_95_22_pad_groupi_n_1066, csa_tree_add_95_22_pad_groupi_n_1067, csa_tree_add_95_22_pad_groupi_n_1068, csa_tree_add_95_22_pad_groupi_n_1069, csa_tree_add_95_22_pad_groupi_n_1070, csa_tree_add_95_22_pad_groupi_n_1071, csa_tree_add_95_22_pad_groupi_n_1072, csa_tree_add_95_22_pad_groupi_n_1073;
  wire csa_tree_add_95_22_pad_groupi_n_1074, csa_tree_add_95_22_pad_groupi_n_1075, csa_tree_add_95_22_pad_groupi_n_1076, csa_tree_add_95_22_pad_groupi_n_1077, csa_tree_add_95_22_pad_groupi_n_1078, csa_tree_add_95_22_pad_groupi_n_1079, csa_tree_add_95_22_pad_groupi_n_1080, csa_tree_add_95_22_pad_groupi_n_1081;
  wire csa_tree_add_95_22_pad_groupi_n_1082, csa_tree_add_95_22_pad_groupi_n_1083, csa_tree_add_95_22_pad_groupi_n_1084, csa_tree_add_95_22_pad_groupi_n_1085, csa_tree_add_95_22_pad_groupi_n_1086, csa_tree_add_95_22_pad_groupi_n_1087, csa_tree_add_95_22_pad_groupi_n_1088, csa_tree_add_95_22_pad_groupi_n_1089;
  wire csa_tree_add_95_22_pad_groupi_n_1090, csa_tree_add_95_22_pad_groupi_n_1091, csa_tree_add_95_22_pad_groupi_n_1092, csa_tree_add_95_22_pad_groupi_n_1093, csa_tree_add_95_22_pad_groupi_n_1094, csa_tree_add_95_22_pad_groupi_n_1095, csa_tree_add_95_22_pad_groupi_n_1096, csa_tree_add_95_22_pad_groupi_n_1097;
  wire csa_tree_add_95_22_pad_groupi_n_1098, csa_tree_add_95_22_pad_groupi_n_1099, csa_tree_add_95_22_pad_groupi_n_1100, csa_tree_add_95_22_pad_groupi_n_1101, csa_tree_add_95_22_pad_groupi_n_1102, csa_tree_add_95_22_pad_groupi_n_1103, csa_tree_add_95_22_pad_groupi_n_1104, csa_tree_add_95_22_pad_groupi_n_1105;
  wire csa_tree_add_95_22_pad_groupi_n_1106, csa_tree_add_95_22_pad_groupi_n_1107, csa_tree_add_95_22_pad_groupi_n_1108, csa_tree_add_95_22_pad_groupi_n_1109, csa_tree_add_95_22_pad_groupi_n_1110, csa_tree_add_95_22_pad_groupi_n_1111, csa_tree_add_95_22_pad_groupi_n_1112, csa_tree_add_95_22_pad_groupi_n_1113;
  wire csa_tree_add_95_22_pad_groupi_n_1114, csa_tree_add_95_22_pad_groupi_n_1115, csa_tree_add_95_22_pad_groupi_n_1116, csa_tree_add_95_22_pad_groupi_n_1117, csa_tree_add_95_22_pad_groupi_n_1118, csa_tree_add_95_22_pad_groupi_n_1119, csa_tree_add_95_22_pad_groupi_n_1120, csa_tree_add_95_22_pad_groupi_n_1121;
  wire csa_tree_add_95_22_pad_groupi_n_1122, csa_tree_add_95_22_pad_groupi_n_1123, csa_tree_add_95_22_pad_groupi_n_1124, csa_tree_add_95_22_pad_groupi_n_1125, csa_tree_add_95_22_pad_groupi_n_1126, csa_tree_add_95_22_pad_groupi_n_1127, csa_tree_add_95_22_pad_groupi_n_1128, csa_tree_add_95_22_pad_groupi_n_1129;
  wire csa_tree_add_95_22_pad_groupi_n_1130, csa_tree_add_95_22_pad_groupi_n_1131, csa_tree_add_95_22_pad_groupi_n_1132, csa_tree_add_95_22_pad_groupi_n_1133, csa_tree_add_95_22_pad_groupi_n_1134, csa_tree_add_95_22_pad_groupi_n_1135, csa_tree_add_95_22_pad_groupi_n_1136, csa_tree_add_95_22_pad_groupi_n_1137;
  wire csa_tree_add_95_22_pad_groupi_n_1138, csa_tree_add_95_22_pad_groupi_n_1139, csa_tree_add_95_22_pad_groupi_n_1140, csa_tree_add_95_22_pad_groupi_n_1141, csa_tree_add_95_22_pad_groupi_n_1142, csa_tree_add_95_22_pad_groupi_n_1143, csa_tree_add_95_22_pad_groupi_n_1144, csa_tree_add_95_22_pad_groupi_n_1145;
  wire csa_tree_add_95_22_pad_groupi_n_1146, csa_tree_add_95_22_pad_groupi_n_1147, csa_tree_add_95_22_pad_groupi_n_1148, csa_tree_add_95_22_pad_groupi_n_1149, csa_tree_add_95_22_pad_groupi_n_1150, csa_tree_add_95_22_pad_groupi_n_1151, csa_tree_add_95_22_pad_groupi_n_1152, csa_tree_add_95_22_pad_groupi_n_1153;
  wire csa_tree_add_95_22_pad_groupi_n_1154, csa_tree_add_95_22_pad_groupi_n_1155, csa_tree_add_95_22_pad_groupi_n_1156, csa_tree_add_95_22_pad_groupi_n_1157, csa_tree_add_95_22_pad_groupi_n_1158, csa_tree_add_95_22_pad_groupi_n_1159, csa_tree_add_95_22_pad_groupi_n_1160, csa_tree_add_95_22_pad_groupi_n_1161;
  wire csa_tree_add_95_22_pad_groupi_n_1162, csa_tree_add_95_22_pad_groupi_n_1163, csa_tree_add_95_22_pad_groupi_n_1164, csa_tree_add_95_22_pad_groupi_n_1165, csa_tree_add_95_22_pad_groupi_n_1166, csa_tree_add_95_22_pad_groupi_n_1167, csa_tree_add_95_22_pad_groupi_n_1168, csa_tree_add_95_22_pad_groupi_n_1169;
  wire csa_tree_add_95_22_pad_groupi_n_1170, csa_tree_add_95_22_pad_groupi_n_1171, csa_tree_add_95_22_pad_groupi_n_1172, csa_tree_add_95_22_pad_groupi_n_1173, csa_tree_add_95_22_pad_groupi_n_1174, csa_tree_add_95_22_pad_groupi_n_1175, csa_tree_add_95_22_pad_groupi_n_1176, csa_tree_add_95_22_pad_groupi_n_1177;
  wire csa_tree_add_95_22_pad_groupi_n_1178, csa_tree_add_95_22_pad_groupi_n_1179, csa_tree_add_95_22_pad_groupi_n_1180, csa_tree_add_95_22_pad_groupi_n_1181, csa_tree_add_95_22_pad_groupi_n_1182, csa_tree_add_95_22_pad_groupi_n_1183, csa_tree_add_95_22_pad_groupi_n_1184, csa_tree_add_95_22_pad_groupi_n_1185;
  wire csa_tree_add_95_22_pad_groupi_n_1186, csa_tree_add_95_22_pad_groupi_n_1187, csa_tree_add_95_22_pad_groupi_n_1188, csa_tree_add_95_22_pad_groupi_n_1189, csa_tree_add_95_22_pad_groupi_n_1190, csa_tree_add_95_22_pad_groupi_n_1191, csa_tree_add_95_22_pad_groupi_n_1192, csa_tree_add_95_22_pad_groupi_n_1193;
  wire csa_tree_add_95_22_pad_groupi_n_1194, csa_tree_add_95_22_pad_groupi_n_1195, csa_tree_add_95_22_pad_groupi_n_1196, csa_tree_add_95_22_pad_groupi_n_1197, csa_tree_add_95_22_pad_groupi_n_1198, csa_tree_add_95_22_pad_groupi_n_1199, csa_tree_add_95_22_pad_groupi_n_1200, csa_tree_add_95_22_pad_groupi_n_1201;
  wire csa_tree_add_95_22_pad_groupi_n_1202, csa_tree_add_95_22_pad_groupi_n_1203, csa_tree_add_95_22_pad_groupi_n_1204, csa_tree_add_95_22_pad_groupi_n_1205, csa_tree_add_95_22_pad_groupi_n_1206, csa_tree_add_95_22_pad_groupi_n_1207, csa_tree_add_95_22_pad_groupi_n_1208, csa_tree_add_95_22_pad_groupi_n_1209;
  wire csa_tree_add_95_22_pad_groupi_n_1210, csa_tree_add_95_22_pad_groupi_n_1211, csa_tree_add_95_22_pad_groupi_n_1212, csa_tree_add_95_22_pad_groupi_n_1213, csa_tree_add_95_22_pad_groupi_n_1214, csa_tree_add_95_22_pad_groupi_n_1215, csa_tree_add_95_22_pad_groupi_n_1216, csa_tree_add_95_22_pad_groupi_n_1217;
  wire csa_tree_add_95_22_pad_groupi_n_1218, csa_tree_add_95_22_pad_groupi_n_1219, csa_tree_add_95_22_pad_groupi_n_1220, csa_tree_add_95_22_pad_groupi_n_1221, csa_tree_add_95_22_pad_groupi_n_1222, csa_tree_add_95_22_pad_groupi_n_1223, csa_tree_add_95_22_pad_groupi_n_1224, csa_tree_add_95_22_pad_groupi_n_1225;
  wire csa_tree_add_95_22_pad_groupi_n_1226, csa_tree_add_95_22_pad_groupi_n_1227, csa_tree_add_95_22_pad_groupi_n_1228, csa_tree_add_95_22_pad_groupi_n_1229, csa_tree_add_95_22_pad_groupi_n_1230, csa_tree_add_95_22_pad_groupi_n_1231, csa_tree_add_95_22_pad_groupi_n_1232, csa_tree_add_95_22_pad_groupi_n_1233;
  wire csa_tree_add_95_22_pad_groupi_n_1234, csa_tree_add_95_22_pad_groupi_n_1235, csa_tree_add_95_22_pad_groupi_n_1236, csa_tree_add_95_22_pad_groupi_n_1237, csa_tree_add_95_22_pad_groupi_n_1238, csa_tree_add_95_22_pad_groupi_n_1239, csa_tree_add_95_22_pad_groupi_n_1240, csa_tree_add_95_22_pad_groupi_n_1241;
  wire csa_tree_add_95_22_pad_groupi_n_1242, csa_tree_add_95_22_pad_groupi_n_1243, csa_tree_add_95_22_pad_groupi_n_1244, csa_tree_add_95_22_pad_groupi_n_1245, csa_tree_add_95_22_pad_groupi_n_1246, csa_tree_add_95_22_pad_groupi_n_1247, csa_tree_add_95_22_pad_groupi_n_1248, csa_tree_add_95_22_pad_groupi_n_1249;
  wire csa_tree_add_95_22_pad_groupi_n_1250, csa_tree_add_95_22_pad_groupi_n_1251, csa_tree_add_95_22_pad_groupi_n_1252, csa_tree_add_95_22_pad_groupi_n_1253, csa_tree_add_95_22_pad_groupi_n_1254, csa_tree_add_95_22_pad_groupi_n_1255, csa_tree_add_95_22_pad_groupi_n_1256, csa_tree_add_95_22_pad_groupi_n_1257;
  wire csa_tree_add_95_22_pad_groupi_n_1258, csa_tree_add_95_22_pad_groupi_n_1259, csa_tree_add_95_22_pad_groupi_n_1260, csa_tree_add_95_22_pad_groupi_n_1261, csa_tree_add_95_22_pad_groupi_n_1262, csa_tree_add_95_22_pad_groupi_n_1263, csa_tree_add_95_22_pad_groupi_n_1264, csa_tree_add_95_22_pad_groupi_n_1265;
  wire csa_tree_add_95_22_pad_groupi_n_1266, csa_tree_add_95_22_pad_groupi_n_1267, csa_tree_add_95_22_pad_groupi_n_1268, csa_tree_add_95_22_pad_groupi_n_1269, csa_tree_add_95_22_pad_groupi_n_1270, csa_tree_add_95_22_pad_groupi_n_1271, csa_tree_add_95_22_pad_groupi_n_1272, csa_tree_add_95_22_pad_groupi_n_1273;
  wire csa_tree_add_95_22_pad_groupi_n_1274, csa_tree_add_95_22_pad_groupi_n_1275, csa_tree_add_95_22_pad_groupi_n_1276, csa_tree_add_95_22_pad_groupi_n_1277, csa_tree_add_95_22_pad_groupi_n_1278, csa_tree_add_95_22_pad_groupi_n_1279, csa_tree_add_95_22_pad_groupi_n_1280, csa_tree_add_95_22_pad_groupi_n_1281;
  wire csa_tree_add_95_22_pad_groupi_n_1282, csa_tree_add_95_22_pad_groupi_n_1283, csa_tree_add_95_22_pad_groupi_n_1284, csa_tree_add_95_22_pad_groupi_n_1285, csa_tree_add_95_22_pad_groupi_n_1286, csa_tree_add_95_22_pad_groupi_n_1287, csa_tree_add_95_22_pad_groupi_n_1288, csa_tree_add_95_22_pad_groupi_n_1289;
  wire csa_tree_add_95_22_pad_groupi_n_1290, csa_tree_add_95_22_pad_groupi_n_1291, csa_tree_add_95_22_pad_groupi_n_1292, csa_tree_add_95_22_pad_groupi_n_1293, csa_tree_add_95_22_pad_groupi_n_1294, csa_tree_add_95_22_pad_groupi_n_1295, csa_tree_add_95_22_pad_groupi_n_1296, csa_tree_add_95_22_pad_groupi_n_1297;
  wire csa_tree_add_95_22_pad_groupi_n_1298, csa_tree_add_95_22_pad_groupi_n_1299, csa_tree_add_95_22_pad_groupi_n_1300, csa_tree_add_95_22_pad_groupi_n_1301, csa_tree_add_95_22_pad_groupi_n_1302, csa_tree_add_95_22_pad_groupi_n_1303, csa_tree_add_95_22_pad_groupi_n_1304, csa_tree_add_95_22_pad_groupi_n_1305;
  wire csa_tree_add_95_22_pad_groupi_n_1306, csa_tree_add_95_22_pad_groupi_n_1307, csa_tree_add_95_22_pad_groupi_n_1308, csa_tree_add_95_22_pad_groupi_n_1309, csa_tree_add_95_22_pad_groupi_n_1310, csa_tree_add_95_22_pad_groupi_n_1311, csa_tree_add_95_22_pad_groupi_n_1312, csa_tree_add_95_22_pad_groupi_n_1313;
  wire csa_tree_add_95_22_pad_groupi_n_1314, csa_tree_add_95_22_pad_groupi_n_1315, csa_tree_add_95_22_pad_groupi_n_1316, csa_tree_add_95_22_pad_groupi_n_1317, csa_tree_add_95_22_pad_groupi_n_1318, csa_tree_add_95_22_pad_groupi_n_1319, csa_tree_add_95_22_pad_groupi_n_1320, csa_tree_add_95_22_pad_groupi_n_1321;
  wire csa_tree_add_95_22_pad_groupi_n_1322, csa_tree_add_95_22_pad_groupi_n_1323, csa_tree_add_95_22_pad_groupi_n_1324, csa_tree_add_95_22_pad_groupi_n_1325, csa_tree_add_95_22_pad_groupi_n_1326, csa_tree_add_95_22_pad_groupi_n_1327, csa_tree_add_95_22_pad_groupi_n_1328, csa_tree_add_95_22_pad_groupi_n_1329;
  wire csa_tree_add_95_22_pad_groupi_n_1330, csa_tree_add_95_22_pad_groupi_n_1331, csa_tree_add_95_22_pad_groupi_n_1332, csa_tree_add_95_22_pad_groupi_n_1333, csa_tree_add_95_22_pad_groupi_n_1334, csa_tree_add_95_22_pad_groupi_n_1335, csa_tree_add_95_22_pad_groupi_n_1336, csa_tree_add_95_22_pad_groupi_n_1337;
  wire csa_tree_add_95_22_pad_groupi_n_1338, csa_tree_add_95_22_pad_groupi_n_1339, csa_tree_add_95_22_pad_groupi_n_1340, csa_tree_add_95_22_pad_groupi_n_1341, csa_tree_add_95_22_pad_groupi_n_1342, csa_tree_add_95_22_pad_groupi_n_1343, csa_tree_add_95_22_pad_groupi_n_1344, csa_tree_add_95_22_pad_groupi_n_1345;
  wire csa_tree_add_95_22_pad_groupi_n_1346, csa_tree_add_95_22_pad_groupi_n_1347, csa_tree_add_95_22_pad_groupi_n_1348, csa_tree_add_95_22_pad_groupi_n_1349, csa_tree_add_95_22_pad_groupi_n_1350, csa_tree_add_95_22_pad_groupi_n_1351, csa_tree_add_95_22_pad_groupi_n_1352, csa_tree_add_95_22_pad_groupi_n_1353;
  wire csa_tree_add_95_22_pad_groupi_n_1354, csa_tree_add_95_22_pad_groupi_n_1355, csa_tree_add_95_22_pad_groupi_n_1356, csa_tree_add_95_22_pad_groupi_n_1357, csa_tree_add_95_22_pad_groupi_n_1358, csa_tree_add_95_22_pad_groupi_n_1359, csa_tree_add_95_22_pad_groupi_n_1360, csa_tree_add_95_22_pad_groupi_n_1361;
  wire csa_tree_add_95_22_pad_groupi_n_1362, csa_tree_add_95_22_pad_groupi_n_1363, csa_tree_add_95_22_pad_groupi_n_1364, csa_tree_add_95_22_pad_groupi_n_1365, csa_tree_add_95_22_pad_groupi_n_1366, csa_tree_add_95_22_pad_groupi_n_1367, csa_tree_add_95_22_pad_groupi_n_1368, csa_tree_add_95_22_pad_groupi_n_1369;
  wire csa_tree_add_95_22_pad_groupi_n_1370, csa_tree_add_95_22_pad_groupi_n_1371, csa_tree_add_95_22_pad_groupi_n_1372, csa_tree_add_95_22_pad_groupi_n_1373, csa_tree_add_95_22_pad_groupi_n_1374, csa_tree_add_95_22_pad_groupi_n_1375, csa_tree_add_95_22_pad_groupi_n_1376, csa_tree_add_95_22_pad_groupi_n_1377;
  wire csa_tree_add_95_22_pad_groupi_n_1378, csa_tree_add_95_22_pad_groupi_n_1379, csa_tree_add_95_22_pad_groupi_n_1380, csa_tree_add_95_22_pad_groupi_n_1381, csa_tree_add_95_22_pad_groupi_n_1382, csa_tree_add_95_22_pad_groupi_n_1383, csa_tree_add_95_22_pad_groupi_n_1384, csa_tree_add_95_22_pad_groupi_n_1385;
  wire csa_tree_add_95_22_pad_groupi_n_1386, csa_tree_add_95_22_pad_groupi_n_1387, csa_tree_add_95_22_pad_groupi_n_1388, csa_tree_add_95_22_pad_groupi_n_1389, csa_tree_add_95_22_pad_groupi_n_1390, csa_tree_add_95_22_pad_groupi_n_1391, csa_tree_add_95_22_pad_groupi_n_1392, csa_tree_add_95_22_pad_groupi_n_1393;
  wire csa_tree_add_95_22_pad_groupi_n_1394, csa_tree_add_95_22_pad_groupi_n_1395, csa_tree_add_95_22_pad_groupi_n_1396, csa_tree_add_95_22_pad_groupi_n_1397, csa_tree_add_95_22_pad_groupi_n_1398, csa_tree_add_95_22_pad_groupi_n_1399, csa_tree_add_95_22_pad_groupi_n_1400, csa_tree_add_95_22_pad_groupi_n_1401;
  wire csa_tree_add_95_22_pad_groupi_n_1402, csa_tree_add_95_22_pad_groupi_n_1403, csa_tree_add_95_22_pad_groupi_n_1404, csa_tree_add_95_22_pad_groupi_n_1405, csa_tree_add_95_22_pad_groupi_n_1406, csa_tree_add_95_22_pad_groupi_n_1407, csa_tree_add_95_22_pad_groupi_n_1408, csa_tree_add_95_22_pad_groupi_n_1409;
  wire csa_tree_add_95_22_pad_groupi_n_1410, csa_tree_add_95_22_pad_groupi_n_1411, csa_tree_add_95_22_pad_groupi_n_1412, csa_tree_add_95_22_pad_groupi_n_1413, csa_tree_add_95_22_pad_groupi_n_1414, csa_tree_add_95_22_pad_groupi_n_1415, csa_tree_add_95_22_pad_groupi_n_1416, csa_tree_add_95_22_pad_groupi_n_1417;
  wire csa_tree_add_95_22_pad_groupi_n_1418, csa_tree_add_95_22_pad_groupi_n_1419, csa_tree_add_95_22_pad_groupi_n_1420, csa_tree_add_95_22_pad_groupi_n_1421, csa_tree_add_95_22_pad_groupi_n_1422, csa_tree_add_95_22_pad_groupi_n_1423, csa_tree_add_95_22_pad_groupi_n_1424, csa_tree_add_95_22_pad_groupi_n_1425;
  wire csa_tree_add_95_22_pad_groupi_n_1426, csa_tree_add_95_22_pad_groupi_n_1427, csa_tree_add_95_22_pad_groupi_n_1428, csa_tree_add_95_22_pad_groupi_n_1429, csa_tree_add_95_22_pad_groupi_n_1430, csa_tree_add_95_22_pad_groupi_n_1431, csa_tree_add_95_22_pad_groupi_n_1432, csa_tree_add_95_22_pad_groupi_n_1433;
  wire csa_tree_add_95_22_pad_groupi_n_1434, csa_tree_add_95_22_pad_groupi_n_1435, csa_tree_add_95_22_pad_groupi_n_1436, csa_tree_add_95_22_pad_groupi_n_1437, csa_tree_add_95_22_pad_groupi_n_1438, csa_tree_add_95_22_pad_groupi_n_1439, csa_tree_add_95_22_pad_groupi_n_1440, csa_tree_add_95_22_pad_groupi_n_1441;
  wire csa_tree_add_95_22_pad_groupi_n_1442, csa_tree_add_95_22_pad_groupi_n_1443, csa_tree_add_95_22_pad_groupi_n_1444, csa_tree_add_95_22_pad_groupi_n_1445, csa_tree_add_95_22_pad_groupi_n_1446, csa_tree_add_95_22_pad_groupi_n_1447, csa_tree_add_95_22_pad_groupi_n_1448, csa_tree_add_95_22_pad_groupi_n_1449;
  wire csa_tree_add_95_22_pad_groupi_n_1450, csa_tree_add_95_22_pad_groupi_n_1451, csa_tree_add_95_22_pad_groupi_n_1452, csa_tree_add_95_22_pad_groupi_n_1453, csa_tree_add_95_22_pad_groupi_n_1454, csa_tree_add_95_22_pad_groupi_n_1455, csa_tree_add_95_22_pad_groupi_n_1456, csa_tree_add_95_22_pad_groupi_n_1457;
  wire csa_tree_add_95_22_pad_groupi_n_1458, csa_tree_add_95_22_pad_groupi_n_1459, csa_tree_add_95_22_pad_groupi_n_1460, csa_tree_add_95_22_pad_groupi_n_1461, csa_tree_add_95_22_pad_groupi_n_1462, csa_tree_add_95_22_pad_groupi_n_1463, csa_tree_add_95_22_pad_groupi_n_1464, csa_tree_add_95_22_pad_groupi_n_1465;
  wire csa_tree_add_95_22_pad_groupi_n_1466, csa_tree_add_95_22_pad_groupi_n_1467, csa_tree_add_95_22_pad_groupi_n_1468, csa_tree_add_95_22_pad_groupi_n_1469, csa_tree_add_95_22_pad_groupi_n_1470, csa_tree_add_95_22_pad_groupi_n_1471, csa_tree_add_95_22_pad_groupi_n_1472, csa_tree_add_95_22_pad_groupi_n_1473;
  wire csa_tree_add_95_22_pad_groupi_n_1474, csa_tree_add_95_22_pad_groupi_n_1475, csa_tree_add_95_22_pad_groupi_n_1476, csa_tree_add_95_22_pad_groupi_n_1477, csa_tree_add_95_22_pad_groupi_n_1478, csa_tree_add_95_22_pad_groupi_n_1479, csa_tree_add_95_22_pad_groupi_n_1480, csa_tree_add_95_22_pad_groupi_n_1481;
  wire csa_tree_add_95_22_pad_groupi_n_1482, csa_tree_add_95_22_pad_groupi_n_1483, csa_tree_add_95_22_pad_groupi_n_1484, csa_tree_add_95_22_pad_groupi_n_1485, csa_tree_add_95_22_pad_groupi_n_1486, csa_tree_add_95_22_pad_groupi_n_1487, csa_tree_add_95_22_pad_groupi_n_1488, csa_tree_add_95_22_pad_groupi_n_1489;
  wire csa_tree_add_95_22_pad_groupi_n_1490, csa_tree_add_95_22_pad_groupi_n_1491, csa_tree_add_95_22_pad_groupi_n_1492, csa_tree_add_95_22_pad_groupi_n_1493, csa_tree_add_95_22_pad_groupi_n_1494, csa_tree_add_95_22_pad_groupi_n_1495, csa_tree_add_95_22_pad_groupi_n_1496, csa_tree_add_95_22_pad_groupi_n_1497;
  wire csa_tree_add_95_22_pad_groupi_n_1498, csa_tree_add_95_22_pad_groupi_n_1499, csa_tree_add_95_22_pad_groupi_n_1500, csa_tree_add_95_22_pad_groupi_n_1501, csa_tree_add_95_22_pad_groupi_n_1502, csa_tree_add_95_22_pad_groupi_n_1503, csa_tree_add_95_22_pad_groupi_n_1505, csa_tree_add_95_22_pad_groupi_n_1506;
  wire csa_tree_add_95_22_pad_groupi_n_1507, csa_tree_add_95_22_pad_groupi_n_1508, csa_tree_add_95_22_pad_groupi_n_1509, csa_tree_add_95_22_pad_groupi_n_1510, csa_tree_add_95_22_pad_groupi_n_1511, csa_tree_add_95_22_pad_groupi_n_1512, csa_tree_add_95_22_pad_groupi_n_1513, csa_tree_add_95_22_pad_groupi_n_1514;
  wire csa_tree_add_95_22_pad_groupi_n_1515, csa_tree_add_95_22_pad_groupi_n_1516, csa_tree_add_95_22_pad_groupi_n_1517, csa_tree_add_95_22_pad_groupi_n_1518, csa_tree_add_95_22_pad_groupi_n_1519, csa_tree_add_95_22_pad_groupi_n_1520, csa_tree_add_95_22_pad_groupi_n_1521, csa_tree_add_95_22_pad_groupi_n_1522;
  wire csa_tree_add_95_22_pad_groupi_n_1523, csa_tree_add_95_22_pad_groupi_n_1524, csa_tree_add_95_22_pad_groupi_n_1525, csa_tree_add_95_22_pad_groupi_n_1526, csa_tree_add_95_22_pad_groupi_n_1527, csa_tree_add_95_22_pad_groupi_n_1529, csa_tree_add_95_22_pad_groupi_n_1530, csa_tree_add_95_22_pad_groupi_n_1532;
  wire csa_tree_add_95_22_pad_groupi_n_1533, csa_tree_add_95_22_pad_groupi_n_1534, csa_tree_add_95_22_pad_groupi_n_1535, csa_tree_add_95_22_pad_groupi_n_1537, csa_tree_add_95_22_pad_groupi_n_1538, csa_tree_add_95_22_pad_groupi_n_1539, csa_tree_add_95_22_pad_groupi_n_1540, csa_tree_add_95_22_pad_groupi_n_1542;
  wire csa_tree_add_95_22_pad_groupi_n_1543, csa_tree_add_95_22_pad_groupi_n_1544, csa_tree_add_95_22_pad_groupi_n_1546, csa_tree_add_95_22_pad_groupi_n_1547, csa_tree_add_95_22_pad_groupi_n_1549, csa_tree_add_95_22_pad_groupi_n_1550, csa_tree_add_95_22_pad_groupi_n_1552, csa_tree_add_95_22_pad_groupi_n_1553;
  wire csa_tree_add_95_22_pad_groupi_n_1555, csa_tree_add_95_22_pad_groupi_n_1556, csa_tree_add_95_22_pad_groupi_n_1558, csa_tree_add_101_22_pad_groupi_n_0, csa_tree_add_101_22_pad_groupi_n_1, csa_tree_add_101_22_pad_groupi_n_3, csa_tree_add_101_22_pad_groupi_n_4, csa_tree_add_101_22_pad_groupi_n_5;
  wire csa_tree_add_101_22_pad_groupi_n_6, csa_tree_add_101_22_pad_groupi_n_12, csa_tree_add_101_22_pad_groupi_n_13, csa_tree_add_101_22_pad_groupi_n_14, csa_tree_add_101_22_pad_groupi_n_15, csa_tree_add_101_22_pad_groupi_n_16, csa_tree_add_101_22_pad_groupi_n_17, csa_tree_add_101_22_pad_groupi_n_18;
  wire csa_tree_add_101_22_pad_groupi_n_19, csa_tree_add_101_22_pad_groupi_n_20, csa_tree_add_101_22_pad_groupi_n_21, csa_tree_add_101_22_pad_groupi_n_22, csa_tree_add_101_22_pad_groupi_n_23, csa_tree_add_101_22_pad_groupi_n_24, csa_tree_add_101_22_pad_groupi_n_25, csa_tree_add_101_22_pad_groupi_n_26;
  wire csa_tree_add_101_22_pad_groupi_n_27, csa_tree_add_101_22_pad_groupi_n_28, csa_tree_add_101_22_pad_groupi_n_29, csa_tree_add_101_22_pad_groupi_n_30, csa_tree_add_101_22_pad_groupi_n_31, csa_tree_add_101_22_pad_groupi_n_32, csa_tree_add_101_22_pad_groupi_n_33, csa_tree_add_101_22_pad_groupi_n_34;
  wire csa_tree_add_101_22_pad_groupi_n_35, csa_tree_add_101_22_pad_groupi_n_36, csa_tree_add_101_22_pad_groupi_n_37, csa_tree_add_101_22_pad_groupi_n_38, csa_tree_add_101_22_pad_groupi_n_39, csa_tree_add_101_22_pad_groupi_n_40, csa_tree_add_101_22_pad_groupi_n_41, csa_tree_add_101_22_pad_groupi_n_42;
  wire csa_tree_add_101_22_pad_groupi_n_43, csa_tree_add_101_22_pad_groupi_n_45, csa_tree_add_101_22_pad_groupi_n_46, csa_tree_add_101_22_pad_groupi_n_47, csa_tree_add_101_22_pad_groupi_n_48, csa_tree_add_101_22_pad_groupi_n_50, csa_tree_add_101_22_pad_groupi_n_51, csa_tree_add_101_22_pad_groupi_n_52;
  wire csa_tree_add_101_22_pad_groupi_n_53, csa_tree_add_101_22_pad_groupi_n_54, csa_tree_add_101_22_pad_groupi_n_55, csa_tree_add_101_22_pad_groupi_n_56, csa_tree_add_101_22_pad_groupi_n_57, csa_tree_add_101_22_pad_groupi_n_58, csa_tree_add_101_22_pad_groupi_n_59, csa_tree_add_101_22_pad_groupi_n_60;
  wire csa_tree_add_101_22_pad_groupi_n_61, csa_tree_add_101_22_pad_groupi_n_62, csa_tree_add_101_22_pad_groupi_n_64, csa_tree_add_101_22_pad_groupi_n_65, csa_tree_add_101_22_pad_groupi_n_66, csa_tree_add_101_22_pad_groupi_n_67, csa_tree_add_101_22_pad_groupi_n_68, csa_tree_add_101_22_pad_groupi_n_69;
  wire csa_tree_add_101_22_pad_groupi_n_70, csa_tree_add_101_22_pad_groupi_n_71, csa_tree_add_101_22_pad_groupi_n_72, csa_tree_add_101_22_pad_groupi_n_73, csa_tree_add_101_22_pad_groupi_n_74, csa_tree_add_101_22_pad_groupi_n_75, csa_tree_add_101_22_pad_groupi_n_76, csa_tree_add_101_22_pad_groupi_n_77;
  wire csa_tree_add_101_22_pad_groupi_n_78, csa_tree_add_101_22_pad_groupi_n_79, csa_tree_add_101_22_pad_groupi_n_80, csa_tree_add_101_22_pad_groupi_n_82, csa_tree_add_101_22_pad_groupi_n_83, csa_tree_add_101_22_pad_groupi_n_84, csa_tree_add_101_22_pad_groupi_n_85, csa_tree_add_101_22_pad_groupi_n_86;
  wire csa_tree_add_101_22_pad_groupi_n_87, csa_tree_add_101_22_pad_groupi_n_88, csa_tree_add_101_22_pad_groupi_n_89, csa_tree_add_101_22_pad_groupi_n_90, csa_tree_add_101_22_pad_groupi_n_91, csa_tree_add_101_22_pad_groupi_n_92, csa_tree_add_101_22_pad_groupi_n_93, csa_tree_add_101_22_pad_groupi_n_94;
  wire csa_tree_add_101_22_pad_groupi_n_95, csa_tree_add_101_22_pad_groupi_n_96, csa_tree_add_101_22_pad_groupi_n_97, csa_tree_add_101_22_pad_groupi_n_98, csa_tree_add_101_22_pad_groupi_n_99, csa_tree_add_101_22_pad_groupi_n_100, csa_tree_add_101_22_pad_groupi_n_101, csa_tree_add_101_22_pad_groupi_n_102;
  wire csa_tree_add_101_22_pad_groupi_n_103, csa_tree_add_101_22_pad_groupi_n_104, csa_tree_add_101_22_pad_groupi_n_105, csa_tree_add_101_22_pad_groupi_n_106, csa_tree_add_101_22_pad_groupi_n_107, csa_tree_add_101_22_pad_groupi_n_108, csa_tree_add_101_22_pad_groupi_n_109, csa_tree_add_101_22_pad_groupi_n_110;
  wire csa_tree_add_101_22_pad_groupi_n_111, csa_tree_add_101_22_pad_groupi_n_112, csa_tree_add_101_22_pad_groupi_n_113, csa_tree_add_101_22_pad_groupi_n_114, csa_tree_add_101_22_pad_groupi_n_115, csa_tree_add_101_22_pad_groupi_n_116, csa_tree_add_101_22_pad_groupi_n_117, csa_tree_add_101_22_pad_groupi_n_118;
  wire csa_tree_add_101_22_pad_groupi_n_119, csa_tree_add_101_22_pad_groupi_n_120, csa_tree_add_101_22_pad_groupi_n_121, csa_tree_add_101_22_pad_groupi_n_122, csa_tree_add_101_22_pad_groupi_n_123, csa_tree_add_101_22_pad_groupi_n_124, csa_tree_add_101_22_pad_groupi_n_125, csa_tree_add_101_22_pad_groupi_n_126;
  wire csa_tree_add_101_22_pad_groupi_n_127, csa_tree_add_101_22_pad_groupi_n_128, csa_tree_add_101_22_pad_groupi_n_129, csa_tree_add_101_22_pad_groupi_n_130, csa_tree_add_101_22_pad_groupi_n_131, csa_tree_add_101_22_pad_groupi_n_132, csa_tree_add_101_22_pad_groupi_n_133, csa_tree_add_101_22_pad_groupi_n_134;
  wire csa_tree_add_101_22_pad_groupi_n_135, csa_tree_add_101_22_pad_groupi_n_136, csa_tree_add_101_22_pad_groupi_n_137, csa_tree_add_101_22_pad_groupi_n_138, csa_tree_add_101_22_pad_groupi_n_139, csa_tree_add_101_22_pad_groupi_n_140, csa_tree_add_101_22_pad_groupi_n_141, csa_tree_add_101_22_pad_groupi_n_142;
  wire csa_tree_add_101_22_pad_groupi_n_143, csa_tree_add_101_22_pad_groupi_n_144, csa_tree_add_101_22_pad_groupi_n_145, csa_tree_add_101_22_pad_groupi_n_146, csa_tree_add_101_22_pad_groupi_n_147, csa_tree_add_101_22_pad_groupi_n_148, csa_tree_add_101_22_pad_groupi_n_149, csa_tree_add_101_22_pad_groupi_n_150;
  wire csa_tree_add_101_22_pad_groupi_n_151, csa_tree_add_101_22_pad_groupi_n_152, csa_tree_add_101_22_pad_groupi_n_153, csa_tree_add_101_22_pad_groupi_n_154, csa_tree_add_101_22_pad_groupi_n_155, csa_tree_add_101_22_pad_groupi_n_158, csa_tree_add_101_22_pad_groupi_n_159, csa_tree_add_101_22_pad_groupi_n_160;
  wire csa_tree_add_101_22_pad_groupi_n_161, csa_tree_add_101_22_pad_groupi_n_162, csa_tree_add_101_22_pad_groupi_n_163, csa_tree_add_101_22_pad_groupi_n_164, csa_tree_add_101_22_pad_groupi_n_165, csa_tree_add_101_22_pad_groupi_n_166, csa_tree_add_101_22_pad_groupi_n_167, csa_tree_add_101_22_pad_groupi_n_168;
  wire csa_tree_add_101_22_pad_groupi_n_169, csa_tree_add_101_22_pad_groupi_n_170, csa_tree_add_101_22_pad_groupi_n_171, csa_tree_add_101_22_pad_groupi_n_172, csa_tree_add_101_22_pad_groupi_n_173, csa_tree_add_101_22_pad_groupi_n_174, csa_tree_add_101_22_pad_groupi_n_175, csa_tree_add_101_22_pad_groupi_n_176;
  wire csa_tree_add_101_22_pad_groupi_n_177, csa_tree_add_101_22_pad_groupi_n_178, csa_tree_add_101_22_pad_groupi_n_179, csa_tree_add_101_22_pad_groupi_n_180, csa_tree_add_101_22_pad_groupi_n_181, csa_tree_add_101_22_pad_groupi_n_182, csa_tree_add_101_22_pad_groupi_n_183, csa_tree_add_101_22_pad_groupi_n_184;
  wire csa_tree_add_101_22_pad_groupi_n_185, csa_tree_add_101_22_pad_groupi_n_186, csa_tree_add_101_22_pad_groupi_n_187, csa_tree_add_101_22_pad_groupi_n_188, csa_tree_add_101_22_pad_groupi_n_189, csa_tree_add_101_22_pad_groupi_n_190, csa_tree_add_101_22_pad_groupi_n_191, csa_tree_add_101_22_pad_groupi_n_192;
  wire csa_tree_add_101_22_pad_groupi_n_193, csa_tree_add_101_22_pad_groupi_n_194, csa_tree_add_101_22_pad_groupi_n_195, csa_tree_add_101_22_pad_groupi_n_196, csa_tree_add_101_22_pad_groupi_n_197, csa_tree_add_101_22_pad_groupi_n_198, csa_tree_add_101_22_pad_groupi_n_200, csa_tree_add_101_22_pad_groupi_n_201;
  wire csa_tree_add_101_22_pad_groupi_n_202, csa_tree_add_101_22_pad_groupi_n_203, csa_tree_add_101_22_pad_groupi_n_204, csa_tree_add_101_22_pad_groupi_n_205, csa_tree_add_101_22_pad_groupi_n_206, csa_tree_add_101_22_pad_groupi_n_207, csa_tree_add_101_22_pad_groupi_n_208, csa_tree_add_101_22_pad_groupi_n_209;
  wire csa_tree_add_101_22_pad_groupi_n_210, csa_tree_add_101_22_pad_groupi_n_211, csa_tree_add_101_22_pad_groupi_n_212, csa_tree_add_101_22_pad_groupi_n_213, csa_tree_add_101_22_pad_groupi_n_214, csa_tree_add_101_22_pad_groupi_n_215, csa_tree_add_101_22_pad_groupi_n_216, csa_tree_add_101_22_pad_groupi_n_217;
  wire csa_tree_add_101_22_pad_groupi_n_218, csa_tree_add_101_22_pad_groupi_n_219, csa_tree_add_101_22_pad_groupi_n_220, csa_tree_add_101_22_pad_groupi_n_221, csa_tree_add_101_22_pad_groupi_n_222, csa_tree_add_101_22_pad_groupi_n_223, csa_tree_add_101_22_pad_groupi_n_224, csa_tree_add_101_22_pad_groupi_n_225;
  wire csa_tree_add_101_22_pad_groupi_n_226, csa_tree_add_101_22_pad_groupi_n_227, csa_tree_add_101_22_pad_groupi_n_228, csa_tree_add_101_22_pad_groupi_n_229, csa_tree_add_101_22_pad_groupi_n_230, csa_tree_add_101_22_pad_groupi_n_231, csa_tree_add_101_22_pad_groupi_n_232, csa_tree_add_101_22_pad_groupi_n_233;
  wire csa_tree_add_101_22_pad_groupi_n_234, csa_tree_add_101_22_pad_groupi_n_235, csa_tree_add_101_22_pad_groupi_n_236, csa_tree_add_101_22_pad_groupi_n_237, csa_tree_add_101_22_pad_groupi_n_238, csa_tree_add_101_22_pad_groupi_n_239, csa_tree_add_101_22_pad_groupi_n_240, csa_tree_add_101_22_pad_groupi_n_241;
  wire csa_tree_add_101_22_pad_groupi_n_242, csa_tree_add_101_22_pad_groupi_n_243, csa_tree_add_101_22_pad_groupi_n_244, csa_tree_add_101_22_pad_groupi_n_245, csa_tree_add_101_22_pad_groupi_n_246, csa_tree_add_101_22_pad_groupi_n_247, csa_tree_add_101_22_pad_groupi_n_248, csa_tree_add_101_22_pad_groupi_n_249;
  wire csa_tree_add_101_22_pad_groupi_n_250, csa_tree_add_101_22_pad_groupi_n_251, csa_tree_add_101_22_pad_groupi_n_252, csa_tree_add_101_22_pad_groupi_n_253, csa_tree_add_101_22_pad_groupi_n_254, csa_tree_add_101_22_pad_groupi_n_255, csa_tree_add_101_22_pad_groupi_n_256, csa_tree_add_101_22_pad_groupi_n_257;
  wire csa_tree_add_101_22_pad_groupi_n_258, csa_tree_add_101_22_pad_groupi_n_259, csa_tree_add_101_22_pad_groupi_n_260, csa_tree_add_101_22_pad_groupi_n_261, csa_tree_add_101_22_pad_groupi_n_262, csa_tree_add_101_22_pad_groupi_n_263, csa_tree_add_101_22_pad_groupi_n_264, csa_tree_add_101_22_pad_groupi_n_265;
  wire csa_tree_add_101_22_pad_groupi_n_266, csa_tree_add_101_22_pad_groupi_n_267, csa_tree_add_101_22_pad_groupi_n_268, csa_tree_add_101_22_pad_groupi_n_269, csa_tree_add_101_22_pad_groupi_n_270, csa_tree_add_101_22_pad_groupi_n_271, csa_tree_add_101_22_pad_groupi_n_272, csa_tree_add_101_22_pad_groupi_n_273;
  wire csa_tree_add_101_22_pad_groupi_n_274, csa_tree_add_101_22_pad_groupi_n_275, csa_tree_add_101_22_pad_groupi_n_276, csa_tree_add_101_22_pad_groupi_n_277, csa_tree_add_101_22_pad_groupi_n_278, csa_tree_add_101_22_pad_groupi_n_279, csa_tree_add_101_22_pad_groupi_n_280, csa_tree_add_101_22_pad_groupi_n_281;
  wire csa_tree_add_101_22_pad_groupi_n_282, csa_tree_add_101_22_pad_groupi_n_283, csa_tree_add_101_22_pad_groupi_n_284, csa_tree_add_101_22_pad_groupi_n_285, csa_tree_add_101_22_pad_groupi_n_286, csa_tree_add_101_22_pad_groupi_n_287, csa_tree_add_101_22_pad_groupi_n_288, csa_tree_add_101_22_pad_groupi_n_289;
  wire csa_tree_add_101_22_pad_groupi_n_290, csa_tree_add_101_22_pad_groupi_n_291, csa_tree_add_101_22_pad_groupi_n_292, csa_tree_add_101_22_pad_groupi_n_293, csa_tree_add_101_22_pad_groupi_n_294, csa_tree_add_101_22_pad_groupi_n_295, csa_tree_add_101_22_pad_groupi_n_296, csa_tree_add_101_22_pad_groupi_n_297;
  wire csa_tree_add_101_22_pad_groupi_n_298, csa_tree_add_101_22_pad_groupi_n_299, csa_tree_add_101_22_pad_groupi_n_300, csa_tree_add_101_22_pad_groupi_n_301, csa_tree_add_101_22_pad_groupi_n_302, csa_tree_add_101_22_pad_groupi_n_303, csa_tree_add_101_22_pad_groupi_n_304, csa_tree_add_101_22_pad_groupi_n_305;
  wire csa_tree_add_101_22_pad_groupi_n_306, csa_tree_add_101_22_pad_groupi_n_307, csa_tree_add_101_22_pad_groupi_n_308, csa_tree_add_101_22_pad_groupi_n_309, csa_tree_add_101_22_pad_groupi_n_310, csa_tree_add_101_22_pad_groupi_n_311, csa_tree_add_101_22_pad_groupi_n_312, csa_tree_add_101_22_pad_groupi_n_313;
  wire csa_tree_add_101_22_pad_groupi_n_314, csa_tree_add_101_22_pad_groupi_n_315, csa_tree_add_101_22_pad_groupi_n_316, csa_tree_add_101_22_pad_groupi_n_317, csa_tree_add_101_22_pad_groupi_n_318, csa_tree_add_101_22_pad_groupi_n_319, csa_tree_add_101_22_pad_groupi_n_320, csa_tree_add_101_22_pad_groupi_n_321;
  wire csa_tree_add_101_22_pad_groupi_n_322, csa_tree_add_101_22_pad_groupi_n_323, csa_tree_add_101_22_pad_groupi_n_324, csa_tree_add_101_22_pad_groupi_n_325, csa_tree_add_101_22_pad_groupi_n_326, csa_tree_add_101_22_pad_groupi_n_327, csa_tree_add_101_22_pad_groupi_n_328, csa_tree_add_101_22_pad_groupi_n_329;
  wire csa_tree_add_101_22_pad_groupi_n_330, csa_tree_add_101_22_pad_groupi_n_331, csa_tree_add_101_22_pad_groupi_n_332, csa_tree_add_101_22_pad_groupi_n_333, csa_tree_add_101_22_pad_groupi_n_334, csa_tree_add_101_22_pad_groupi_n_335, csa_tree_add_101_22_pad_groupi_n_336, csa_tree_add_101_22_pad_groupi_n_337;
  wire csa_tree_add_101_22_pad_groupi_n_338, csa_tree_add_101_22_pad_groupi_n_339, csa_tree_add_101_22_pad_groupi_n_340, csa_tree_add_101_22_pad_groupi_n_341, csa_tree_add_101_22_pad_groupi_n_342, csa_tree_add_101_22_pad_groupi_n_343, csa_tree_add_101_22_pad_groupi_n_344, csa_tree_add_101_22_pad_groupi_n_345;
  wire csa_tree_add_101_22_pad_groupi_n_346, csa_tree_add_101_22_pad_groupi_n_347, csa_tree_add_101_22_pad_groupi_n_348, csa_tree_add_101_22_pad_groupi_n_349, csa_tree_add_101_22_pad_groupi_n_350, csa_tree_add_101_22_pad_groupi_n_351, csa_tree_add_101_22_pad_groupi_n_352, csa_tree_add_101_22_pad_groupi_n_353;
  wire csa_tree_add_101_22_pad_groupi_n_354, csa_tree_add_101_22_pad_groupi_n_355, csa_tree_add_101_22_pad_groupi_n_356, csa_tree_add_101_22_pad_groupi_n_357, csa_tree_add_101_22_pad_groupi_n_358, csa_tree_add_101_22_pad_groupi_n_359, csa_tree_add_101_22_pad_groupi_n_361, csa_tree_add_101_22_pad_groupi_n_362;
  wire csa_tree_add_101_22_pad_groupi_n_363, csa_tree_add_101_22_pad_groupi_n_364, csa_tree_add_101_22_pad_groupi_n_365, csa_tree_add_101_22_pad_groupi_n_366, csa_tree_add_101_22_pad_groupi_n_367, csa_tree_add_101_22_pad_groupi_n_368, csa_tree_add_101_22_pad_groupi_n_369, csa_tree_add_101_22_pad_groupi_n_370;
  wire csa_tree_add_101_22_pad_groupi_n_371, csa_tree_add_101_22_pad_groupi_n_372, csa_tree_add_101_22_pad_groupi_n_373, csa_tree_add_101_22_pad_groupi_n_374, csa_tree_add_101_22_pad_groupi_n_375, csa_tree_add_101_22_pad_groupi_n_376, csa_tree_add_101_22_pad_groupi_n_377, csa_tree_add_101_22_pad_groupi_n_378;
  wire csa_tree_add_101_22_pad_groupi_n_379, csa_tree_add_101_22_pad_groupi_n_380, csa_tree_add_101_22_pad_groupi_n_381, csa_tree_add_101_22_pad_groupi_n_382, csa_tree_add_101_22_pad_groupi_n_383, csa_tree_add_101_22_pad_groupi_n_384, csa_tree_add_101_22_pad_groupi_n_385, csa_tree_add_101_22_pad_groupi_n_386;
  wire csa_tree_add_101_22_pad_groupi_n_387, csa_tree_add_101_22_pad_groupi_n_388, csa_tree_add_101_22_pad_groupi_n_389, csa_tree_add_101_22_pad_groupi_n_390, csa_tree_add_101_22_pad_groupi_n_391, csa_tree_add_101_22_pad_groupi_n_392, csa_tree_add_101_22_pad_groupi_n_393, csa_tree_add_101_22_pad_groupi_n_394;
  wire csa_tree_add_101_22_pad_groupi_n_395, csa_tree_add_101_22_pad_groupi_n_396, csa_tree_add_101_22_pad_groupi_n_397, csa_tree_add_101_22_pad_groupi_n_398, csa_tree_add_101_22_pad_groupi_n_399, csa_tree_add_101_22_pad_groupi_n_401, csa_tree_add_101_22_pad_groupi_n_402, csa_tree_add_101_22_pad_groupi_n_403;
  wire csa_tree_add_101_22_pad_groupi_n_404, csa_tree_add_101_22_pad_groupi_n_406, csa_tree_add_101_22_pad_groupi_n_409, csa_tree_add_101_22_pad_groupi_n_410, csa_tree_add_101_22_pad_groupi_n_411, csa_tree_add_101_22_pad_groupi_n_412, csa_tree_add_101_22_pad_groupi_n_413, csa_tree_add_101_22_pad_groupi_n_414;
  wire csa_tree_add_101_22_pad_groupi_n_415, csa_tree_add_101_22_pad_groupi_n_416, csa_tree_add_101_22_pad_groupi_n_417, csa_tree_add_101_22_pad_groupi_n_418, csa_tree_add_101_22_pad_groupi_n_419, csa_tree_add_101_22_pad_groupi_n_420, csa_tree_add_101_22_pad_groupi_n_421, csa_tree_add_101_22_pad_groupi_n_422;
  wire csa_tree_add_101_22_pad_groupi_n_423, csa_tree_add_101_22_pad_groupi_n_424, csa_tree_add_101_22_pad_groupi_n_425, csa_tree_add_101_22_pad_groupi_n_426, csa_tree_add_101_22_pad_groupi_n_427, csa_tree_add_101_22_pad_groupi_n_428, csa_tree_add_101_22_pad_groupi_n_429, csa_tree_add_101_22_pad_groupi_n_430;
  wire csa_tree_add_101_22_pad_groupi_n_431, csa_tree_add_101_22_pad_groupi_n_432, csa_tree_add_101_22_pad_groupi_n_433, csa_tree_add_101_22_pad_groupi_n_434, csa_tree_add_101_22_pad_groupi_n_435, csa_tree_add_101_22_pad_groupi_n_438, csa_tree_add_101_22_pad_groupi_n_439, csa_tree_add_101_22_pad_groupi_n_445;
  wire csa_tree_add_101_22_pad_groupi_n_455, csa_tree_add_101_22_pad_groupi_n_456, csa_tree_add_101_22_pad_groupi_n_457, csa_tree_add_101_22_pad_groupi_n_458, csa_tree_add_101_22_pad_groupi_n_459, csa_tree_add_101_22_pad_groupi_n_460, csa_tree_add_101_22_pad_groupi_n_461, csa_tree_add_101_22_pad_groupi_n_462;
  wire csa_tree_add_101_22_pad_groupi_n_463, csa_tree_add_101_22_pad_groupi_n_464, csa_tree_add_101_22_pad_groupi_n_465, csa_tree_add_101_22_pad_groupi_n_466, csa_tree_add_101_22_pad_groupi_n_467, csa_tree_add_101_22_pad_groupi_n_468, csa_tree_add_101_22_pad_groupi_n_469, csa_tree_add_101_22_pad_groupi_n_470;
  wire csa_tree_add_101_22_pad_groupi_n_471, csa_tree_add_101_22_pad_groupi_n_472, csa_tree_add_101_22_pad_groupi_n_473, csa_tree_add_101_22_pad_groupi_n_474, csa_tree_add_101_22_pad_groupi_n_475, csa_tree_add_101_22_pad_groupi_n_476, csa_tree_add_101_22_pad_groupi_n_477, csa_tree_add_101_22_pad_groupi_n_478;
  wire csa_tree_add_101_22_pad_groupi_n_479, csa_tree_add_101_22_pad_groupi_n_480, csa_tree_add_101_22_pad_groupi_n_481, csa_tree_add_101_22_pad_groupi_n_482, csa_tree_add_101_22_pad_groupi_n_483, csa_tree_add_101_22_pad_groupi_n_484, csa_tree_add_101_22_pad_groupi_n_485, csa_tree_add_101_22_pad_groupi_n_486;
  wire csa_tree_add_101_22_pad_groupi_n_487, csa_tree_add_101_22_pad_groupi_n_488, csa_tree_add_101_22_pad_groupi_n_489, csa_tree_add_101_22_pad_groupi_n_490, csa_tree_add_101_22_pad_groupi_n_491, csa_tree_add_101_22_pad_groupi_n_492, csa_tree_add_101_22_pad_groupi_n_493, csa_tree_add_101_22_pad_groupi_n_494;
  wire csa_tree_add_101_22_pad_groupi_n_495, csa_tree_add_101_22_pad_groupi_n_496, csa_tree_add_101_22_pad_groupi_n_497, csa_tree_add_101_22_pad_groupi_n_498, csa_tree_add_101_22_pad_groupi_n_499, csa_tree_add_101_22_pad_groupi_n_500, csa_tree_add_101_22_pad_groupi_n_501, csa_tree_add_101_22_pad_groupi_n_502;
  wire csa_tree_add_101_22_pad_groupi_n_503, csa_tree_add_101_22_pad_groupi_n_504, csa_tree_add_101_22_pad_groupi_n_505, csa_tree_add_101_22_pad_groupi_n_506, csa_tree_add_101_22_pad_groupi_n_507, csa_tree_add_101_22_pad_groupi_n_508, csa_tree_add_101_22_pad_groupi_n_509, csa_tree_add_101_22_pad_groupi_n_510;
  wire csa_tree_add_101_22_pad_groupi_n_511, csa_tree_add_101_22_pad_groupi_n_512, csa_tree_add_101_22_pad_groupi_n_513, csa_tree_add_101_22_pad_groupi_n_514, csa_tree_add_101_22_pad_groupi_n_515, csa_tree_add_101_22_pad_groupi_n_516, csa_tree_add_101_22_pad_groupi_n_517, csa_tree_add_101_22_pad_groupi_n_518;
  wire csa_tree_add_101_22_pad_groupi_n_519, csa_tree_add_101_22_pad_groupi_n_520, csa_tree_add_101_22_pad_groupi_n_521, csa_tree_add_101_22_pad_groupi_n_522, csa_tree_add_101_22_pad_groupi_n_523, csa_tree_add_101_22_pad_groupi_n_524, csa_tree_add_101_22_pad_groupi_n_525, csa_tree_add_101_22_pad_groupi_n_526;
  wire csa_tree_add_101_22_pad_groupi_n_527, csa_tree_add_101_22_pad_groupi_n_528, csa_tree_add_101_22_pad_groupi_n_529, csa_tree_add_101_22_pad_groupi_n_530, csa_tree_add_101_22_pad_groupi_n_531, csa_tree_add_101_22_pad_groupi_n_532, csa_tree_add_101_22_pad_groupi_n_533, csa_tree_add_101_22_pad_groupi_n_534;
  wire csa_tree_add_101_22_pad_groupi_n_535, csa_tree_add_101_22_pad_groupi_n_536, csa_tree_add_101_22_pad_groupi_n_537, csa_tree_add_101_22_pad_groupi_n_538, csa_tree_add_101_22_pad_groupi_n_539, csa_tree_add_101_22_pad_groupi_n_540, csa_tree_add_101_22_pad_groupi_n_541, csa_tree_add_101_22_pad_groupi_n_542;
  wire csa_tree_add_101_22_pad_groupi_n_543, csa_tree_add_101_22_pad_groupi_n_544, csa_tree_add_101_22_pad_groupi_n_545, csa_tree_add_101_22_pad_groupi_n_546, csa_tree_add_101_22_pad_groupi_n_547, csa_tree_add_101_22_pad_groupi_n_548, csa_tree_add_101_22_pad_groupi_n_549, csa_tree_add_101_22_pad_groupi_n_550;
  wire csa_tree_add_101_22_pad_groupi_n_551, csa_tree_add_101_22_pad_groupi_n_552, csa_tree_add_101_22_pad_groupi_n_553, csa_tree_add_101_22_pad_groupi_n_554, csa_tree_add_101_22_pad_groupi_n_555, csa_tree_add_101_22_pad_groupi_n_556, csa_tree_add_101_22_pad_groupi_n_557, csa_tree_add_101_22_pad_groupi_n_559;
  wire csa_tree_add_101_22_pad_groupi_n_561, csa_tree_add_101_22_pad_groupi_n_562, csa_tree_add_101_22_pad_groupi_n_563, csa_tree_add_101_22_pad_groupi_n_564, csa_tree_add_101_22_pad_groupi_n_565, csa_tree_add_101_22_pad_groupi_n_566, csa_tree_add_101_22_pad_groupi_n_567, csa_tree_add_101_22_pad_groupi_n_568;
  wire csa_tree_add_101_22_pad_groupi_n_569, csa_tree_add_101_22_pad_groupi_n_570, csa_tree_add_101_22_pad_groupi_n_572, csa_tree_add_101_22_pad_groupi_n_573, csa_tree_add_101_22_pad_groupi_n_574, csa_tree_add_101_22_pad_groupi_n_575, csa_tree_add_101_22_pad_groupi_n_576, csa_tree_add_101_22_pad_groupi_n_577;
  wire csa_tree_add_101_22_pad_groupi_n_578, csa_tree_add_101_22_pad_groupi_n_579, csa_tree_add_101_22_pad_groupi_n_580, csa_tree_add_101_22_pad_groupi_n_581, csa_tree_add_101_22_pad_groupi_n_582, csa_tree_add_101_22_pad_groupi_n_583, csa_tree_add_101_22_pad_groupi_n_584, csa_tree_add_101_22_pad_groupi_n_586;
  wire csa_tree_add_101_22_pad_groupi_n_587, csa_tree_add_101_22_pad_groupi_n_588, csa_tree_add_101_22_pad_groupi_n_589, csa_tree_add_101_22_pad_groupi_n_590, csa_tree_add_101_22_pad_groupi_n_591, csa_tree_add_101_22_pad_groupi_n_592, csa_tree_add_101_22_pad_groupi_n_593, csa_tree_add_101_22_pad_groupi_n_594;
  wire csa_tree_add_101_22_pad_groupi_n_595, csa_tree_add_101_22_pad_groupi_n_598, csa_tree_add_101_22_pad_groupi_n_599, csa_tree_add_101_22_pad_groupi_n_600, csa_tree_add_101_22_pad_groupi_n_601, csa_tree_add_101_22_pad_groupi_n_602, csa_tree_add_101_22_pad_groupi_n_603, csa_tree_add_101_22_pad_groupi_n_604;
  wire csa_tree_add_101_22_pad_groupi_n_605, csa_tree_add_101_22_pad_groupi_n_606, csa_tree_add_101_22_pad_groupi_n_607, csa_tree_add_101_22_pad_groupi_n_608, csa_tree_add_101_22_pad_groupi_n_609, csa_tree_add_101_22_pad_groupi_n_610, csa_tree_add_101_22_pad_groupi_n_611, csa_tree_add_101_22_pad_groupi_n_612;
  wire csa_tree_add_101_22_pad_groupi_n_613, csa_tree_add_101_22_pad_groupi_n_614, csa_tree_add_101_22_pad_groupi_n_615, csa_tree_add_101_22_pad_groupi_n_616, csa_tree_add_101_22_pad_groupi_n_617, csa_tree_add_101_22_pad_groupi_n_618, csa_tree_add_101_22_pad_groupi_n_619, csa_tree_add_101_22_pad_groupi_n_620;
  wire csa_tree_add_101_22_pad_groupi_n_621, csa_tree_add_101_22_pad_groupi_n_622, csa_tree_add_101_22_pad_groupi_n_623, csa_tree_add_101_22_pad_groupi_n_624, csa_tree_add_101_22_pad_groupi_n_625, csa_tree_add_101_22_pad_groupi_n_626, csa_tree_add_101_22_pad_groupi_n_627, csa_tree_add_101_22_pad_groupi_n_628;
  wire csa_tree_add_101_22_pad_groupi_n_629, csa_tree_add_101_22_pad_groupi_n_630, csa_tree_add_101_22_pad_groupi_n_631, csa_tree_add_101_22_pad_groupi_n_633, csa_tree_add_101_22_pad_groupi_n_634, csa_tree_add_101_22_pad_groupi_n_635, csa_tree_add_101_22_pad_groupi_n_637, csa_tree_add_101_22_pad_groupi_n_638;
  wire csa_tree_add_101_22_pad_groupi_n_639, csa_tree_add_101_22_pad_groupi_n_640, csa_tree_add_101_22_pad_groupi_n_641, csa_tree_add_101_22_pad_groupi_n_642, csa_tree_add_101_22_pad_groupi_n_643, csa_tree_add_101_22_pad_groupi_n_644, csa_tree_add_101_22_pad_groupi_n_645, csa_tree_add_101_22_pad_groupi_n_646;
  wire csa_tree_add_101_22_pad_groupi_n_647, csa_tree_add_101_22_pad_groupi_n_648, csa_tree_add_101_22_pad_groupi_n_649, csa_tree_add_101_22_pad_groupi_n_650, csa_tree_add_101_22_pad_groupi_n_651, csa_tree_add_101_22_pad_groupi_n_652, csa_tree_add_101_22_pad_groupi_n_653, csa_tree_add_101_22_pad_groupi_n_654;
  wire csa_tree_add_101_22_pad_groupi_n_655, csa_tree_add_101_22_pad_groupi_n_656, csa_tree_add_101_22_pad_groupi_n_657, csa_tree_add_101_22_pad_groupi_n_658, csa_tree_add_101_22_pad_groupi_n_659, csa_tree_add_101_22_pad_groupi_n_660, csa_tree_add_101_22_pad_groupi_n_661, csa_tree_add_101_22_pad_groupi_n_662;
  wire csa_tree_add_101_22_pad_groupi_n_663, csa_tree_add_101_22_pad_groupi_n_664, csa_tree_add_101_22_pad_groupi_n_665, csa_tree_add_101_22_pad_groupi_n_666, csa_tree_add_101_22_pad_groupi_n_667, csa_tree_add_101_22_pad_groupi_n_668, csa_tree_add_101_22_pad_groupi_n_669, csa_tree_add_101_22_pad_groupi_n_670;
  wire csa_tree_add_101_22_pad_groupi_n_671, csa_tree_add_101_22_pad_groupi_n_672, csa_tree_add_101_22_pad_groupi_n_673, csa_tree_add_101_22_pad_groupi_n_674, csa_tree_add_101_22_pad_groupi_n_675, csa_tree_add_101_22_pad_groupi_n_676, csa_tree_add_101_22_pad_groupi_n_677, csa_tree_add_101_22_pad_groupi_n_678;
  wire csa_tree_add_101_22_pad_groupi_n_679, csa_tree_add_101_22_pad_groupi_n_680, csa_tree_add_101_22_pad_groupi_n_681, csa_tree_add_101_22_pad_groupi_n_682, csa_tree_add_101_22_pad_groupi_n_683, csa_tree_add_101_22_pad_groupi_n_684, csa_tree_add_101_22_pad_groupi_n_685, csa_tree_add_101_22_pad_groupi_n_686;
  wire csa_tree_add_101_22_pad_groupi_n_688, csa_tree_add_101_22_pad_groupi_n_689, csa_tree_add_101_22_pad_groupi_n_690, csa_tree_add_101_22_pad_groupi_n_691, csa_tree_add_101_22_pad_groupi_n_692, csa_tree_add_101_22_pad_groupi_n_693, csa_tree_add_101_22_pad_groupi_n_694, csa_tree_add_101_22_pad_groupi_n_695;
  wire csa_tree_add_101_22_pad_groupi_n_696, csa_tree_add_101_22_pad_groupi_n_697, csa_tree_add_101_22_pad_groupi_n_698, csa_tree_add_101_22_pad_groupi_n_699, csa_tree_add_101_22_pad_groupi_n_700, csa_tree_add_101_22_pad_groupi_n_702, csa_tree_add_101_22_pad_groupi_n_703, csa_tree_add_101_22_pad_groupi_n_704;
  wire csa_tree_add_101_22_pad_groupi_n_705, csa_tree_add_101_22_pad_groupi_n_706, csa_tree_add_101_22_pad_groupi_n_707, csa_tree_add_101_22_pad_groupi_n_708, csa_tree_add_101_22_pad_groupi_n_709, csa_tree_add_101_22_pad_groupi_n_710, csa_tree_add_101_22_pad_groupi_n_711, csa_tree_add_101_22_pad_groupi_n_712;
  wire csa_tree_add_101_22_pad_groupi_n_713, csa_tree_add_101_22_pad_groupi_n_714, csa_tree_add_101_22_pad_groupi_n_715, csa_tree_add_101_22_pad_groupi_n_716, csa_tree_add_101_22_pad_groupi_n_717, csa_tree_add_101_22_pad_groupi_n_718, csa_tree_add_101_22_pad_groupi_n_719, csa_tree_add_101_22_pad_groupi_n_720;
  wire csa_tree_add_101_22_pad_groupi_n_721, csa_tree_add_101_22_pad_groupi_n_722, csa_tree_add_101_22_pad_groupi_n_723, csa_tree_add_101_22_pad_groupi_n_724, csa_tree_add_101_22_pad_groupi_n_725, csa_tree_add_101_22_pad_groupi_n_726, csa_tree_add_101_22_pad_groupi_n_727, csa_tree_add_101_22_pad_groupi_n_728;
  wire csa_tree_add_101_22_pad_groupi_n_729, csa_tree_add_101_22_pad_groupi_n_730, csa_tree_add_101_22_pad_groupi_n_731, csa_tree_add_101_22_pad_groupi_n_732, csa_tree_add_101_22_pad_groupi_n_733, csa_tree_add_101_22_pad_groupi_n_734, csa_tree_add_101_22_pad_groupi_n_735, csa_tree_add_101_22_pad_groupi_n_736;
  wire csa_tree_add_101_22_pad_groupi_n_737, csa_tree_add_101_22_pad_groupi_n_738, csa_tree_add_101_22_pad_groupi_n_739, csa_tree_add_101_22_pad_groupi_n_740, csa_tree_add_101_22_pad_groupi_n_741, csa_tree_add_101_22_pad_groupi_n_742, csa_tree_add_101_22_pad_groupi_n_743, csa_tree_add_101_22_pad_groupi_n_744;
  wire csa_tree_add_101_22_pad_groupi_n_745, csa_tree_add_101_22_pad_groupi_n_746, csa_tree_add_101_22_pad_groupi_n_747, csa_tree_add_101_22_pad_groupi_n_748, csa_tree_add_101_22_pad_groupi_n_749, csa_tree_add_101_22_pad_groupi_n_750, csa_tree_add_101_22_pad_groupi_n_751, csa_tree_add_101_22_pad_groupi_n_752;
  wire csa_tree_add_101_22_pad_groupi_n_753, csa_tree_add_101_22_pad_groupi_n_754, csa_tree_add_101_22_pad_groupi_n_755, csa_tree_add_101_22_pad_groupi_n_756, csa_tree_add_101_22_pad_groupi_n_757, csa_tree_add_101_22_pad_groupi_n_758, csa_tree_add_101_22_pad_groupi_n_759, csa_tree_add_101_22_pad_groupi_n_760;
  wire csa_tree_add_101_22_pad_groupi_n_761, csa_tree_add_101_22_pad_groupi_n_762, csa_tree_add_101_22_pad_groupi_n_763, csa_tree_add_101_22_pad_groupi_n_764, csa_tree_add_101_22_pad_groupi_n_765, csa_tree_add_101_22_pad_groupi_n_766, csa_tree_add_101_22_pad_groupi_n_767, csa_tree_add_101_22_pad_groupi_n_768;
  wire csa_tree_add_101_22_pad_groupi_n_769, csa_tree_add_101_22_pad_groupi_n_770, csa_tree_add_101_22_pad_groupi_n_771, csa_tree_add_101_22_pad_groupi_n_772, csa_tree_add_101_22_pad_groupi_n_773, csa_tree_add_101_22_pad_groupi_n_774, csa_tree_add_101_22_pad_groupi_n_775, csa_tree_add_101_22_pad_groupi_n_776;
  wire csa_tree_add_101_22_pad_groupi_n_777, csa_tree_add_101_22_pad_groupi_n_778, csa_tree_add_101_22_pad_groupi_n_779, csa_tree_add_101_22_pad_groupi_n_780, csa_tree_add_101_22_pad_groupi_n_781, csa_tree_add_101_22_pad_groupi_n_782, csa_tree_add_101_22_pad_groupi_n_783, csa_tree_add_101_22_pad_groupi_n_784;
  wire csa_tree_add_101_22_pad_groupi_n_785, csa_tree_add_101_22_pad_groupi_n_786, csa_tree_add_101_22_pad_groupi_n_787, csa_tree_add_101_22_pad_groupi_n_788, csa_tree_add_101_22_pad_groupi_n_789, csa_tree_add_101_22_pad_groupi_n_790, csa_tree_add_101_22_pad_groupi_n_791, csa_tree_add_101_22_pad_groupi_n_792;
  wire csa_tree_add_101_22_pad_groupi_n_793, csa_tree_add_101_22_pad_groupi_n_794, csa_tree_add_101_22_pad_groupi_n_795, csa_tree_add_101_22_pad_groupi_n_796, csa_tree_add_101_22_pad_groupi_n_797, csa_tree_add_101_22_pad_groupi_n_798, csa_tree_add_101_22_pad_groupi_n_799, csa_tree_add_101_22_pad_groupi_n_800;
  wire csa_tree_add_101_22_pad_groupi_n_801, csa_tree_add_101_22_pad_groupi_n_802, csa_tree_add_101_22_pad_groupi_n_803, csa_tree_add_101_22_pad_groupi_n_804, csa_tree_add_101_22_pad_groupi_n_805, csa_tree_add_101_22_pad_groupi_n_806, csa_tree_add_101_22_pad_groupi_n_807, csa_tree_add_101_22_pad_groupi_n_808;
  wire csa_tree_add_101_22_pad_groupi_n_809, csa_tree_add_101_22_pad_groupi_n_810, csa_tree_add_101_22_pad_groupi_n_811, csa_tree_add_101_22_pad_groupi_n_812, csa_tree_add_101_22_pad_groupi_n_813, csa_tree_add_101_22_pad_groupi_n_814, csa_tree_add_101_22_pad_groupi_n_815, csa_tree_add_101_22_pad_groupi_n_816;
  wire csa_tree_add_101_22_pad_groupi_n_817, csa_tree_add_101_22_pad_groupi_n_818, csa_tree_add_101_22_pad_groupi_n_819, csa_tree_add_101_22_pad_groupi_n_820, csa_tree_add_101_22_pad_groupi_n_821, csa_tree_add_101_22_pad_groupi_n_822, csa_tree_add_101_22_pad_groupi_n_823, csa_tree_add_101_22_pad_groupi_n_824;
  wire csa_tree_add_101_22_pad_groupi_n_825, csa_tree_add_101_22_pad_groupi_n_826, csa_tree_add_101_22_pad_groupi_n_827, csa_tree_add_101_22_pad_groupi_n_828, csa_tree_add_101_22_pad_groupi_n_829, csa_tree_add_101_22_pad_groupi_n_830, csa_tree_add_101_22_pad_groupi_n_831, csa_tree_add_101_22_pad_groupi_n_832;
  wire csa_tree_add_101_22_pad_groupi_n_833, csa_tree_add_101_22_pad_groupi_n_834, csa_tree_add_101_22_pad_groupi_n_835, csa_tree_add_101_22_pad_groupi_n_836, csa_tree_add_101_22_pad_groupi_n_837, csa_tree_add_101_22_pad_groupi_n_838, csa_tree_add_101_22_pad_groupi_n_839, csa_tree_add_101_22_pad_groupi_n_840;
  wire csa_tree_add_101_22_pad_groupi_n_841, csa_tree_add_101_22_pad_groupi_n_842, csa_tree_add_101_22_pad_groupi_n_843, csa_tree_add_101_22_pad_groupi_n_844, csa_tree_add_101_22_pad_groupi_n_845, csa_tree_add_101_22_pad_groupi_n_846, csa_tree_add_101_22_pad_groupi_n_847, csa_tree_add_101_22_pad_groupi_n_848;
  wire csa_tree_add_101_22_pad_groupi_n_849, csa_tree_add_101_22_pad_groupi_n_851, csa_tree_add_101_22_pad_groupi_n_852, csa_tree_add_101_22_pad_groupi_n_853, csa_tree_add_101_22_pad_groupi_n_854, csa_tree_add_101_22_pad_groupi_n_855, csa_tree_add_101_22_pad_groupi_n_856, csa_tree_add_101_22_pad_groupi_n_857;
  wire csa_tree_add_101_22_pad_groupi_n_858, csa_tree_add_101_22_pad_groupi_n_859, csa_tree_add_101_22_pad_groupi_n_860, csa_tree_add_101_22_pad_groupi_n_861, csa_tree_add_101_22_pad_groupi_n_862, csa_tree_add_101_22_pad_groupi_n_863, csa_tree_add_101_22_pad_groupi_n_864, csa_tree_add_101_22_pad_groupi_n_865;
  wire csa_tree_add_101_22_pad_groupi_n_866, csa_tree_add_101_22_pad_groupi_n_867, csa_tree_add_101_22_pad_groupi_n_868, csa_tree_add_101_22_pad_groupi_n_869, csa_tree_add_101_22_pad_groupi_n_870, csa_tree_add_101_22_pad_groupi_n_871, csa_tree_add_101_22_pad_groupi_n_872, csa_tree_add_101_22_pad_groupi_n_873;
  wire csa_tree_add_101_22_pad_groupi_n_874, csa_tree_add_101_22_pad_groupi_n_875, csa_tree_add_101_22_pad_groupi_n_876, csa_tree_add_101_22_pad_groupi_n_877, csa_tree_add_101_22_pad_groupi_n_878, csa_tree_add_101_22_pad_groupi_n_879, csa_tree_add_101_22_pad_groupi_n_880, csa_tree_add_101_22_pad_groupi_n_881;
  wire csa_tree_add_101_22_pad_groupi_n_882, csa_tree_add_101_22_pad_groupi_n_883, csa_tree_add_101_22_pad_groupi_n_884, csa_tree_add_101_22_pad_groupi_n_885, csa_tree_add_101_22_pad_groupi_n_886, csa_tree_add_101_22_pad_groupi_n_887, csa_tree_add_101_22_pad_groupi_n_888, csa_tree_add_101_22_pad_groupi_n_889;
  wire csa_tree_add_101_22_pad_groupi_n_890, csa_tree_add_101_22_pad_groupi_n_891, csa_tree_add_101_22_pad_groupi_n_892, csa_tree_add_101_22_pad_groupi_n_893, csa_tree_add_101_22_pad_groupi_n_894, csa_tree_add_101_22_pad_groupi_n_895, csa_tree_add_101_22_pad_groupi_n_896, csa_tree_add_101_22_pad_groupi_n_897;
  wire csa_tree_add_101_22_pad_groupi_n_898, csa_tree_add_101_22_pad_groupi_n_899, csa_tree_add_101_22_pad_groupi_n_900, csa_tree_add_101_22_pad_groupi_n_901, csa_tree_add_101_22_pad_groupi_n_902, csa_tree_add_101_22_pad_groupi_n_903, csa_tree_add_101_22_pad_groupi_n_904, csa_tree_add_101_22_pad_groupi_n_905;
  wire csa_tree_add_101_22_pad_groupi_n_906, csa_tree_add_101_22_pad_groupi_n_907, csa_tree_add_101_22_pad_groupi_n_908, csa_tree_add_101_22_pad_groupi_n_909, csa_tree_add_101_22_pad_groupi_n_910, csa_tree_add_101_22_pad_groupi_n_911, csa_tree_add_101_22_pad_groupi_n_912, csa_tree_add_101_22_pad_groupi_n_913;
  wire csa_tree_add_101_22_pad_groupi_n_914, csa_tree_add_101_22_pad_groupi_n_915, csa_tree_add_101_22_pad_groupi_n_916, csa_tree_add_101_22_pad_groupi_n_917, csa_tree_add_101_22_pad_groupi_n_918, csa_tree_add_101_22_pad_groupi_n_919, csa_tree_add_101_22_pad_groupi_n_920, csa_tree_add_101_22_pad_groupi_n_921;
  wire csa_tree_add_101_22_pad_groupi_n_922, csa_tree_add_101_22_pad_groupi_n_923, csa_tree_add_101_22_pad_groupi_n_924, csa_tree_add_101_22_pad_groupi_n_925, csa_tree_add_101_22_pad_groupi_n_926, csa_tree_add_101_22_pad_groupi_n_927, csa_tree_add_101_22_pad_groupi_n_928, csa_tree_add_101_22_pad_groupi_n_929;
  wire csa_tree_add_101_22_pad_groupi_n_930, csa_tree_add_101_22_pad_groupi_n_931, csa_tree_add_101_22_pad_groupi_n_932, csa_tree_add_101_22_pad_groupi_n_933, csa_tree_add_101_22_pad_groupi_n_934, csa_tree_add_101_22_pad_groupi_n_935, csa_tree_add_101_22_pad_groupi_n_936, csa_tree_add_101_22_pad_groupi_n_937;
  wire csa_tree_add_101_22_pad_groupi_n_938, csa_tree_add_101_22_pad_groupi_n_939, csa_tree_add_101_22_pad_groupi_n_940, csa_tree_add_101_22_pad_groupi_n_941, csa_tree_add_101_22_pad_groupi_n_942, csa_tree_add_101_22_pad_groupi_n_943, csa_tree_add_101_22_pad_groupi_n_944, csa_tree_add_101_22_pad_groupi_n_945;
  wire csa_tree_add_101_22_pad_groupi_n_946, csa_tree_add_101_22_pad_groupi_n_947, csa_tree_add_101_22_pad_groupi_n_948, csa_tree_add_101_22_pad_groupi_n_949, csa_tree_add_101_22_pad_groupi_n_950, csa_tree_add_101_22_pad_groupi_n_951, csa_tree_add_101_22_pad_groupi_n_952, csa_tree_add_101_22_pad_groupi_n_953;
  wire csa_tree_add_101_22_pad_groupi_n_954, csa_tree_add_101_22_pad_groupi_n_955, csa_tree_add_101_22_pad_groupi_n_956, csa_tree_add_101_22_pad_groupi_n_957, csa_tree_add_101_22_pad_groupi_n_958, csa_tree_add_101_22_pad_groupi_n_959, csa_tree_add_101_22_pad_groupi_n_960, csa_tree_add_101_22_pad_groupi_n_961;
  wire csa_tree_add_101_22_pad_groupi_n_962, csa_tree_add_101_22_pad_groupi_n_963, csa_tree_add_101_22_pad_groupi_n_964, csa_tree_add_101_22_pad_groupi_n_965, csa_tree_add_101_22_pad_groupi_n_966, csa_tree_add_101_22_pad_groupi_n_967, csa_tree_add_101_22_pad_groupi_n_968, csa_tree_add_101_22_pad_groupi_n_969;
  wire csa_tree_add_101_22_pad_groupi_n_970, csa_tree_add_101_22_pad_groupi_n_971, csa_tree_add_101_22_pad_groupi_n_972, csa_tree_add_101_22_pad_groupi_n_973, csa_tree_add_101_22_pad_groupi_n_974, csa_tree_add_101_22_pad_groupi_n_975, csa_tree_add_101_22_pad_groupi_n_976, csa_tree_add_101_22_pad_groupi_n_977;
  wire csa_tree_add_101_22_pad_groupi_n_978, csa_tree_add_101_22_pad_groupi_n_979, csa_tree_add_101_22_pad_groupi_n_980, csa_tree_add_101_22_pad_groupi_n_981, csa_tree_add_101_22_pad_groupi_n_982, csa_tree_add_101_22_pad_groupi_n_983, csa_tree_add_101_22_pad_groupi_n_984, csa_tree_add_101_22_pad_groupi_n_985;
  wire csa_tree_add_101_22_pad_groupi_n_986, csa_tree_add_101_22_pad_groupi_n_987, csa_tree_add_101_22_pad_groupi_n_988, csa_tree_add_101_22_pad_groupi_n_989, csa_tree_add_101_22_pad_groupi_n_990, csa_tree_add_101_22_pad_groupi_n_991, csa_tree_add_101_22_pad_groupi_n_992, csa_tree_add_101_22_pad_groupi_n_993;
  wire csa_tree_add_101_22_pad_groupi_n_994, csa_tree_add_101_22_pad_groupi_n_995, csa_tree_add_101_22_pad_groupi_n_996, csa_tree_add_101_22_pad_groupi_n_997, csa_tree_add_101_22_pad_groupi_n_998, csa_tree_add_101_22_pad_groupi_n_999, csa_tree_add_101_22_pad_groupi_n_1000, csa_tree_add_101_22_pad_groupi_n_1001;
  wire csa_tree_add_101_22_pad_groupi_n_1002, csa_tree_add_101_22_pad_groupi_n_1003, csa_tree_add_101_22_pad_groupi_n_1004, csa_tree_add_101_22_pad_groupi_n_1005, csa_tree_add_101_22_pad_groupi_n_1006, csa_tree_add_101_22_pad_groupi_n_1007, csa_tree_add_101_22_pad_groupi_n_1008, csa_tree_add_101_22_pad_groupi_n_1009;
  wire csa_tree_add_101_22_pad_groupi_n_1010, csa_tree_add_101_22_pad_groupi_n_1011, csa_tree_add_101_22_pad_groupi_n_1012, csa_tree_add_101_22_pad_groupi_n_1013, csa_tree_add_101_22_pad_groupi_n_1014, csa_tree_add_101_22_pad_groupi_n_1015, csa_tree_add_101_22_pad_groupi_n_1016, csa_tree_add_101_22_pad_groupi_n_1017;
  wire csa_tree_add_101_22_pad_groupi_n_1018, csa_tree_add_101_22_pad_groupi_n_1019, csa_tree_add_101_22_pad_groupi_n_1020, csa_tree_add_101_22_pad_groupi_n_1021, csa_tree_add_101_22_pad_groupi_n_1022, csa_tree_add_101_22_pad_groupi_n_1023, csa_tree_add_101_22_pad_groupi_n_1024, csa_tree_add_101_22_pad_groupi_n_1025;
  wire csa_tree_add_101_22_pad_groupi_n_1026, csa_tree_add_101_22_pad_groupi_n_1027, csa_tree_add_101_22_pad_groupi_n_1028, csa_tree_add_101_22_pad_groupi_n_1029, csa_tree_add_101_22_pad_groupi_n_1030, csa_tree_add_101_22_pad_groupi_n_1031, csa_tree_add_101_22_pad_groupi_n_1032, csa_tree_add_101_22_pad_groupi_n_1033;
  wire csa_tree_add_101_22_pad_groupi_n_1034, csa_tree_add_101_22_pad_groupi_n_1035, csa_tree_add_101_22_pad_groupi_n_1036, csa_tree_add_101_22_pad_groupi_n_1037, csa_tree_add_101_22_pad_groupi_n_1038, csa_tree_add_101_22_pad_groupi_n_1039, csa_tree_add_101_22_pad_groupi_n_1040, csa_tree_add_101_22_pad_groupi_n_1041;
  wire csa_tree_add_101_22_pad_groupi_n_1042, csa_tree_add_101_22_pad_groupi_n_1043, csa_tree_add_101_22_pad_groupi_n_1044, csa_tree_add_101_22_pad_groupi_n_1045, csa_tree_add_101_22_pad_groupi_n_1046, csa_tree_add_101_22_pad_groupi_n_1047, csa_tree_add_101_22_pad_groupi_n_1048, csa_tree_add_101_22_pad_groupi_n_1049;
  wire csa_tree_add_101_22_pad_groupi_n_1050, csa_tree_add_101_22_pad_groupi_n_1051, csa_tree_add_101_22_pad_groupi_n_1052, csa_tree_add_101_22_pad_groupi_n_1053, csa_tree_add_101_22_pad_groupi_n_1054, csa_tree_add_101_22_pad_groupi_n_1055, csa_tree_add_101_22_pad_groupi_n_1056, csa_tree_add_101_22_pad_groupi_n_1057;
  wire csa_tree_add_101_22_pad_groupi_n_1058, csa_tree_add_101_22_pad_groupi_n_1059, csa_tree_add_101_22_pad_groupi_n_1060, csa_tree_add_101_22_pad_groupi_n_1061, csa_tree_add_101_22_pad_groupi_n_1062, csa_tree_add_101_22_pad_groupi_n_1063, csa_tree_add_101_22_pad_groupi_n_1064, csa_tree_add_101_22_pad_groupi_n_1065;
  wire csa_tree_add_101_22_pad_groupi_n_1066, csa_tree_add_101_22_pad_groupi_n_1067, csa_tree_add_101_22_pad_groupi_n_1068, csa_tree_add_101_22_pad_groupi_n_1069, csa_tree_add_101_22_pad_groupi_n_1070, csa_tree_add_101_22_pad_groupi_n_1071, csa_tree_add_101_22_pad_groupi_n_1072, csa_tree_add_101_22_pad_groupi_n_1073;
  wire csa_tree_add_101_22_pad_groupi_n_1074, csa_tree_add_101_22_pad_groupi_n_1075, csa_tree_add_101_22_pad_groupi_n_1076, csa_tree_add_101_22_pad_groupi_n_1077, csa_tree_add_101_22_pad_groupi_n_1078, csa_tree_add_101_22_pad_groupi_n_1079, csa_tree_add_101_22_pad_groupi_n_1080, csa_tree_add_101_22_pad_groupi_n_1081;
  wire csa_tree_add_101_22_pad_groupi_n_1082, csa_tree_add_101_22_pad_groupi_n_1083, csa_tree_add_101_22_pad_groupi_n_1084, csa_tree_add_101_22_pad_groupi_n_1085, csa_tree_add_101_22_pad_groupi_n_1086, csa_tree_add_101_22_pad_groupi_n_1087, csa_tree_add_101_22_pad_groupi_n_1088, csa_tree_add_101_22_pad_groupi_n_1089;
  wire csa_tree_add_101_22_pad_groupi_n_1090, csa_tree_add_101_22_pad_groupi_n_1091, csa_tree_add_101_22_pad_groupi_n_1092, csa_tree_add_101_22_pad_groupi_n_1093, csa_tree_add_101_22_pad_groupi_n_1094, csa_tree_add_101_22_pad_groupi_n_1095, csa_tree_add_101_22_pad_groupi_n_1096, csa_tree_add_101_22_pad_groupi_n_1097;
  wire csa_tree_add_101_22_pad_groupi_n_1098, csa_tree_add_101_22_pad_groupi_n_1099, csa_tree_add_101_22_pad_groupi_n_1100, csa_tree_add_101_22_pad_groupi_n_1101, csa_tree_add_101_22_pad_groupi_n_1102, csa_tree_add_101_22_pad_groupi_n_1103, csa_tree_add_101_22_pad_groupi_n_1104, csa_tree_add_101_22_pad_groupi_n_1105;
  wire csa_tree_add_101_22_pad_groupi_n_1106, csa_tree_add_101_22_pad_groupi_n_1107, csa_tree_add_101_22_pad_groupi_n_1108, csa_tree_add_101_22_pad_groupi_n_1109, csa_tree_add_101_22_pad_groupi_n_1110, csa_tree_add_101_22_pad_groupi_n_1111, csa_tree_add_101_22_pad_groupi_n_1112, csa_tree_add_101_22_pad_groupi_n_1113;
  wire csa_tree_add_101_22_pad_groupi_n_1114, csa_tree_add_101_22_pad_groupi_n_1115, csa_tree_add_101_22_pad_groupi_n_1116, csa_tree_add_101_22_pad_groupi_n_1117, csa_tree_add_101_22_pad_groupi_n_1118, csa_tree_add_101_22_pad_groupi_n_1119, csa_tree_add_101_22_pad_groupi_n_1120, csa_tree_add_101_22_pad_groupi_n_1121;
  wire csa_tree_add_101_22_pad_groupi_n_1122, csa_tree_add_101_22_pad_groupi_n_1123, csa_tree_add_101_22_pad_groupi_n_1124, csa_tree_add_101_22_pad_groupi_n_1125, csa_tree_add_101_22_pad_groupi_n_1126, csa_tree_add_101_22_pad_groupi_n_1127, csa_tree_add_101_22_pad_groupi_n_1128, csa_tree_add_101_22_pad_groupi_n_1129;
  wire csa_tree_add_101_22_pad_groupi_n_1130, csa_tree_add_101_22_pad_groupi_n_1131, csa_tree_add_101_22_pad_groupi_n_1132, csa_tree_add_101_22_pad_groupi_n_1133, csa_tree_add_101_22_pad_groupi_n_1134, csa_tree_add_101_22_pad_groupi_n_1135, csa_tree_add_101_22_pad_groupi_n_1136, csa_tree_add_101_22_pad_groupi_n_1137;
  wire csa_tree_add_101_22_pad_groupi_n_1138, csa_tree_add_101_22_pad_groupi_n_1139, csa_tree_add_101_22_pad_groupi_n_1140, csa_tree_add_101_22_pad_groupi_n_1141, csa_tree_add_101_22_pad_groupi_n_1142, csa_tree_add_101_22_pad_groupi_n_1143, csa_tree_add_101_22_pad_groupi_n_1144, csa_tree_add_101_22_pad_groupi_n_1145;
  wire csa_tree_add_101_22_pad_groupi_n_1146, csa_tree_add_101_22_pad_groupi_n_1147, csa_tree_add_101_22_pad_groupi_n_1148, csa_tree_add_101_22_pad_groupi_n_1149, csa_tree_add_101_22_pad_groupi_n_1150, csa_tree_add_101_22_pad_groupi_n_1151, csa_tree_add_101_22_pad_groupi_n_1152, csa_tree_add_101_22_pad_groupi_n_1153;
  wire csa_tree_add_101_22_pad_groupi_n_1154, csa_tree_add_101_22_pad_groupi_n_1155, csa_tree_add_101_22_pad_groupi_n_1156, csa_tree_add_101_22_pad_groupi_n_1157, csa_tree_add_101_22_pad_groupi_n_1158, csa_tree_add_101_22_pad_groupi_n_1159, csa_tree_add_101_22_pad_groupi_n_1160, csa_tree_add_101_22_pad_groupi_n_1161;
  wire csa_tree_add_101_22_pad_groupi_n_1162, csa_tree_add_101_22_pad_groupi_n_1163, csa_tree_add_101_22_pad_groupi_n_1164, csa_tree_add_101_22_pad_groupi_n_1165, csa_tree_add_101_22_pad_groupi_n_1166, csa_tree_add_101_22_pad_groupi_n_1167, csa_tree_add_101_22_pad_groupi_n_1168, csa_tree_add_101_22_pad_groupi_n_1169;
  wire csa_tree_add_101_22_pad_groupi_n_1170, csa_tree_add_101_22_pad_groupi_n_1171, csa_tree_add_101_22_pad_groupi_n_1172, csa_tree_add_101_22_pad_groupi_n_1173, csa_tree_add_101_22_pad_groupi_n_1174, csa_tree_add_101_22_pad_groupi_n_1175, csa_tree_add_101_22_pad_groupi_n_1176, csa_tree_add_101_22_pad_groupi_n_1177;
  wire csa_tree_add_101_22_pad_groupi_n_1178, csa_tree_add_101_22_pad_groupi_n_1179, csa_tree_add_101_22_pad_groupi_n_1180, csa_tree_add_101_22_pad_groupi_n_1181, csa_tree_add_101_22_pad_groupi_n_1182, csa_tree_add_101_22_pad_groupi_n_1183, csa_tree_add_101_22_pad_groupi_n_1184, csa_tree_add_101_22_pad_groupi_n_1185;
  wire csa_tree_add_101_22_pad_groupi_n_1186, csa_tree_add_101_22_pad_groupi_n_1187, csa_tree_add_101_22_pad_groupi_n_1188, csa_tree_add_101_22_pad_groupi_n_1189, csa_tree_add_101_22_pad_groupi_n_1190, csa_tree_add_101_22_pad_groupi_n_1191, csa_tree_add_101_22_pad_groupi_n_1192, csa_tree_add_101_22_pad_groupi_n_1193;
  wire csa_tree_add_101_22_pad_groupi_n_1194, csa_tree_add_101_22_pad_groupi_n_1195, csa_tree_add_101_22_pad_groupi_n_1196, csa_tree_add_101_22_pad_groupi_n_1197, csa_tree_add_101_22_pad_groupi_n_1198, csa_tree_add_101_22_pad_groupi_n_1199, csa_tree_add_101_22_pad_groupi_n_1200, csa_tree_add_101_22_pad_groupi_n_1201;
  wire csa_tree_add_101_22_pad_groupi_n_1202, csa_tree_add_101_22_pad_groupi_n_1203, csa_tree_add_101_22_pad_groupi_n_1204, csa_tree_add_101_22_pad_groupi_n_1205, csa_tree_add_101_22_pad_groupi_n_1206, csa_tree_add_101_22_pad_groupi_n_1207, csa_tree_add_101_22_pad_groupi_n_1208, csa_tree_add_101_22_pad_groupi_n_1209;
  wire csa_tree_add_101_22_pad_groupi_n_1210, csa_tree_add_101_22_pad_groupi_n_1211, csa_tree_add_101_22_pad_groupi_n_1212, csa_tree_add_101_22_pad_groupi_n_1213, csa_tree_add_101_22_pad_groupi_n_1214, csa_tree_add_101_22_pad_groupi_n_1215, csa_tree_add_101_22_pad_groupi_n_1216, csa_tree_add_101_22_pad_groupi_n_1217;
  wire csa_tree_add_101_22_pad_groupi_n_1218, csa_tree_add_101_22_pad_groupi_n_1219, csa_tree_add_101_22_pad_groupi_n_1220, csa_tree_add_101_22_pad_groupi_n_1221, csa_tree_add_101_22_pad_groupi_n_1222, csa_tree_add_101_22_pad_groupi_n_1223, csa_tree_add_101_22_pad_groupi_n_1224, csa_tree_add_101_22_pad_groupi_n_1225;
  wire csa_tree_add_101_22_pad_groupi_n_1226, csa_tree_add_101_22_pad_groupi_n_1227, csa_tree_add_101_22_pad_groupi_n_1228, csa_tree_add_101_22_pad_groupi_n_1229, csa_tree_add_101_22_pad_groupi_n_1230, csa_tree_add_101_22_pad_groupi_n_1231, csa_tree_add_101_22_pad_groupi_n_1232, csa_tree_add_101_22_pad_groupi_n_1233;
  wire csa_tree_add_101_22_pad_groupi_n_1234, csa_tree_add_101_22_pad_groupi_n_1235, csa_tree_add_101_22_pad_groupi_n_1236, csa_tree_add_101_22_pad_groupi_n_1237, csa_tree_add_101_22_pad_groupi_n_1238, csa_tree_add_101_22_pad_groupi_n_1239, csa_tree_add_101_22_pad_groupi_n_1240, csa_tree_add_101_22_pad_groupi_n_1241;
  wire csa_tree_add_101_22_pad_groupi_n_1242, csa_tree_add_101_22_pad_groupi_n_1243, csa_tree_add_101_22_pad_groupi_n_1244, csa_tree_add_101_22_pad_groupi_n_1245, csa_tree_add_101_22_pad_groupi_n_1246, csa_tree_add_101_22_pad_groupi_n_1247, csa_tree_add_101_22_pad_groupi_n_1248, csa_tree_add_101_22_pad_groupi_n_1249;
  wire csa_tree_add_101_22_pad_groupi_n_1250, csa_tree_add_101_22_pad_groupi_n_1251, csa_tree_add_101_22_pad_groupi_n_1252, csa_tree_add_101_22_pad_groupi_n_1253, csa_tree_add_101_22_pad_groupi_n_1254, csa_tree_add_101_22_pad_groupi_n_1255, csa_tree_add_101_22_pad_groupi_n_1256, csa_tree_add_101_22_pad_groupi_n_1257;
  wire csa_tree_add_101_22_pad_groupi_n_1258, csa_tree_add_101_22_pad_groupi_n_1259, csa_tree_add_101_22_pad_groupi_n_1260, csa_tree_add_101_22_pad_groupi_n_1261, csa_tree_add_101_22_pad_groupi_n_1262, csa_tree_add_101_22_pad_groupi_n_1263, csa_tree_add_101_22_pad_groupi_n_1264, csa_tree_add_101_22_pad_groupi_n_1265;
  wire csa_tree_add_101_22_pad_groupi_n_1266, csa_tree_add_101_22_pad_groupi_n_1267, csa_tree_add_101_22_pad_groupi_n_1268, csa_tree_add_101_22_pad_groupi_n_1269, csa_tree_add_101_22_pad_groupi_n_1270, csa_tree_add_101_22_pad_groupi_n_1271, csa_tree_add_101_22_pad_groupi_n_1272, csa_tree_add_101_22_pad_groupi_n_1273;
  wire csa_tree_add_101_22_pad_groupi_n_1274, csa_tree_add_101_22_pad_groupi_n_1275, csa_tree_add_101_22_pad_groupi_n_1276, csa_tree_add_101_22_pad_groupi_n_1277, csa_tree_add_101_22_pad_groupi_n_1278, csa_tree_add_101_22_pad_groupi_n_1279, csa_tree_add_101_22_pad_groupi_n_1280, csa_tree_add_101_22_pad_groupi_n_1281;
  wire csa_tree_add_101_22_pad_groupi_n_1282, csa_tree_add_101_22_pad_groupi_n_1283, csa_tree_add_101_22_pad_groupi_n_1284, csa_tree_add_101_22_pad_groupi_n_1285, csa_tree_add_101_22_pad_groupi_n_1286, csa_tree_add_101_22_pad_groupi_n_1287, csa_tree_add_101_22_pad_groupi_n_1288, csa_tree_add_101_22_pad_groupi_n_1289;
  wire csa_tree_add_101_22_pad_groupi_n_1290, csa_tree_add_101_22_pad_groupi_n_1291, csa_tree_add_101_22_pad_groupi_n_1292, csa_tree_add_101_22_pad_groupi_n_1293, csa_tree_add_101_22_pad_groupi_n_1294, csa_tree_add_101_22_pad_groupi_n_1295, csa_tree_add_101_22_pad_groupi_n_1296, csa_tree_add_101_22_pad_groupi_n_1297;
  wire csa_tree_add_101_22_pad_groupi_n_1298, csa_tree_add_101_22_pad_groupi_n_1299, csa_tree_add_101_22_pad_groupi_n_1300, csa_tree_add_101_22_pad_groupi_n_1301, csa_tree_add_101_22_pad_groupi_n_1302, csa_tree_add_101_22_pad_groupi_n_1303, csa_tree_add_101_22_pad_groupi_n_1304, csa_tree_add_101_22_pad_groupi_n_1305;
  wire csa_tree_add_101_22_pad_groupi_n_1306, csa_tree_add_101_22_pad_groupi_n_1307, csa_tree_add_101_22_pad_groupi_n_1308, csa_tree_add_101_22_pad_groupi_n_1309, csa_tree_add_101_22_pad_groupi_n_1310, csa_tree_add_101_22_pad_groupi_n_1311, csa_tree_add_101_22_pad_groupi_n_1312, csa_tree_add_101_22_pad_groupi_n_1313;
  wire csa_tree_add_101_22_pad_groupi_n_1314, csa_tree_add_101_22_pad_groupi_n_1315, csa_tree_add_101_22_pad_groupi_n_1316, csa_tree_add_101_22_pad_groupi_n_1317, csa_tree_add_101_22_pad_groupi_n_1318, csa_tree_add_101_22_pad_groupi_n_1319, csa_tree_add_101_22_pad_groupi_n_1320, csa_tree_add_101_22_pad_groupi_n_1321;
  wire csa_tree_add_101_22_pad_groupi_n_1322, csa_tree_add_101_22_pad_groupi_n_1323, csa_tree_add_101_22_pad_groupi_n_1324, csa_tree_add_101_22_pad_groupi_n_1325, csa_tree_add_101_22_pad_groupi_n_1326, csa_tree_add_101_22_pad_groupi_n_1327, csa_tree_add_101_22_pad_groupi_n_1328, csa_tree_add_101_22_pad_groupi_n_1329;
  wire csa_tree_add_101_22_pad_groupi_n_1330, csa_tree_add_101_22_pad_groupi_n_1331, csa_tree_add_101_22_pad_groupi_n_1332, csa_tree_add_101_22_pad_groupi_n_1333, csa_tree_add_101_22_pad_groupi_n_1334, csa_tree_add_101_22_pad_groupi_n_1335, csa_tree_add_101_22_pad_groupi_n_1336, csa_tree_add_101_22_pad_groupi_n_1337;
  wire csa_tree_add_101_22_pad_groupi_n_1338, csa_tree_add_101_22_pad_groupi_n_1339, csa_tree_add_101_22_pad_groupi_n_1340, csa_tree_add_101_22_pad_groupi_n_1341, csa_tree_add_101_22_pad_groupi_n_1342, csa_tree_add_101_22_pad_groupi_n_1343, csa_tree_add_101_22_pad_groupi_n_1344, csa_tree_add_101_22_pad_groupi_n_1345;
  wire csa_tree_add_101_22_pad_groupi_n_1346, csa_tree_add_101_22_pad_groupi_n_1347, csa_tree_add_101_22_pad_groupi_n_1348, csa_tree_add_101_22_pad_groupi_n_1349, csa_tree_add_101_22_pad_groupi_n_1350, csa_tree_add_101_22_pad_groupi_n_1351, csa_tree_add_101_22_pad_groupi_n_1352, csa_tree_add_101_22_pad_groupi_n_1353;
  wire csa_tree_add_101_22_pad_groupi_n_1354, csa_tree_add_101_22_pad_groupi_n_1355, csa_tree_add_101_22_pad_groupi_n_1356, csa_tree_add_101_22_pad_groupi_n_1357, csa_tree_add_101_22_pad_groupi_n_1358, csa_tree_add_101_22_pad_groupi_n_1359, csa_tree_add_101_22_pad_groupi_n_1360, csa_tree_add_101_22_pad_groupi_n_1361;
  wire csa_tree_add_101_22_pad_groupi_n_1362, csa_tree_add_101_22_pad_groupi_n_1363, csa_tree_add_101_22_pad_groupi_n_1364, csa_tree_add_101_22_pad_groupi_n_1365, csa_tree_add_101_22_pad_groupi_n_1366, csa_tree_add_101_22_pad_groupi_n_1367, csa_tree_add_101_22_pad_groupi_n_1368, csa_tree_add_101_22_pad_groupi_n_1369;
  wire csa_tree_add_101_22_pad_groupi_n_1370, csa_tree_add_101_22_pad_groupi_n_1371, csa_tree_add_101_22_pad_groupi_n_1372, csa_tree_add_101_22_pad_groupi_n_1373, csa_tree_add_101_22_pad_groupi_n_1374, csa_tree_add_101_22_pad_groupi_n_1375, csa_tree_add_101_22_pad_groupi_n_1376, csa_tree_add_101_22_pad_groupi_n_1377;
  wire csa_tree_add_101_22_pad_groupi_n_1378, csa_tree_add_101_22_pad_groupi_n_1379, csa_tree_add_101_22_pad_groupi_n_1380, csa_tree_add_101_22_pad_groupi_n_1381, csa_tree_add_101_22_pad_groupi_n_1382, csa_tree_add_101_22_pad_groupi_n_1383, csa_tree_add_101_22_pad_groupi_n_1384, csa_tree_add_101_22_pad_groupi_n_1385;
  wire csa_tree_add_101_22_pad_groupi_n_1386, csa_tree_add_101_22_pad_groupi_n_1387, csa_tree_add_101_22_pad_groupi_n_1388, csa_tree_add_101_22_pad_groupi_n_1389, csa_tree_add_101_22_pad_groupi_n_1390, csa_tree_add_101_22_pad_groupi_n_1391, csa_tree_add_101_22_pad_groupi_n_1392, csa_tree_add_101_22_pad_groupi_n_1393;
  wire csa_tree_add_101_22_pad_groupi_n_1394, csa_tree_add_101_22_pad_groupi_n_1395, csa_tree_add_101_22_pad_groupi_n_1396, csa_tree_add_101_22_pad_groupi_n_1397, csa_tree_add_101_22_pad_groupi_n_1398, csa_tree_add_101_22_pad_groupi_n_1399, csa_tree_add_101_22_pad_groupi_n_1400, csa_tree_add_101_22_pad_groupi_n_1401;
  wire csa_tree_add_101_22_pad_groupi_n_1402, csa_tree_add_101_22_pad_groupi_n_1403, csa_tree_add_101_22_pad_groupi_n_1404, csa_tree_add_101_22_pad_groupi_n_1405, csa_tree_add_101_22_pad_groupi_n_1406, csa_tree_add_101_22_pad_groupi_n_1407, csa_tree_add_101_22_pad_groupi_n_1408, csa_tree_add_101_22_pad_groupi_n_1409;
  wire csa_tree_add_101_22_pad_groupi_n_1410, csa_tree_add_101_22_pad_groupi_n_1411, csa_tree_add_101_22_pad_groupi_n_1412, csa_tree_add_101_22_pad_groupi_n_1413, csa_tree_add_101_22_pad_groupi_n_1414, csa_tree_add_101_22_pad_groupi_n_1415, csa_tree_add_101_22_pad_groupi_n_1416, csa_tree_add_101_22_pad_groupi_n_1417;
  wire csa_tree_add_101_22_pad_groupi_n_1418, csa_tree_add_101_22_pad_groupi_n_1419, csa_tree_add_101_22_pad_groupi_n_1420, csa_tree_add_101_22_pad_groupi_n_1421, csa_tree_add_101_22_pad_groupi_n_1422, csa_tree_add_101_22_pad_groupi_n_1423, csa_tree_add_101_22_pad_groupi_n_1424, csa_tree_add_101_22_pad_groupi_n_1425;
  wire csa_tree_add_101_22_pad_groupi_n_1426, csa_tree_add_101_22_pad_groupi_n_1427, csa_tree_add_101_22_pad_groupi_n_1428, csa_tree_add_101_22_pad_groupi_n_1429, csa_tree_add_101_22_pad_groupi_n_1430, csa_tree_add_101_22_pad_groupi_n_1431, csa_tree_add_101_22_pad_groupi_n_1432, csa_tree_add_101_22_pad_groupi_n_1433;
  wire csa_tree_add_101_22_pad_groupi_n_1434, csa_tree_add_101_22_pad_groupi_n_1435, csa_tree_add_101_22_pad_groupi_n_1436, csa_tree_add_101_22_pad_groupi_n_1437, csa_tree_add_101_22_pad_groupi_n_1438, csa_tree_add_101_22_pad_groupi_n_1439, csa_tree_add_101_22_pad_groupi_n_1440, csa_tree_add_101_22_pad_groupi_n_1441;
  wire csa_tree_add_101_22_pad_groupi_n_1442, csa_tree_add_101_22_pad_groupi_n_1443, csa_tree_add_101_22_pad_groupi_n_1444, csa_tree_add_101_22_pad_groupi_n_1445, csa_tree_add_101_22_pad_groupi_n_1446, csa_tree_add_101_22_pad_groupi_n_1447, csa_tree_add_101_22_pad_groupi_n_1448, csa_tree_add_101_22_pad_groupi_n_1449;
  wire csa_tree_add_101_22_pad_groupi_n_1450, csa_tree_add_101_22_pad_groupi_n_1451, csa_tree_add_101_22_pad_groupi_n_1452, csa_tree_add_101_22_pad_groupi_n_1453, csa_tree_add_101_22_pad_groupi_n_1454, csa_tree_add_101_22_pad_groupi_n_1455, csa_tree_add_101_22_pad_groupi_n_1456, csa_tree_add_101_22_pad_groupi_n_1457;
  wire csa_tree_add_101_22_pad_groupi_n_1458, csa_tree_add_101_22_pad_groupi_n_1459, csa_tree_add_101_22_pad_groupi_n_1460, csa_tree_add_101_22_pad_groupi_n_1461, csa_tree_add_101_22_pad_groupi_n_1462, csa_tree_add_101_22_pad_groupi_n_1463, csa_tree_add_101_22_pad_groupi_n_1464, csa_tree_add_101_22_pad_groupi_n_1465;
  wire csa_tree_add_101_22_pad_groupi_n_1466, csa_tree_add_101_22_pad_groupi_n_1467, csa_tree_add_101_22_pad_groupi_n_1468, csa_tree_add_101_22_pad_groupi_n_1469, csa_tree_add_101_22_pad_groupi_n_1470, csa_tree_add_101_22_pad_groupi_n_1471, csa_tree_add_101_22_pad_groupi_n_1472, csa_tree_add_101_22_pad_groupi_n_1473;
  wire csa_tree_add_101_22_pad_groupi_n_1474, csa_tree_add_101_22_pad_groupi_n_1475, csa_tree_add_101_22_pad_groupi_n_1476, csa_tree_add_101_22_pad_groupi_n_1477, csa_tree_add_101_22_pad_groupi_n_1478, csa_tree_add_101_22_pad_groupi_n_1479, csa_tree_add_101_22_pad_groupi_n_1480, csa_tree_add_101_22_pad_groupi_n_1481;
  wire csa_tree_add_101_22_pad_groupi_n_1482, csa_tree_add_101_22_pad_groupi_n_1483, csa_tree_add_101_22_pad_groupi_n_1484, csa_tree_add_101_22_pad_groupi_n_1485, csa_tree_add_101_22_pad_groupi_n_1486, csa_tree_add_101_22_pad_groupi_n_1487, csa_tree_add_101_22_pad_groupi_n_1488, csa_tree_add_101_22_pad_groupi_n_1489;
  wire csa_tree_add_101_22_pad_groupi_n_1490, csa_tree_add_101_22_pad_groupi_n_1491, csa_tree_add_101_22_pad_groupi_n_1492, csa_tree_add_101_22_pad_groupi_n_1493, csa_tree_add_101_22_pad_groupi_n_1494, csa_tree_add_101_22_pad_groupi_n_1495, csa_tree_add_101_22_pad_groupi_n_1496, csa_tree_add_101_22_pad_groupi_n_1497;
  wire csa_tree_add_101_22_pad_groupi_n_1498, csa_tree_add_101_22_pad_groupi_n_1499, csa_tree_add_101_22_pad_groupi_n_1500, csa_tree_add_101_22_pad_groupi_n_1501, csa_tree_add_101_22_pad_groupi_n_1502, csa_tree_add_101_22_pad_groupi_n_1503, csa_tree_add_101_22_pad_groupi_n_1505, csa_tree_add_101_22_pad_groupi_n_1506;
  wire csa_tree_add_101_22_pad_groupi_n_1507, csa_tree_add_101_22_pad_groupi_n_1508, csa_tree_add_101_22_pad_groupi_n_1509, csa_tree_add_101_22_pad_groupi_n_1510, csa_tree_add_101_22_pad_groupi_n_1511, csa_tree_add_101_22_pad_groupi_n_1512, csa_tree_add_101_22_pad_groupi_n_1513, csa_tree_add_101_22_pad_groupi_n_1514;
  wire csa_tree_add_101_22_pad_groupi_n_1515, csa_tree_add_101_22_pad_groupi_n_1516, csa_tree_add_101_22_pad_groupi_n_1517, csa_tree_add_101_22_pad_groupi_n_1518, csa_tree_add_101_22_pad_groupi_n_1519, csa_tree_add_101_22_pad_groupi_n_1520, csa_tree_add_101_22_pad_groupi_n_1521, csa_tree_add_101_22_pad_groupi_n_1522;
  wire csa_tree_add_101_22_pad_groupi_n_1523, csa_tree_add_101_22_pad_groupi_n_1524, csa_tree_add_101_22_pad_groupi_n_1525, csa_tree_add_101_22_pad_groupi_n_1526, csa_tree_add_101_22_pad_groupi_n_1527, csa_tree_add_101_22_pad_groupi_n_1529, csa_tree_add_101_22_pad_groupi_n_1530, csa_tree_add_101_22_pad_groupi_n_1532;
  wire csa_tree_add_101_22_pad_groupi_n_1533, csa_tree_add_101_22_pad_groupi_n_1534, csa_tree_add_101_22_pad_groupi_n_1535, csa_tree_add_101_22_pad_groupi_n_1537, csa_tree_add_101_22_pad_groupi_n_1538, csa_tree_add_101_22_pad_groupi_n_1539, csa_tree_add_101_22_pad_groupi_n_1540, csa_tree_add_101_22_pad_groupi_n_1542;
  wire csa_tree_add_101_22_pad_groupi_n_1543, csa_tree_add_101_22_pad_groupi_n_1544, csa_tree_add_101_22_pad_groupi_n_1546, csa_tree_add_101_22_pad_groupi_n_1547, csa_tree_add_101_22_pad_groupi_n_1549, csa_tree_add_101_22_pad_groupi_n_1550, csa_tree_add_101_22_pad_groupi_n_1552, csa_tree_add_101_22_pad_groupi_n_1553;
  wire csa_tree_add_101_22_pad_groupi_n_1555, csa_tree_add_101_22_pad_groupi_n_1556, csa_tree_add_101_22_pad_groupi_n_1558, csa_tree_add_107_22_pad_groupi_n_0, csa_tree_add_107_22_pad_groupi_n_1, csa_tree_add_107_22_pad_groupi_n_3, csa_tree_add_107_22_pad_groupi_n_4, csa_tree_add_107_22_pad_groupi_n_5;
  wire csa_tree_add_107_22_pad_groupi_n_6, csa_tree_add_107_22_pad_groupi_n_12, csa_tree_add_107_22_pad_groupi_n_13, csa_tree_add_107_22_pad_groupi_n_14, csa_tree_add_107_22_pad_groupi_n_15, csa_tree_add_107_22_pad_groupi_n_16, csa_tree_add_107_22_pad_groupi_n_17, csa_tree_add_107_22_pad_groupi_n_18;
  wire csa_tree_add_107_22_pad_groupi_n_19, csa_tree_add_107_22_pad_groupi_n_20, csa_tree_add_107_22_pad_groupi_n_21, csa_tree_add_107_22_pad_groupi_n_22, csa_tree_add_107_22_pad_groupi_n_23, csa_tree_add_107_22_pad_groupi_n_24, csa_tree_add_107_22_pad_groupi_n_25, csa_tree_add_107_22_pad_groupi_n_26;
  wire csa_tree_add_107_22_pad_groupi_n_27, csa_tree_add_107_22_pad_groupi_n_28, csa_tree_add_107_22_pad_groupi_n_29, csa_tree_add_107_22_pad_groupi_n_30, csa_tree_add_107_22_pad_groupi_n_31, csa_tree_add_107_22_pad_groupi_n_32, csa_tree_add_107_22_pad_groupi_n_33, csa_tree_add_107_22_pad_groupi_n_34;
  wire csa_tree_add_107_22_pad_groupi_n_35, csa_tree_add_107_22_pad_groupi_n_36, csa_tree_add_107_22_pad_groupi_n_37, csa_tree_add_107_22_pad_groupi_n_38, csa_tree_add_107_22_pad_groupi_n_39, csa_tree_add_107_22_pad_groupi_n_40, csa_tree_add_107_22_pad_groupi_n_41, csa_tree_add_107_22_pad_groupi_n_42;
  wire csa_tree_add_107_22_pad_groupi_n_43, csa_tree_add_107_22_pad_groupi_n_45, csa_tree_add_107_22_pad_groupi_n_46, csa_tree_add_107_22_pad_groupi_n_47, csa_tree_add_107_22_pad_groupi_n_48, csa_tree_add_107_22_pad_groupi_n_50, csa_tree_add_107_22_pad_groupi_n_51, csa_tree_add_107_22_pad_groupi_n_52;
  wire csa_tree_add_107_22_pad_groupi_n_53, csa_tree_add_107_22_pad_groupi_n_54, csa_tree_add_107_22_pad_groupi_n_55, csa_tree_add_107_22_pad_groupi_n_56, csa_tree_add_107_22_pad_groupi_n_57, csa_tree_add_107_22_pad_groupi_n_58, csa_tree_add_107_22_pad_groupi_n_59, csa_tree_add_107_22_pad_groupi_n_60;
  wire csa_tree_add_107_22_pad_groupi_n_61, csa_tree_add_107_22_pad_groupi_n_62, csa_tree_add_107_22_pad_groupi_n_64, csa_tree_add_107_22_pad_groupi_n_65, csa_tree_add_107_22_pad_groupi_n_66, csa_tree_add_107_22_pad_groupi_n_67, csa_tree_add_107_22_pad_groupi_n_68, csa_tree_add_107_22_pad_groupi_n_69;
  wire csa_tree_add_107_22_pad_groupi_n_70, csa_tree_add_107_22_pad_groupi_n_71, csa_tree_add_107_22_pad_groupi_n_72, csa_tree_add_107_22_pad_groupi_n_73, csa_tree_add_107_22_pad_groupi_n_74, csa_tree_add_107_22_pad_groupi_n_75, csa_tree_add_107_22_pad_groupi_n_76, csa_tree_add_107_22_pad_groupi_n_77;
  wire csa_tree_add_107_22_pad_groupi_n_78, csa_tree_add_107_22_pad_groupi_n_79, csa_tree_add_107_22_pad_groupi_n_80, csa_tree_add_107_22_pad_groupi_n_82, csa_tree_add_107_22_pad_groupi_n_83, csa_tree_add_107_22_pad_groupi_n_84, csa_tree_add_107_22_pad_groupi_n_85, csa_tree_add_107_22_pad_groupi_n_86;
  wire csa_tree_add_107_22_pad_groupi_n_87, csa_tree_add_107_22_pad_groupi_n_88, csa_tree_add_107_22_pad_groupi_n_89, csa_tree_add_107_22_pad_groupi_n_90, csa_tree_add_107_22_pad_groupi_n_91, csa_tree_add_107_22_pad_groupi_n_92, csa_tree_add_107_22_pad_groupi_n_93, csa_tree_add_107_22_pad_groupi_n_94;
  wire csa_tree_add_107_22_pad_groupi_n_95, csa_tree_add_107_22_pad_groupi_n_96, csa_tree_add_107_22_pad_groupi_n_97, csa_tree_add_107_22_pad_groupi_n_98, csa_tree_add_107_22_pad_groupi_n_99, csa_tree_add_107_22_pad_groupi_n_100, csa_tree_add_107_22_pad_groupi_n_101, csa_tree_add_107_22_pad_groupi_n_102;
  wire csa_tree_add_107_22_pad_groupi_n_103, csa_tree_add_107_22_pad_groupi_n_104, csa_tree_add_107_22_pad_groupi_n_105, csa_tree_add_107_22_pad_groupi_n_106, csa_tree_add_107_22_pad_groupi_n_107, csa_tree_add_107_22_pad_groupi_n_108, csa_tree_add_107_22_pad_groupi_n_109, csa_tree_add_107_22_pad_groupi_n_110;
  wire csa_tree_add_107_22_pad_groupi_n_111, csa_tree_add_107_22_pad_groupi_n_112, csa_tree_add_107_22_pad_groupi_n_113, csa_tree_add_107_22_pad_groupi_n_114, csa_tree_add_107_22_pad_groupi_n_115, csa_tree_add_107_22_pad_groupi_n_116, csa_tree_add_107_22_pad_groupi_n_117, csa_tree_add_107_22_pad_groupi_n_118;
  wire csa_tree_add_107_22_pad_groupi_n_119, csa_tree_add_107_22_pad_groupi_n_120, csa_tree_add_107_22_pad_groupi_n_121, csa_tree_add_107_22_pad_groupi_n_122, csa_tree_add_107_22_pad_groupi_n_123, csa_tree_add_107_22_pad_groupi_n_124, csa_tree_add_107_22_pad_groupi_n_125, csa_tree_add_107_22_pad_groupi_n_126;
  wire csa_tree_add_107_22_pad_groupi_n_127, csa_tree_add_107_22_pad_groupi_n_128, csa_tree_add_107_22_pad_groupi_n_129, csa_tree_add_107_22_pad_groupi_n_130, csa_tree_add_107_22_pad_groupi_n_131, csa_tree_add_107_22_pad_groupi_n_132, csa_tree_add_107_22_pad_groupi_n_133, csa_tree_add_107_22_pad_groupi_n_134;
  wire csa_tree_add_107_22_pad_groupi_n_135, csa_tree_add_107_22_pad_groupi_n_136, csa_tree_add_107_22_pad_groupi_n_137, csa_tree_add_107_22_pad_groupi_n_138, csa_tree_add_107_22_pad_groupi_n_139, csa_tree_add_107_22_pad_groupi_n_140, csa_tree_add_107_22_pad_groupi_n_141, csa_tree_add_107_22_pad_groupi_n_142;
  wire csa_tree_add_107_22_pad_groupi_n_143, csa_tree_add_107_22_pad_groupi_n_144, csa_tree_add_107_22_pad_groupi_n_145, csa_tree_add_107_22_pad_groupi_n_146, csa_tree_add_107_22_pad_groupi_n_147, csa_tree_add_107_22_pad_groupi_n_148, csa_tree_add_107_22_pad_groupi_n_149, csa_tree_add_107_22_pad_groupi_n_150;
  wire csa_tree_add_107_22_pad_groupi_n_151, csa_tree_add_107_22_pad_groupi_n_152, csa_tree_add_107_22_pad_groupi_n_153, csa_tree_add_107_22_pad_groupi_n_154, csa_tree_add_107_22_pad_groupi_n_155, csa_tree_add_107_22_pad_groupi_n_158, csa_tree_add_107_22_pad_groupi_n_159, csa_tree_add_107_22_pad_groupi_n_160;
  wire csa_tree_add_107_22_pad_groupi_n_161, csa_tree_add_107_22_pad_groupi_n_162, csa_tree_add_107_22_pad_groupi_n_163, csa_tree_add_107_22_pad_groupi_n_164, csa_tree_add_107_22_pad_groupi_n_165, csa_tree_add_107_22_pad_groupi_n_166, csa_tree_add_107_22_pad_groupi_n_167, csa_tree_add_107_22_pad_groupi_n_168;
  wire csa_tree_add_107_22_pad_groupi_n_169, csa_tree_add_107_22_pad_groupi_n_170, csa_tree_add_107_22_pad_groupi_n_171, csa_tree_add_107_22_pad_groupi_n_172, csa_tree_add_107_22_pad_groupi_n_173, csa_tree_add_107_22_pad_groupi_n_174, csa_tree_add_107_22_pad_groupi_n_175, csa_tree_add_107_22_pad_groupi_n_176;
  wire csa_tree_add_107_22_pad_groupi_n_177, csa_tree_add_107_22_pad_groupi_n_178, csa_tree_add_107_22_pad_groupi_n_179, csa_tree_add_107_22_pad_groupi_n_180, csa_tree_add_107_22_pad_groupi_n_181, csa_tree_add_107_22_pad_groupi_n_182, csa_tree_add_107_22_pad_groupi_n_183, csa_tree_add_107_22_pad_groupi_n_184;
  wire csa_tree_add_107_22_pad_groupi_n_185, csa_tree_add_107_22_pad_groupi_n_186, csa_tree_add_107_22_pad_groupi_n_187, csa_tree_add_107_22_pad_groupi_n_188, csa_tree_add_107_22_pad_groupi_n_189, csa_tree_add_107_22_pad_groupi_n_190, csa_tree_add_107_22_pad_groupi_n_191, csa_tree_add_107_22_pad_groupi_n_192;
  wire csa_tree_add_107_22_pad_groupi_n_193, csa_tree_add_107_22_pad_groupi_n_194, csa_tree_add_107_22_pad_groupi_n_195, csa_tree_add_107_22_pad_groupi_n_196, csa_tree_add_107_22_pad_groupi_n_197, csa_tree_add_107_22_pad_groupi_n_198, csa_tree_add_107_22_pad_groupi_n_200, csa_tree_add_107_22_pad_groupi_n_201;
  wire csa_tree_add_107_22_pad_groupi_n_202, csa_tree_add_107_22_pad_groupi_n_203, csa_tree_add_107_22_pad_groupi_n_204, csa_tree_add_107_22_pad_groupi_n_205, csa_tree_add_107_22_pad_groupi_n_206, csa_tree_add_107_22_pad_groupi_n_207, csa_tree_add_107_22_pad_groupi_n_208, csa_tree_add_107_22_pad_groupi_n_209;
  wire csa_tree_add_107_22_pad_groupi_n_210, csa_tree_add_107_22_pad_groupi_n_211, csa_tree_add_107_22_pad_groupi_n_212, csa_tree_add_107_22_pad_groupi_n_213, csa_tree_add_107_22_pad_groupi_n_214, csa_tree_add_107_22_pad_groupi_n_215, csa_tree_add_107_22_pad_groupi_n_216, csa_tree_add_107_22_pad_groupi_n_217;
  wire csa_tree_add_107_22_pad_groupi_n_218, csa_tree_add_107_22_pad_groupi_n_219, csa_tree_add_107_22_pad_groupi_n_220, csa_tree_add_107_22_pad_groupi_n_221, csa_tree_add_107_22_pad_groupi_n_222, csa_tree_add_107_22_pad_groupi_n_223, csa_tree_add_107_22_pad_groupi_n_224, csa_tree_add_107_22_pad_groupi_n_225;
  wire csa_tree_add_107_22_pad_groupi_n_226, csa_tree_add_107_22_pad_groupi_n_227, csa_tree_add_107_22_pad_groupi_n_228, csa_tree_add_107_22_pad_groupi_n_229, csa_tree_add_107_22_pad_groupi_n_230, csa_tree_add_107_22_pad_groupi_n_231, csa_tree_add_107_22_pad_groupi_n_232, csa_tree_add_107_22_pad_groupi_n_233;
  wire csa_tree_add_107_22_pad_groupi_n_234, csa_tree_add_107_22_pad_groupi_n_235, csa_tree_add_107_22_pad_groupi_n_236, csa_tree_add_107_22_pad_groupi_n_237, csa_tree_add_107_22_pad_groupi_n_238, csa_tree_add_107_22_pad_groupi_n_239, csa_tree_add_107_22_pad_groupi_n_240, csa_tree_add_107_22_pad_groupi_n_241;
  wire csa_tree_add_107_22_pad_groupi_n_242, csa_tree_add_107_22_pad_groupi_n_243, csa_tree_add_107_22_pad_groupi_n_244, csa_tree_add_107_22_pad_groupi_n_245, csa_tree_add_107_22_pad_groupi_n_246, csa_tree_add_107_22_pad_groupi_n_247, csa_tree_add_107_22_pad_groupi_n_248, csa_tree_add_107_22_pad_groupi_n_249;
  wire csa_tree_add_107_22_pad_groupi_n_250, csa_tree_add_107_22_pad_groupi_n_251, csa_tree_add_107_22_pad_groupi_n_252, csa_tree_add_107_22_pad_groupi_n_253, csa_tree_add_107_22_pad_groupi_n_254, csa_tree_add_107_22_pad_groupi_n_255, csa_tree_add_107_22_pad_groupi_n_256, csa_tree_add_107_22_pad_groupi_n_257;
  wire csa_tree_add_107_22_pad_groupi_n_258, csa_tree_add_107_22_pad_groupi_n_259, csa_tree_add_107_22_pad_groupi_n_260, csa_tree_add_107_22_pad_groupi_n_261, csa_tree_add_107_22_pad_groupi_n_262, csa_tree_add_107_22_pad_groupi_n_263, csa_tree_add_107_22_pad_groupi_n_264, csa_tree_add_107_22_pad_groupi_n_265;
  wire csa_tree_add_107_22_pad_groupi_n_266, csa_tree_add_107_22_pad_groupi_n_267, csa_tree_add_107_22_pad_groupi_n_268, csa_tree_add_107_22_pad_groupi_n_269, csa_tree_add_107_22_pad_groupi_n_270, csa_tree_add_107_22_pad_groupi_n_271, csa_tree_add_107_22_pad_groupi_n_272, csa_tree_add_107_22_pad_groupi_n_273;
  wire csa_tree_add_107_22_pad_groupi_n_274, csa_tree_add_107_22_pad_groupi_n_275, csa_tree_add_107_22_pad_groupi_n_276, csa_tree_add_107_22_pad_groupi_n_277, csa_tree_add_107_22_pad_groupi_n_278, csa_tree_add_107_22_pad_groupi_n_279, csa_tree_add_107_22_pad_groupi_n_280, csa_tree_add_107_22_pad_groupi_n_281;
  wire csa_tree_add_107_22_pad_groupi_n_282, csa_tree_add_107_22_pad_groupi_n_283, csa_tree_add_107_22_pad_groupi_n_284, csa_tree_add_107_22_pad_groupi_n_285, csa_tree_add_107_22_pad_groupi_n_286, csa_tree_add_107_22_pad_groupi_n_287, csa_tree_add_107_22_pad_groupi_n_288, csa_tree_add_107_22_pad_groupi_n_289;
  wire csa_tree_add_107_22_pad_groupi_n_290, csa_tree_add_107_22_pad_groupi_n_291, csa_tree_add_107_22_pad_groupi_n_292, csa_tree_add_107_22_pad_groupi_n_293, csa_tree_add_107_22_pad_groupi_n_294, csa_tree_add_107_22_pad_groupi_n_295, csa_tree_add_107_22_pad_groupi_n_296, csa_tree_add_107_22_pad_groupi_n_297;
  wire csa_tree_add_107_22_pad_groupi_n_298, csa_tree_add_107_22_pad_groupi_n_299, csa_tree_add_107_22_pad_groupi_n_300, csa_tree_add_107_22_pad_groupi_n_301, csa_tree_add_107_22_pad_groupi_n_302, csa_tree_add_107_22_pad_groupi_n_303, csa_tree_add_107_22_pad_groupi_n_304, csa_tree_add_107_22_pad_groupi_n_305;
  wire csa_tree_add_107_22_pad_groupi_n_306, csa_tree_add_107_22_pad_groupi_n_307, csa_tree_add_107_22_pad_groupi_n_308, csa_tree_add_107_22_pad_groupi_n_309, csa_tree_add_107_22_pad_groupi_n_310, csa_tree_add_107_22_pad_groupi_n_311, csa_tree_add_107_22_pad_groupi_n_312, csa_tree_add_107_22_pad_groupi_n_313;
  wire csa_tree_add_107_22_pad_groupi_n_314, csa_tree_add_107_22_pad_groupi_n_315, csa_tree_add_107_22_pad_groupi_n_316, csa_tree_add_107_22_pad_groupi_n_317, csa_tree_add_107_22_pad_groupi_n_318, csa_tree_add_107_22_pad_groupi_n_319, csa_tree_add_107_22_pad_groupi_n_320, csa_tree_add_107_22_pad_groupi_n_321;
  wire csa_tree_add_107_22_pad_groupi_n_322, csa_tree_add_107_22_pad_groupi_n_323, csa_tree_add_107_22_pad_groupi_n_324, csa_tree_add_107_22_pad_groupi_n_325, csa_tree_add_107_22_pad_groupi_n_326, csa_tree_add_107_22_pad_groupi_n_327, csa_tree_add_107_22_pad_groupi_n_328, csa_tree_add_107_22_pad_groupi_n_329;
  wire csa_tree_add_107_22_pad_groupi_n_330, csa_tree_add_107_22_pad_groupi_n_331, csa_tree_add_107_22_pad_groupi_n_332, csa_tree_add_107_22_pad_groupi_n_333, csa_tree_add_107_22_pad_groupi_n_334, csa_tree_add_107_22_pad_groupi_n_335, csa_tree_add_107_22_pad_groupi_n_336, csa_tree_add_107_22_pad_groupi_n_337;
  wire csa_tree_add_107_22_pad_groupi_n_338, csa_tree_add_107_22_pad_groupi_n_339, csa_tree_add_107_22_pad_groupi_n_340, csa_tree_add_107_22_pad_groupi_n_341, csa_tree_add_107_22_pad_groupi_n_342, csa_tree_add_107_22_pad_groupi_n_343, csa_tree_add_107_22_pad_groupi_n_344, csa_tree_add_107_22_pad_groupi_n_345;
  wire csa_tree_add_107_22_pad_groupi_n_346, csa_tree_add_107_22_pad_groupi_n_347, csa_tree_add_107_22_pad_groupi_n_348, csa_tree_add_107_22_pad_groupi_n_349, csa_tree_add_107_22_pad_groupi_n_350, csa_tree_add_107_22_pad_groupi_n_351, csa_tree_add_107_22_pad_groupi_n_352, csa_tree_add_107_22_pad_groupi_n_353;
  wire csa_tree_add_107_22_pad_groupi_n_354, csa_tree_add_107_22_pad_groupi_n_355, csa_tree_add_107_22_pad_groupi_n_356, csa_tree_add_107_22_pad_groupi_n_357, csa_tree_add_107_22_pad_groupi_n_358, csa_tree_add_107_22_pad_groupi_n_359, csa_tree_add_107_22_pad_groupi_n_361, csa_tree_add_107_22_pad_groupi_n_362;
  wire csa_tree_add_107_22_pad_groupi_n_363, csa_tree_add_107_22_pad_groupi_n_364, csa_tree_add_107_22_pad_groupi_n_365, csa_tree_add_107_22_pad_groupi_n_366, csa_tree_add_107_22_pad_groupi_n_367, csa_tree_add_107_22_pad_groupi_n_368, csa_tree_add_107_22_pad_groupi_n_369, csa_tree_add_107_22_pad_groupi_n_370;
  wire csa_tree_add_107_22_pad_groupi_n_371, csa_tree_add_107_22_pad_groupi_n_372, csa_tree_add_107_22_pad_groupi_n_373, csa_tree_add_107_22_pad_groupi_n_374, csa_tree_add_107_22_pad_groupi_n_375, csa_tree_add_107_22_pad_groupi_n_376, csa_tree_add_107_22_pad_groupi_n_377, csa_tree_add_107_22_pad_groupi_n_378;
  wire csa_tree_add_107_22_pad_groupi_n_379, csa_tree_add_107_22_pad_groupi_n_380, csa_tree_add_107_22_pad_groupi_n_381, csa_tree_add_107_22_pad_groupi_n_382, csa_tree_add_107_22_pad_groupi_n_383, csa_tree_add_107_22_pad_groupi_n_384, csa_tree_add_107_22_pad_groupi_n_385, csa_tree_add_107_22_pad_groupi_n_386;
  wire csa_tree_add_107_22_pad_groupi_n_387, csa_tree_add_107_22_pad_groupi_n_388, csa_tree_add_107_22_pad_groupi_n_389, csa_tree_add_107_22_pad_groupi_n_390, csa_tree_add_107_22_pad_groupi_n_391, csa_tree_add_107_22_pad_groupi_n_392, csa_tree_add_107_22_pad_groupi_n_393, csa_tree_add_107_22_pad_groupi_n_394;
  wire csa_tree_add_107_22_pad_groupi_n_395, csa_tree_add_107_22_pad_groupi_n_396, csa_tree_add_107_22_pad_groupi_n_397, csa_tree_add_107_22_pad_groupi_n_398, csa_tree_add_107_22_pad_groupi_n_399, csa_tree_add_107_22_pad_groupi_n_401, csa_tree_add_107_22_pad_groupi_n_402, csa_tree_add_107_22_pad_groupi_n_403;
  wire csa_tree_add_107_22_pad_groupi_n_404, csa_tree_add_107_22_pad_groupi_n_406, csa_tree_add_107_22_pad_groupi_n_409, csa_tree_add_107_22_pad_groupi_n_410, csa_tree_add_107_22_pad_groupi_n_411, csa_tree_add_107_22_pad_groupi_n_412, csa_tree_add_107_22_pad_groupi_n_413, csa_tree_add_107_22_pad_groupi_n_414;
  wire csa_tree_add_107_22_pad_groupi_n_415, csa_tree_add_107_22_pad_groupi_n_416, csa_tree_add_107_22_pad_groupi_n_417, csa_tree_add_107_22_pad_groupi_n_418, csa_tree_add_107_22_pad_groupi_n_419, csa_tree_add_107_22_pad_groupi_n_420, csa_tree_add_107_22_pad_groupi_n_421, csa_tree_add_107_22_pad_groupi_n_422;
  wire csa_tree_add_107_22_pad_groupi_n_423, csa_tree_add_107_22_pad_groupi_n_424, csa_tree_add_107_22_pad_groupi_n_425, csa_tree_add_107_22_pad_groupi_n_426, csa_tree_add_107_22_pad_groupi_n_427, csa_tree_add_107_22_pad_groupi_n_428, csa_tree_add_107_22_pad_groupi_n_429, csa_tree_add_107_22_pad_groupi_n_430;
  wire csa_tree_add_107_22_pad_groupi_n_431, csa_tree_add_107_22_pad_groupi_n_432, csa_tree_add_107_22_pad_groupi_n_433, csa_tree_add_107_22_pad_groupi_n_434, csa_tree_add_107_22_pad_groupi_n_435, csa_tree_add_107_22_pad_groupi_n_438, csa_tree_add_107_22_pad_groupi_n_439, csa_tree_add_107_22_pad_groupi_n_445;
  wire csa_tree_add_107_22_pad_groupi_n_455, csa_tree_add_107_22_pad_groupi_n_456, csa_tree_add_107_22_pad_groupi_n_457, csa_tree_add_107_22_pad_groupi_n_458, csa_tree_add_107_22_pad_groupi_n_459, csa_tree_add_107_22_pad_groupi_n_460, csa_tree_add_107_22_pad_groupi_n_461, csa_tree_add_107_22_pad_groupi_n_462;
  wire csa_tree_add_107_22_pad_groupi_n_463, csa_tree_add_107_22_pad_groupi_n_464, csa_tree_add_107_22_pad_groupi_n_465, csa_tree_add_107_22_pad_groupi_n_466, csa_tree_add_107_22_pad_groupi_n_467, csa_tree_add_107_22_pad_groupi_n_468, csa_tree_add_107_22_pad_groupi_n_469, csa_tree_add_107_22_pad_groupi_n_470;
  wire csa_tree_add_107_22_pad_groupi_n_471, csa_tree_add_107_22_pad_groupi_n_472, csa_tree_add_107_22_pad_groupi_n_473, csa_tree_add_107_22_pad_groupi_n_474, csa_tree_add_107_22_pad_groupi_n_475, csa_tree_add_107_22_pad_groupi_n_476, csa_tree_add_107_22_pad_groupi_n_477, csa_tree_add_107_22_pad_groupi_n_478;
  wire csa_tree_add_107_22_pad_groupi_n_479, csa_tree_add_107_22_pad_groupi_n_480, csa_tree_add_107_22_pad_groupi_n_481, csa_tree_add_107_22_pad_groupi_n_482, csa_tree_add_107_22_pad_groupi_n_483, csa_tree_add_107_22_pad_groupi_n_484, csa_tree_add_107_22_pad_groupi_n_485, csa_tree_add_107_22_pad_groupi_n_486;
  wire csa_tree_add_107_22_pad_groupi_n_487, csa_tree_add_107_22_pad_groupi_n_488, csa_tree_add_107_22_pad_groupi_n_489, csa_tree_add_107_22_pad_groupi_n_490, csa_tree_add_107_22_pad_groupi_n_491, csa_tree_add_107_22_pad_groupi_n_492, csa_tree_add_107_22_pad_groupi_n_493, csa_tree_add_107_22_pad_groupi_n_494;
  wire csa_tree_add_107_22_pad_groupi_n_495, csa_tree_add_107_22_pad_groupi_n_496, csa_tree_add_107_22_pad_groupi_n_497, csa_tree_add_107_22_pad_groupi_n_498, csa_tree_add_107_22_pad_groupi_n_499, csa_tree_add_107_22_pad_groupi_n_500, csa_tree_add_107_22_pad_groupi_n_501, csa_tree_add_107_22_pad_groupi_n_502;
  wire csa_tree_add_107_22_pad_groupi_n_503, csa_tree_add_107_22_pad_groupi_n_504, csa_tree_add_107_22_pad_groupi_n_505, csa_tree_add_107_22_pad_groupi_n_506, csa_tree_add_107_22_pad_groupi_n_507, csa_tree_add_107_22_pad_groupi_n_508, csa_tree_add_107_22_pad_groupi_n_509, csa_tree_add_107_22_pad_groupi_n_510;
  wire csa_tree_add_107_22_pad_groupi_n_511, csa_tree_add_107_22_pad_groupi_n_512, csa_tree_add_107_22_pad_groupi_n_513, csa_tree_add_107_22_pad_groupi_n_514, csa_tree_add_107_22_pad_groupi_n_515, csa_tree_add_107_22_pad_groupi_n_516, csa_tree_add_107_22_pad_groupi_n_517, csa_tree_add_107_22_pad_groupi_n_518;
  wire csa_tree_add_107_22_pad_groupi_n_519, csa_tree_add_107_22_pad_groupi_n_520, csa_tree_add_107_22_pad_groupi_n_521, csa_tree_add_107_22_pad_groupi_n_522, csa_tree_add_107_22_pad_groupi_n_523, csa_tree_add_107_22_pad_groupi_n_524, csa_tree_add_107_22_pad_groupi_n_525, csa_tree_add_107_22_pad_groupi_n_526;
  wire csa_tree_add_107_22_pad_groupi_n_527, csa_tree_add_107_22_pad_groupi_n_528, csa_tree_add_107_22_pad_groupi_n_529, csa_tree_add_107_22_pad_groupi_n_530, csa_tree_add_107_22_pad_groupi_n_531, csa_tree_add_107_22_pad_groupi_n_532, csa_tree_add_107_22_pad_groupi_n_533, csa_tree_add_107_22_pad_groupi_n_534;
  wire csa_tree_add_107_22_pad_groupi_n_535, csa_tree_add_107_22_pad_groupi_n_536, csa_tree_add_107_22_pad_groupi_n_537, csa_tree_add_107_22_pad_groupi_n_538, csa_tree_add_107_22_pad_groupi_n_539, csa_tree_add_107_22_pad_groupi_n_540, csa_tree_add_107_22_pad_groupi_n_541, csa_tree_add_107_22_pad_groupi_n_542;
  wire csa_tree_add_107_22_pad_groupi_n_543, csa_tree_add_107_22_pad_groupi_n_544, csa_tree_add_107_22_pad_groupi_n_545, csa_tree_add_107_22_pad_groupi_n_546, csa_tree_add_107_22_pad_groupi_n_547, csa_tree_add_107_22_pad_groupi_n_548, csa_tree_add_107_22_pad_groupi_n_549, csa_tree_add_107_22_pad_groupi_n_550;
  wire csa_tree_add_107_22_pad_groupi_n_551, csa_tree_add_107_22_pad_groupi_n_552, csa_tree_add_107_22_pad_groupi_n_553, csa_tree_add_107_22_pad_groupi_n_554, csa_tree_add_107_22_pad_groupi_n_555, csa_tree_add_107_22_pad_groupi_n_556, csa_tree_add_107_22_pad_groupi_n_557, csa_tree_add_107_22_pad_groupi_n_559;
  wire csa_tree_add_107_22_pad_groupi_n_561, csa_tree_add_107_22_pad_groupi_n_562, csa_tree_add_107_22_pad_groupi_n_563, csa_tree_add_107_22_pad_groupi_n_564, csa_tree_add_107_22_pad_groupi_n_565, csa_tree_add_107_22_pad_groupi_n_566, csa_tree_add_107_22_pad_groupi_n_567, csa_tree_add_107_22_pad_groupi_n_568;
  wire csa_tree_add_107_22_pad_groupi_n_569, csa_tree_add_107_22_pad_groupi_n_570, csa_tree_add_107_22_pad_groupi_n_572, csa_tree_add_107_22_pad_groupi_n_573, csa_tree_add_107_22_pad_groupi_n_574, csa_tree_add_107_22_pad_groupi_n_575, csa_tree_add_107_22_pad_groupi_n_576, csa_tree_add_107_22_pad_groupi_n_577;
  wire csa_tree_add_107_22_pad_groupi_n_578, csa_tree_add_107_22_pad_groupi_n_579, csa_tree_add_107_22_pad_groupi_n_580, csa_tree_add_107_22_pad_groupi_n_581, csa_tree_add_107_22_pad_groupi_n_582, csa_tree_add_107_22_pad_groupi_n_583, csa_tree_add_107_22_pad_groupi_n_584, csa_tree_add_107_22_pad_groupi_n_586;
  wire csa_tree_add_107_22_pad_groupi_n_587, csa_tree_add_107_22_pad_groupi_n_588, csa_tree_add_107_22_pad_groupi_n_589, csa_tree_add_107_22_pad_groupi_n_590, csa_tree_add_107_22_pad_groupi_n_591, csa_tree_add_107_22_pad_groupi_n_592, csa_tree_add_107_22_pad_groupi_n_593, csa_tree_add_107_22_pad_groupi_n_594;
  wire csa_tree_add_107_22_pad_groupi_n_595, csa_tree_add_107_22_pad_groupi_n_598, csa_tree_add_107_22_pad_groupi_n_599, csa_tree_add_107_22_pad_groupi_n_600, csa_tree_add_107_22_pad_groupi_n_601, csa_tree_add_107_22_pad_groupi_n_602, csa_tree_add_107_22_pad_groupi_n_603, csa_tree_add_107_22_pad_groupi_n_604;
  wire csa_tree_add_107_22_pad_groupi_n_605, csa_tree_add_107_22_pad_groupi_n_606, csa_tree_add_107_22_pad_groupi_n_607, csa_tree_add_107_22_pad_groupi_n_608, csa_tree_add_107_22_pad_groupi_n_609, csa_tree_add_107_22_pad_groupi_n_610, csa_tree_add_107_22_pad_groupi_n_611, csa_tree_add_107_22_pad_groupi_n_612;
  wire csa_tree_add_107_22_pad_groupi_n_613, csa_tree_add_107_22_pad_groupi_n_614, csa_tree_add_107_22_pad_groupi_n_615, csa_tree_add_107_22_pad_groupi_n_616, csa_tree_add_107_22_pad_groupi_n_617, csa_tree_add_107_22_pad_groupi_n_618, csa_tree_add_107_22_pad_groupi_n_619, csa_tree_add_107_22_pad_groupi_n_620;
  wire csa_tree_add_107_22_pad_groupi_n_621, csa_tree_add_107_22_pad_groupi_n_622, csa_tree_add_107_22_pad_groupi_n_623, csa_tree_add_107_22_pad_groupi_n_624, csa_tree_add_107_22_pad_groupi_n_625, csa_tree_add_107_22_pad_groupi_n_626, csa_tree_add_107_22_pad_groupi_n_627, csa_tree_add_107_22_pad_groupi_n_628;
  wire csa_tree_add_107_22_pad_groupi_n_629, csa_tree_add_107_22_pad_groupi_n_630, csa_tree_add_107_22_pad_groupi_n_631, csa_tree_add_107_22_pad_groupi_n_633, csa_tree_add_107_22_pad_groupi_n_634, csa_tree_add_107_22_pad_groupi_n_635, csa_tree_add_107_22_pad_groupi_n_637, csa_tree_add_107_22_pad_groupi_n_638;
  wire csa_tree_add_107_22_pad_groupi_n_639, csa_tree_add_107_22_pad_groupi_n_640, csa_tree_add_107_22_pad_groupi_n_641, csa_tree_add_107_22_pad_groupi_n_642, csa_tree_add_107_22_pad_groupi_n_643, csa_tree_add_107_22_pad_groupi_n_644, csa_tree_add_107_22_pad_groupi_n_645, csa_tree_add_107_22_pad_groupi_n_646;
  wire csa_tree_add_107_22_pad_groupi_n_647, csa_tree_add_107_22_pad_groupi_n_648, csa_tree_add_107_22_pad_groupi_n_649, csa_tree_add_107_22_pad_groupi_n_650, csa_tree_add_107_22_pad_groupi_n_651, csa_tree_add_107_22_pad_groupi_n_652, csa_tree_add_107_22_pad_groupi_n_653, csa_tree_add_107_22_pad_groupi_n_654;
  wire csa_tree_add_107_22_pad_groupi_n_655, csa_tree_add_107_22_pad_groupi_n_656, csa_tree_add_107_22_pad_groupi_n_657, csa_tree_add_107_22_pad_groupi_n_658, csa_tree_add_107_22_pad_groupi_n_659, csa_tree_add_107_22_pad_groupi_n_660, csa_tree_add_107_22_pad_groupi_n_661, csa_tree_add_107_22_pad_groupi_n_662;
  wire csa_tree_add_107_22_pad_groupi_n_663, csa_tree_add_107_22_pad_groupi_n_664, csa_tree_add_107_22_pad_groupi_n_665, csa_tree_add_107_22_pad_groupi_n_666, csa_tree_add_107_22_pad_groupi_n_667, csa_tree_add_107_22_pad_groupi_n_668, csa_tree_add_107_22_pad_groupi_n_669, csa_tree_add_107_22_pad_groupi_n_670;
  wire csa_tree_add_107_22_pad_groupi_n_671, csa_tree_add_107_22_pad_groupi_n_672, csa_tree_add_107_22_pad_groupi_n_673, csa_tree_add_107_22_pad_groupi_n_674, csa_tree_add_107_22_pad_groupi_n_675, csa_tree_add_107_22_pad_groupi_n_676, csa_tree_add_107_22_pad_groupi_n_677, csa_tree_add_107_22_pad_groupi_n_678;
  wire csa_tree_add_107_22_pad_groupi_n_679, csa_tree_add_107_22_pad_groupi_n_680, csa_tree_add_107_22_pad_groupi_n_681, csa_tree_add_107_22_pad_groupi_n_682, csa_tree_add_107_22_pad_groupi_n_683, csa_tree_add_107_22_pad_groupi_n_684, csa_tree_add_107_22_pad_groupi_n_685, csa_tree_add_107_22_pad_groupi_n_686;
  wire csa_tree_add_107_22_pad_groupi_n_688, csa_tree_add_107_22_pad_groupi_n_689, csa_tree_add_107_22_pad_groupi_n_690, csa_tree_add_107_22_pad_groupi_n_691, csa_tree_add_107_22_pad_groupi_n_692, csa_tree_add_107_22_pad_groupi_n_693, csa_tree_add_107_22_pad_groupi_n_694, csa_tree_add_107_22_pad_groupi_n_695;
  wire csa_tree_add_107_22_pad_groupi_n_696, csa_tree_add_107_22_pad_groupi_n_697, csa_tree_add_107_22_pad_groupi_n_698, csa_tree_add_107_22_pad_groupi_n_699, csa_tree_add_107_22_pad_groupi_n_700, csa_tree_add_107_22_pad_groupi_n_702, csa_tree_add_107_22_pad_groupi_n_703, csa_tree_add_107_22_pad_groupi_n_704;
  wire csa_tree_add_107_22_pad_groupi_n_705, csa_tree_add_107_22_pad_groupi_n_706, csa_tree_add_107_22_pad_groupi_n_707, csa_tree_add_107_22_pad_groupi_n_708, csa_tree_add_107_22_pad_groupi_n_709, csa_tree_add_107_22_pad_groupi_n_710, csa_tree_add_107_22_pad_groupi_n_711, csa_tree_add_107_22_pad_groupi_n_712;
  wire csa_tree_add_107_22_pad_groupi_n_713, csa_tree_add_107_22_pad_groupi_n_714, csa_tree_add_107_22_pad_groupi_n_715, csa_tree_add_107_22_pad_groupi_n_716, csa_tree_add_107_22_pad_groupi_n_717, csa_tree_add_107_22_pad_groupi_n_718, csa_tree_add_107_22_pad_groupi_n_719, csa_tree_add_107_22_pad_groupi_n_720;
  wire csa_tree_add_107_22_pad_groupi_n_721, csa_tree_add_107_22_pad_groupi_n_722, csa_tree_add_107_22_pad_groupi_n_723, csa_tree_add_107_22_pad_groupi_n_724, csa_tree_add_107_22_pad_groupi_n_725, csa_tree_add_107_22_pad_groupi_n_726, csa_tree_add_107_22_pad_groupi_n_727, csa_tree_add_107_22_pad_groupi_n_728;
  wire csa_tree_add_107_22_pad_groupi_n_729, csa_tree_add_107_22_pad_groupi_n_730, csa_tree_add_107_22_pad_groupi_n_731, csa_tree_add_107_22_pad_groupi_n_732, csa_tree_add_107_22_pad_groupi_n_733, csa_tree_add_107_22_pad_groupi_n_734, csa_tree_add_107_22_pad_groupi_n_735, csa_tree_add_107_22_pad_groupi_n_736;
  wire csa_tree_add_107_22_pad_groupi_n_737, csa_tree_add_107_22_pad_groupi_n_738, csa_tree_add_107_22_pad_groupi_n_739, csa_tree_add_107_22_pad_groupi_n_740, csa_tree_add_107_22_pad_groupi_n_741, csa_tree_add_107_22_pad_groupi_n_742, csa_tree_add_107_22_pad_groupi_n_743, csa_tree_add_107_22_pad_groupi_n_744;
  wire csa_tree_add_107_22_pad_groupi_n_745, csa_tree_add_107_22_pad_groupi_n_746, csa_tree_add_107_22_pad_groupi_n_747, csa_tree_add_107_22_pad_groupi_n_748, csa_tree_add_107_22_pad_groupi_n_749, csa_tree_add_107_22_pad_groupi_n_750, csa_tree_add_107_22_pad_groupi_n_751, csa_tree_add_107_22_pad_groupi_n_752;
  wire csa_tree_add_107_22_pad_groupi_n_753, csa_tree_add_107_22_pad_groupi_n_754, csa_tree_add_107_22_pad_groupi_n_755, csa_tree_add_107_22_pad_groupi_n_756, csa_tree_add_107_22_pad_groupi_n_757, csa_tree_add_107_22_pad_groupi_n_758, csa_tree_add_107_22_pad_groupi_n_759, csa_tree_add_107_22_pad_groupi_n_760;
  wire csa_tree_add_107_22_pad_groupi_n_761, csa_tree_add_107_22_pad_groupi_n_762, csa_tree_add_107_22_pad_groupi_n_763, csa_tree_add_107_22_pad_groupi_n_764, csa_tree_add_107_22_pad_groupi_n_765, csa_tree_add_107_22_pad_groupi_n_766, csa_tree_add_107_22_pad_groupi_n_767, csa_tree_add_107_22_pad_groupi_n_768;
  wire csa_tree_add_107_22_pad_groupi_n_769, csa_tree_add_107_22_pad_groupi_n_770, csa_tree_add_107_22_pad_groupi_n_771, csa_tree_add_107_22_pad_groupi_n_772, csa_tree_add_107_22_pad_groupi_n_773, csa_tree_add_107_22_pad_groupi_n_774, csa_tree_add_107_22_pad_groupi_n_775, csa_tree_add_107_22_pad_groupi_n_776;
  wire csa_tree_add_107_22_pad_groupi_n_777, csa_tree_add_107_22_pad_groupi_n_778, csa_tree_add_107_22_pad_groupi_n_779, csa_tree_add_107_22_pad_groupi_n_780, csa_tree_add_107_22_pad_groupi_n_781, csa_tree_add_107_22_pad_groupi_n_782, csa_tree_add_107_22_pad_groupi_n_783, csa_tree_add_107_22_pad_groupi_n_784;
  wire csa_tree_add_107_22_pad_groupi_n_785, csa_tree_add_107_22_pad_groupi_n_786, csa_tree_add_107_22_pad_groupi_n_787, csa_tree_add_107_22_pad_groupi_n_788, csa_tree_add_107_22_pad_groupi_n_789, csa_tree_add_107_22_pad_groupi_n_790, csa_tree_add_107_22_pad_groupi_n_791, csa_tree_add_107_22_pad_groupi_n_792;
  wire csa_tree_add_107_22_pad_groupi_n_793, csa_tree_add_107_22_pad_groupi_n_794, csa_tree_add_107_22_pad_groupi_n_795, csa_tree_add_107_22_pad_groupi_n_796, csa_tree_add_107_22_pad_groupi_n_797, csa_tree_add_107_22_pad_groupi_n_798, csa_tree_add_107_22_pad_groupi_n_799, csa_tree_add_107_22_pad_groupi_n_800;
  wire csa_tree_add_107_22_pad_groupi_n_801, csa_tree_add_107_22_pad_groupi_n_802, csa_tree_add_107_22_pad_groupi_n_803, csa_tree_add_107_22_pad_groupi_n_804, csa_tree_add_107_22_pad_groupi_n_805, csa_tree_add_107_22_pad_groupi_n_806, csa_tree_add_107_22_pad_groupi_n_807, csa_tree_add_107_22_pad_groupi_n_808;
  wire csa_tree_add_107_22_pad_groupi_n_809, csa_tree_add_107_22_pad_groupi_n_810, csa_tree_add_107_22_pad_groupi_n_811, csa_tree_add_107_22_pad_groupi_n_812, csa_tree_add_107_22_pad_groupi_n_813, csa_tree_add_107_22_pad_groupi_n_814, csa_tree_add_107_22_pad_groupi_n_815, csa_tree_add_107_22_pad_groupi_n_816;
  wire csa_tree_add_107_22_pad_groupi_n_817, csa_tree_add_107_22_pad_groupi_n_818, csa_tree_add_107_22_pad_groupi_n_819, csa_tree_add_107_22_pad_groupi_n_820, csa_tree_add_107_22_pad_groupi_n_821, csa_tree_add_107_22_pad_groupi_n_822, csa_tree_add_107_22_pad_groupi_n_823, csa_tree_add_107_22_pad_groupi_n_824;
  wire csa_tree_add_107_22_pad_groupi_n_825, csa_tree_add_107_22_pad_groupi_n_826, csa_tree_add_107_22_pad_groupi_n_827, csa_tree_add_107_22_pad_groupi_n_828, csa_tree_add_107_22_pad_groupi_n_829, csa_tree_add_107_22_pad_groupi_n_830, csa_tree_add_107_22_pad_groupi_n_831, csa_tree_add_107_22_pad_groupi_n_832;
  wire csa_tree_add_107_22_pad_groupi_n_833, csa_tree_add_107_22_pad_groupi_n_834, csa_tree_add_107_22_pad_groupi_n_835, csa_tree_add_107_22_pad_groupi_n_836, csa_tree_add_107_22_pad_groupi_n_837, csa_tree_add_107_22_pad_groupi_n_838, csa_tree_add_107_22_pad_groupi_n_839, csa_tree_add_107_22_pad_groupi_n_840;
  wire csa_tree_add_107_22_pad_groupi_n_841, csa_tree_add_107_22_pad_groupi_n_842, csa_tree_add_107_22_pad_groupi_n_843, csa_tree_add_107_22_pad_groupi_n_844, csa_tree_add_107_22_pad_groupi_n_845, csa_tree_add_107_22_pad_groupi_n_846, csa_tree_add_107_22_pad_groupi_n_847, csa_tree_add_107_22_pad_groupi_n_848;
  wire csa_tree_add_107_22_pad_groupi_n_849, csa_tree_add_107_22_pad_groupi_n_851, csa_tree_add_107_22_pad_groupi_n_852, csa_tree_add_107_22_pad_groupi_n_853, csa_tree_add_107_22_pad_groupi_n_854, csa_tree_add_107_22_pad_groupi_n_855, csa_tree_add_107_22_pad_groupi_n_856, csa_tree_add_107_22_pad_groupi_n_857;
  wire csa_tree_add_107_22_pad_groupi_n_858, csa_tree_add_107_22_pad_groupi_n_859, csa_tree_add_107_22_pad_groupi_n_860, csa_tree_add_107_22_pad_groupi_n_861, csa_tree_add_107_22_pad_groupi_n_862, csa_tree_add_107_22_pad_groupi_n_863, csa_tree_add_107_22_pad_groupi_n_864, csa_tree_add_107_22_pad_groupi_n_865;
  wire csa_tree_add_107_22_pad_groupi_n_866, csa_tree_add_107_22_pad_groupi_n_867, csa_tree_add_107_22_pad_groupi_n_868, csa_tree_add_107_22_pad_groupi_n_869, csa_tree_add_107_22_pad_groupi_n_870, csa_tree_add_107_22_pad_groupi_n_871, csa_tree_add_107_22_pad_groupi_n_872, csa_tree_add_107_22_pad_groupi_n_873;
  wire csa_tree_add_107_22_pad_groupi_n_874, csa_tree_add_107_22_pad_groupi_n_875, csa_tree_add_107_22_pad_groupi_n_876, csa_tree_add_107_22_pad_groupi_n_877, csa_tree_add_107_22_pad_groupi_n_878, csa_tree_add_107_22_pad_groupi_n_879, csa_tree_add_107_22_pad_groupi_n_880, csa_tree_add_107_22_pad_groupi_n_881;
  wire csa_tree_add_107_22_pad_groupi_n_882, csa_tree_add_107_22_pad_groupi_n_883, csa_tree_add_107_22_pad_groupi_n_884, csa_tree_add_107_22_pad_groupi_n_885, csa_tree_add_107_22_pad_groupi_n_886, csa_tree_add_107_22_pad_groupi_n_887, csa_tree_add_107_22_pad_groupi_n_888, csa_tree_add_107_22_pad_groupi_n_889;
  wire csa_tree_add_107_22_pad_groupi_n_890, csa_tree_add_107_22_pad_groupi_n_891, csa_tree_add_107_22_pad_groupi_n_892, csa_tree_add_107_22_pad_groupi_n_893, csa_tree_add_107_22_pad_groupi_n_894, csa_tree_add_107_22_pad_groupi_n_895, csa_tree_add_107_22_pad_groupi_n_896, csa_tree_add_107_22_pad_groupi_n_897;
  wire csa_tree_add_107_22_pad_groupi_n_898, csa_tree_add_107_22_pad_groupi_n_899, csa_tree_add_107_22_pad_groupi_n_900, csa_tree_add_107_22_pad_groupi_n_901, csa_tree_add_107_22_pad_groupi_n_902, csa_tree_add_107_22_pad_groupi_n_903, csa_tree_add_107_22_pad_groupi_n_904, csa_tree_add_107_22_pad_groupi_n_905;
  wire csa_tree_add_107_22_pad_groupi_n_906, csa_tree_add_107_22_pad_groupi_n_907, csa_tree_add_107_22_pad_groupi_n_908, csa_tree_add_107_22_pad_groupi_n_909, csa_tree_add_107_22_pad_groupi_n_910, csa_tree_add_107_22_pad_groupi_n_911, csa_tree_add_107_22_pad_groupi_n_912, csa_tree_add_107_22_pad_groupi_n_913;
  wire csa_tree_add_107_22_pad_groupi_n_914, csa_tree_add_107_22_pad_groupi_n_915, csa_tree_add_107_22_pad_groupi_n_916, csa_tree_add_107_22_pad_groupi_n_917, csa_tree_add_107_22_pad_groupi_n_918, csa_tree_add_107_22_pad_groupi_n_919, csa_tree_add_107_22_pad_groupi_n_920, csa_tree_add_107_22_pad_groupi_n_921;
  wire csa_tree_add_107_22_pad_groupi_n_922, csa_tree_add_107_22_pad_groupi_n_923, csa_tree_add_107_22_pad_groupi_n_924, csa_tree_add_107_22_pad_groupi_n_925, csa_tree_add_107_22_pad_groupi_n_926, csa_tree_add_107_22_pad_groupi_n_927, csa_tree_add_107_22_pad_groupi_n_928, csa_tree_add_107_22_pad_groupi_n_929;
  wire csa_tree_add_107_22_pad_groupi_n_930, csa_tree_add_107_22_pad_groupi_n_931, csa_tree_add_107_22_pad_groupi_n_932, csa_tree_add_107_22_pad_groupi_n_933, csa_tree_add_107_22_pad_groupi_n_934, csa_tree_add_107_22_pad_groupi_n_935, csa_tree_add_107_22_pad_groupi_n_936, csa_tree_add_107_22_pad_groupi_n_937;
  wire csa_tree_add_107_22_pad_groupi_n_938, csa_tree_add_107_22_pad_groupi_n_939, csa_tree_add_107_22_pad_groupi_n_940, csa_tree_add_107_22_pad_groupi_n_941, csa_tree_add_107_22_pad_groupi_n_942, csa_tree_add_107_22_pad_groupi_n_943, csa_tree_add_107_22_pad_groupi_n_944, csa_tree_add_107_22_pad_groupi_n_945;
  wire csa_tree_add_107_22_pad_groupi_n_946, csa_tree_add_107_22_pad_groupi_n_947, csa_tree_add_107_22_pad_groupi_n_948, csa_tree_add_107_22_pad_groupi_n_949, csa_tree_add_107_22_pad_groupi_n_950, csa_tree_add_107_22_pad_groupi_n_951, csa_tree_add_107_22_pad_groupi_n_952, csa_tree_add_107_22_pad_groupi_n_953;
  wire csa_tree_add_107_22_pad_groupi_n_954, csa_tree_add_107_22_pad_groupi_n_955, csa_tree_add_107_22_pad_groupi_n_956, csa_tree_add_107_22_pad_groupi_n_957, csa_tree_add_107_22_pad_groupi_n_958, csa_tree_add_107_22_pad_groupi_n_959, csa_tree_add_107_22_pad_groupi_n_960, csa_tree_add_107_22_pad_groupi_n_961;
  wire csa_tree_add_107_22_pad_groupi_n_962, csa_tree_add_107_22_pad_groupi_n_963, csa_tree_add_107_22_pad_groupi_n_964, csa_tree_add_107_22_pad_groupi_n_965, csa_tree_add_107_22_pad_groupi_n_966, csa_tree_add_107_22_pad_groupi_n_967, csa_tree_add_107_22_pad_groupi_n_968, csa_tree_add_107_22_pad_groupi_n_969;
  wire csa_tree_add_107_22_pad_groupi_n_970, csa_tree_add_107_22_pad_groupi_n_971, csa_tree_add_107_22_pad_groupi_n_972, csa_tree_add_107_22_pad_groupi_n_973, csa_tree_add_107_22_pad_groupi_n_974, csa_tree_add_107_22_pad_groupi_n_975, csa_tree_add_107_22_pad_groupi_n_976, csa_tree_add_107_22_pad_groupi_n_977;
  wire csa_tree_add_107_22_pad_groupi_n_978, csa_tree_add_107_22_pad_groupi_n_979, csa_tree_add_107_22_pad_groupi_n_980, csa_tree_add_107_22_pad_groupi_n_981, csa_tree_add_107_22_pad_groupi_n_982, csa_tree_add_107_22_pad_groupi_n_983, csa_tree_add_107_22_pad_groupi_n_984, csa_tree_add_107_22_pad_groupi_n_985;
  wire csa_tree_add_107_22_pad_groupi_n_986, csa_tree_add_107_22_pad_groupi_n_987, csa_tree_add_107_22_pad_groupi_n_988, csa_tree_add_107_22_pad_groupi_n_989, csa_tree_add_107_22_pad_groupi_n_990, csa_tree_add_107_22_pad_groupi_n_991, csa_tree_add_107_22_pad_groupi_n_992, csa_tree_add_107_22_pad_groupi_n_993;
  wire csa_tree_add_107_22_pad_groupi_n_994, csa_tree_add_107_22_pad_groupi_n_995, csa_tree_add_107_22_pad_groupi_n_996, csa_tree_add_107_22_pad_groupi_n_997, csa_tree_add_107_22_pad_groupi_n_998, csa_tree_add_107_22_pad_groupi_n_999, csa_tree_add_107_22_pad_groupi_n_1000, csa_tree_add_107_22_pad_groupi_n_1001;
  wire csa_tree_add_107_22_pad_groupi_n_1002, csa_tree_add_107_22_pad_groupi_n_1003, csa_tree_add_107_22_pad_groupi_n_1004, csa_tree_add_107_22_pad_groupi_n_1005, csa_tree_add_107_22_pad_groupi_n_1006, csa_tree_add_107_22_pad_groupi_n_1007, csa_tree_add_107_22_pad_groupi_n_1008, csa_tree_add_107_22_pad_groupi_n_1009;
  wire csa_tree_add_107_22_pad_groupi_n_1010, csa_tree_add_107_22_pad_groupi_n_1011, csa_tree_add_107_22_pad_groupi_n_1012, csa_tree_add_107_22_pad_groupi_n_1013, csa_tree_add_107_22_pad_groupi_n_1014, csa_tree_add_107_22_pad_groupi_n_1015, csa_tree_add_107_22_pad_groupi_n_1016, csa_tree_add_107_22_pad_groupi_n_1017;
  wire csa_tree_add_107_22_pad_groupi_n_1018, csa_tree_add_107_22_pad_groupi_n_1019, csa_tree_add_107_22_pad_groupi_n_1020, csa_tree_add_107_22_pad_groupi_n_1021, csa_tree_add_107_22_pad_groupi_n_1022, csa_tree_add_107_22_pad_groupi_n_1023, csa_tree_add_107_22_pad_groupi_n_1024, csa_tree_add_107_22_pad_groupi_n_1025;
  wire csa_tree_add_107_22_pad_groupi_n_1026, csa_tree_add_107_22_pad_groupi_n_1027, csa_tree_add_107_22_pad_groupi_n_1028, csa_tree_add_107_22_pad_groupi_n_1029, csa_tree_add_107_22_pad_groupi_n_1030, csa_tree_add_107_22_pad_groupi_n_1031, csa_tree_add_107_22_pad_groupi_n_1032, csa_tree_add_107_22_pad_groupi_n_1033;
  wire csa_tree_add_107_22_pad_groupi_n_1034, csa_tree_add_107_22_pad_groupi_n_1035, csa_tree_add_107_22_pad_groupi_n_1036, csa_tree_add_107_22_pad_groupi_n_1037, csa_tree_add_107_22_pad_groupi_n_1038, csa_tree_add_107_22_pad_groupi_n_1039, csa_tree_add_107_22_pad_groupi_n_1040, csa_tree_add_107_22_pad_groupi_n_1041;
  wire csa_tree_add_107_22_pad_groupi_n_1042, csa_tree_add_107_22_pad_groupi_n_1043, csa_tree_add_107_22_pad_groupi_n_1044, csa_tree_add_107_22_pad_groupi_n_1045, csa_tree_add_107_22_pad_groupi_n_1046, csa_tree_add_107_22_pad_groupi_n_1047, csa_tree_add_107_22_pad_groupi_n_1048, csa_tree_add_107_22_pad_groupi_n_1049;
  wire csa_tree_add_107_22_pad_groupi_n_1050, csa_tree_add_107_22_pad_groupi_n_1051, csa_tree_add_107_22_pad_groupi_n_1052, csa_tree_add_107_22_pad_groupi_n_1053, csa_tree_add_107_22_pad_groupi_n_1054, csa_tree_add_107_22_pad_groupi_n_1055, csa_tree_add_107_22_pad_groupi_n_1056, csa_tree_add_107_22_pad_groupi_n_1057;
  wire csa_tree_add_107_22_pad_groupi_n_1058, csa_tree_add_107_22_pad_groupi_n_1059, csa_tree_add_107_22_pad_groupi_n_1060, csa_tree_add_107_22_pad_groupi_n_1061, csa_tree_add_107_22_pad_groupi_n_1062, csa_tree_add_107_22_pad_groupi_n_1063, csa_tree_add_107_22_pad_groupi_n_1064, csa_tree_add_107_22_pad_groupi_n_1065;
  wire csa_tree_add_107_22_pad_groupi_n_1066, csa_tree_add_107_22_pad_groupi_n_1067, csa_tree_add_107_22_pad_groupi_n_1068, csa_tree_add_107_22_pad_groupi_n_1069, csa_tree_add_107_22_pad_groupi_n_1070, csa_tree_add_107_22_pad_groupi_n_1071, csa_tree_add_107_22_pad_groupi_n_1072, csa_tree_add_107_22_pad_groupi_n_1073;
  wire csa_tree_add_107_22_pad_groupi_n_1074, csa_tree_add_107_22_pad_groupi_n_1075, csa_tree_add_107_22_pad_groupi_n_1076, csa_tree_add_107_22_pad_groupi_n_1077, csa_tree_add_107_22_pad_groupi_n_1078, csa_tree_add_107_22_pad_groupi_n_1079, csa_tree_add_107_22_pad_groupi_n_1080, csa_tree_add_107_22_pad_groupi_n_1081;
  wire csa_tree_add_107_22_pad_groupi_n_1082, csa_tree_add_107_22_pad_groupi_n_1083, csa_tree_add_107_22_pad_groupi_n_1084, csa_tree_add_107_22_pad_groupi_n_1085, csa_tree_add_107_22_pad_groupi_n_1086, csa_tree_add_107_22_pad_groupi_n_1087, csa_tree_add_107_22_pad_groupi_n_1088, csa_tree_add_107_22_pad_groupi_n_1089;
  wire csa_tree_add_107_22_pad_groupi_n_1090, csa_tree_add_107_22_pad_groupi_n_1091, csa_tree_add_107_22_pad_groupi_n_1092, csa_tree_add_107_22_pad_groupi_n_1093, csa_tree_add_107_22_pad_groupi_n_1094, csa_tree_add_107_22_pad_groupi_n_1095, csa_tree_add_107_22_pad_groupi_n_1096, csa_tree_add_107_22_pad_groupi_n_1097;
  wire csa_tree_add_107_22_pad_groupi_n_1098, csa_tree_add_107_22_pad_groupi_n_1099, csa_tree_add_107_22_pad_groupi_n_1100, csa_tree_add_107_22_pad_groupi_n_1101, csa_tree_add_107_22_pad_groupi_n_1102, csa_tree_add_107_22_pad_groupi_n_1103, csa_tree_add_107_22_pad_groupi_n_1104, csa_tree_add_107_22_pad_groupi_n_1105;
  wire csa_tree_add_107_22_pad_groupi_n_1106, csa_tree_add_107_22_pad_groupi_n_1107, csa_tree_add_107_22_pad_groupi_n_1108, csa_tree_add_107_22_pad_groupi_n_1109, csa_tree_add_107_22_pad_groupi_n_1110, csa_tree_add_107_22_pad_groupi_n_1111, csa_tree_add_107_22_pad_groupi_n_1112, csa_tree_add_107_22_pad_groupi_n_1113;
  wire csa_tree_add_107_22_pad_groupi_n_1114, csa_tree_add_107_22_pad_groupi_n_1115, csa_tree_add_107_22_pad_groupi_n_1116, csa_tree_add_107_22_pad_groupi_n_1117, csa_tree_add_107_22_pad_groupi_n_1118, csa_tree_add_107_22_pad_groupi_n_1119, csa_tree_add_107_22_pad_groupi_n_1120, csa_tree_add_107_22_pad_groupi_n_1121;
  wire csa_tree_add_107_22_pad_groupi_n_1122, csa_tree_add_107_22_pad_groupi_n_1123, csa_tree_add_107_22_pad_groupi_n_1124, csa_tree_add_107_22_pad_groupi_n_1125, csa_tree_add_107_22_pad_groupi_n_1126, csa_tree_add_107_22_pad_groupi_n_1127, csa_tree_add_107_22_pad_groupi_n_1128, csa_tree_add_107_22_pad_groupi_n_1129;
  wire csa_tree_add_107_22_pad_groupi_n_1130, csa_tree_add_107_22_pad_groupi_n_1131, csa_tree_add_107_22_pad_groupi_n_1132, csa_tree_add_107_22_pad_groupi_n_1133, csa_tree_add_107_22_pad_groupi_n_1134, csa_tree_add_107_22_pad_groupi_n_1135, csa_tree_add_107_22_pad_groupi_n_1136, csa_tree_add_107_22_pad_groupi_n_1137;
  wire csa_tree_add_107_22_pad_groupi_n_1138, csa_tree_add_107_22_pad_groupi_n_1139, csa_tree_add_107_22_pad_groupi_n_1140, csa_tree_add_107_22_pad_groupi_n_1141, csa_tree_add_107_22_pad_groupi_n_1142, csa_tree_add_107_22_pad_groupi_n_1143, csa_tree_add_107_22_pad_groupi_n_1144, csa_tree_add_107_22_pad_groupi_n_1145;
  wire csa_tree_add_107_22_pad_groupi_n_1146, csa_tree_add_107_22_pad_groupi_n_1147, csa_tree_add_107_22_pad_groupi_n_1148, csa_tree_add_107_22_pad_groupi_n_1149, csa_tree_add_107_22_pad_groupi_n_1150, csa_tree_add_107_22_pad_groupi_n_1151, csa_tree_add_107_22_pad_groupi_n_1152, csa_tree_add_107_22_pad_groupi_n_1153;
  wire csa_tree_add_107_22_pad_groupi_n_1154, csa_tree_add_107_22_pad_groupi_n_1155, csa_tree_add_107_22_pad_groupi_n_1156, csa_tree_add_107_22_pad_groupi_n_1157, csa_tree_add_107_22_pad_groupi_n_1158, csa_tree_add_107_22_pad_groupi_n_1159, csa_tree_add_107_22_pad_groupi_n_1160, csa_tree_add_107_22_pad_groupi_n_1161;
  wire csa_tree_add_107_22_pad_groupi_n_1162, csa_tree_add_107_22_pad_groupi_n_1163, csa_tree_add_107_22_pad_groupi_n_1164, csa_tree_add_107_22_pad_groupi_n_1165, csa_tree_add_107_22_pad_groupi_n_1166, csa_tree_add_107_22_pad_groupi_n_1167, csa_tree_add_107_22_pad_groupi_n_1168, csa_tree_add_107_22_pad_groupi_n_1169;
  wire csa_tree_add_107_22_pad_groupi_n_1170, csa_tree_add_107_22_pad_groupi_n_1171, csa_tree_add_107_22_pad_groupi_n_1172, csa_tree_add_107_22_pad_groupi_n_1173, csa_tree_add_107_22_pad_groupi_n_1174, csa_tree_add_107_22_pad_groupi_n_1175, csa_tree_add_107_22_pad_groupi_n_1176, csa_tree_add_107_22_pad_groupi_n_1177;
  wire csa_tree_add_107_22_pad_groupi_n_1178, csa_tree_add_107_22_pad_groupi_n_1179, csa_tree_add_107_22_pad_groupi_n_1180, csa_tree_add_107_22_pad_groupi_n_1181, csa_tree_add_107_22_pad_groupi_n_1182, csa_tree_add_107_22_pad_groupi_n_1183, csa_tree_add_107_22_pad_groupi_n_1184, csa_tree_add_107_22_pad_groupi_n_1185;
  wire csa_tree_add_107_22_pad_groupi_n_1186, csa_tree_add_107_22_pad_groupi_n_1187, csa_tree_add_107_22_pad_groupi_n_1188, csa_tree_add_107_22_pad_groupi_n_1189, csa_tree_add_107_22_pad_groupi_n_1190, csa_tree_add_107_22_pad_groupi_n_1191, csa_tree_add_107_22_pad_groupi_n_1192, csa_tree_add_107_22_pad_groupi_n_1193;
  wire csa_tree_add_107_22_pad_groupi_n_1194, csa_tree_add_107_22_pad_groupi_n_1195, csa_tree_add_107_22_pad_groupi_n_1196, csa_tree_add_107_22_pad_groupi_n_1197, csa_tree_add_107_22_pad_groupi_n_1198, csa_tree_add_107_22_pad_groupi_n_1199, csa_tree_add_107_22_pad_groupi_n_1200, csa_tree_add_107_22_pad_groupi_n_1201;
  wire csa_tree_add_107_22_pad_groupi_n_1202, csa_tree_add_107_22_pad_groupi_n_1203, csa_tree_add_107_22_pad_groupi_n_1204, csa_tree_add_107_22_pad_groupi_n_1205, csa_tree_add_107_22_pad_groupi_n_1206, csa_tree_add_107_22_pad_groupi_n_1207, csa_tree_add_107_22_pad_groupi_n_1208, csa_tree_add_107_22_pad_groupi_n_1209;
  wire csa_tree_add_107_22_pad_groupi_n_1210, csa_tree_add_107_22_pad_groupi_n_1211, csa_tree_add_107_22_pad_groupi_n_1212, csa_tree_add_107_22_pad_groupi_n_1213, csa_tree_add_107_22_pad_groupi_n_1214, csa_tree_add_107_22_pad_groupi_n_1215, csa_tree_add_107_22_pad_groupi_n_1216, csa_tree_add_107_22_pad_groupi_n_1217;
  wire csa_tree_add_107_22_pad_groupi_n_1218, csa_tree_add_107_22_pad_groupi_n_1219, csa_tree_add_107_22_pad_groupi_n_1220, csa_tree_add_107_22_pad_groupi_n_1221, csa_tree_add_107_22_pad_groupi_n_1222, csa_tree_add_107_22_pad_groupi_n_1223, csa_tree_add_107_22_pad_groupi_n_1224, csa_tree_add_107_22_pad_groupi_n_1225;
  wire csa_tree_add_107_22_pad_groupi_n_1226, csa_tree_add_107_22_pad_groupi_n_1227, csa_tree_add_107_22_pad_groupi_n_1228, csa_tree_add_107_22_pad_groupi_n_1229, csa_tree_add_107_22_pad_groupi_n_1230, csa_tree_add_107_22_pad_groupi_n_1231, csa_tree_add_107_22_pad_groupi_n_1232, csa_tree_add_107_22_pad_groupi_n_1233;
  wire csa_tree_add_107_22_pad_groupi_n_1234, csa_tree_add_107_22_pad_groupi_n_1235, csa_tree_add_107_22_pad_groupi_n_1236, csa_tree_add_107_22_pad_groupi_n_1237, csa_tree_add_107_22_pad_groupi_n_1238, csa_tree_add_107_22_pad_groupi_n_1239, csa_tree_add_107_22_pad_groupi_n_1240, csa_tree_add_107_22_pad_groupi_n_1241;
  wire csa_tree_add_107_22_pad_groupi_n_1242, csa_tree_add_107_22_pad_groupi_n_1243, csa_tree_add_107_22_pad_groupi_n_1244, csa_tree_add_107_22_pad_groupi_n_1245, csa_tree_add_107_22_pad_groupi_n_1246, csa_tree_add_107_22_pad_groupi_n_1247, csa_tree_add_107_22_pad_groupi_n_1248, csa_tree_add_107_22_pad_groupi_n_1249;
  wire csa_tree_add_107_22_pad_groupi_n_1250, csa_tree_add_107_22_pad_groupi_n_1251, csa_tree_add_107_22_pad_groupi_n_1252, csa_tree_add_107_22_pad_groupi_n_1253, csa_tree_add_107_22_pad_groupi_n_1254, csa_tree_add_107_22_pad_groupi_n_1255, csa_tree_add_107_22_pad_groupi_n_1256, csa_tree_add_107_22_pad_groupi_n_1257;
  wire csa_tree_add_107_22_pad_groupi_n_1258, csa_tree_add_107_22_pad_groupi_n_1259, csa_tree_add_107_22_pad_groupi_n_1260, csa_tree_add_107_22_pad_groupi_n_1261, csa_tree_add_107_22_pad_groupi_n_1262, csa_tree_add_107_22_pad_groupi_n_1263, csa_tree_add_107_22_pad_groupi_n_1264, csa_tree_add_107_22_pad_groupi_n_1265;
  wire csa_tree_add_107_22_pad_groupi_n_1266, csa_tree_add_107_22_pad_groupi_n_1267, csa_tree_add_107_22_pad_groupi_n_1268, csa_tree_add_107_22_pad_groupi_n_1269, csa_tree_add_107_22_pad_groupi_n_1270, csa_tree_add_107_22_pad_groupi_n_1271, csa_tree_add_107_22_pad_groupi_n_1272, csa_tree_add_107_22_pad_groupi_n_1273;
  wire csa_tree_add_107_22_pad_groupi_n_1274, csa_tree_add_107_22_pad_groupi_n_1275, csa_tree_add_107_22_pad_groupi_n_1276, csa_tree_add_107_22_pad_groupi_n_1277, csa_tree_add_107_22_pad_groupi_n_1278, csa_tree_add_107_22_pad_groupi_n_1279, csa_tree_add_107_22_pad_groupi_n_1280, csa_tree_add_107_22_pad_groupi_n_1281;
  wire csa_tree_add_107_22_pad_groupi_n_1282, csa_tree_add_107_22_pad_groupi_n_1283, csa_tree_add_107_22_pad_groupi_n_1284, csa_tree_add_107_22_pad_groupi_n_1285, csa_tree_add_107_22_pad_groupi_n_1286, csa_tree_add_107_22_pad_groupi_n_1287, csa_tree_add_107_22_pad_groupi_n_1288, csa_tree_add_107_22_pad_groupi_n_1289;
  wire csa_tree_add_107_22_pad_groupi_n_1290, csa_tree_add_107_22_pad_groupi_n_1291, csa_tree_add_107_22_pad_groupi_n_1292, csa_tree_add_107_22_pad_groupi_n_1293, csa_tree_add_107_22_pad_groupi_n_1294, csa_tree_add_107_22_pad_groupi_n_1295, csa_tree_add_107_22_pad_groupi_n_1296, csa_tree_add_107_22_pad_groupi_n_1297;
  wire csa_tree_add_107_22_pad_groupi_n_1298, csa_tree_add_107_22_pad_groupi_n_1299, csa_tree_add_107_22_pad_groupi_n_1300, csa_tree_add_107_22_pad_groupi_n_1301, csa_tree_add_107_22_pad_groupi_n_1302, csa_tree_add_107_22_pad_groupi_n_1303, csa_tree_add_107_22_pad_groupi_n_1304, csa_tree_add_107_22_pad_groupi_n_1305;
  wire csa_tree_add_107_22_pad_groupi_n_1306, csa_tree_add_107_22_pad_groupi_n_1307, csa_tree_add_107_22_pad_groupi_n_1308, csa_tree_add_107_22_pad_groupi_n_1309, csa_tree_add_107_22_pad_groupi_n_1310, csa_tree_add_107_22_pad_groupi_n_1311, csa_tree_add_107_22_pad_groupi_n_1312, csa_tree_add_107_22_pad_groupi_n_1313;
  wire csa_tree_add_107_22_pad_groupi_n_1314, csa_tree_add_107_22_pad_groupi_n_1315, csa_tree_add_107_22_pad_groupi_n_1316, csa_tree_add_107_22_pad_groupi_n_1317, csa_tree_add_107_22_pad_groupi_n_1318, csa_tree_add_107_22_pad_groupi_n_1319, csa_tree_add_107_22_pad_groupi_n_1320, csa_tree_add_107_22_pad_groupi_n_1321;
  wire csa_tree_add_107_22_pad_groupi_n_1322, csa_tree_add_107_22_pad_groupi_n_1323, csa_tree_add_107_22_pad_groupi_n_1324, csa_tree_add_107_22_pad_groupi_n_1325, csa_tree_add_107_22_pad_groupi_n_1326, csa_tree_add_107_22_pad_groupi_n_1327, csa_tree_add_107_22_pad_groupi_n_1328, csa_tree_add_107_22_pad_groupi_n_1329;
  wire csa_tree_add_107_22_pad_groupi_n_1330, csa_tree_add_107_22_pad_groupi_n_1331, csa_tree_add_107_22_pad_groupi_n_1332, csa_tree_add_107_22_pad_groupi_n_1333, csa_tree_add_107_22_pad_groupi_n_1334, csa_tree_add_107_22_pad_groupi_n_1335, csa_tree_add_107_22_pad_groupi_n_1336, csa_tree_add_107_22_pad_groupi_n_1337;
  wire csa_tree_add_107_22_pad_groupi_n_1338, csa_tree_add_107_22_pad_groupi_n_1339, csa_tree_add_107_22_pad_groupi_n_1340, csa_tree_add_107_22_pad_groupi_n_1341, csa_tree_add_107_22_pad_groupi_n_1342, csa_tree_add_107_22_pad_groupi_n_1343, csa_tree_add_107_22_pad_groupi_n_1344, csa_tree_add_107_22_pad_groupi_n_1345;
  wire csa_tree_add_107_22_pad_groupi_n_1346, csa_tree_add_107_22_pad_groupi_n_1347, csa_tree_add_107_22_pad_groupi_n_1348, csa_tree_add_107_22_pad_groupi_n_1349, csa_tree_add_107_22_pad_groupi_n_1350, csa_tree_add_107_22_pad_groupi_n_1351, csa_tree_add_107_22_pad_groupi_n_1352, csa_tree_add_107_22_pad_groupi_n_1353;
  wire csa_tree_add_107_22_pad_groupi_n_1354, csa_tree_add_107_22_pad_groupi_n_1355, csa_tree_add_107_22_pad_groupi_n_1356, csa_tree_add_107_22_pad_groupi_n_1357, csa_tree_add_107_22_pad_groupi_n_1358, csa_tree_add_107_22_pad_groupi_n_1359, csa_tree_add_107_22_pad_groupi_n_1360, csa_tree_add_107_22_pad_groupi_n_1361;
  wire csa_tree_add_107_22_pad_groupi_n_1362, csa_tree_add_107_22_pad_groupi_n_1363, csa_tree_add_107_22_pad_groupi_n_1364, csa_tree_add_107_22_pad_groupi_n_1365, csa_tree_add_107_22_pad_groupi_n_1366, csa_tree_add_107_22_pad_groupi_n_1367, csa_tree_add_107_22_pad_groupi_n_1368, csa_tree_add_107_22_pad_groupi_n_1369;
  wire csa_tree_add_107_22_pad_groupi_n_1370, csa_tree_add_107_22_pad_groupi_n_1371, csa_tree_add_107_22_pad_groupi_n_1372, csa_tree_add_107_22_pad_groupi_n_1373, csa_tree_add_107_22_pad_groupi_n_1374, csa_tree_add_107_22_pad_groupi_n_1375, csa_tree_add_107_22_pad_groupi_n_1376, csa_tree_add_107_22_pad_groupi_n_1377;
  wire csa_tree_add_107_22_pad_groupi_n_1378, csa_tree_add_107_22_pad_groupi_n_1379, csa_tree_add_107_22_pad_groupi_n_1380, csa_tree_add_107_22_pad_groupi_n_1381, csa_tree_add_107_22_pad_groupi_n_1382, csa_tree_add_107_22_pad_groupi_n_1383, csa_tree_add_107_22_pad_groupi_n_1384, csa_tree_add_107_22_pad_groupi_n_1385;
  wire csa_tree_add_107_22_pad_groupi_n_1386, csa_tree_add_107_22_pad_groupi_n_1387, csa_tree_add_107_22_pad_groupi_n_1388, csa_tree_add_107_22_pad_groupi_n_1389, csa_tree_add_107_22_pad_groupi_n_1390, csa_tree_add_107_22_pad_groupi_n_1391, csa_tree_add_107_22_pad_groupi_n_1392, csa_tree_add_107_22_pad_groupi_n_1393;
  wire csa_tree_add_107_22_pad_groupi_n_1394, csa_tree_add_107_22_pad_groupi_n_1395, csa_tree_add_107_22_pad_groupi_n_1396, csa_tree_add_107_22_pad_groupi_n_1397, csa_tree_add_107_22_pad_groupi_n_1398, csa_tree_add_107_22_pad_groupi_n_1399, csa_tree_add_107_22_pad_groupi_n_1400, csa_tree_add_107_22_pad_groupi_n_1401;
  wire csa_tree_add_107_22_pad_groupi_n_1402, csa_tree_add_107_22_pad_groupi_n_1403, csa_tree_add_107_22_pad_groupi_n_1404, csa_tree_add_107_22_pad_groupi_n_1405, csa_tree_add_107_22_pad_groupi_n_1406, csa_tree_add_107_22_pad_groupi_n_1407, csa_tree_add_107_22_pad_groupi_n_1408, csa_tree_add_107_22_pad_groupi_n_1409;
  wire csa_tree_add_107_22_pad_groupi_n_1410, csa_tree_add_107_22_pad_groupi_n_1411, csa_tree_add_107_22_pad_groupi_n_1412, csa_tree_add_107_22_pad_groupi_n_1413, csa_tree_add_107_22_pad_groupi_n_1414, csa_tree_add_107_22_pad_groupi_n_1415, csa_tree_add_107_22_pad_groupi_n_1416, csa_tree_add_107_22_pad_groupi_n_1417;
  wire csa_tree_add_107_22_pad_groupi_n_1418, csa_tree_add_107_22_pad_groupi_n_1419, csa_tree_add_107_22_pad_groupi_n_1420, csa_tree_add_107_22_pad_groupi_n_1421, csa_tree_add_107_22_pad_groupi_n_1422, csa_tree_add_107_22_pad_groupi_n_1423, csa_tree_add_107_22_pad_groupi_n_1424, csa_tree_add_107_22_pad_groupi_n_1425;
  wire csa_tree_add_107_22_pad_groupi_n_1426, csa_tree_add_107_22_pad_groupi_n_1427, csa_tree_add_107_22_pad_groupi_n_1428, csa_tree_add_107_22_pad_groupi_n_1429, csa_tree_add_107_22_pad_groupi_n_1430, csa_tree_add_107_22_pad_groupi_n_1431, csa_tree_add_107_22_pad_groupi_n_1432, csa_tree_add_107_22_pad_groupi_n_1433;
  wire csa_tree_add_107_22_pad_groupi_n_1434, csa_tree_add_107_22_pad_groupi_n_1435, csa_tree_add_107_22_pad_groupi_n_1436, csa_tree_add_107_22_pad_groupi_n_1437, csa_tree_add_107_22_pad_groupi_n_1438, csa_tree_add_107_22_pad_groupi_n_1439, csa_tree_add_107_22_pad_groupi_n_1440, csa_tree_add_107_22_pad_groupi_n_1441;
  wire csa_tree_add_107_22_pad_groupi_n_1442, csa_tree_add_107_22_pad_groupi_n_1443, csa_tree_add_107_22_pad_groupi_n_1444, csa_tree_add_107_22_pad_groupi_n_1445, csa_tree_add_107_22_pad_groupi_n_1446, csa_tree_add_107_22_pad_groupi_n_1447, csa_tree_add_107_22_pad_groupi_n_1448, csa_tree_add_107_22_pad_groupi_n_1449;
  wire csa_tree_add_107_22_pad_groupi_n_1450, csa_tree_add_107_22_pad_groupi_n_1451, csa_tree_add_107_22_pad_groupi_n_1452, csa_tree_add_107_22_pad_groupi_n_1453, csa_tree_add_107_22_pad_groupi_n_1454, csa_tree_add_107_22_pad_groupi_n_1455, csa_tree_add_107_22_pad_groupi_n_1456, csa_tree_add_107_22_pad_groupi_n_1457;
  wire csa_tree_add_107_22_pad_groupi_n_1458, csa_tree_add_107_22_pad_groupi_n_1459, csa_tree_add_107_22_pad_groupi_n_1460, csa_tree_add_107_22_pad_groupi_n_1461, csa_tree_add_107_22_pad_groupi_n_1462, csa_tree_add_107_22_pad_groupi_n_1463, csa_tree_add_107_22_pad_groupi_n_1464, csa_tree_add_107_22_pad_groupi_n_1465;
  wire csa_tree_add_107_22_pad_groupi_n_1466, csa_tree_add_107_22_pad_groupi_n_1467, csa_tree_add_107_22_pad_groupi_n_1468, csa_tree_add_107_22_pad_groupi_n_1469, csa_tree_add_107_22_pad_groupi_n_1470, csa_tree_add_107_22_pad_groupi_n_1471, csa_tree_add_107_22_pad_groupi_n_1472, csa_tree_add_107_22_pad_groupi_n_1473;
  wire csa_tree_add_107_22_pad_groupi_n_1474, csa_tree_add_107_22_pad_groupi_n_1475, csa_tree_add_107_22_pad_groupi_n_1476, csa_tree_add_107_22_pad_groupi_n_1477, csa_tree_add_107_22_pad_groupi_n_1478, csa_tree_add_107_22_pad_groupi_n_1479, csa_tree_add_107_22_pad_groupi_n_1480, csa_tree_add_107_22_pad_groupi_n_1481;
  wire csa_tree_add_107_22_pad_groupi_n_1482, csa_tree_add_107_22_pad_groupi_n_1483, csa_tree_add_107_22_pad_groupi_n_1484, csa_tree_add_107_22_pad_groupi_n_1485, csa_tree_add_107_22_pad_groupi_n_1486, csa_tree_add_107_22_pad_groupi_n_1487, csa_tree_add_107_22_pad_groupi_n_1488, csa_tree_add_107_22_pad_groupi_n_1489;
  wire csa_tree_add_107_22_pad_groupi_n_1490, csa_tree_add_107_22_pad_groupi_n_1491, csa_tree_add_107_22_pad_groupi_n_1492, csa_tree_add_107_22_pad_groupi_n_1493, csa_tree_add_107_22_pad_groupi_n_1494, csa_tree_add_107_22_pad_groupi_n_1495, csa_tree_add_107_22_pad_groupi_n_1496, csa_tree_add_107_22_pad_groupi_n_1497;
  wire csa_tree_add_107_22_pad_groupi_n_1498, csa_tree_add_107_22_pad_groupi_n_1499, csa_tree_add_107_22_pad_groupi_n_1500, csa_tree_add_107_22_pad_groupi_n_1501, csa_tree_add_107_22_pad_groupi_n_1502, csa_tree_add_107_22_pad_groupi_n_1503, csa_tree_add_107_22_pad_groupi_n_1505, csa_tree_add_107_22_pad_groupi_n_1506;
  wire csa_tree_add_107_22_pad_groupi_n_1507, csa_tree_add_107_22_pad_groupi_n_1508, csa_tree_add_107_22_pad_groupi_n_1509, csa_tree_add_107_22_pad_groupi_n_1510, csa_tree_add_107_22_pad_groupi_n_1511, csa_tree_add_107_22_pad_groupi_n_1512, csa_tree_add_107_22_pad_groupi_n_1513, csa_tree_add_107_22_pad_groupi_n_1514;
  wire csa_tree_add_107_22_pad_groupi_n_1515, csa_tree_add_107_22_pad_groupi_n_1516, csa_tree_add_107_22_pad_groupi_n_1517, csa_tree_add_107_22_pad_groupi_n_1518, csa_tree_add_107_22_pad_groupi_n_1519, csa_tree_add_107_22_pad_groupi_n_1520, csa_tree_add_107_22_pad_groupi_n_1521, csa_tree_add_107_22_pad_groupi_n_1522;
  wire csa_tree_add_107_22_pad_groupi_n_1523, csa_tree_add_107_22_pad_groupi_n_1524, csa_tree_add_107_22_pad_groupi_n_1525, csa_tree_add_107_22_pad_groupi_n_1526, csa_tree_add_107_22_pad_groupi_n_1527, csa_tree_add_107_22_pad_groupi_n_1529, csa_tree_add_107_22_pad_groupi_n_1530, csa_tree_add_107_22_pad_groupi_n_1532;
  wire csa_tree_add_107_22_pad_groupi_n_1533, csa_tree_add_107_22_pad_groupi_n_1534, csa_tree_add_107_22_pad_groupi_n_1535, csa_tree_add_107_22_pad_groupi_n_1537, csa_tree_add_107_22_pad_groupi_n_1538, csa_tree_add_107_22_pad_groupi_n_1539, csa_tree_add_107_22_pad_groupi_n_1540, csa_tree_add_107_22_pad_groupi_n_1542;
  wire csa_tree_add_107_22_pad_groupi_n_1543, csa_tree_add_107_22_pad_groupi_n_1544, csa_tree_add_107_22_pad_groupi_n_1546, csa_tree_add_107_22_pad_groupi_n_1547, csa_tree_add_107_22_pad_groupi_n_1549, csa_tree_add_107_22_pad_groupi_n_1550, csa_tree_add_107_22_pad_groupi_n_1552, csa_tree_add_107_22_pad_groupi_n_1553;
  wire csa_tree_add_107_22_pad_groupi_n_1555, csa_tree_add_107_22_pad_groupi_n_1556, csa_tree_add_107_22_pad_groupi_n_1558, csa_tree_add_110_49_pad_groupi_n_0, csa_tree_add_110_49_pad_groupi_n_1, csa_tree_add_110_49_pad_groupi_n_4, csa_tree_add_110_49_pad_groupi_n_5, csa_tree_add_110_49_pad_groupi_n_6;
  wire csa_tree_add_110_49_pad_groupi_n_7, csa_tree_add_110_49_pad_groupi_n_8, csa_tree_add_110_49_pad_groupi_n_9, csa_tree_add_110_49_pad_groupi_n_10, csa_tree_add_110_49_pad_groupi_n_11, csa_tree_add_110_49_pad_groupi_n_12, csa_tree_add_110_49_pad_groupi_n_13, csa_tree_add_110_49_pad_groupi_n_14;
  wire csa_tree_add_110_49_pad_groupi_n_15, csa_tree_add_110_49_pad_groupi_n_16, csa_tree_add_110_49_pad_groupi_n_17, csa_tree_add_110_49_pad_groupi_n_18, csa_tree_add_110_49_pad_groupi_n_19, csa_tree_add_110_49_pad_groupi_n_20, csa_tree_add_110_49_pad_groupi_n_21, csa_tree_add_110_49_pad_groupi_n_22;
  wire csa_tree_add_110_49_pad_groupi_n_23, csa_tree_add_110_49_pad_groupi_n_24, csa_tree_add_110_49_pad_groupi_n_25, csa_tree_add_110_49_pad_groupi_n_26, csa_tree_add_110_49_pad_groupi_n_27, csa_tree_add_110_49_pad_groupi_n_28, csa_tree_add_110_49_pad_groupi_n_29, csa_tree_add_110_49_pad_groupi_n_30;
  wire csa_tree_add_110_49_pad_groupi_n_31, csa_tree_add_110_49_pad_groupi_n_32, csa_tree_add_110_49_pad_groupi_n_33, csa_tree_add_110_49_pad_groupi_n_34, csa_tree_add_110_49_pad_groupi_n_35, csa_tree_add_110_49_pad_groupi_n_36, csa_tree_add_110_49_pad_groupi_n_37, csa_tree_add_110_49_pad_groupi_n_38;
  wire csa_tree_add_110_49_pad_groupi_n_39, csa_tree_add_110_49_pad_groupi_n_40, csa_tree_add_110_49_pad_groupi_n_41, csa_tree_add_110_49_pad_groupi_n_42, csa_tree_add_110_49_pad_groupi_n_43, csa_tree_add_110_49_pad_groupi_n_44, csa_tree_add_110_49_pad_groupi_n_45, csa_tree_add_110_49_pad_groupi_n_46;
  wire csa_tree_add_110_49_pad_groupi_n_47, csa_tree_add_110_49_pad_groupi_n_48, csa_tree_add_110_49_pad_groupi_n_49, csa_tree_add_110_49_pad_groupi_n_50, csa_tree_add_110_49_pad_groupi_n_51, csa_tree_add_110_49_pad_groupi_n_52, csa_tree_add_110_49_pad_groupi_n_53, csa_tree_add_110_49_pad_groupi_n_54;
  wire csa_tree_add_110_49_pad_groupi_n_55, csa_tree_add_110_49_pad_groupi_n_56, csa_tree_add_110_49_pad_groupi_n_57, csa_tree_add_110_49_pad_groupi_n_58, csa_tree_add_110_49_pad_groupi_n_59, csa_tree_add_110_49_pad_groupi_n_60, csa_tree_add_110_49_pad_groupi_n_61, csa_tree_add_110_49_pad_groupi_n_62;
  wire csa_tree_add_110_49_pad_groupi_n_63, csa_tree_add_110_49_pad_groupi_n_64, csa_tree_add_110_49_pad_groupi_n_65, csa_tree_add_110_49_pad_groupi_n_66, csa_tree_add_110_49_pad_groupi_n_67, csa_tree_add_110_49_pad_groupi_n_68, csa_tree_add_110_49_pad_groupi_n_69, csa_tree_add_110_49_pad_groupi_n_70;
  wire csa_tree_add_110_49_pad_groupi_n_71, csa_tree_add_110_49_pad_groupi_n_72, csa_tree_add_110_49_pad_groupi_n_73, csa_tree_add_110_49_pad_groupi_n_74, csa_tree_add_110_49_pad_groupi_n_75, csa_tree_add_110_49_pad_groupi_n_76, csa_tree_add_110_49_pad_groupi_n_77, csa_tree_add_110_49_pad_groupi_n_78;
  wire csa_tree_add_110_49_pad_groupi_n_79, csa_tree_add_110_49_pad_groupi_n_80, csa_tree_add_110_49_pad_groupi_n_81, csa_tree_add_110_49_pad_groupi_n_82, csa_tree_add_110_49_pad_groupi_n_83, csa_tree_add_110_49_pad_groupi_n_84, csa_tree_add_110_49_pad_groupi_n_85, csa_tree_add_110_49_pad_groupi_n_86;
  wire csa_tree_add_110_49_pad_groupi_n_87, csa_tree_add_110_49_pad_groupi_n_88, csa_tree_add_110_49_pad_groupi_n_89, csa_tree_add_110_49_pad_groupi_n_90, csa_tree_add_110_49_pad_groupi_n_91, csa_tree_add_110_49_pad_groupi_n_92, csa_tree_add_110_49_pad_groupi_n_93, csa_tree_add_110_49_pad_groupi_n_94;
  wire csa_tree_add_110_49_pad_groupi_n_95, csa_tree_add_110_49_pad_groupi_n_96, csa_tree_add_110_49_pad_groupi_n_97, csa_tree_add_110_49_pad_groupi_n_98, csa_tree_add_110_49_pad_groupi_n_99, csa_tree_add_110_49_pad_groupi_n_100, csa_tree_add_110_49_pad_groupi_n_101, csa_tree_add_110_49_pad_groupi_n_102;
  wire csa_tree_add_110_49_pad_groupi_n_103, csa_tree_add_110_49_pad_groupi_n_104, csa_tree_add_110_49_pad_groupi_n_105, csa_tree_add_110_49_pad_groupi_n_106, csa_tree_add_110_49_pad_groupi_n_107, csa_tree_add_110_49_pad_groupi_n_108, csa_tree_add_110_49_pad_groupi_n_109, csa_tree_add_110_49_pad_groupi_n_110;
  wire csa_tree_add_110_49_pad_groupi_n_111, csa_tree_add_110_49_pad_groupi_n_112, csa_tree_add_110_49_pad_groupi_n_113, csa_tree_add_110_49_pad_groupi_n_114, csa_tree_add_110_49_pad_groupi_n_115, csa_tree_add_110_49_pad_groupi_n_116, csa_tree_add_110_49_pad_groupi_n_117, csa_tree_add_110_49_pad_groupi_n_118;
  wire csa_tree_add_110_49_pad_groupi_n_119, csa_tree_add_110_49_pad_groupi_n_120, csa_tree_add_110_49_pad_groupi_n_121, csa_tree_add_110_49_pad_groupi_n_122, csa_tree_add_110_49_pad_groupi_n_123, csa_tree_add_110_49_pad_groupi_n_124, csa_tree_add_110_49_pad_groupi_n_125, csa_tree_add_110_49_pad_groupi_n_126;
  wire csa_tree_add_110_49_pad_groupi_n_127, csa_tree_add_110_49_pad_groupi_n_128, csa_tree_add_110_49_pad_groupi_n_129, csa_tree_add_110_49_pad_groupi_n_130, csa_tree_add_110_49_pad_groupi_n_131, csa_tree_add_110_49_pad_groupi_n_132, csa_tree_add_110_49_pad_groupi_n_133, csa_tree_add_110_49_pad_groupi_n_134;
  wire csa_tree_add_110_49_pad_groupi_n_135, csa_tree_add_110_49_pad_groupi_n_136, csa_tree_add_110_49_pad_groupi_n_137, csa_tree_add_110_49_pad_groupi_n_138, csa_tree_add_110_49_pad_groupi_n_139, csa_tree_add_110_49_pad_groupi_n_140, csa_tree_add_110_49_pad_groupi_n_141, csa_tree_add_110_49_pad_groupi_n_142;
  wire csa_tree_add_110_49_pad_groupi_n_143, csa_tree_add_110_49_pad_groupi_n_144, csa_tree_add_110_49_pad_groupi_n_145, csa_tree_add_110_49_pad_groupi_n_146, csa_tree_add_110_49_pad_groupi_n_147, csa_tree_add_110_49_pad_groupi_n_148, csa_tree_add_110_49_pad_groupi_n_149, csa_tree_add_110_49_pad_groupi_n_150;
  wire csa_tree_add_110_49_pad_groupi_n_151, csa_tree_add_110_49_pad_groupi_n_152, csa_tree_add_110_49_pad_groupi_n_153, csa_tree_add_110_49_pad_groupi_n_154, csa_tree_add_110_49_pad_groupi_n_155, csa_tree_add_110_49_pad_groupi_n_156, csa_tree_add_110_49_pad_groupi_n_157, csa_tree_add_110_49_pad_groupi_n_158;
  wire csa_tree_add_110_49_pad_groupi_n_159, csa_tree_add_110_49_pad_groupi_n_160, csa_tree_add_110_49_pad_groupi_n_161, csa_tree_add_110_49_pad_groupi_n_162, csa_tree_add_110_49_pad_groupi_n_163, csa_tree_add_110_49_pad_groupi_n_164, csa_tree_add_110_49_pad_groupi_n_165, csa_tree_add_110_49_pad_groupi_n_166;
  wire csa_tree_add_110_49_pad_groupi_n_167, csa_tree_add_110_49_pad_groupi_n_168, csa_tree_add_110_49_pad_groupi_n_169, csa_tree_add_110_49_pad_groupi_n_170, csa_tree_add_110_49_pad_groupi_n_171, csa_tree_add_110_49_pad_groupi_n_172, csa_tree_add_110_49_pad_groupi_n_173, csa_tree_add_110_49_pad_groupi_n_174;
  wire csa_tree_add_110_49_pad_groupi_n_175, csa_tree_add_110_49_pad_groupi_n_176, csa_tree_add_110_49_pad_groupi_n_177, csa_tree_add_110_49_pad_groupi_n_178, csa_tree_add_110_49_pad_groupi_n_179, csa_tree_add_110_49_pad_groupi_n_180, csa_tree_add_110_49_pad_groupi_n_181, csa_tree_add_110_49_pad_groupi_n_182;
  wire csa_tree_add_110_49_pad_groupi_n_183, csa_tree_add_110_49_pad_groupi_n_184, csa_tree_add_110_49_pad_groupi_n_185, csa_tree_add_110_49_pad_groupi_n_186, csa_tree_add_110_49_pad_groupi_n_187, csa_tree_add_110_49_pad_groupi_n_188, csa_tree_add_110_49_pad_groupi_n_189, csa_tree_add_110_49_pad_groupi_n_190;
  wire csa_tree_add_110_49_pad_groupi_n_191, csa_tree_add_110_49_pad_groupi_n_192, csa_tree_add_110_49_pad_groupi_n_193, csa_tree_add_110_49_pad_groupi_n_194, csa_tree_add_110_49_pad_groupi_n_195, csa_tree_add_110_49_pad_groupi_n_196, csa_tree_add_110_49_pad_groupi_n_197, csa_tree_add_110_49_pad_groupi_n_198;
  wire csa_tree_add_110_49_pad_groupi_n_199, csa_tree_add_110_49_pad_groupi_n_200, csa_tree_add_110_49_pad_groupi_n_201, csa_tree_add_110_49_pad_groupi_n_202, csa_tree_add_110_49_pad_groupi_n_203, csa_tree_add_110_49_pad_groupi_n_204, csa_tree_add_110_49_pad_groupi_n_205, csa_tree_add_110_49_pad_groupi_n_206;
  wire csa_tree_add_110_49_pad_groupi_n_207, csa_tree_add_110_49_pad_groupi_n_208, csa_tree_add_110_49_pad_groupi_n_209, csa_tree_add_110_49_pad_groupi_n_210, csa_tree_add_110_49_pad_groupi_n_211, csa_tree_add_110_49_pad_groupi_n_212, csa_tree_add_110_49_pad_groupi_n_213, csa_tree_add_110_49_pad_groupi_n_214;
  wire csa_tree_add_110_49_pad_groupi_n_215, csa_tree_add_110_49_pad_groupi_n_216, csa_tree_add_110_49_pad_groupi_n_217, csa_tree_add_110_49_pad_groupi_n_218, csa_tree_add_110_49_pad_groupi_n_219, csa_tree_add_110_49_pad_groupi_n_220, csa_tree_add_110_49_pad_groupi_n_221, csa_tree_add_110_49_pad_groupi_n_222;
  wire csa_tree_add_110_49_pad_groupi_n_223, csa_tree_add_110_49_pad_groupi_n_224, csa_tree_add_110_49_pad_groupi_n_225, csa_tree_add_110_49_pad_groupi_n_226, csa_tree_add_110_49_pad_groupi_n_227, csa_tree_add_110_49_pad_groupi_n_228, csa_tree_add_110_49_pad_groupi_n_229, csa_tree_add_110_49_pad_groupi_n_230;
  wire csa_tree_add_110_49_pad_groupi_n_231, csa_tree_add_110_49_pad_groupi_n_232, csa_tree_add_110_49_pad_groupi_n_233, csa_tree_add_110_49_pad_groupi_n_234, csa_tree_add_110_49_pad_groupi_n_235, csa_tree_add_110_49_pad_groupi_n_236, csa_tree_add_110_49_pad_groupi_n_237, csa_tree_add_110_49_pad_groupi_n_238;
  wire csa_tree_add_110_49_pad_groupi_n_239, csa_tree_add_110_49_pad_groupi_n_240, csa_tree_add_110_49_pad_groupi_n_241, csa_tree_add_110_49_pad_groupi_n_242, csa_tree_add_110_49_pad_groupi_n_243, csa_tree_add_110_49_pad_groupi_n_244, csa_tree_add_110_49_pad_groupi_n_245, csa_tree_add_110_49_pad_groupi_n_246;
  wire csa_tree_add_110_49_pad_groupi_n_247, csa_tree_add_110_49_pad_groupi_n_248, csa_tree_add_110_49_pad_groupi_n_249, csa_tree_add_110_49_pad_groupi_n_250, csa_tree_add_110_49_pad_groupi_n_251, csa_tree_add_110_49_pad_groupi_n_252, csa_tree_add_110_49_pad_groupi_n_253, csa_tree_add_110_49_pad_groupi_n_254;
  wire csa_tree_add_110_49_pad_groupi_n_255, csa_tree_add_110_49_pad_groupi_n_256, csa_tree_add_110_49_pad_groupi_n_257, csa_tree_add_110_49_pad_groupi_n_258, csa_tree_add_110_49_pad_groupi_n_259, csa_tree_add_110_49_pad_groupi_n_260, csa_tree_add_110_49_pad_groupi_n_261, csa_tree_add_110_49_pad_groupi_n_262;
  wire csa_tree_add_110_49_pad_groupi_n_263, csa_tree_add_110_49_pad_groupi_n_264, csa_tree_add_110_49_pad_groupi_n_265, csa_tree_add_110_49_pad_groupi_n_266, csa_tree_add_110_49_pad_groupi_n_267, csa_tree_add_110_49_pad_groupi_n_268, csa_tree_add_110_49_pad_groupi_n_269, csa_tree_add_110_49_pad_groupi_n_270;
  wire csa_tree_add_110_49_pad_groupi_n_271, csa_tree_add_110_49_pad_groupi_n_272, csa_tree_add_110_49_pad_groupi_n_273, csa_tree_add_110_49_pad_groupi_n_274, csa_tree_add_110_49_pad_groupi_n_275, csa_tree_add_110_49_pad_groupi_n_276, csa_tree_add_110_49_pad_groupi_n_277, csa_tree_add_110_49_pad_groupi_n_278;
  wire csa_tree_add_110_49_pad_groupi_n_279, csa_tree_add_110_49_pad_groupi_n_280, csa_tree_add_110_49_pad_groupi_n_281, csa_tree_add_110_49_pad_groupi_n_282, csa_tree_add_110_49_pad_groupi_n_283, csa_tree_add_110_49_pad_groupi_n_284, csa_tree_add_110_49_pad_groupi_n_285, csa_tree_add_110_49_pad_groupi_n_286;
  wire csa_tree_add_110_49_pad_groupi_n_287, csa_tree_add_110_49_pad_groupi_n_289, csa_tree_add_110_49_pad_groupi_n_290, csa_tree_add_110_49_pad_groupi_n_291, csa_tree_add_110_49_pad_groupi_n_292, csa_tree_add_110_49_pad_groupi_n_293, csa_tree_add_110_49_pad_groupi_n_294, csa_tree_add_110_49_pad_groupi_n_295;
  wire csa_tree_add_110_49_pad_groupi_n_296, csa_tree_add_110_49_pad_groupi_n_297, csa_tree_add_110_49_pad_groupi_n_298, csa_tree_add_110_49_pad_groupi_n_299, csa_tree_add_110_49_pad_groupi_n_300, csa_tree_add_110_49_pad_groupi_n_301, csa_tree_add_110_49_pad_groupi_n_302, csa_tree_add_110_49_pad_groupi_n_303;
  wire csa_tree_add_110_49_pad_groupi_n_304, csa_tree_add_110_49_pad_groupi_n_305, csa_tree_add_110_49_pad_groupi_n_306, csa_tree_add_110_49_pad_groupi_n_307, csa_tree_add_110_49_pad_groupi_n_308, csa_tree_add_110_49_pad_groupi_n_309, csa_tree_add_110_49_pad_groupi_n_310, csa_tree_add_110_49_pad_groupi_n_311;
  wire csa_tree_add_110_49_pad_groupi_n_312, csa_tree_add_110_49_pad_groupi_n_313, csa_tree_add_110_49_pad_groupi_n_314, csa_tree_add_110_49_pad_groupi_n_315, csa_tree_add_110_49_pad_groupi_n_316, csa_tree_add_110_49_pad_groupi_n_317, csa_tree_add_110_49_pad_groupi_n_318, csa_tree_add_110_49_pad_groupi_n_319;
  wire csa_tree_add_110_49_pad_groupi_n_320, csa_tree_add_110_49_pad_groupi_n_321, csa_tree_add_110_49_pad_groupi_n_322, csa_tree_add_110_49_pad_groupi_n_323, csa_tree_add_110_49_pad_groupi_n_324, csa_tree_add_110_49_pad_groupi_n_325, csa_tree_add_110_49_pad_groupi_n_326, csa_tree_add_110_49_pad_groupi_n_327;
  wire csa_tree_add_110_49_pad_groupi_n_328, csa_tree_add_110_49_pad_groupi_n_329, csa_tree_add_110_49_pad_groupi_n_330, csa_tree_add_110_49_pad_groupi_n_331, csa_tree_add_110_49_pad_groupi_n_332, csa_tree_add_110_49_pad_groupi_n_333, csa_tree_add_110_49_pad_groupi_n_334, csa_tree_add_110_49_pad_groupi_n_335;
  wire csa_tree_add_110_49_pad_groupi_n_336, csa_tree_add_110_49_pad_groupi_n_337, csa_tree_add_110_49_pad_groupi_n_338, csa_tree_add_110_49_pad_groupi_n_339, csa_tree_add_110_49_pad_groupi_n_340, csa_tree_add_110_49_pad_groupi_n_341, csa_tree_add_110_49_pad_groupi_n_342, csa_tree_add_110_49_pad_groupi_n_343;
  wire csa_tree_add_110_49_pad_groupi_n_344, csa_tree_add_110_49_pad_groupi_n_345, csa_tree_add_110_49_pad_groupi_n_346, csa_tree_add_110_49_pad_groupi_n_347, csa_tree_add_110_49_pad_groupi_n_348, csa_tree_add_110_49_pad_groupi_n_349, csa_tree_add_110_49_pad_groupi_n_350, csa_tree_add_110_49_pad_groupi_n_351;
  wire csa_tree_add_110_49_pad_groupi_n_352, csa_tree_add_110_49_pad_groupi_n_353, csa_tree_add_110_49_pad_groupi_n_354, csa_tree_add_110_49_pad_groupi_n_355, csa_tree_add_110_49_pad_groupi_n_356, csa_tree_add_110_49_pad_groupi_n_357, csa_tree_add_110_49_pad_groupi_n_358, csa_tree_add_110_49_pad_groupi_n_359;
  wire csa_tree_add_110_49_pad_groupi_n_360, csa_tree_add_110_49_pad_groupi_n_361, csa_tree_add_110_49_pad_groupi_n_362, csa_tree_add_110_49_pad_groupi_n_363, csa_tree_add_110_49_pad_groupi_n_364, csa_tree_add_110_49_pad_groupi_n_365, csa_tree_add_110_49_pad_groupi_n_366, csa_tree_add_110_49_pad_groupi_n_367;
  wire csa_tree_add_110_49_pad_groupi_n_368, csa_tree_add_110_49_pad_groupi_n_369, csa_tree_add_110_49_pad_groupi_n_370, csa_tree_add_110_49_pad_groupi_n_371, csa_tree_add_110_49_pad_groupi_n_372, csa_tree_add_110_49_pad_groupi_n_373, csa_tree_add_110_49_pad_groupi_n_374, csa_tree_add_110_49_pad_groupi_n_375;
  wire csa_tree_add_110_49_pad_groupi_n_376, csa_tree_add_110_49_pad_groupi_n_377, csa_tree_add_110_49_pad_groupi_n_378, csa_tree_add_110_49_pad_groupi_n_379, csa_tree_add_110_49_pad_groupi_n_380, csa_tree_add_110_49_pad_groupi_n_381, csa_tree_add_110_49_pad_groupi_n_382, csa_tree_add_110_49_pad_groupi_n_383;
  wire csa_tree_add_110_49_pad_groupi_n_384, csa_tree_add_110_49_pad_groupi_n_385, csa_tree_add_110_49_pad_groupi_n_386, csa_tree_add_110_49_pad_groupi_n_387, csa_tree_add_110_49_pad_groupi_n_388, csa_tree_add_110_49_pad_groupi_n_389, csa_tree_add_110_49_pad_groupi_n_390, csa_tree_add_110_49_pad_groupi_n_391;
  wire csa_tree_add_110_49_pad_groupi_n_392, csa_tree_add_110_49_pad_groupi_n_393, csa_tree_add_110_49_pad_groupi_n_394, csa_tree_add_110_49_pad_groupi_n_395, csa_tree_add_110_49_pad_groupi_n_396, csa_tree_add_110_49_pad_groupi_n_397, csa_tree_add_110_49_pad_groupi_n_398, csa_tree_add_110_49_pad_groupi_n_399;
  wire csa_tree_add_110_49_pad_groupi_n_400, csa_tree_add_110_49_pad_groupi_n_401, csa_tree_add_110_49_pad_groupi_n_402, csa_tree_add_110_49_pad_groupi_n_403, csa_tree_add_110_49_pad_groupi_n_404, csa_tree_add_110_49_pad_groupi_n_405, csa_tree_add_110_49_pad_groupi_n_406, csa_tree_add_110_49_pad_groupi_n_407;
  wire csa_tree_add_110_49_pad_groupi_n_408, csa_tree_add_110_49_pad_groupi_n_409, csa_tree_add_110_49_pad_groupi_n_410, csa_tree_add_110_49_pad_groupi_n_411, csa_tree_add_110_49_pad_groupi_n_412, csa_tree_add_110_49_pad_groupi_n_413, csa_tree_add_110_49_pad_groupi_n_414, csa_tree_add_110_49_pad_groupi_n_415;
  wire csa_tree_add_110_49_pad_groupi_n_416, csa_tree_add_110_49_pad_groupi_n_417, csa_tree_add_110_49_pad_groupi_n_418, csa_tree_add_110_49_pad_groupi_n_419, csa_tree_add_110_49_pad_groupi_n_420, csa_tree_add_110_49_pad_groupi_n_421, csa_tree_add_110_49_pad_groupi_n_422, csa_tree_add_110_49_pad_groupi_n_423;
  wire csa_tree_add_110_49_pad_groupi_n_424, csa_tree_add_110_49_pad_groupi_n_425, csa_tree_add_110_49_pad_groupi_n_426, csa_tree_add_110_49_pad_groupi_n_427, csa_tree_add_110_49_pad_groupi_n_428, csa_tree_add_110_49_pad_groupi_n_429, csa_tree_add_110_49_pad_groupi_n_430, csa_tree_add_110_49_pad_groupi_n_431;
  wire csa_tree_add_110_49_pad_groupi_n_432, csa_tree_add_110_49_pad_groupi_n_433, csa_tree_add_110_49_pad_groupi_n_434, csa_tree_add_110_49_pad_groupi_n_435, csa_tree_add_110_49_pad_groupi_n_436, csa_tree_add_110_49_pad_groupi_n_437, csa_tree_add_110_49_pad_groupi_n_438, csa_tree_add_110_49_pad_groupi_n_439;
  wire csa_tree_add_110_49_pad_groupi_n_440, csa_tree_add_110_49_pad_groupi_n_441, csa_tree_add_110_49_pad_groupi_n_442, csa_tree_add_110_49_pad_groupi_n_443, csa_tree_add_110_49_pad_groupi_n_444, csa_tree_add_110_49_pad_groupi_n_445, csa_tree_add_110_49_pad_groupi_n_446, csa_tree_add_110_49_pad_groupi_n_447;
  wire csa_tree_add_110_49_pad_groupi_n_448, csa_tree_add_110_49_pad_groupi_n_449, csa_tree_add_110_49_pad_groupi_n_450, csa_tree_add_110_49_pad_groupi_n_451, csa_tree_add_110_49_pad_groupi_n_452, csa_tree_add_110_49_pad_groupi_n_453, csa_tree_add_110_49_pad_groupi_n_454, csa_tree_add_110_49_pad_groupi_n_455;
  wire csa_tree_add_110_49_pad_groupi_n_456, csa_tree_add_110_49_pad_groupi_n_457, csa_tree_add_110_49_pad_groupi_n_458, csa_tree_add_110_49_pad_groupi_n_459, csa_tree_add_110_49_pad_groupi_n_460, csa_tree_add_110_49_pad_groupi_n_461, csa_tree_add_110_49_pad_groupi_n_462, csa_tree_add_110_49_pad_groupi_n_463;
  wire csa_tree_add_110_49_pad_groupi_n_464, csa_tree_add_110_49_pad_groupi_n_465, csa_tree_add_110_49_pad_groupi_n_466, csa_tree_add_110_49_pad_groupi_n_467, csa_tree_add_110_49_pad_groupi_n_468, csa_tree_add_110_49_pad_groupi_n_469, csa_tree_add_110_49_pad_groupi_n_470, csa_tree_add_110_49_pad_groupi_n_471;
  wire csa_tree_add_110_49_pad_groupi_n_472, csa_tree_add_110_49_pad_groupi_n_473, csa_tree_add_110_49_pad_groupi_n_474, csa_tree_add_110_49_pad_groupi_n_475, csa_tree_add_110_49_pad_groupi_n_476, csa_tree_add_110_49_pad_groupi_n_477, csa_tree_add_110_49_pad_groupi_n_478, csa_tree_add_110_49_pad_groupi_n_479;
  wire csa_tree_add_110_49_pad_groupi_n_480, csa_tree_add_110_49_pad_groupi_n_481, csa_tree_add_110_49_pad_groupi_n_482, csa_tree_add_110_49_pad_groupi_n_483, csa_tree_add_110_49_pad_groupi_n_484, csa_tree_add_110_49_pad_groupi_n_485, csa_tree_add_110_49_pad_groupi_n_486, csa_tree_add_110_49_pad_groupi_n_487;
  wire csa_tree_add_110_49_pad_groupi_n_488, csa_tree_add_110_49_pad_groupi_n_489, csa_tree_add_110_49_pad_groupi_n_490, csa_tree_add_110_49_pad_groupi_n_491, csa_tree_add_110_49_pad_groupi_n_492, csa_tree_add_110_49_pad_groupi_n_493, csa_tree_add_110_49_pad_groupi_n_494, csa_tree_add_110_49_pad_groupi_n_495;
  wire csa_tree_add_110_49_pad_groupi_n_496, csa_tree_add_110_49_pad_groupi_n_497, csa_tree_add_110_49_pad_groupi_n_498, csa_tree_add_110_49_pad_groupi_n_499, csa_tree_add_110_49_pad_groupi_n_500, csa_tree_add_110_49_pad_groupi_n_501, csa_tree_add_110_49_pad_groupi_n_502, csa_tree_add_110_49_pad_groupi_n_503;
  wire csa_tree_add_110_49_pad_groupi_n_504, csa_tree_add_110_49_pad_groupi_n_505, csa_tree_add_110_49_pad_groupi_n_506, csa_tree_add_110_49_pad_groupi_n_507, csa_tree_add_110_49_pad_groupi_n_508, csa_tree_add_110_49_pad_groupi_n_509, csa_tree_add_110_49_pad_groupi_n_510, csa_tree_add_110_49_pad_groupi_n_511;
  wire csa_tree_add_110_49_pad_groupi_n_512, csa_tree_add_110_49_pad_groupi_n_513, csa_tree_add_110_49_pad_groupi_n_514, csa_tree_add_110_49_pad_groupi_n_515, csa_tree_add_110_49_pad_groupi_n_516, csa_tree_add_110_49_pad_groupi_n_517, csa_tree_add_110_49_pad_groupi_n_518, csa_tree_add_110_49_pad_groupi_n_519;
  wire csa_tree_add_110_49_pad_groupi_n_520, csa_tree_add_110_49_pad_groupi_n_521, csa_tree_add_110_49_pad_groupi_n_522, csa_tree_add_110_49_pad_groupi_n_523, csa_tree_add_110_49_pad_groupi_n_524, csa_tree_add_110_49_pad_groupi_n_525, csa_tree_add_110_49_pad_groupi_n_526, csa_tree_add_110_49_pad_groupi_n_527;
  wire csa_tree_add_110_49_pad_groupi_n_528, csa_tree_add_110_49_pad_groupi_n_529, csa_tree_add_110_49_pad_groupi_n_530, csa_tree_add_110_49_pad_groupi_n_531, csa_tree_add_110_49_pad_groupi_n_532, csa_tree_add_110_49_pad_groupi_n_533, csa_tree_add_110_49_pad_groupi_n_534, csa_tree_add_110_49_pad_groupi_n_535;
  wire csa_tree_add_110_49_pad_groupi_n_536, csa_tree_add_110_49_pad_groupi_n_537, csa_tree_add_110_49_pad_groupi_n_538, csa_tree_add_110_49_pad_groupi_n_539, csa_tree_add_110_49_pad_groupi_n_540, csa_tree_add_110_49_pad_groupi_n_541, csa_tree_add_110_49_pad_groupi_n_542, csa_tree_add_110_49_pad_groupi_n_543;
  wire csa_tree_add_110_49_pad_groupi_n_544, csa_tree_add_110_49_pad_groupi_n_545, csa_tree_add_110_49_pad_groupi_n_546, csa_tree_add_110_49_pad_groupi_n_547, csa_tree_add_110_49_pad_groupi_n_548, csa_tree_add_110_49_pad_groupi_n_549, csa_tree_add_110_49_pad_groupi_n_550, csa_tree_add_110_49_pad_groupi_n_551;
  wire csa_tree_add_110_49_pad_groupi_n_552, csa_tree_add_110_49_pad_groupi_n_553, csa_tree_add_110_49_pad_groupi_n_554, csa_tree_add_110_49_pad_groupi_n_555, csa_tree_add_110_49_pad_groupi_n_556, csa_tree_add_110_49_pad_groupi_n_557, csa_tree_add_110_49_pad_groupi_n_558, csa_tree_add_110_49_pad_groupi_n_559;
  wire csa_tree_add_110_49_pad_groupi_n_560, csa_tree_add_110_49_pad_groupi_n_561, csa_tree_add_110_49_pad_groupi_n_562, csa_tree_add_110_49_pad_groupi_n_563, csa_tree_add_110_49_pad_groupi_n_564, csa_tree_add_110_49_pad_groupi_n_565, csa_tree_add_110_49_pad_groupi_n_566, csa_tree_add_110_49_pad_groupi_n_567;
  wire csa_tree_add_110_49_pad_groupi_n_568, csa_tree_add_110_49_pad_groupi_n_569, csa_tree_add_110_49_pad_groupi_n_570, csa_tree_add_110_49_pad_groupi_n_571, csa_tree_add_110_49_pad_groupi_n_572, csa_tree_add_110_49_pad_groupi_n_573, csa_tree_add_110_49_pad_groupi_n_574, csa_tree_add_110_49_pad_groupi_n_575;
  wire csa_tree_add_110_49_pad_groupi_n_576, csa_tree_add_110_49_pad_groupi_n_577, csa_tree_add_110_49_pad_groupi_n_578, csa_tree_add_110_49_pad_groupi_n_579, csa_tree_add_110_49_pad_groupi_n_580, csa_tree_add_110_49_pad_groupi_n_581, csa_tree_add_110_49_pad_groupi_n_582, csa_tree_add_110_49_pad_groupi_n_583;
  wire csa_tree_add_110_49_pad_groupi_n_584, csa_tree_add_110_49_pad_groupi_n_585, csa_tree_add_110_49_pad_groupi_n_586, csa_tree_add_110_49_pad_groupi_n_587, csa_tree_add_110_49_pad_groupi_n_588, csa_tree_add_110_49_pad_groupi_n_589, csa_tree_add_110_49_pad_groupi_n_590, csa_tree_add_110_49_pad_groupi_n_591;
  wire csa_tree_add_110_49_pad_groupi_n_592, csa_tree_add_110_49_pad_groupi_n_593, csa_tree_add_110_49_pad_groupi_n_594, csa_tree_add_110_49_pad_groupi_n_595, csa_tree_add_110_49_pad_groupi_n_596, csa_tree_add_110_49_pad_groupi_n_597, csa_tree_add_110_49_pad_groupi_n_598, csa_tree_add_110_49_pad_groupi_n_599;
  wire csa_tree_add_110_49_pad_groupi_n_600, csa_tree_add_110_49_pad_groupi_n_601, csa_tree_add_110_49_pad_groupi_n_602, csa_tree_add_110_49_pad_groupi_n_603, csa_tree_add_110_49_pad_groupi_n_604, csa_tree_add_110_49_pad_groupi_n_605, csa_tree_add_110_49_pad_groupi_n_606, csa_tree_add_110_49_pad_groupi_n_607;
  wire csa_tree_add_110_49_pad_groupi_n_608, csa_tree_add_110_49_pad_groupi_n_609, csa_tree_add_110_49_pad_groupi_n_610, csa_tree_add_110_49_pad_groupi_n_611, csa_tree_add_110_49_pad_groupi_n_612, csa_tree_add_110_49_pad_groupi_n_613, csa_tree_add_110_49_pad_groupi_n_614, csa_tree_add_110_49_pad_groupi_n_615;
  wire csa_tree_add_110_49_pad_groupi_n_616, csa_tree_add_110_49_pad_groupi_n_617, csa_tree_add_110_49_pad_groupi_n_618, csa_tree_add_110_49_pad_groupi_n_619, csa_tree_add_110_49_pad_groupi_n_620, csa_tree_add_110_49_pad_groupi_n_621, csa_tree_add_110_49_pad_groupi_n_622, csa_tree_add_110_49_pad_groupi_n_623;
  wire csa_tree_add_110_49_pad_groupi_n_624, csa_tree_add_110_49_pad_groupi_n_625, csa_tree_add_110_49_pad_groupi_n_626, csa_tree_add_110_49_pad_groupi_n_627, csa_tree_add_110_49_pad_groupi_n_628, csa_tree_add_110_49_pad_groupi_n_629, csa_tree_add_110_49_pad_groupi_n_630, csa_tree_add_110_49_pad_groupi_n_631;
  wire csa_tree_add_110_49_pad_groupi_n_632, csa_tree_add_110_49_pad_groupi_n_633, csa_tree_add_110_49_pad_groupi_n_634, csa_tree_add_110_49_pad_groupi_n_635, csa_tree_add_110_49_pad_groupi_n_636, csa_tree_add_110_49_pad_groupi_n_637, csa_tree_add_110_49_pad_groupi_n_638, csa_tree_add_110_49_pad_groupi_n_639;
  wire csa_tree_add_110_49_pad_groupi_n_640, csa_tree_add_110_49_pad_groupi_n_641, csa_tree_add_110_49_pad_groupi_n_642, csa_tree_add_110_49_pad_groupi_n_643, csa_tree_add_110_49_pad_groupi_n_644, csa_tree_add_110_49_pad_groupi_n_645, csa_tree_add_110_49_pad_groupi_n_646, csa_tree_add_110_49_pad_groupi_n_647;
  wire csa_tree_add_110_49_pad_groupi_n_648, csa_tree_add_110_49_pad_groupi_n_649, csa_tree_add_110_49_pad_groupi_n_650, csa_tree_add_110_49_pad_groupi_n_651, csa_tree_add_110_49_pad_groupi_n_652, csa_tree_add_110_49_pad_groupi_n_653, csa_tree_add_110_49_pad_groupi_n_654, csa_tree_add_110_49_pad_groupi_n_655;
  wire csa_tree_add_110_49_pad_groupi_n_656, csa_tree_add_110_49_pad_groupi_n_657, csa_tree_add_110_49_pad_groupi_n_658, csa_tree_add_110_49_pad_groupi_n_659, csa_tree_add_110_49_pad_groupi_n_660, csa_tree_add_110_49_pad_groupi_n_661, csa_tree_add_110_49_pad_groupi_n_662, csa_tree_add_110_49_pad_groupi_n_663;
  wire csa_tree_add_110_49_pad_groupi_n_664, csa_tree_add_110_49_pad_groupi_n_665, csa_tree_add_110_49_pad_groupi_n_666, csa_tree_add_110_49_pad_groupi_n_667, csa_tree_add_110_49_pad_groupi_n_668, csa_tree_add_110_49_pad_groupi_n_669, csa_tree_add_110_49_pad_groupi_n_670, csa_tree_add_110_49_pad_groupi_n_671;
  wire csa_tree_add_110_49_pad_groupi_n_672, csa_tree_add_110_49_pad_groupi_n_673, csa_tree_add_110_49_pad_groupi_n_674, csa_tree_add_110_49_pad_groupi_n_675, csa_tree_add_110_49_pad_groupi_n_676, csa_tree_add_110_49_pad_groupi_n_677, csa_tree_add_110_49_pad_groupi_n_678, csa_tree_add_110_49_pad_groupi_n_679;
  wire csa_tree_add_110_49_pad_groupi_n_680, csa_tree_add_110_49_pad_groupi_n_681, csa_tree_add_110_49_pad_groupi_n_682, csa_tree_add_110_49_pad_groupi_n_683, csa_tree_add_110_49_pad_groupi_n_684, csa_tree_add_110_49_pad_groupi_n_685, csa_tree_add_110_49_pad_groupi_n_686, csa_tree_add_110_49_pad_groupi_n_687;
  wire csa_tree_add_110_49_pad_groupi_n_688, csa_tree_add_110_49_pad_groupi_n_689, csa_tree_add_110_49_pad_groupi_n_690, csa_tree_add_110_49_pad_groupi_n_691, csa_tree_add_110_49_pad_groupi_n_692, csa_tree_add_110_49_pad_groupi_n_693, csa_tree_add_110_49_pad_groupi_n_694, csa_tree_add_110_49_pad_groupi_n_695;
  wire csa_tree_add_110_49_pad_groupi_n_696, csa_tree_add_110_49_pad_groupi_n_697, csa_tree_add_110_49_pad_groupi_n_698, csa_tree_add_110_49_pad_groupi_n_699, csa_tree_add_110_49_pad_groupi_n_700, csa_tree_add_110_49_pad_groupi_n_701, csa_tree_add_110_49_pad_groupi_n_702, csa_tree_add_110_49_pad_groupi_n_703;
  wire csa_tree_add_110_49_pad_groupi_n_704, csa_tree_add_110_49_pad_groupi_n_705, csa_tree_add_110_49_pad_groupi_n_706, csa_tree_add_110_49_pad_groupi_n_707, csa_tree_add_110_49_pad_groupi_n_708, csa_tree_add_110_49_pad_groupi_n_709, csa_tree_add_110_49_pad_groupi_n_710, csa_tree_add_110_49_pad_groupi_n_711;
  wire csa_tree_add_110_49_pad_groupi_n_712, csa_tree_add_110_49_pad_groupi_n_713, csa_tree_add_110_49_pad_groupi_n_714, csa_tree_add_110_49_pad_groupi_n_715, csa_tree_add_110_49_pad_groupi_n_716, csa_tree_add_110_49_pad_groupi_n_717, csa_tree_add_110_49_pad_groupi_n_718, csa_tree_add_110_49_pad_groupi_n_719;
  wire csa_tree_add_110_49_pad_groupi_n_720, csa_tree_add_110_49_pad_groupi_n_721, csa_tree_add_110_49_pad_groupi_n_722, csa_tree_add_110_49_pad_groupi_n_723, csa_tree_add_110_49_pad_groupi_n_724, csa_tree_add_110_49_pad_groupi_n_725, csa_tree_add_110_49_pad_groupi_n_726, csa_tree_add_110_49_pad_groupi_n_727;
  wire csa_tree_add_110_49_pad_groupi_n_728, csa_tree_add_110_49_pad_groupi_n_729, csa_tree_add_110_49_pad_groupi_n_730, csa_tree_add_110_49_pad_groupi_n_731, csa_tree_add_110_49_pad_groupi_n_732, csa_tree_add_110_49_pad_groupi_n_733, csa_tree_add_110_49_pad_groupi_n_734, csa_tree_add_110_49_pad_groupi_n_735;
  wire csa_tree_add_110_49_pad_groupi_n_736, csa_tree_add_110_49_pad_groupi_n_737, csa_tree_add_110_49_pad_groupi_n_738, csa_tree_add_110_49_pad_groupi_n_739, csa_tree_add_110_49_pad_groupi_n_740, csa_tree_add_110_49_pad_groupi_n_741, csa_tree_add_110_49_pad_groupi_n_742, csa_tree_add_110_49_pad_groupi_n_743;
  wire csa_tree_add_110_49_pad_groupi_n_744, csa_tree_add_110_49_pad_groupi_n_745, csa_tree_add_110_49_pad_groupi_n_746, csa_tree_add_110_49_pad_groupi_n_747, csa_tree_add_110_49_pad_groupi_n_748, csa_tree_add_110_49_pad_groupi_n_749, csa_tree_add_110_49_pad_groupi_n_750, csa_tree_add_110_49_pad_groupi_n_751;
  wire csa_tree_add_110_49_pad_groupi_n_752, csa_tree_add_110_49_pad_groupi_n_753, csa_tree_add_110_49_pad_groupi_n_754, csa_tree_add_110_49_pad_groupi_n_755, csa_tree_add_110_49_pad_groupi_n_756, csa_tree_add_110_49_pad_groupi_n_757, csa_tree_add_110_49_pad_groupi_n_758, csa_tree_add_110_49_pad_groupi_n_759;
  wire csa_tree_add_110_49_pad_groupi_n_760, csa_tree_add_110_49_pad_groupi_n_761, csa_tree_add_110_49_pad_groupi_n_762, csa_tree_add_110_49_pad_groupi_n_763, csa_tree_add_110_49_pad_groupi_n_764, csa_tree_add_110_49_pad_groupi_n_765, csa_tree_add_110_49_pad_groupi_n_766, csa_tree_add_110_49_pad_groupi_n_767;
  wire csa_tree_add_110_49_pad_groupi_n_768, csa_tree_add_110_49_pad_groupi_n_769, csa_tree_add_110_49_pad_groupi_n_770, csa_tree_add_110_49_pad_groupi_n_771, csa_tree_add_110_49_pad_groupi_n_772, csa_tree_add_110_49_pad_groupi_n_773, csa_tree_add_110_49_pad_groupi_n_774, csa_tree_add_110_49_pad_groupi_n_775;
  wire csa_tree_add_110_49_pad_groupi_n_776, csa_tree_add_110_49_pad_groupi_n_777, csa_tree_add_110_49_pad_groupi_n_778, csa_tree_add_110_49_pad_groupi_n_779, csa_tree_add_110_49_pad_groupi_n_780, csa_tree_add_110_49_pad_groupi_n_781, csa_tree_add_110_49_pad_groupi_n_782, csa_tree_add_110_49_pad_groupi_n_783;
  wire csa_tree_add_110_49_pad_groupi_n_784, csa_tree_add_110_49_pad_groupi_n_785, csa_tree_add_110_49_pad_groupi_n_786, csa_tree_add_110_49_pad_groupi_n_787, csa_tree_add_110_49_pad_groupi_n_788, csa_tree_add_110_49_pad_groupi_n_789, csa_tree_add_110_49_pad_groupi_n_790, csa_tree_add_110_49_pad_groupi_n_791;
  wire csa_tree_add_110_49_pad_groupi_n_792, csa_tree_add_110_49_pad_groupi_n_793, csa_tree_add_110_49_pad_groupi_n_794, csa_tree_add_110_49_pad_groupi_n_795, csa_tree_add_110_49_pad_groupi_n_796, csa_tree_add_110_49_pad_groupi_n_797, csa_tree_add_110_49_pad_groupi_n_798, csa_tree_add_110_49_pad_groupi_n_799;
  wire csa_tree_add_110_49_pad_groupi_n_800, csa_tree_add_110_49_pad_groupi_n_801, csa_tree_add_110_49_pad_groupi_n_802, csa_tree_add_110_49_pad_groupi_n_803, csa_tree_add_110_49_pad_groupi_n_804, csa_tree_add_110_49_pad_groupi_n_805, csa_tree_add_110_49_pad_groupi_n_806, csa_tree_add_110_49_pad_groupi_n_807;
  wire csa_tree_add_110_49_pad_groupi_n_808, csa_tree_add_110_49_pad_groupi_n_809, csa_tree_add_110_49_pad_groupi_n_810, csa_tree_add_110_49_pad_groupi_n_811, csa_tree_add_110_49_pad_groupi_n_812, csa_tree_add_110_49_pad_groupi_n_813, csa_tree_add_110_49_pad_groupi_n_814, csa_tree_add_110_49_pad_groupi_n_815;
  wire csa_tree_add_110_49_pad_groupi_n_816, csa_tree_add_110_49_pad_groupi_n_817, csa_tree_add_110_49_pad_groupi_n_818, csa_tree_add_110_49_pad_groupi_n_819, csa_tree_add_110_49_pad_groupi_n_820, csa_tree_add_110_49_pad_groupi_n_821, csa_tree_add_110_49_pad_groupi_n_822, csa_tree_add_110_49_pad_groupi_n_823;
  wire csa_tree_add_110_49_pad_groupi_n_824, csa_tree_add_110_49_pad_groupi_n_825, csa_tree_add_110_49_pad_groupi_n_826, csa_tree_add_110_49_pad_groupi_n_827, csa_tree_add_110_49_pad_groupi_n_828, csa_tree_add_110_49_pad_groupi_n_829, csa_tree_add_110_49_pad_groupi_n_830, csa_tree_add_110_49_pad_groupi_n_831;
  wire csa_tree_add_110_49_pad_groupi_n_832, csa_tree_add_110_49_pad_groupi_n_833, csa_tree_add_110_49_pad_groupi_n_834, csa_tree_add_110_49_pad_groupi_n_835, csa_tree_add_110_49_pad_groupi_n_836, csa_tree_add_110_49_pad_groupi_n_837, csa_tree_add_110_49_pad_groupi_n_838, csa_tree_add_110_49_pad_groupi_n_839;
  wire csa_tree_add_110_49_pad_groupi_n_840, csa_tree_add_110_49_pad_groupi_n_841, csa_tree_add_110_49_pad_groupi_n_842, csa_tree_add_110_49_pad_groupi_n_843, csa_tree_add_110_49_pad_groupi_n_844, csa_tree_add_110_49_pad_groupi_n_845, csa_tree_add_110_49_pad_groupi_n_846, csa_tree_add_110_49_pad_groupi_n_847;
  wire csa_tree_add_110_49_pad_groupi_n_848, csa_tree_add_110_49_pad_groupi_n_849, csa_tree_add_110_49_pad_groupi_n_850, csa_tree_add_110_49_pad_groupi_n_851, csa_tree_add_110_49_pad_groupi_n_852, csa_tree_add_110_49_pad_groupi_n_853, csa_tree_add_110_49_pad_groupi_n_854, csa_tree_add_110_49_pad_groupi_n_855;
  wire csa_tree_add_110_49_pad_groupi_n_856, csa_tree_add_110_49_pad_groupi_n_857, csa_tree_add_110_49_pad_groupi_n_858, csa_tree_add_110_49_pad_groupi_n_859, csa_tree_add_110_49_pad_groupi_n_860, csa_tree_add_110_49_pad_groupi_n_861, csa_tree_add_110_49_pad_groupi_n_862, csa_tree_add_110_49_pad_groupi_n_863;
  wire csa_tree_add_110_49_pad_groupi_n_864, csa_tree_add_110_49_pad_groupi_n_865, csa_tree_add_110_49_pad_groupi_n_866, csa_tree_add_110_49_pad_groupi_n_867, csa_tree_add_110_49_pad_groupi_n_868, csa_tree_add_110_49_pad_groupi_n_869, csa_tree_add_110_49_pad_groupi_n_870, csa_tree_add_110_49_pad_groupi_n_871;
  wire csa_tree_add_110_49_pad_groupi_n_872, csa_tree_add_110_49_pad_groupi_n_873, csa_tree_add_110_49_pad_groupi_n_874, csa_tree_add_110_49_pad_groupi_n_875, csa_tree_add_110_49_pad_groupi_n_876, csa_tree_add_110_49_pad_groupi_n_877, csa_tree_add_110_49_pad_groupi_n_878, csa_tree_add_110_49_pad_groupi_n_879;
  wire csa_tree_add_110_49_pad_groupi_n_880, csa_tree_add_110_49_pad_groupi_n_881, csa_tree_add_110_49_pad_groupi_n_882, csa_tree_add_110_49_pad_groupi_n_883, csa_tree_add_110_49_pad_groupi_n_884, csa_tree_add_110_49_pad_groupi_n_885, csa_tree_add_110_49_pad_groupi_n_886, csa_tree_add_110_49_pad_groupi_n_887;
  wire csa_tree_add_110_49_pad_groupi_n_888, csa_tree_add_110_49_pad_groupi_n_889, csa_tree_add_110_49_pad_groupi_n_890, csa_tree_add_110_49_pad_groupi_n_891, csa_tree_add_110_49_pad_groupi_n_892, csa_tree_add_110_49_pad_groupi_n_893, csa_tree_add_110_49_pad_groupi_n_894, csa_tree_add_110_49_pad_groupi_n_895;
  wire csa_tree_add_110_49_pad_groupi_n_896, csa_tree_add_110_49_pad_groupi_n_897, csa_tree_add_110_49_pad_groupi_n_898, csa_tree_add_110_49_pad_groupi_n_899, csa_tree_add_110_49_pad_groupi_n_900, csa_tree_add_110_49_pad_groupi_n_901, csa_tree_add_110_49_pad_groupi_n_902, csa_tree_add_110_49_pad_groupi_n_903;
  wire csa_tree_add_110_49_pad_groupi_n_904, csa_tree_add_110_49_pad_groupi_n_905, csa_tree_add_110_49_pad_groupi_n_906, csa_tree_add_110_49_pad_groupi_n_907, csa_tree_add_110_49_pad_groupi_n_908, csa_tree_add_110_49_pad_groupi_n_909, csa_tree_add_110_49_pad_groupi_n_910, csa_tree_add_110_49_pad_groupi_n_911;
  wire csa_tree_add_110_49_pad_groupi_n_912, csa_tree_add_110_49_pad_groupi_n_913, csa_tree_add_110_49_pad_groupi_n_914, csa_tree_add_110_49_pad_groupi_n_915, csa_tree_add_110_49_pad_groupi_n_916, csa_tree_add_110_49_pad_groupi_n_917, csa_tree_add_110_49_pad_groupi_n_918, csa_tree_add_110_49_pad_groupi_n_919;
  wire csa_tree_add_110_49_pad_groupi_n_920, csa_tree_add_110_49_pad_groupi_n_921, csa_tree_add_110_49_pad_groupi_n_922, csa_tree_add_110_49_pad_groupi_n_923, csa_tree_add_110_49_pad_groupi_n_924, csa_tree_add_110_49_pad_groupi_n_925, csa_tree_add_110_49_pad_groupi_n_926, csa_tree_add_110_49_pad_groupi_n_927;
  wire csa_tree_add_110_49_pad_groupi_n_928, csa_tree_add_110_49_pad_groupi_n_929, csa_tree_add_110_49_pad_groupi_n_930, csa_tree_add_110_49_pad_groupi_n_931, csa_tree_add_110_49_pad_groupi_n_932, csa_tree_add_110_49_pad_groupi_n_933, csa_tree_add_110_49_pad_groupi_n_934, csa_tree_add_110_49_pad_groupi_n_935;
  wire csa_tree_add_110_49_pad_groupi_n_936, csa_tree_add_110_49_pad_groupi_n_937, csa_tree_add_110_49_pad_groupi_n_938, csa_tree_add_110_49_pad_groupi_n_939, csa_tree_add_110_49_pad_groupi_n_940, csa_tree_add_110_49_pad_groupi_n_941, csa_tree_add_110_49_pad_groupi_n_942, csa_tree_add_110_49_pad_groupi_n_943;
  wire csa_tree_add_110_49_pad_groupi_n_944, csa_tree_add_110_49_pad_groupi_n_945, csa_tree_add_110_49_pad_groupi_n_946, csa_tree_add_110_49_pad_groupi_n_947, csa_tree_add_110_49_pad_groupi_n_948, csa_tree_add_110_49_pad_groupi_n_949, csa_tree_add_110_49_pad_groupi_n_950, csa_tree_add_110_49_pad_groupi_n_951;
  wire csa_tree_add_110_49_pad_groupi_n_952, csa_tree_add_110_49_pad_groupi_n_953, csa_tree_add_110_49_pad_groupi_n_954, csa_tree_add_110_49_pad_groupi_n_955, csa_tree_add_110_49_pad_groupi_n_956, csa_tree_add_110_49_pad_groupi_n_957, csa_tree_add_110_49_pad_groupi_n_958, csa_tree_add_110_49_pad_groupi_n_959;
  wire csa_tree_add_110_49_pad_groupi_n_960, csa_tree_add_110_49_pad_groupi_n_961, csa_tree_add_110_49_pad_groupi_n_962, csa_tree_add_110_49_pad_groupi_n_963, csa_tree_add_110_49_pad_groupi_n_964, csa_tree_add_110_49_pad_groupi_n_965, csa_tree_add_110_49_pad_groupi_n_966, csa_tree_add_110_49_pad_groupi_n_967;
  wire csa_tree_add_110_49_pad_groupi_n_968, csa_tree_add_110_49_pad_groupi_n_969, csa_tree_add_110_49_pad_groupi_n_970, csa_tree_add_110_49_pad_groupi_n_971, csa_tree_add_110_49_pad_groupi_n_972, csa_tree_add_110_49_pad_groupi_n_973, csa_tree_add_110_49_pad_groupi_n_974, csa_tree_add_110_49_pad_groupi_n_975;
  wire csa_tree_add_110_49_pad_groupi_n_976, csa_tree_add_110_49_pad_groupi_n_977, csa_tree_add_110_49_pad_groupi_n_978, csa_tree_add_110_49_pad_groupi_n_979, csa_tree_add_110_49_pad_groupi_n_980, csa_tree_add_110_49_pad_groupi_n_981, csa_tree_add_110_49_pad_groupi_n_982, csa_tree_add_110_49_pad_groupi_n_983;
  wire csa_tree_add_110_49_pad_groupi_n_984, csa_tree_add_110_49_pad_groupi_n_985, csa_tree_add_110_49_pad_groupi_n_986, csa_tree_add_110_49_pad_groupi_n_987, csa_tree_add_110_49_pad_groupi_n_988, csa_tree_add_110_49_pad_groupi_n_989, csa_tree_add_110_49_pad_groupi_n_990, csa_tree_add_110_49_pad_groupi_n_991;
  wire csa_tree_add_110_49_pad_groupi_n_992, csa_tree_add_110_49_pad_groupi_n_993, csa_tree_add_110_49_pad_groupi_n_994, csa_tree_add_110_49_pad_groupi_n_995, csa_tree_add_110_49_pad_groupi_n_996, csa_tree_add_110_49_pad_groupi_n_997, csa_tree_add_110_49_pad_groupi_n_998, csa_tree_add_110_49_pad_groupi_n_999;
  wire csa_tree_add_110_49_pad_groupi_n_1000, csa_tree_add_110_49_pad_groupi_n_1001, csa_tree_add_110_49_pad_groupi_n_1002, csa_tree_add_110_49_pad_groupi_n_1003, csa_tree_add_110_49_pad_groupi_n_1004, csa_tree_add_110_49_pad_groupi_n_1005, csa_tree_add_110_49_pad_groupi_n_1006, csa_tree_add_110_49_pad_groupi_n_1007;
  wire csa_tree_add_110_49_pad_groupi_n_1008, csa_tree_add_110_49_pad_groupi_n_1009, csa_tree_add_110_49_pad_groupi_n_1010, csa_tree_add_110_49_pad_groupi_n_1011, csa_tree_add_110_49_pad_groupi_n_1012, csa_tree_add_110_49_pad_groupi_n_1013, csa_tree_add_110_49_pad_groupi_n_1014, csa_tree_add_110_49_pad_groupi_n_1015;
  wire csa_tree_add_110_49_pad_groupi_n_1016, csa_tree_add_110_49_pad_groupi_n_1017, csa_tree_add_110_49_pad_groupi_n_1018, csa_tree_add_110_49_pad_groupi_n_1019, csa_tree_add_110_49_pad_groupi_n_1020, csa_tree_add_110_49_pad_groupi_n_1021, csa_tree_add_110_49_pad_groupi_n_1022, csa_tree_add_110_49_pad_groupi_n_1023;
  wire csa_tree_add_110_49_pad_groupi_n_1024, csa_tree_add_110_49_pad_groupi_n_1025, csa_tree_add_110_49_pad_groupi_n_1026, csa_tree_add_110_49_pad_groupi_n_1027, csa_tree_add_110_49_pad_groupi_n_1028, csa_tree_add_110_49_pad_groupi_n_1029, csa_tree_add_110_49_pad_groupi_n_1030, csa_tree_add_110_49_pad_groupi_n_1031;
  wire csa_tree_add_110_49_pad_groupi_n_1032, csa_tree_add_110_49_pad_groupi_n_1033, csa_tree_add_110_49_pad_groupi_n_1034, csa_tree_add_110_49_pad_groupi_n_1035, csa_tree_add_110_49_pad_groupi_n_1036, csa_tree_add_110_49_pad_groupi_n_1037, csa_tree_add_110_49_pad_groupi_n_1038, csa_tree_add_110_49_pad_groupi_n_1039;
  wire csa_tree_add_110_49_pad_groupi_n_1040, csa_tree_add_110_49_pad_groupi_n_1041, csa_tree_add_110_49_pad_groupi_n_1042, csa_tree_add_110_49_pad_groupi_n_1043, csa_tree_add_110_49_pad_groupi_n_1044, csa_tree_add_110_49_pad_groupi_n_1045, csa_tree_add_110_49_pad_groupi_n_1046, csa_tree_add_110_49_pad_groupi_n_1047;
  wire csa_tree_add_110_49_pad_groupi_n_1048, csa_tree_add_110_49_pad_groupi_n_1049, csa_tree_add_110_49_pad_groupi_n_1050, csa_tree_add_110_49_pad_groupi_n_1051, csa_tree_add_110_49_pad_groupi_n_1052, csa_tree_add_110_49_pad_groupi_n_1053, csa_tree_add_110_49_pad_groupi_n_1054, csa_tree_add_110_49_pad_groupi_n_1055;
  wire csa_tree_add_110_49_pad_groupi_n_1056, csa_tree_add_110_49_pad_groupi_n_1057, csa_tree_add_110_49_pad_groupi_n_1058, csa_tree_add_110_49_pad_groupi_n_1059, csa_tree_add_110_49_pad_groupi_n_1060, csa_tree_add_110_49_pad_groupi_n_1061, csa_tree_add_110_49_pad_groupi_n_1062, csa_tree_add_110_49_pad_groupi_n_1063;
  wire csa_tree_add_110_49_pad_groupi_n_1064, csa_tree_add_110_49_pad_groupi_n_1065, csa_tree_add_110_49_pad_groupi_n_1066, csa_tree_add_110_49_pad_groupi_n_1067, csa_tree_add_110_49_pad_groupi_n_1068, csa_tree_add_110_49_pad_groupi_n_1069, csa_tree_add_110_49_pad_groupi_n_1070, csa_tree_add_110_49_pad_groupi_n_1071;
  wire csa_tree_add_110_49_pad_groupi_n_1072, csa_tree_add_110_49_pad_groupi_n_1073, csa_tree_add_110_49_pad_groupi_n_1074, csa_tree_add_110_49_pad_groupi_n_1075, csa_tree_add_110_49_pad_groupi_n_1076, csa_tree_add_110_49_pad_groupi_n_1077, csa_tree_add_110_49_pad_groupi_n_1078, csa_tree_add_110_49_pad_groupi_n_1079;
  wire csa_tree_add_110_49_pad_groupi_n_1080, csa_tree_add_110_49_pad_groupi_n_1081, csa_tree_add_110_49_pad_groupi_n_1082, csa_tree_add_110_49_pad_groupi_n_1083, csa_tree_add_110_49_pad_groupi_n_1084, csa_tree_add_110_49_pad_groupi_n_1085, csa_tree_add_110_49_pad_groupi_n_1086, csa_tree_add_110_49_pad_groupi_n_1087;
  wire csa_tree_add_110_49_pad_groupi_n_1088, csa_tree_add_110_49_pad_groupi_n_1089, csa_tree_add_110_49_pad_groupi_n_1090, csa_tree_add_110_49_pad_groupi_n_1091, csa_tree_add_110_49_pad_groupi_n_1092, csa_tree_add_110_49_pad_groupi_n_1093, csa_tree_add_110_49_pad_groupi_n_1094, csa_tree_add_110_49_pad_groupi_n_1095;
  wire csa_tree_add_110_49_pad_groupi_n_1096, csa_tree_add_110_49_pad_groupi_n_1097, csa_tree_add_110_49_pad_groupi_n_1098, csa_tree_add_110_49_pad_groupi_n_1099, csa_tree_add_110_49_pad_groupi_n_1100, csa_tree_add_110_49_pad_groupi_n_1101, csa_tree_add_110_49_pad_groupi_n_1102, csa_tree_add_110_49_pad_groupi_n_1103;
  wire csa_tree_add_110_49_pad_groupi_n_1104, csa_tree_add_110_49_pad_groupi_n_1105, csa_tree_add_110_49_pad_groupi_n_1106, csa_tree_add_110_49_pad_groupi_n_1107, csa_tree_add_110_49_pad_groupi_n_1108, csa_tree_add_110_49_pad_groupi_n_1109, csa_tree_add_110_49_pad_groupi_n_1110, csa_tree_add_110_49_pad_groupi_n_1111;
  wire csa_tree_add_110_49_pad_groupi_n_1112, csa_tree_add_110_49_pad_groupi_n_1113, csa_tree_add_110_49_pad_groupi_n_1114, csa_tree_add_110_49_pad_groupi_n_1115, csa_tree_add_110_49_pad_groupi_n_1116, csa_tree_add_110_49_pad_groupi_n_1117, csa_tree_add_110_49_pad_groupi_n_1118, csa_tree_add_110_49_pad_groupi_n_1119;
  wire csa_tree_add_110_49_pad_groupi_n_1120, csa_tree_add_110_49_pad_groupi_n_1121, csa_tree_add_110_49_pad_groupi_n_1122, csa_tree_add_110_49_pad_groupi_n_1123, csa_tree_add_110_49_pad_groupi_n_1124, csa_tree_add_110_49_pad_groupi_n_1125, csa_tree_add_110_49_pad_groupi_n_1126, csa_tree_add_110_49_pad_groupi_n_1127;
  wire csa_tree_add_110_49_pad_groupi_n_1128, csa_tree_add_110_49_pad_groupi_n_1129, csa_tree_add_110_49_pad_groupi_n_1130, csa_tree_add_110_49_pad_groupi_n_1131, csa_tree_add_110_49_pad_groupi_n_1132, csa_tree_add_110_49_pad_groupi_n_1133, csa_tree_add_110_49_pad_groupi_n_1134, csa_tree_add_110_49_pad_groupi_n_1135;
  wire csa_tree_add_110_49_pad_groupi_n_1136, csa_tree_add_110_49_pad_groupi_n_1137, csa_tree_add_110_49_pad_groupi_n_1138, csa_tree_add_110_49_pad_groupi_n_1139, csa_tree_add_110_49_pad_groupi_n_1140, csa_tree_add_110_49_pad_groupi_n_1141, csa_tree_add_110_49_pad_groupi_n_1142, csa_tree_add_110_49_pad_groupi_n_1143;
  wire csa_tree_add_110_49_pad_groupi_n_1144, csa_tree_add_110_49_pad_groupi_n_1145, csa_tree_add_110_49_pad_groupi_n_1146, csa_tree_add_110_49_pad_groupi_n_1147, csa_tree_add_110_49_pad_groupi_n_1148, csa_tree_add_110_49_pad_groupi_n_1149, csa_tree_add_110_49_pad_groupi_n_1150, csa_tree_add_110_49_pad_groupi_n_1151;
  wire csa_tree_add_110_49_pad_groupi_n_1152, csa_tree_add_110_49_pad_groupi_n_1153, csa_tree_add_110_49_pad_groupi_n_1154, csa_tree_add_110_49_pad_groupi_n_1155, csa_tree_add_110_49_pad_groupi_n_1156, csa_tree_add_110_49_pad_groupi_n_1157, csa_tree_add_110_49_pad_groupi_n_1158, csa_tree_add_110_49_pad_groupi_n_1159;
  wire csa_tree_add_110_49_pad_groupi_n_1160, csa_tree_add_110_49_pad_groupi_n_1161, csa_tree_add_110_49_pad_groupi_n_1162, csa_tree_add_110_49_pad_groupi_n_1163, csa_tree_add_110_49_pad_groupi_n_1164, csa_tree_add_110_49_pad_groupi_n_1165, csa_tree_add_110_49_pad_groupi_n_1166, csa_tree_add_110_49_pad_groupi_n_1167;
  wire csa_tree_add_110_49_pad_groupi_n_1168, csa_tree_add_110_49_pad_groupi_n_1169, csa_tree_add_110_49_pad_groupi_n_1170, csa_tree_add_110_49_pad_groupi_n_1171, csa_tree_add_110_49_pad_groupi_n_1172, csa_tree_add_110_49_pad_groupi_n_1173, csa_tree_add_110_49_pad_groupi_n_1174, csa_tree_add_110_49_pad_groupi_n_1175;
  wire csa_tree_add_110_49_pad_groupi_n_1176, csa_tree_add_110_49_pad_groupi_n_1177, csa_tree_add_110_49_pad_groupi_n_1178, csa_tree_add_110_49_pad_groupi_n_1179, csa_tree_add_110_49_pad_groupi_n_1180, csa_tree_add_110_49_pad_groupi_n_1181, csa_tree_add_110_49_pad_groupi_n_1182, csa_tree_add_110_49_pad_groupi_n_1183;
  wire csa_tree_add_110_49_pad_groupi_n_1184, csa_tree_add_110_49_pad_groupi_n_1185, csa_tree_add_110_49_pad_groupi_n_1186, csa_tree_add_110_49_pad_groupi_n_1187, csa_tree_add_110_49_pad_groupi_n_1188, csa_tree_add_110_49_pad_groupi_n_1189, csa_tree_add_110_49_pad_groupi_n_1190, csa_tree_add_110_49_pad_groupi_n_1191;
  wire csa_tree_add_110_49_pad_groupi_n_1192, csa_tree_add_110_49_pad_groupi_n_1193, csa_tree_add_110_49_pad_groupi_n_1194, csa_tree_add_110_49_pad_groupi_n_1195, csa_tree_add_110_49_pad_groupi_n_1196, csa_tree_add_110_49_pad_groupi_n_1197, csa_tree_add_110_49_pad_groupi_n_1198, csa_tree_add_110_49_pad_groupi_n_1199;
  wire csa_tree_add_110_49_pad_groupi_n_1200, csa_tree_add_110_49_pad_groupi_n_1201, csa_tree_add_110_49_pad_groupi_n_1202, csa_tree_add_110_49_pad_groupi_n_1203, csa_tree_add_110_49_pad_groupi_n_1204, csa_tree_add_110_49_pad_groupi_n_1205, csa_tree_add_110_49_pad_groupi_n_1206, csa_tree_add_110_49_pad_groupi_n_1207;
  wire csa_tree_add_110_49_pad_groupi_n_1208, csa_tree_add_110_49_pad_groupi_n_1209, csa_tree_add_110_49_pad_groupi_n_1210, csa_tree_add_110_49_pad_groupi_n_1211, csa_tree_add_110_49_pad_groupi_n_1212, csa_tree_add_110_49_pad_groupi_n_1213, csa_tree_add_110_49_pad_groupi_n_1214, csa_tree_add_110_49_pad_groupi_n_1215;
  wire csa_tree_add_110_49_pad_groupi_n_1216, csa_tree_add_110_49_pad_groupi_n_1217, csa_tree_add_110_49_pad_groupi_n_1218, csa_tree_add_110_49_pad_groupi_n_1219, csa_tree_add_110_49_pad_groupi_n_1220, csa_tree_add_110_49_pad_groupi_n_1221, csa_tree_add_110_49_pad_groupi_n_1222, csa_tree_add_110_49_pad_groupi_n_1223;
  wire csa_tree_add_110_49_pad_groupi_n_1224, csa_tree_add_110_49_pad_groupi_n_1225, csa_tree_add_110_49_pad_groupi_n_1226, csa_tree_add_110_49_pad_groupi_n_1227, csa_tree_add_110_49_pad_groupi_n_1228, csa_tree_add_110_49_pad_groupi_n_1229, csa_tree_add_110_49_pad_groupi_n_1230, csa_tree_add_110_49_pad_groupi_n_1231;
  wire csa_tree_add_110_49_pad_groupi_n_1232, csa_tree_add_110_49_pad_groupi_n_1233, csa_tree_add_110_49_pad_groupi_n_1234, csa_tree_add_110_49_pad_groupi_n_1235, csa_tree_add_110_49_pad_groupi_n_1236, csa_tree_add_110_49_pad_groupi_n_1237, csa_tree_add_110_49_pad_groupi_n_1238, csa_tree_add_110_49_pad_groupi_n_1239;
  wire csa_tree_add_110_49_pad_groupi_n_1240, csa_tree_add_110_49_pad_groupi_n_1241, csa_tree_add_110_49_pad_groupi_n_1242, csa_tree_add_110_49_pad_groupi_n_1243, csa_tree_add_110_49_pad_groupi_n_1244, csa_tree_add_110_49_pad_groupi_n_1245, csa_tree_add_110_49_pad_groupi_n_1246, csa_tree_add_110_49_pad_groupi_n_1247;
  wire csa_tree_add_110_49_pad_groupi_n_1248, csa_tree_add_110_49_pad_groupi_n_1249, csa_tree_add_110_49_pad_groupi_n_1250, csa_tree_add_110_49_pad_groupi_n_1251, csa_tree_add_110_49_pad_groupi_n_1252, csa_tree_add_110_49_pad_groupi_n_1253, csa_tree_add_110_49_pad_groupi_n_1254, csa_tree_add_110_49_pad_groupi_n_1255;
  wire csa_tree_add_110_49_pad_groupi_n_1256, csa_tree_add_110_49_pad_groupi_n_1257, csa_tree_add_110_49_pad_groupi_n_1258, csa_tree_add_110_49_pad_groupi_n_1259, csa_tree_add_110_49_pad_groupi_n_1260, csa_tree_add_110_49_pad_groupi_n_1261, csa_tree_add_110_49_pad_groupi_n_1262, csa_tree_add_110_49_pad_groupi_n_1263;
  wire csa_tree_add_110_49_pad_groupi_n_1264, csa_tree_add_110_49_pad_groupi_n_1265, csa_tree_add_110_49_pad_groupi_n_1266, csa_tree_add_110_49_pad_groupi_n_1267, csa_tree_add_110_49_pad_groupi_n_1268, csa_tree_add_110_49_pad_groupi_n_1269, csa_tree_add_110_49_pad_groupi_n_1270, csa_tree_add_110_49_pad_groupi_n_1271;
  wire csa_tree_add_110_49_pad_groupi_n_1272, csa_tree_add_110_49_pad_groupi_n_1273, csa_tree_add_110_49_pad_groupi_n_1274, csa_tree_add_110_49_pad_groupi_n_1275, csa_tree_add_110_49_pad_groupi_n_1276, csa_tree_add_110_49_pad_groupi_n_1277, csa_tree_add_110_49_pad_groupi_n_1278, csa_tree_add_110_49_pad_groupi_n_1279;
  wire csa_tree_add_110_49_pad_groupi_n_1280, csa_tree_add_110_49_pad_groupi_n_1281, csa_tree_add_110_49_pad_groupi_n_1282, csa_tree_add_110_49_pad_groupi_n_1283, csa_tree_add_110_49_pad_groupi_n_1284, csa_tree_add_110_49_pad_groupi_n_1285, csa_tree_add_110_49_pad_groupi_n_1286, csa_tree_add_110_49_pad_groupi_n_1287;
  wire csa_tree_add_110_49_pad_groupi_n_1288, csa_tree_add_110_49_pad_groupi_n_1289, csa_tree_add_110_49_pad_groupi_n_1290, csa_tree_add_110_49_pad_groupi_n_1291, csa_tree_add_110_49_pad_groupi_n_1292, csa_tree_add_110_49_pad_groupi_n_1293, csa_tree_add_110_49_pad_groupi_n_1294, csa_tree_add_110_49_pad_groupi_n_1295;
  wire csa_tree_add_110_49_pad_groupi_n_1296, csa_tree_add_110_49_pad_groupi_n_1297, csa_tree_add_110_49_pad_groupi_n_1298, csa_tree_add_110_49_pad_groupi_n_1299, csa_tree_add_110_49_pad_groupi_n_1300, csa_tree_add_110_49_pad_groupi_n_1301, csa_tree_add_110_49_pad_groupi_n_1302, csa_tree_add_110_49_pad_groupi_n_1303;
  wire csa_tree_add_110_49_pad_groupi_n_1304, csa_tree_add_110_49_pad_groupi_n_1305, csa_tree_add_110_49_pad_groupi_n_1306, csa_tree_add_110_49_pad_groupi_n_1307, csa_tree_add_110_49_pad_groupi_n_1308, csa_tree_add_110_49_pad_groupi_n_1309, csa_tree_add_110_49_pad_groupi_n_1310, csa_tree_add_110_49_pad_groupi_n_1311;
  wire csa_tree_add_110_49_pad_groupi_n_1312, csa_tree_add_110_49_pad_groupi_n_1313, csa_tree_add_110_49_pad_groupi_n_1314, csa_tree_add_110_49_pad_groupi_n_1315, csa_tree_add_110_49_pad_groupi_n_1316, csa_tree_add_110_49_pad_groupi_n_1317, csa_tree_add_110_49_pad_groupi_n_1318, csa_tree_add_110_49_pad_groupi_n_1319;
  wire csa_tree_add_110_49_pad_groupi_n_1320, csa_tree_add_110_49_pad_groupi_n_1321, csa_tree_add_110_49_pad_groupi_n_1322, csa_tree_add_110_49_pad_groupi_n_1323, csa_tree_add_110_49_pad_groupi_n_1324, csa_tree_add_110_49_pad_groupi_n_1325, csa_tree_add_110_49_pad_groupi_n_1326, csa_tree_add_110_49_pad_groupi_n_1327;
  wire csa_tree_add_110_49_pad_groupi_n_1328, csa_tree_add_110_49_pad_groupi_n_1329, csa_tree_add_110_49_pad_groupi_n_1330, csa_tree_add_110_49_pad_groupi_n_1331, csa_tree_add_110_49_pad_groupi_n_1332, csa_tree_add_110_49_pad_groupi_n_1333, csa_tree_add_110_49_pad_groupi_n_1334, csa_tree_add_110_49_pad_groupi_n_1335;
  wire csa_tree_add_110_49_pad_groupi_n_1336, csa_tree_add_110_49_pad_groupi_n_1337, csa_tree_add_110_49_pad_groupi_n_1338, csa_tree_add_110_49_pad_groupi_n_1339, csa_tree_add_110_49_pad_groupi_n_1340, csa_tree_add_110_49_pad_groupi_n_1341, csa_tree_add_110_49_pad_groupi_n_1342, csa_tree_add_110_49_pad_groupi_n_1343;
  wire csa_tree_add_110_49_pad_groupi_n_1344, csa_tree_add_110_49_pad_groupi_n_1345, csa_tree_add_110_49_pad_groupi_n_1346, csa_tree_add_110_49_pad_groupi_n_1347, csa_tree_add_110_49_pad_groupi_n_1348, csa_tree_add_110_49_pad_groupi_n_1349, csa_tree_add_110_49_pad_groupi_n_1350, csa_tree_add_110_49_pad_groupi_n_1351;
  wire csa_tree_add_110_49_pad_groupi_n_1352, csa_tree_add_110_49_pad_groupi_n_1353, csa_tree_add_110_49_pad_groupi_n_1354, csa_tree_add_110_49_pad_groupi_n_1355, csa_tree_add_110_49_pad_groupi_n_1356, csa_tree_add_110_49_pad_groupi_n_1357, csa_tree_add_110_49_pad_groupi_n_1358, csa_tree_add_110_49_pad_groupi_n_1359;
  wire csa_tree_add_110_49_pad_groupi_n_1360, csa_tree_add_110_49_pad_groupi_n_1361, csa_tree_add_110_49_pad_groupi_n_1362, csa_tree_add_110_49_pad_groupi_n_1363, csa_tree_add_110_49_pad_groupi_n_1364, csa_tree_add_110_49_pad_groupi_n_1365, csa_tree_add_110_49_pad_groupi_n_1366, csa_tree_add_110_49_pad_groupi_n_1367;
  wire csa_tree_add_110_49_pad_groupi_n_1368, csa_tree_add_110_49_pad_groupi_n_1369, csa_tree_add_110_49_pad_groupi_n_1370, csa_tree_add_110_49_pad_groupi_n_1371, csa_tree_add_110_49_pad_groupi_n_1372, csa_tree_add_110_49_pad_groupi_n_1373, csa_tree_add_110_49_pad_groupi_n_1374, csa_tree_add_110_49_pad_groupi_n_1375;
  wire csa_tree_add_110_49_pad_groupi_n_1376, csa_tree_add_110_49_pad_groupi_n_1377, csa_tree_add_110_49_pad_groupi_n_1378, csa_tree_add_110_49_pad_groupi_n_1379, csa_tree_add_110_49_pad_groupi_n_1380, csa_tree_add_110_49_pad_groupi_n_1381, csa_tree_add_110_49_pad_groupi_n_1382, csa_tree_add_110_49_pad_groupi_n_1383;
  wire csa_tree_add_110_49_pad_groupi_n_1384, csa_tree_add_110_49_pad_groupi_n_1385, csa_tree_add_110_49_pad_groupi_n_1386, csa_tree_add_110_49_pad_groupi_n_1387, csa_tree_add_110_49_pad_groupi_n_1388, csa_tree_add_110_49_pad_groupi_n_1389, csa_tree_add_110_49_pad_groupi_n_1390, csa_tree_add_110_49_pad_groupi_n_1391;
  wire csa_tree_add_110_49_pad_groupi_n_1392, csa_tree_add_110_49_pad_groupi_n_1393, csa_tree_add_110_49_pad_groupi_n_1394, csa_tree_add_110_49_pad_groupi_n_1395, csa_tree_add_110_49_pad_groupi_n_1396, csa_tree_add_110_49_pad_groupi_n_1397, csa_tree_add_110_49_pad_groupi_n_1398, csa_tree_add_110_49_pad_groupi_n_1399;
  wire csa_tree_add_110_49_pad_groupi_n_1400, csa_tree_add_110_49_pad_groupi_n_1401, csa_tree_add_110_49_pad_groupi_n_1402, csa_tree_add_110_49_pad_groupi_n_1403, csa_tree_add_110_49_pad_groupi_n_1404, csa_tree_add_110_49_pad_groupi_n_1405, csa_tree_add_110_49_pad_groupi_n_1406, csa_tree_add_110_49_pad_groupi_n_1407;
  wire csa_tree_add_110_49_pad_groupi_n_1408, csa_tree_add_110_49_pad_groupi_n_1409, csa_tree_add_110_49_pad_groupi_n_1410, csa_tree_add_110_49_pad_groupi_n_1411, csa_tree_add_110_49_pad_groupi_n_1412, csa_tree_add_110_49_pad_groupi_n_1413, csa_tree_add_110_49_pad_groupi_n_1414, csa_tree_add_110_49_pad_groupi_n_1415;
  wire csa_tree_add_110_49_pad_groupi_n_1416, csa_tree_add_110_49_pad_groupi_n_1417, csa_tree_add_110_49_pad_groupi_n_1418, csa_tree_add_110_49_pad_groupi_n_1419, csa_tree_add_110_49_pad_groupi_n_1420, csa_tree_add_110_49_pad_groupi_n_1421, csa_tree_add_110_49_pad_groupi_n_1422, csa_tree_add_110_49_pad_groupi_n_1423;
  wire csa_tree_add_110_49_pad_groupi_n_1424, csa_tree_add_110_49_pad_groupi_n_1425, csa_tree_add_110_49_pad_groupi_n_1426, csa_tree_add_110_49_pad_groupi_n_1427, csa_tree_add_110_49_pad_groupi_n_1428, csa_tree_add_110_49_pad_groupi_n_1429, csa_tree_add_110_49_pad_groupi_n_1430, csa_tree_add_110_49_pad_groupi_n_1431;
  wire csa_tree_add_110_49_pad_groupi_n_1432, csa_tree_add_110_49_pad_groupi_n_1433, csa_tree_add_110_49_pad_groupi_n_1434, csa_tree_add_110_49_pad_groupi_n_1435, csa_tree_add_110_49_pad_groupi_n_1436, csa_tree_add_110_49_pad_groupi_n_1437, csa_tree_add_110_49_pad_groupi_n_1438, csa_tree_add_110_49_pad_groupi_n_1439;
  wire csa_tree_add_110_49_pad_groupi_n_1440, csa_tree_add_110_49_pad_groupi_n_1441, csa_tree_add_110_49_pad_groupi_n_1442, csa_tree_add_110_49_pad_groupi_n_1443, csa_tree_add_110_49_pad_groupi_n_1444, csa_tree_add_110_49_pad_groupi_n_1445, csa_tree_add_110_49_pad_groupi_n_1446, csa_tree_add_110_49_pad_groupi_n_1447;
  wire csa_tree_add_110_49_pad_groupi_n_1448, csa_tree_add_110_49_pad_groupi_n_1449, csa_tree_add_110_49_pad_groupi_n_1450, csa_tree_add_110_49_pad_groupi_n_1451, csa_tree_add_110_49_pad_groupi_n_1452, csa_tree_add_110_49_pad_groupi_n_1453, csa_tree_add_110_49_pad_groupi_n_1454, csa_tree_add_110_49_pad_groupi_n_1455;
  wire csa_tree_add_110_49_pad_groupi_n_1456, csa_tree_add_110_49_pad_groupi_n_1457, csa_tree_add_110_49_pad_groupi_n_1458, csa_tree_add_110_49_pad_groupi_n_1459, csa_tree_add_110_49_pad_groupi_n_1460, csa_tree_add_110_49_pad_groupi_n_1461, csa_tree_add_110_49_pad_groupi_n_1462, csa_tree_add_110_49_pad_groupi_n_1463;
  wire csa_tree_add_110_49_pad_groupi_n_1464, csa_tree_add_110_49_pad_groupi_n_1465, csa_tree_add_110_49_pad_groupi_n_1466, csa_tree_add_110_49_pad_groupi_n_1467, csa_tree_add_110_49_pad_groupi_n_1468, csa_tree_add_110_49_pad_groupi_n_1469, csa_tree_add_110_49_pad_groupi_n_1470, csa_tree_add_110_49_pad_groupi_n_1471;
  wire csa_tree_add_110_49_pad_groupi_n_1472, csa_tree_add_110_49_pad_groupi_n_1473, csa_tree_add_110_49_pad_groupi_n_1474, csa_tree_add_110_49_pad_groupi_n_1475, csa_tree_add_110_49_pad_groupi_n_1476, csa_tree_add_110_49_pad_groupi_n_1477, csa_tree_add_110_49_pad_groupi_n_1478, csa_tree_add_110_49_pad_groupi_n_1479;
  wire csa_tree_add_110_49_pad_groupi_n_1480, csa_tree_add_110_49_pad_groupi_n_1481, csa_tree_add_110_49_pad_groupi_n_1482, csa_tree_add_110_49_pad_groupi_n_1483, csa_tree_add_110_49_pad_groupi_n_1484, csa_tree_add_110_49_pad_groupi_n_1485, csa_tree_add_110_49_pad_groupi_n_1487, csa_tree_add_110_49_pad_groupi_n_1488;
  wire csa_tree_add_110_49_pad_groupi_n_1489, csa_tree_add_110_49_pad_groupi_n_1490, csa_tree_add_110_49_pad_groupi_n_1491, csa_tree_add_110_49_pad_groupi_n_1492, csa_tree_add_110_49_pad_groupi_n_1493, csa_tree_add_110_49_pad_groupi_n_1494, csa_tree_add_110_49_pad_groupi_n_1495, csa_tree_add_110_49_pad_groupi_n_1496;
  wire csa_tree_add_110_49_pad_groupi_n_1497, csa_tree_add_110_49_pad_groupi_n_1498, csa_tree_add_110_49_pad_groupi_n_1499, csa_tree_add_110_49_pad_groupi_n_1500, csa_tree_add_110_49_pad_groupi_n_1501, csa_tree_add_110_49_pad_groupi_n_1502, csa_tree_add_110_49_pad_groupi_n_1503, csa_tree_add_110_49_pad_groupi_n_1504;
  wire csa_tree_add_110_49_pad_groupi_n_1505, csa_tree_add_110_49_pad_groupi_n_1506, csa_tree_add_110_49_pad_groupi_n_1507, csa_tree_add_110_49_pad_groupi_n_1508, csa_tree_add_110_49_pad_groupi_n_1510, csa_tree_add_110_49_pad_groupi_n_1511, csa_tree_add_110_49_pad_groupi_n_1512, csa_tree_add_110_49_pad_groupi_n_1513;
  wire csa_tree_add_110_49_pad_groupi_n_1514, csa_tree_add_110_49_pad_groupi_n_1515, csa_tree_add_110_49_pad_groupi_n_1516, csa_tree_add_110_49_pad_groupi_n_1517, csa_tree_add_110_49_pad_groupi_n_1518, csa_tree_add_110_49_pad_groupi_n_1519, csa_tree_add_110_49_pad_groupi_n_1521, csa_tree_add_110_49_pad_groupi_n_1522;
  wire csa_tree_add_110_49_pad_groupi_n_1524, csa_tree_add_110_49_pad_groupi_n_1525, csa_tree_add_110_49_pad_groupi_n_1527, csa_tree_add_110_49_pad_groupi_n_1528, csa_tree_add_110_49_pad_groupi_n_1530, csa_tree_add_110_49_pad_groupi_n_1531, csa_tree_add_110_49_pad_groupi_n_1533, csa_tree_add_110_49_pad_groupi_n_1534;
  wire csa_tree_add_110_49_pad_groupi_n_1536, csa_tree_add_110_49_pad_groupi_n_1537, csa_tree_add_110_49_pad_groupi_n_1539, csa_tree_add_110_49_pad_groupi_n_1540, csa_tree_add_110_49_pad_groupi_n_1542, csa_tree_add_110_49_pad_groupi_n_1543, csa_tree_add_110_49_pad_groupi_n_1545, csa_tree_add_110_49_pad_groupi_n_1546;
  wire csa_tree_add_110_49_pad_groupi_n_1548, csa_tree_add_110_49_pad_groupi_n_1549, csa_tree_add_110_49_pad_groupi_n_1550, csa_tree_add_110_49_pad_groupi_n_1551, csa_tree_add_110_49_pad_groupi_n_1552, csa_tree_add_110_49_pad_groupi_n_1553, csa_tree_add_110_49_pad_groupi_n_1555, csa_tree_add_117_21_pad_groupi_n_0;
  wire csa_tree_add_117_21_pad_groupi_n_1, csa_tree_add_117_21_pad_groupi_n_2, csa_tree_add_117_21_pad_groupi_n_3, csa_tree_add_117_21_pad_groupi_n_4, csa_tree_add_117_21_pad_groupi_n_5, csa_tree_add_117_21_pad_groupi_n_6, csa_tree_add_117_21_pad_groupi_n_7, csa_tree_add_117_21_pad_groupi_n_8;
  wire csa_tree_add_117_21_pad_groupi_n_9, csa_tree_add_117_21_pad_groupi_n_10, csa_tree_add_117_21_pad_groupi_n_11, csa_tree_add_117_21_pad_groupi_n_12, csa_tree_add_117_21_pad_groupi_n_13, csa_tree_add_117_21_pad_groupi_n_14, csa_tree_add_117_21_pad_groupi_n_15, csa_tree_add_117_21_pad_groupi_n_16;
  wire csa_tree_add_117_21_pad_groupi_n_17, csa_tree_add_117_21_pad_groupi_n_18, csa_tree_add_117_21_pad_groupi_n_19, csa_tree_add_117_21_pad_groupi_n_20, csa_tree_add_117_21_pad_groupi_n_21, csa_tree_add_117_21_pad_groupi_n_22, csa_tree_add_117_21_pad_groupi_n_23, csa_tree_add_117_21_pad_groupi_n_24;
  wire csa_tree_add_117_21_pad_groupi_n_25, csa_tree_add_117_21_pad_groupi_n_26, csa_tree_add_117_21_pad_groupi_n_27, csa_tree_add_117_21_pad_groupi_n_28, csa_tree_add_117_21_pad_groupi_n_29, csa_tree_add_117_21_pad_groupi_n_30, csa_tree_add_117_21_pad_groupi_n_31, csa_tree_add_117_21_pad_groupi_n_32;
  wire csa_tree_add_117_21_pad_groupi_n_33, csa_tree_add_117_21_pad_groupi_n_34, csa_tree_add_117_21_pad_groupi_n_35, csa_tree_add_117_21_pad_groupi_n_36, csa_tree_add_117_21_pad_groupi_n_37, csa_tree_add_117_21_pad_groupi_n_38, csa_tree_add_117_21_pad_groupi_n_39, csa_tree_add_117_21_pad_groupi_n_40;
  wire csa_tree_add_117_21_pad_groupi_n_41, csa_tree_add_117_21_pad_groupi_n_42, csa_tree_add_117_21_pad_groupi_n_43, csa_tree_add_117_21_pad_groupi_n_44, csa_tree_add_117_21_pad_groupi_n_45, csa_tree_add_117_21_pad_groupi_n_46, csa_tree_add_117_21_pad_groupi_n_47, csa_tree_add_117_21_pad_groupi_n_48;
  wire csa_tree_add_117_21_pad_groupi_n_49, csa_tree_add_117_21_pad_groupi_n_50, csa_tree_add_117_21_pad_groupi_n_51, csa_tree_add_117_21_pad_groupi_n_52, csa_tree_add_117_21_pad_groupi_n_53, csa_tree_add_117_21_pad_groupi_n_54, csa_tree_add_117_21_pad_groupi_n_55, csa_tree_add_117_21_pad_groupi_n_56;
  wire csa_tree_add_117_21_pad_groupi_n_57, csa_tree_add_117_21_pad_groupi_n_58, csa_tree_add_117_21_pad_groupi_n_59, csa_tree_add_117_21_pad_groupi_n_60, csa_tree_add_117_21_pad_groupi_n_61, csa_tree_add_117_21_pad_groupi_n_62, csa_tree_add_117_21_pad_groupi_n_63, csa_tree_add_117_21_pad_groupi_n_64;
  wire csa_tree_add_117_21_pad_groupi_n_65, csa_tree_add_117_21_pad_groupi_n_66, csa_tree_add_117_21_pad_groupi_n_67, csa_tree_add_117_21_pad_groupi_n_68, csa_tree_add_117_21_pad_groupi_n_69, csa_tree_add_117_21_pad_groupi_n_70, csa_tree_add_117_21_pad_groupi_n_71, csa_tree_add_117_21_pad_groupi_n_72;
  wire csa_tree_add_117_21_pad_groupi_n_73, csa_tree_add_117_21_pad_groupi_n_74, csa_tree_add_117_21_pad_groupi_n_75, csa_tree_add_117_21_pad_groupi_n_76, csa_tree_add_117_21_pad_groupi_n_77, csa_tree_add_117_21_pad_groupi_n_78, csa_tree_add_117_21_pad_groupi_n_79, csa_tree_add_117_21_pad_groupi_n_80;
  wire csa_tree_add_117_21_pad_groupi_n_81, csa_tree_add_117_21_pad_groupi_n_82, csa_tree_add_117_21_pad_groupi_n_83, csa_tree_add_117_21_pad_groupi_n_84, csa_tree_add_117_21_pad_groupi_n_85, csa_tree_add_117_21_pad_groupi_n_86, csa_tree_add_117_21_pad_groupi_n_87, csa_tree_add_117_21_pad_groupi_n_88;
  wire csa_tree_add_117_21_pad_groupi_n_89, csa_tree_add_117_21_pad_groupi_n_90, csa_tree_add_117_21_pad_groupi_n_91, csa_tree_add_117_21_pad_groupi_n_92, csa_tree_add_117_21_pad_groupi_n_93, csa_tree_add_117_21_pad_groupi_n_94, csa_tree_add_117_21_pad_groupi_n_95, csa_tree_add_117_21_pad_groupi_n_96;
  wire csa_tree_add_117_21_pad_groupi_n_97, csa_tree_add_117_21_pad_groupi_n_98, csa_tree_add_117_21_pad_groupi_n_99, csa_tree_add_117_21_pad_groupi_n_100, csa_tree_add_117_21_pad_groupi_n_101, csa_tree_add_117_21_pad_groupi_n_102, csa_tree_add_117_21_pad_groupi_n_103, csa_tree_add_117_21_pad_groupi_n_104;
  wire csa_tree_add_117_21_pad_groupi_n_105, csa_tree_add_117_21_pad_groupi_n_106, csa_tree_add_117_21_pad_groupi_n_107, csa_tree_add_117_21_pad_groupi_n_108, csa_tree_add_117_21_pad_groupi_n_109, csa_tree_add_117_21_pad_groupi_n_110, csa_tree_add_117_21_pad_groupi_n_111, csa_tree_add_117_21_pad_groupi_n_112;
  wire csa_tree_add_117_21_pad_groupi_n_116, csa_tree_add_117_21_pad_groupi_n_117, csa_tree_add_117_21_pad_groupi_n_118, csa_tree_add_117_21_pad_groupi_n_119, csa_tree_add_117_21_pad_groupi_n_120, csa_tree_add_117_21_pad_groupi_n_121, csa_tree_add_117_21_pad_groupi_n_122, csa_tree_add_117_21_pad_groupi_n_123;
  wire csa_tree_add_117_21_pad_groupi_n_124, csa_tree_add_117_21_pad_groupi_n_125, csa_tree_add_117_21_pad_groupi_n_126, csa_tree_add_117_21_pad_groupi_n_127, csa_tree_add_117_21_pad_groupi_n_128, csa_tree_add_117_21_pad_groupi_n_129, csa_tree_add_117_21_pad_groupi_n_130, csa_tree_add_117_21_pad_groupi_n_131;
  wire csa_tree_add_117_21_pad_groupi_n_132, csa_tree_add_117_21_pad_groupi_n_133, csa_tree_add_117_21_pad_groupi_n_134, csa_tree_add_117_21_pad_groupi_n_135, csa_tree_add_117_21_pad_groupi_n_136, csa_tree_add_117_21_pad_groupi_n_137, csa_tree_add_117_21_pad_groupi_n_138, csa_tree_add_117_21_pad_groupi_n_139;
  wire csa_tree_add_117_21_pad_groupi_n_140, csa_tree_add_117_21_pad_groupi_n_141, csa_tree_add_117_21_pad_groupi_n_142, csa_tree_add_117_21_pad_groupi_n_143, csa_tree_add_117_21_pad_groupi_n_144, csa_tree_add_117_21_pad_groupi_n_145, csa_tree_add_117_21_pad_groupi_n_146, csa_tree_add_117_21_pad_groupi_n_147;
  wire csa_tree_add_117_21_pad_groupi_n_148, csa_tree_add_117_21_pad_groupi_n_149, csa_tree_add_117_21_pad_groupi_n_150, csa_tree_add_117_21_pad_groupi_n_151, csa_tree_add_117_21_pad_groupi_n_152, csa_tree_add_117_21_pad_groupi_n_153, csa_tree_add_117_21_pad_groupi_n_154, csa_tree_add_117_21_pad_groupi_n_155;
  wire csa_tree_add_117_21_pad_groupi_n_156, csa_tree_add_117_21_pad_groupi_n_157, csa_tree_add_117_21_pad_groupi_n_158, csa_tree_add_117_21_pad_groupi_n_159, csa_tree_add_117_21_pad_groupi_n_160, csa_tree_add_117_21_pad_groupi_n_161, csa_tree_add_117_21_pad_groupi_n_162, csa_tree_add_117_21_pad_groupi_n_163;
  wire csa_tree_add_117_21_pad_groupi_n_164, csa_tree_add_117_21_pad_groupi_n_165, csa_tree_add_117_21_pad_groupi_n_166, csa_tree_add_117_21_pad_groupi_n_167, csa_tree_add_117_21_pad_groupi_n_168, csa_tree_add_117_21_pad_groupi_n_169, csa_tree_add_117_21_pad_groupi_n_170, csa_tree_add_117_21_pad_groupi_n_171;
  wire csa_tree_add_117_21_pad_groupi_n_172, csa_tree_add_117_21_pad_groupi_n_173, csa_tree_add_117_21_pad_groupi_n_174, csa_tree_add_117_21_pad_groupi_n_175, csa_tree_add_117_21_pad_groupi_n_176, csa_tree_add_117_21_pad_groupi_n_177, csa_tree_add_117_21_pad_groupi_n_178, csa_tree_add_117_21_pad_groupi_n_179;
  wire csa_tree_add_117_21_pad_groupi_n_180, csa_tree_add_117_21_pad_groupi_n_181, csa_tree_add_117_21_pad_groupi_n_182, csa_tree_add_117_21_pad_groupi_n_183, csa_tree_add_117_21_pad_groupi_n_184, csa_tree_add_117_21_pad_groupi_n_185, csa_tree_add_117_21_pad_groupi_n_186, csa_tree_add_117_21_pad_groupi_n_187;
  wire csa_tree_add_117_21_pad_groupi_n_188, csa_tree_add_117_21_pad_groupi_n_189, csa_tree_add_117_21_pad_groupi_n_190, csa_tree_add_117_21_pad_groupi_n_191, csa_tree_add_117_21_pad_groupi_n_192, csa_tree_add_117_21_pad_groupi_n_193, csa_tree_add_117_21_pad_groupi_n_194, csa_tree_add_117_21_pad_groupi_n_195;
  wire csa_tree_add_117_21_pad_groupi_n_196, csa_tree_add_117_21_pad_groupi_n_197, csa_tree_add_117_21_pad_groupi_n_198, csa_tree_add_117_21_pad_groupi_n_199, csa_tree_add_117_21_pad_groupi_n_200, csa_tree_add_117_21_pad_groupi_n_201, csa_tree_add_117_21_pad_groupi_n_202, csa_tree_add_117_21_pad_groupi_n_203;
  wire csa_tree_add_117_21_pad_groupi_n_204, csa_tree_add_117_21_pad_groupi_n_205, csa_tree_add_117_21_pad_groupi_n_206, csa_tree_add_117_21_pad_groupi_n_207, csa_tree_add_117_21_pad_groupi_n_208, csa_tree_add_117_21_pad_groupi_n_209, csa_tree_add_117_21_pad_groupi_n_210, csa_tree_add_117_21_pad_groupi_n_211;
  wire csa_tree_add_117_21_pad_groupi_n_213, csa_tree_add_117_21_pad_groupi_n_214, csa_tree_add_117_21_pad_groupi_n_215, csa_tree_add_117_21_pad_groupi_n_216, csa_tree_add_117_21_pad_groupi_n_217, csa_tree_add_117_21_pad_groupi_n_218, csa_tree_add_117_21_pad_groupi_n_219, csa_tree_add_117_21_pad_groupi_n_220;
  wire csa_tree_add_117_21_pad_groupi_n_221, csa_tree_add_117_21_pad_groupi_n_222, csa_tree_add_117_21_pad_groupi_n_223, csa_tree_add_117_21_pad_groupi_n_224, csa_tree_add_117_21_pad_groupi_n_225, csa_tree_add_117_21_pad_groupi_n_226, csa_tree_add_117_21_pad_groupi_n_227, csa_tree_add_117_21_pad_groupi_n_228;
  wire csa_tree_add_117_21_pad_groupi_n_229, csa_tree_add_117_21_pad_groupi_n_231, csa_tree_add_117_21_pad_groupi_n_232, csa_tree_add_117_21_pad_groupi_n_233, csa_tree_add_117_21_pad_groupi_n_234, csa_tree_add_117_21_pad_groupi_n_235, csa_tree_add_117_21_pad_groupi_n_236, csa_tree_add_117_21_pad_groupi_n_237;
  wire csa_tree_add_117_21_pad_groupi_n_238, csa_tree_add_117_21_pad_groupi_n_239, csa_tree_add_117_21_pad_groupi_n_240, csa_tree_add_117_21_pad_groupi_n_241, csa_tree_add_117_21_pad_groupi_n_243, csa_tree_add_117_21_pad_groupi_n_245, csa_tree_add_117_21_pad_groupi_n_246, csa_tree_add_117_21_pad_groupi_n_247;
  wire csa_tree_add_117_21_pad_groupi_n_248, csa_tree_add_117_21_pad_groupi_n_249, csa_tree_add_117_21_pad_groupi_n_250, csa_tree_add_117_21_pad_groupi_n_254, csa_tree_add_117_21_pad_groupi_n_255, csa_tree_add_117_21_pad_groupi_n_256, csa_tree_add_117_21_pad_groupi_n_257, csa_tree_add_117_21_pad_groupi_n_258;
  wire csa_tree_add_117_21_pad_groupi_n_259, csa_tree_add_117_21_pad_groupi_n_260, csa_tree_add_117_21_pad_groupi_n_261, csa_tree_add_117_21_pad_groupi_n_262, csa_tree_add_117_21_pad_groupi_n_263, csa_tree_add_117_21_pad_groupi_n_264, csa_tree_add_117_21_pad_groupi_n_265, csa_tree_add_117_21_pad_groupi_n_266;
  wire csa_tree_add_117_21_pad_groupi_n_267, csa_tree_add_117_21_pad_groupi_n_268, csa_tree_add_117_21_pad_groupi_n_269, csa_tree_add_117_21_pad_groupi_n_271, csa_tree_add_117_21_pad_groupi_n_272, csa_tree_add_117_21_pad_groupi_n_273, csa_tree_add_117_21_pad_groupi_n_274, csa_tree_add_117_21_pad_groupi_n_275;
  wire csa_tree_add_117_21_pad_groupi_n_276, csa_tree_add_117_21_pad_groupi_n_277, csa_tree_add_117_21_pad_groupi_n_278, csa_tree_add_117_21_pad_groupi_n_279, csa_tree_add_117_21_pad_groupi_n_281, csa_tree_add_117_21_pad_groupi_n_283, csa_tree_add_117_21_pad_groupi_n_284, csa_tree_add_117_21_pad_groupi_n_285;
  wire csa_tree_add_117_21_pad_groupi_n_286, csa_tree_add_117_21_pad_groupi_n_287, csa_tree_add_117_21_pad_groupi_n_288, csa_tree_add_117_21_pad_groupi_n_289, csa_tree_add_117_21_pad_groupi_n_290, csa_tree_add_117_21_pad_groupi_n_291, csa_tree_add_117_21_pad_groupi_n_292, csa_tree_add_117_21_pad_groupi_n_293;
  wire csa_tree_add_117_21_pad_groupi_n_294, csa_tree_add_117_21_pad_groupi_n_295, csa_tree_add_117_21_pad_groupi_n_296, csa_tree_add_117_21_pad_groupi_n_297, csa_tree_add_117_21_pad_groupi_n_298, csa_tree_add_117_21_pad_groupi_n_299, csa_tree_add_117_21_pad_groupi_n_300, csa_tree_add_117_21_pad_groupi_n_301;
  wire csa_tree_add_117_21_pad_groupi_n_302, csa_tree_add_117_21_pad_groupi_n_303, csa_tree_add_117_21_pad_groupi_n_304, csa_tree_add_117_21_pad_groupi_n_305, csa_tree_add_117_21_pad_groupi_n_306, csa_tree_add_117_21_pad_groupi_n_307, csa_tree_add_117_21_pad_groupi_n_308, csa_tree_add_117_21_pad_groupi_n_309;
  wire csa_tree_add_117_21_pad_groupi_n_310, csa_tree_add_117_21_pad_groupi_n_312, csa_tree_add_117_21_pad_groupi_n_313, csa_tree_add_117_21_pad_groupi_n_314, csa_tree_add_117_21_pad_groupi_n_315, csa_tree_add_117_21_pad_groupi_n_316, csa_tree_add_117_21_pad_groupi_n_317, csa_tree_add_117_21_pad_groupi_n_318;
  wire csa_tree_add_117_21_pad_groupi_n_319, csa_tree_add_117_21_pad_groupi_n_320, csa_tree_add_117_21_pad_groupi_n_323, csa_tree_add_117_21_pad_groupi_n_324, csa_tree_add_117_21_pad_groupi_n_325, csa_tree_add_117_21_pad_groupi_n_326, csa_tree_add_117_21_pad_groupi_n_327, csa_tree_add_117_21_pad_groupi_n_328;
  wire csa_tree_add_117_21_pad_groupi_n_329, csa_tree_add_117_21_pad_groupi_n_330, csa_tree_add_117_21_pad_groupi_n_331, csa_tree_add_117_21_pad_groupi_n_332, csa_tree_add_117_21_pad_groupi_n_333, csa_tree_add_117_21_pad_groupi_n_334, csa_tree_add_117_21_pad_groupi_n_335, csa_tree_add_117_21_pad_groupi_n_336;
  wire csa_tree_add_117_21_pad_groupi_n_337, csa_tree_add_117_21_pad_groupi_n_338, csa_tree_add_117_21_pad_groupi_n_339, csa_tree_add_117_21_pad_groupi_n_340, csa_tree_add_117_21_pad_groupi_n_341, csa_tree_add_117_21_pad_groupi_n_342, csa_tree_add_117_21_pad_groupi_n_343, csa_tree_add_117_21_pad_groupi_n_344;
  wire csa_tree_add_117_21_pad_groupi_n_345, csa_tree_add_117_21_pad_groupi_n_346, csa_tree_add_117_21_pad_groupi_n_347, csa_tree_add_117_21_pad_groupi_n_348, csa_tree_add_117_21_pad_groupi_n_349, csa_tree_add_117_21_pad_groupi_n_350, csa_tree_add_117_21_pad_groupi_n_352, csa_tree_add_117_21_pad_groupi_n_353;
  wire csa_tree_add_117_21_pad_groupi_n_354, csa_tree_add_117_21_pad_groupi_n_355, csa_tree_add_117_21_pad_groupi_n_356, csa_tree_add_117_21_pad_groupi_n_357, csa_tree_add_117_21_pad_groupi_n_358, csa_tree_add_117_21_pad_groupi_n_359, csa_tree_add_117_21_pad_groupi_n_360, csa_tree_add_117_21_pad_groupi_n_361;
  wire csa_tree_add_117_21_pad_groupi_n_362, csa_tree_add_117_21_pad_groupi_n_363, csa_tree_add_117_21_pad_groupi_n_364, csa_tree_add_117_21_pad_groupi_n_365, csa_tree_add_117_21_pad_groupi_n_366, csa_tree_add_117_21_pad_groupi_n_367, csa_tree_add_117_21_pad_groupi_n_368, csa_tree_add_117_21_pad_groupi_n_369;
  wire csa_tree_add_117_21_pad_groupi_n_370, csa_tree_add_117_21_pad_groupi_n_371, csa_tree_add_117_21_pad_groupi_n_372, csa_tree_add_117_21_pad_groupi_n_373, csa_tree_add_117_21_pad_groupi_n_374, csa_tree_add_117_21_pad_groupi_n_375, csa_tree_add_117_21_pad_groupi_n_376, csa_tree_add_117_21_pad_groupi_n_377;
  wire csa_tree_add_117_21_pad_groupi_n_378, csa_tree_add_117_21_pad_groupi_n_379, csa_tree_add_117_21_pad_groupi_n_380, csa_tree_add_117_21_pad_groupi_n_381, csa_tree_add_117_21_pad_groupi_n_382, csa_tree_add_117_21_pad_groupi_n_383, csa_tree_add_117_21_pad_groupi_n_384, csa_tree_add_117_21_pad_groupi_n_385;
  wire csa_tree_add_117_21_pad_groupi_n_386, csa_tree_add_117_21_pad_groupi_n_387, csa_tree_add_117_21_pad_groupi_n_388, csa_tree_add_117_21_pad_groupi_n_389, csa_tree_add_117_21_pad_groupi_n_390, csa_tree_add_117_21_pad_groupi_n_391, csa_tree_add_117_21_pad_groupi_n_392, csa_tree_add_117_21_pad_groupi_n_394;
  wire csa_tree_add_117_21_pad_groupi_n_395, csa_tree_add_117_21_pad_groupi_n_396, csa_tree_add_117_21_pad_groupi_n_397, csa_tree_add_117_21_pad_groupi_n_398, csa_tree_add_117_21_pad_groupi_n_399, csa_tree_add_117_21_pad_groupi_n_400, csa_tree_add_117_21_pad_groupi_n_401, csa_tree_add_117_21_pad_groupi_n_402;
  wire csa_tree_add_117_21_pad_groupi_n_403, csa_tree_add_117_21_pad_groupi_n_404, csa_tree_add_117_21_pad_groupi_n_405, csa_tree_add_117_21_pad_groupi_n_406, csa_tree_add_117_21_pad_groupi_n_407, csa_tree_add_117_21_pad_groupi_n_408, csa_tree_add_117_21_pad_groupi_n_409, csa_tree_add_117_21_pad_groupi_n_410;
  wire csa_tree_add_117_21_pad_groupi_n_411, csa_tree_add_117_21_pad_groupi_n_412, csa_tree_add_117_21_pad_groupi_n_413, csa_tree_add_117_21_pad_groupi_n_414, csa_tree_add_117_21_pad_groupi_n_415, csa_tree_add_117_21_pad_groupi_n_416, csa_tree_add_117_21_pad_groupi_n_417, csa_tree_add_117_21_pad_groupi_n_418;
  wire csa_tree_add_117_21_pad_groupi_n_419, csa_tree_add_117_21_pad_groupi_n_420, csa_tree_add_117_21_pad_groupi_n_421, csa_tree_add_117_21_pad_groupi_n_422, csa_tree_add_117_21_pad_groupi_n_423, csa_tree_add_117_21_pad_groupi_n_424, csa_tree_add_117_21_pad_groupi_n_425, csa_tree_add_117_21_pad_groupi_n_426;
  wire csa_tree_add_117_21_pad_groupi_n_427, csa_tree_add_117_21_pad_groupi_n_428, csa_tree_add_117_21_pad_groupi_n_429, csa_tree_add_117_21_pad_groupi_n_430, csa_tree_add_117_21_pad_groupi_n_431, csa_tree_add_117_21_pad_groupi_n_432, csa_tree_add_117_21_pad_groupi_n_433, csa_tree_add_117_21_pad_groupi_n_434;
  wire csa_tree_add_117_21_pad_groupi_n_435, csa_tree_add_117_21_pad_groupi_n_436, csa_tree_add_117_21_pad_groupi_n_437, csa_tree_add_117_21_pad_groupi_n_438, csa_tree_add_117_21_pad_groupi_n_439, csa_tree_add_117_21_pad_groupi_n_440, csa_tree_add_117_21_pad_groupi_n_441, csa_tree_add_117_21_pad_groupi_n_442;
  wire csa_tree_add_117_21_pad_groupi_n_443, csa_tree_add_117_21_pad_groupi_n_444, csa_tree_add_117_21_pad_groupi_n_445, csa_tree_add_117_21_pad_groupi_n_446, csa_tree_add_117_21_pad_groupi_n_447, csa_tree_add_117_21_pad_groupi_n_448, csa_tree_add_117_21_pad_groupi_n_449, csa_tree_add_117_21_pad_groupi_n_450;
  wire csa_tree_add_117_21_pad_groupi_n_451, csa_tree_add_117_21_pad_groupi_n_452, csa_tree_add_117_21_pad_groupi_n_456, csa_tree_add_117_21_pad_groupi_n_467, csa_tree_add_117_21_pad_groupi_n_468, csa_tree_add_117_21_pad_groupi_n_469, csa_tree_add_117_21_pad_groupi_n_470, csa_tree_add_117_21_pad_groupi_n_471;
  wire csa_tree_add_117_21_pad_groupi_n_472, csa_tree_add_117_21_pad_groupi_n_473, csa_tree_add_117_21_pad_groupi_n_474, csa_tree_add_117_21_pad_groupi_n_476, csa_tree_add_117_21_pad_groupi_n_477, csa_tree_add_117_21_pad_groupi_n_478, csa_tree_add_117_21_pad_groupi_n_479, csa_tree_add_117_21_pad_groupi_n_480;
  wire csa_tree_add_117_21_pad_groupi_n_481, csa_tree_add_117_21_pad_groupi_n_482, csa_tree_add_117_21_pad_groupi_n_483, csa_tree_add_117_21_pad_groupi_n_484, csa_tree_add_117_21_pad_groupi_n_485, csa_tree_add_117_21_pad_groupi_n_486, csa_tree_add_117_21_pad_groupi_n_487, csa_tree_add_117_21_pad_groupi_n_488;
  wire csa_tree_add_117_21_pad_groupi_n_489, csa_tree_add_117_21_pad_groupi_n_490, csa_tree_add_117_21_pad_groupi_n_491, csa_tree_add_117_21_pad_groupi_n_492, csa_tree_add_117_21_pad_groupi_n_493, csa_tree_add_117_21_pad_groupi_n_494, csa_tree_add_117_21_pad_groupi_n_495, csa_tree_add_117_21_pad_groupi_n_496;
  wire csa_tree_add_117_21_pad_groupi_n_497, csa_tree_add_117_21_pad_groupi_n_498, csa_tree_add_117_21_pad_groupi_n_499, csa_tree_add_117_21_pad_groupi_n_500, csa_tree_add_117_21_pad_groupi_n_501, csa_tree_add_117_21_pad_groupi_n_502, csa_tree_add_117_21_pad_groupi_n_503, csa_tree_add_117_21_pad_groupi_n_504;
  wire csa_tree_add_117_21_pad_groupi_n_505, csa_tree_add_117_21_pad_groupi_n_506, csa_tree_add_117_21_pad_groupi_n_507, csa_tree_add_117_21_pad_groupi_n_508, csa_tree_add_117_21_pad_groupi_n_509, csa_tree_add_117_21_pad_groupi_n_510, csa_tree_add_117_21_pad_groupi_n_511, csa_tree_add_117_21_pad_groupi_n_512;
  wire csa_tree_add_117_21_pad_groupi_n_513, csa_tree_add_117_21_pad_groupi_n_514, csa_tree_add_117_21_pad_groupi_n_515, csa_tree_add_117_21_pad_groupi_n_516, csa_tree_add_117_21_pad_groupi_n_517, csa_tree_add_117_21_pad_groupi_n_518, csa_tree_add_117_21_pad_groupi_n_519, csa_tree_add_117_21_pad_groupi_n_520;
  wire csa_tree_add_117_21_pad_groupi_n_521, csa_tree_add_117_21_pad_groupi_n_522, csa_tree_add_117_21_pad_groupi_n_523, csa_tree_add_117_21_pad_groupi_n_524, csa_tree_add_117_21_pad_groupi_n_525, csa_tree_add_117_21_pad_groupi_n_526, csa_tree_add_117_21_pad_groupi_n_527, csa_tree_add_117_21_pad_groupi_n_528;
  wire csa_tree_add_117_21_pad_groupi_n_529, csa_tree_add_117_21_pad_groupi_n_530, csa_tree_add_117_21_pad_groupi_n_531, csa_tree_add_117_21_pad_groupi_n_532, csa_tree_add_117_21_pad_groupi_n_533, csa_tree_add_117_21_pad_groupi_n_534, csa_tree_add_117_21_pad_groupi_n_535, csa_tree_add_117_21_pad_groupi_n_536;
  wire csa_tree_add_117_21_pad_groupi_n_537, csa_tree_add_117_21_pad_groupi_n_538, csa_tree_add_117_21_pad_groupi_n_539, csa_tree_add_117_21_pad_groupi_n_540, csa_tree_add_117_21_pad_groupi_n_541, csa_tree_add_117_21_pad_groupi_n_542, csa_tree_add_117_21_pad_groupi_n_543, csa_tree_add_117_21_pad_groupi_n_544;
  wire csa_tree_add_117_21_pad_groupi_n_545, csa_tree_add_117_21_pad_groupi_n_546, csa_tree_add_117_21_pad_groupi_n_547, csa_tree_add_117_21_pad_groupi_n_548, csa_tree_add_117_21_pad_groupi_n_549, csa_tree_add_117_21_pad_groupi_n_550, csa_tree_add_117_21_pad_groupi_n_551, csa_tree_add_117_21_pad_groupi_n_552;
  wire csa_tree_add_117_21_pad_groupi_n_553, csa_tree_add_117_21_pad_groupi_n_554, csa_tree_add_117_21_pad_groupi_n_555, csa_tree_add_117_21_pad_groupi_n_556, csa_tree_add_117_21_pad_groupi_n_557, csa_tree_add_117_21_pad_groupi_n_558, csa_tree_add_117_21_pad_groupi_n_559, csa_tree_add_117_21_pad_groupi_n_560;
  wire csa_tree_add_117_21_pad_groupi_n_561, csa_tree_add_117_21_pad_groupi_n_562, csa_tree_add_117_21_pad_groupi_n_563, csa_tree_add_117_21_pad_groupi_n_564, csa_tree_add_117_21_pad_groupi_n_565, csa_tree_add_117_21_pad_groupi_n_566, csa_tree_add_117_21_pad_groupi_n_567, csa_tree_add_117_21_pad_groupi_n_568;
  wire csa_tree_add_117_21_pad_groupi_n_569, csa_tree_add_117_21_pad_groupi_n_570, csa_tree_add_117_21_pad_groupi_n_571, csa_tree_add_117_21_pad_groupi_n_572, csa_tree_add_117_21_pad_groupi_n_573, csa_tree_add_117_21_pad_groupi_n_574, csa_tree_add_117_21_pad_groupi_n_575, csa_tree_add_117_21_pad_groupi_n_576;
  wire csa_tree_add_117_21_pad_groupi_n_577, csa_tree_add_117_21_pad_groupi_n_578, csa_tree_add_117_21_pad_groupi_n_579, csa_tree_add_117_21_pad_groupi_n_580, csa_tree_add_117_21_pad_groupi_n_581, csa_tree_add_117_21_pad_groupi_n_582, csa_tree_add_117_21_pad_groupi_n_583, csa_tree_add_117_21_pad_groupi_n_584;
  wire csa_tree_add_117_21_pad_groupi_n_585, csa_tree_add_117_21_pad_groupi_n_586, csa_tree_add_117_21_pad_groupi_n_587, csa_tree_add_117_21_pad_groupi_n_588, csa_tree_add_117_21_pad_groupi_n_589, csa_tree_add_117_21_pad_groupi_n_590, csa_tree_add_117_21_pad_groupi_n_591, csa_tree_add_117_21_pad_groupi_n_592;
  wire csa_tree_add_117_21_pad_groupi_n_593, csa_tree_add_117_21_pad_groupi_n_594, csa_tree_add_117_21_pad_groupi_n_595, csa_tree_add_117_21_pad_groupi_n_596, csa_tree_add_117_21_pad_groupi_n_597, csa_tree_add_117_21_pad_groupi_n_598, csa_tree_add_117_21_pad_groupi_n_599, csa_tree_add_117_21_pad_groupi_n_600;
  wire csa_tree_add_117_21_pad_groupi_n_601, csa_tree_add_117_21_pad_groupi_n_602, csa_tree_add_117_21_pad_groupi_n_603, csa_tree_add_117_21_pad_groupi_n_604, csa_tree_add_117_21_pad_groupi_n_605, csa_tree_add_117_21_pad_groupi_n_606, csa_tree_add_117_21_pad_groupi_n_607, csa_tree_add_117_21_pad_groupi_n_608;
  wire csa_tree_add_117_21_pad_groupi_n_609, csa_tree_add_117_21_pad_groupi_n_610, csa_tree_add_117_21_pad_groupi_n_611, csa_tree_add_117_21_pad_groupi_n_612, csa_tree_add_117_21_pad_groupi_n_613, csa_tree_add_117_21_pad_groupi_n_614, csa_tree_add_117_21_pad_groupi_n_615, csa_tree_add_117_21_pad_groupi_n_616;
  wire csa_tree_add_117_21_pad_groupi_n_617, csa_tree_add_117_21_pad_groupi_n_618, csa_tree_add_117_21_pad_groupi_n_619, csa_tree_add_117_21_pad_groupi_n_620, csa_tree_add_117_21_pad_groupi_n_621, csa_tree_add_117_21_pad_groupi_n_622, csa_tree_add_117_21_pad_groupi_n_623, csa_tree_add_117_21_pad_groupi_n_624;
  wire csa_tree_add_117_21_pad_groupi_n_625, csa_tree_add_117_21_pad_groupi_n_626, csa_tree_add_117_21_pad_groupi_n_627, csa_tree_add_117_21_pad_groupi_n_628, csa_tree_add_117_21_pad_groupi_n_629, csa_tree_add_117_21_pad_groupi_n_630, csa_tree_add_117_21_pad_groupi_n_631, csa_tree_add_117_21_pad_groupi_n_632;
  wire csa_tree_add_117_21_pad_groupi_n_633, csa_tree_add_117_21_pad_groupi_n_634, csa_tree_add_117_21_pad_groupi_n_635, csa_tree_add_117_21_pad_groupi_n_636, csa_tree_add_117_21_pad_groupi_n_637, csa_tree_add_117_21_pad_groupi_n_638, csa_tree_add_117_21_pad_groupi_n_639, csa_tree_add_117_21_pad_groupi_n_640;
  wire csa_tree_add_117_21_pad_groupi_n_641, csa_tree_add_117_21_pad_groupi_n_642, csa_tree_add_117_21_pad_groupi_n_643, csa_tree_add_117_21_pad_groupi_n_644, csa_tree_add_117_21_pad_groupi_n_645, csa_tree_add_117_21_pad_groupi_n_646, csa_tree_add_117_21_pad_groupi_n_647, csa_tree_add_117_21_pad_groupi_n_648;
  wire csa_tree_add_117_21_pad_groupi_n_649, csa_tree_add_117_21_pad_groupi_n_650, csa_tree_add_117_21_pad_groupi_n_651, csa_tree_add_117_21_pad_groupi_n_652, csa_tree_add_117_21_pad_groupi_n_653, csa_tree_add_117_21_pad_groupi_n_654, csa_tree_add_117_21_pad_groupi_n_655, csa_tree_add_117_21_pad_groupi_n_656;
  wire csa_tree_add_117_21_pad_groupi_n_657, csa_tree_add_117_21_pad_groupi_n_658, csa_tree_add_117_21_pad_groupi_n_659, csa_tree_add_117_21_pad_groupi_n_660, csa_tree_add_117_21_pad_groupi_n_661, csa_tree_add_117_21_pad_groupi_n_662, csa_tree_add_117_21_pad_groupi_n_663, csa_tree_add_117_21_pad_groupi_n_664;
  wire csa_tree_add_117_21_pad_groupi_n_665, csa_tree_add_117_21_pad_groupi_n_666, csa_tree_add_117_21_pad_groupi_n_667, csa_tree_add_117_21_pad_groupi_n_668, csa_tree_add_117_21_pad_groupi_n_669, csa_tree_add_117_21_pad_groupi_n_670, csa_tree_add_117_21_pad_groupi_n_671, csa_tree_add_117_21_pad_groupi_n_672;
  wire csa_tree_add_117_21_pad_groupi_n_673, csa_tree_add_117_21_pad_groupi_n_674, csa_tree_add_117_21_pad_groupi_n_675, csa_tree_add_117_21_pad_groupi_n_676, csa_tree_add_117_21_pad_groupi_n_677, csa_tree_add_117_21_pad_groupi_n_678, csa_tree_add_117_21_pad_groupi_n_679, csa_tree_add_117_21_pad_groupi_n_680;
  wire csa_tree_add_117_21_pad_groupi_n_681, csa_tree_add_117_21_pad_groupi_n_682, csa_tree_add_117_21_pad_groupi_n_683, csa_tree_add_117_21_pad_groupi_n_684, csa_tree_add_117_21_pad_groupi_n_685, csa_tree_add_117_21_pad_groupi_n_686, csa_tree_add_117_21_pad_groupi_n_687, csa_tree_add_117_21_pad_groupi_n_688;
  wire csa_tree_add_117_21_pad_groupi_n_689, csa_tree_add_117_21_pad_groupi_n_690, csa_tree_add_117_21_pad_groupi_n_691, csa_tree_add_117_21_pad_groupi_n_692, csa_tree_add_117_21_pad_groupi_n_693, csa_tree_add_117_21_pad_groupi_n_694, csa_tree_add_117_21_pad_groupi_n_695, csa_tree_add_117_21_pad_groupi_n_696;
  wire csa_tree_add_117_21_pad_groupi_n_697, csa_tree_add_117_21_pad_groupi_n_698, csa_tree_add_117_21_pad_groupi_n_699, csa_tree_add_117_21_pad_groupi_n_700, csa_tree_add_117_21_pad_groupi_n_701, csa_tree_add_117_21_pad_groupi_n_702, csa_tree_add_117_21_pad_groupi_n_703, csa_tree_add_117_21_pad_groupi_n_704;
  wire csa_tree_add_117_21_pad_groupi_n_705, csa_tree_add_117_21_pad_groupi_n_706, csa_tree_add_117_21_pad_groupi_n_707, csa_tree_add_117_21_pad_groupi_n_708, csa_tree_add_117_21_pad_groupi_n_709, csa_tree_add_117_21_pad_groupi_n_710, csa_tree_add_117_21_pad_groupi_n_711, csa_tree_add_117_21_pad_groupi_n_712;
  wire csa_tree_add_117_21_pad_groupi_n_713, csa_tree_add_117_21_pad_groupi_n_714, csa_tree_add_117_21_pad_groupi_n_715, csa_tree_add_117_21_pad_groupi_n_716, csa_tree_add_117_21_pad_groupi_n_717, csa_tree_add_117_21_pad_groupi_n_718, csa_tree_add_117_21_pad_groupi_n_719, csa_tree_add_117_21_pad_groupi_n_720;
  wire csa_tree_add_117_21_pad_groupi_n_721, csa_tree_add_117_21_pad_groupi_n_722, csa_tree_add_117_21_pad_groupi_n_723, csa_tree_add_117_21_pad_groupi_n_724, csa_tree_add_117_21_pad_groupi_n_725, csa_tree_add_117_21_pad_groupi_n_726, csa_tree_add_117_21_pad_groupi_n_727, csa_tree_add_117_21_pad_groupi_n_728;
  wire csa_tree_add_117_21_pad_groupi_n_729, csa_tree_add_117_21_pad_groupi_n_730, csa_tree_add_117_21_pad_groupi_n_731, csa_tree_add_117_21_pad_groupi_n_732, csa_tree_add_117_21_pad_groupi_n_733, csa_tree_add_117_21_pad_groupi_n_734, csa_tree_add_117_21_pad_groupi_n_735, csa_tree_add_117_21_pad_groupi_n_736;
  wire csa_tree_add_117_21_pad_groupi_n_737, csa_tree_add_117_21_pad_groupi_n_738, csa_tree_add_117_21_pad_groupi_n_739, csa_tree_add_117_21_pad_groupi_n_740, csa_tree_add_117_21_pad_groupi_n_741, csa_tree_add_117_21_pad_groupi_n_742, csa_tree_add_117_21_pad_groupi_n_743, csa_tree_add_117_21_pad_groupi_n_744;
  wire csa_tree_add_117_21_pad_groupi_n_745, csa_tree_add_117_21_pad_groupi_n_746, csa_tree_add_117_21_pad_groupi_n_747, csa_tree_add_117_21_pad_groupi_n_748, csa_tree_add_117_21_pad_groupi_n_749, csa_tree_add_117_21_pad_groupi_n_750, csa_tree_add_117_21_pad_groupi_n_751, csa_tree_add_117_21_pad_groupi_n_752;
  wire csa_tree_add_117_21_pad_groupi_n_753, csa_tree_add_117_21_pad_groupi_n_754, csa_tree_add_117_21_pad_groupi_n_755, csa_tree_add_117_21_pad_groupi_n_756, csa_tree_add_117_21_pad_groupi_n_757, csa_tree_add_117_21_pad_groupi_n_758, csa_tree_add_117_21_pad_groupi_n_759, csa_tree_add_117_21_pad_groupi_n_760;
  wire csa_tree_add_117_21_pad_groupi_n_761, csa_tree_add_117_21_pad_groupi_n_762, csa_tree_add_117_21_pad_groupi_n_763, csa_tree_add_117_21_pad_groupi_n_764, csa_tree_add_117_21_pad_groupi_n_765, csa_tree_add_117_21_pad_groupi_n_766, csa_tree_add_117_21_pad_groupi_n_767, csa_tree_add_117_21_pad_groupi_n_768;
  wire csa_tree_add_117_21_pad_groupi_n_769, csa_tree_add_117_21_pad_groupi_n_770, csa_tree_add_117_21_pad_groupi_n_771, csa_tree_add_117_21_pad_groupi_n_772, csa_tree_add_117_21_pad_groupi_n_773, csa_tree_add_117_21_pad_groupi_n_774, csa_tree_add_117_21_pad_groupi_n_775, csa_tree_add_117_21_pad_groupi_n_776;
  wire csa_tree_add_117_21_pad_groupi_n_777, csa_tree_add_117_21_pad_groupi_n_778, csa_tree_add_117_21_pad_groupi_n_779, csa_tree_add_117_21_pad_groupi_n_780, csa_tree_add_117_21_pad_groupi_n_781, csa_tree_add_117_21_pad_groupi_n_782, csa_tree_add_117_21_pad_groupi_n_783, csa_tree_add_117_21_pad_groupi_n_784;
  wire csa_tree_add_117_21_pad_groupi_n_785, csa_tree_add_117_21_pad_groupi_n_786, csa_tree_add_117_21_pad_groupi_n_787, csa_tree_add_117_21_pad_groupi_n_788, csa_tree_add_117_21_pad_groupi_n_789, csa_tree_add_117_21_pad_groupi_n_790, csa_tree_add_117_21_pad_groupi_n_791, csa_tree_add_117_21_pad_groupi_n_792;
  wire csa_tree_add_117_21_pad_groupi_n_793, csa_tree_add_117_21_pad_groupi_n_794, csa_tree_add_117_21_pad_groupi_n_795, csa_tree_add_117_21_pad_groupi_n_796, csa_tree_add_117_21_pad_groupi_n_797, csa_tree_add_117_21_pad_groupi_n_798, csa_tree_add_117_21_pad_groupi_n_799, csa_tree_add_117_21_pad_groupi_n_800;
  wire csa_tree_add_117_21_pad_groupi_n_801, csa_tree_add_117_21_pad_groupi_n_802, csa_tree_add_117_21_pad_groupi_n_803, csa_tree_add_117_21_pad_groupi_n_804, csa_tree_add_117_21_pad_groupi_n_805, csa_tree_add_117_21_pad_groupi_n_806, csa_tree_add_117_21_pad_groupi_n_807, csa_tree_add_117_21_pad_groupi_n_808;
  wire csa_tree_add_117_21_pad_groupi_n_809, csa_tree_add_117_21_pad_groupi_n_810, csa_tree_add_117_21_pad_groupi_n_811, csa_tree_add_117_21_pad_groupi_n_812, csa_tree_add_117_21_pad_groupi_n_813, csa_tree_add_117_21_pad_groupi_n_814, csa_tree_add_117_21_pad_groupi_n_815, csa_tree_add_117_21_pad_groupi_n_816;
  wire csa_tree_add_117_21_pad_groupi_n_817, csa_tree_add_117_21_pad_groupi_n_818, csa_tree_add_117_21_pad_groupi_n_819, csa_tree_add_117_21_pad_groupi_n_820, csa_tree_add_117_21_pad_groupi_n_821, csa_tree_add_117_21_pad_groupi_n_822, csa_tree_add_117_21_pad_groupi_n_823, csa_tree_add_117_21_pad_groupi_n_824;
  wire csa_tree_add_117_21_pad_groupi_n_825, csa_tree_add_117_21_pad_groupi_n_826, csa_tree_add_117_21_pad_groupi_n_827, csa_tree_add_117_21_pad_groupi_n_828, csa_tree_add_117_21_pad_groupi_n_829, csa_tree_add_117_21_pad_groupi_n_830, csa_tree_add_117_21_pad_groupi_n_831, csa_tree_add_117_21_pad_groupi_n_832;
  wire csa_tree_add_117_21_pad_groupi_n_833, csa_tree_add_117_21_pad_groupi_n_834, csa_tree_add_117_21_pad_groupi_n_835, csa_tree_add_117_21_pad_groupi_n_836, csa_tree_add_117_21_pad_groupi_n_837, csa_tree_add_117_21_pad_groupi_n_838, csa_tree_add_117_21_pad_groupi_n_839, csa_tree_add_117_21_pad_groupi_n_840;
  wire csa_tree_add_117_21_pad_groupi_n_841, csa_tree_add_117_21_pad_groupi_n_842, csa_tree_add_117_21_pad_groupi_n_843, csa_tree_add_117_21_pad_groupi_n_844, csa_tree_add_117_21_pad_groupi_n_845, csa_tree_add_117_21_pad_groupi_n_846, csa_tree_add_117_21_pad_groupi_n_847, csa_tree_add_117_21_pad_groupi_n_848;
  wire csa_tree_add_117_21_pad_groupi_n_849, csa_tree_add_117_21_pad_groupi_n_850, csa_tree_add_117_21_pad_groupi_n_851, csa_tree_add_117_21_pad_groupi_n_852, csa_tree_add_117_21_pad_groupi_n_853, csa_tree_add_117_21_pad_groupi_n_854, csa_tree_add_117_21_pad_groupi_n_855, csa_tree_add_117_21_pad_groupi_n_856;
  wire csa_tree_add_117_21_pad_groupi_n_857, csa_tree_add_117_21_pad_groupi_n_858, csa_tree_add_117_21_pad_groupi_n_859, csa_tree_add_117_21_pad_groupi_n_860, csa_tree_add_117_21_pad_groupi_n_861, csa_tree_add_117_21_pad_groupi_n_862, csa_tree_add_117_21_pad_groupi_n_863, csa_tree_add_117_21_pad_groupi_n_864;
  wire csa_tree_add_117_21_pad_groupi_n_865, csa_tree_add_117_21_pad_groupi_n_866, csa_tree_add_117_21_pad_groupi_n_867, csa_tree_add_117_21_pad_groupi_n_868, csa_tree_add_117_21_pad_groupi_n_869, csa_tree_add_117_21_pad_groupi_n_870, csa_tree_add_117_21_pad_groupi_n_871, csa_tree_add_117_21_pad_groupi_n_872;
  wire csa_tree_add_117_21_pad_groupi_n_873, csa_tree_add_117_21_pad_groupi_n_874, csa_tree_add_117_21_pad_groupi_n_875, csa_tree_add_117_21_pad_groupi_n_876, csa_tree_add_117_21_pad_groupi_n_877, csa_tree_add_117_21_pad_groupi_n_878, csa_tree_add_117_21_pad_groupi_n_879, csa_tree_add_117_21_pad_groupi_n_880;
  wire csa_tree_add_117_21_pad_groupi_n_881, csa_tree_add_117_21_pad_groupi_n_882, csa_tree_add_117_21_pad_groupi_n_883, csa_tree_add_117_21_pad_groupi_n_884, csa_tree_add_117_21_pad_groupi_n_885, csa_tree_add_117_21_pad_groupi_n_886, csa_tree_add_117_21_pad_groupi_n_887, csa_tree_add_117_21_pad_groupi_n_888;
  wire csa_tree_add_117_21_pad_groupi_n_889, csa_tree_add_117_21_pad_groupi_n_890, csa_tree_add_117_21_pad_groupi_n_891, csa_tree_add_117_21_pad_groupi_n_892, csa_tree_add_117_21_pad_groupi_n_893, csa_tree_add_117_21_pad_groupi_n_894, csa_tree_add_117_21_pad_groupi_n_895, csa_tree_add_117_21_pad_groupi_n_896;
  wire csa_tree_add_117_21_pad_groupi_n_897, csa_tree_add_117_21_pad_groupi_n_898, csa_tree_add_117_21_pad_groupi_n_899, csa_tree_add_117_21_pad_groupi_n_900, csa_tree_add_117_21_pad_groupi_n_901, csa_tree_add_117_21_pad_groupi_n_902, csa_tree_add_117_21_pad_groupi_n_903, csa_tree_add_117_21_pad_groupi_n_904;
  wire csa_tree_add_117_21_pad_groupi_n_905, csa_tree_add_117_21_pad_groupi_n_906, csa_tree_add_117_21_pad_groupi_n_907, csa_tree_add_117_21_pad_groupi_n_908, csa_tree_add_117_21_pad_groupi_n_909, csa_tree_add_117_21_pad_groupi_n_910, csa_tree_add_117_21_pad_groupi_n_911, csa_tree_add_117_21_pad_groupi_n_912;
  wire csa_tree_add_117_21_pad_groupi_n_913, csa_tree_add_117_21_pad_groupi_n_914, csa_tree_add_117_21_pad_groupi_n_915, csa_tree_add_117_21_pad_groupi_n_916, csa_tree_add_117_21_pad_groupi_n_917, csa_tree_add_117_21_pad_groupi_n_918, csa_tree_add_117_21_pad_groupi_n_919, csa_tree_add_117_21_pad_groupi_n_920;
  wire csa_tree_add_117_21_pad_groupi_n_921, csa_tree_add_117_21_pad_groupi_n_922, csa_tree_add_117_21_pad_groupi_n_923, csa_tree_add_117_21_pad_groupi_n_924, csa_tree_add_117_21_pad_groupi_n_925, csa_tree_add_117_21_pad_groupi_n_926, csa_tree_add_117_21_pad_groupi_n_927, csa_tree_add_117_21_pad_groupi_n_928;
  wire csa_tree_add_117_21_pad_groupi_n_929, csa_tree_add_117_21_pad_groupi_n_930, csa_tree_add_117_21_pad_groupi_n_931, csa_tree_add_117_21_pad_groupi_n_932, csa_tree_add_117_21_pad_groupi_n_933, csa_tree_add_117_21_pad_groupi_n_934, csa_tree_add_117_21_pad_groupi_n_935, csa_tree_add_117_21_pad_groupi_n_936;
  wire csa_tree_add_117_21_pad_groupi_n_937, csa_tree_add_117_21_pad_groupi_n_938, csa_tree_add_117_21_pad_groupi_n_939, csa_tree_add_117_21_pad_groupi_n_940, csa_tree_add_117_21_pad_groupi_n_941, csa_tree_add_117_21_pad_groupi_n_942, csa_tree_add_117_21_pad_groupi_n_943, csa_tree_add_117_21_pad_groupi_n_944;
  wire csa_tree_add_117_21_pad_groupi_n_945, csa_tree_add_117_21_pad_groupi_n_946, csa_tree_add_117_21_pad_groupi_n_947, csa_tree_add_117_21_pad_groupi_n_948, csa_tree_add_117_21_pad_groupi_n_949, csa_tree_add_117_21_pad_groupi_n_950, csa_tree_add_117_21_pad_groupi_n_951, csa_tree_add_117_21_pad_groupi_n_952;
  wire csa_tree_add_117_21_pad_groupi_n_953, csa_tree_add_117_21_pad_groupi_n_954, csa_tree_add_117_21_pad_groupi_n_955, csa_tree_add_117_21_pad_groupi_n_956, csa_tree_add_117_21_pad_groupi_n_957, csa_tree_add_117_21_pad_groupi_n_958, csa_tree_add_117_21_pad_groupi_n_959, csa_tree_add_117_21_pad_groupi_n_960;
  wire csa_tree_add_117_21_pad_groupi_n_961, csa_tree_add_117_21_pad_groupi_n_962, csa_tree_add_117_21_pad_groupi_n_963, csa_tree_add_117_21_pad_groupi_n_964, csa_tree_add_117_21_pad_groupi_n_965, csa_tree_add_117_21_pad_groupi_n_966, csa_tree_add_117_21_pad_groupi_n_967, csa_tree_add_117_21_pad_groupi_n_968;
  wire csa_tree_add_117_21_pad_groupi_n_969, csa_tree_add_117_21_pad_groupi_n_970, csa_tree_add_117_21_pad_groupi_n_971, csa_tree_add_117_21_pad_groupi_n_972, csa_tree_add_117_21_pad_groupi_n_973, csa_tree_add_117_21_pad_groupi_n_974, csa_tree_add_117_21_pad_groupi_n_975, csa_tree_add_117_21_pad_groupi_n_976;
  wire csa_tree_add_117_21_pad_groupi_n_977, csa_tree_add_117_21_pad_groupi_n_978, csa_tree_add_117_21_pad_groupi_n_979, csa_tree_add_117_21_pad_groupi_n_980, csa_tree_add_117_21_pad_groupi_n_981, csa_tree_add_117_21_pad_groupi_n_982, csa_tree_add_117_21_pad_groupi_n_983, csa_tree_add_117_21_pad_groupi_n_984;
  wire csa_tree_add_117_21_pad_groupi_n_985, csa_tree_add_117_21_pad_groupi_n_986, csa_tree_add_117_21_pad_groupi_n_987, csa_tree_add_117_21_pad_groupi_n_988, csa_tree_add_117_21_pad_groupi_n_989, csa_tree_add_117_21_pad_groupi_n_990, csa_tree_add_117_21_pad_groupi_n_991, csa_tree_add_117_21_pad_groupi_n_992;
  wire csa_tree_add_117_21_pad_groupi_n_993, csa_tree_add_117_21_pad_groupi_n_994, csa_tree_add_117_21_pad_groupi_n_995, csa_tree_add_117_21_pad_groupi_n_996, csa_tree_add_117_21_pad_groupi_n_997, csa_tree_add_117_21_pad_groupi_n_998, csa_tree_add_117_21_pad_groupi_n_999, csa_tree_add_117_21_pad_groupi_n_1000;
  wire csa_tree_add_117_21_pad_groupi_n_1001, csa_tree_add_117_21_pad_groupi_n_1002, csa_tree_add_117_21_pad_groupi_n_1003, csa_tree_add_117_21_pad_groupi_n_1004, csa_tree_add_117_21_pad_groupi_n_1005, csa_tree_add_117_21_pad_groupi_n_1006, csa_tree_add_117_21_pad_groupi_n_1007, csa_tree_add_117_21_pad_groupi_n_1008;
  wire csa_tree_add_117_21_pad_groupi_n_1009, csa_tree_add_117_21_pad_groupi_n_1010, csa_tree_add_117_21_pad_groupi_n_1011, csa_tree_add_117_21_pad_groupi_n_1012, csa_tree_add_117_21_pad_groupi_n_1013, csa_tree_add_117_21_pad_groupi_n_1014, csa_tree_add_117_21_pad_groupi_n_1015, csa_tree_add_117_21_pad_groupi_n_1016;
  wire csa_tree_add_117_21_pad_groupi_n_1017, csa_tree_add_117_21_pad_groupi_n_1018, csa_tree_add_117_21_pad_groupi_n_1019, csa_tree_add_117_21_pad_groupi_n_1020, csa_tree_add_117_21_pad_groupi_n_1021, csa_tree_add_117_21_pad_groupi_n_1022, csa_tree_add_117_21_pad_groupi_n_1023, csa_tree_add_117_21_pad_groupi_n_1024;
  wire csa_tree_add_117_21_pad_groupi_n_1025, csa_tree_add_117_21_pad_groupi_n_1026, csa_tree_add_117_21_pad_groupi_n_1027, csa_tree_add_117_21_pad_groupi_n_1028, csa_tree_add_117_21_pad_groupi_n_1029, csa_tree_add_117_21_pad_groupi_n_1030, csa_tree_add_117_21_pad_groupi_n_1031, csa_tree_add_117_21_pad_groupi_n_1032;
  wire csa_tree_add_117_21_pad_groupi_n_1033, csa_tree_add_117_21_pad_groupi_n_1034, csa_tree_add_117_21_pad_groupi_n_1035, csa_tree_add_117_21_pad_groupi_n_1036, csa_tree_add_117_21_pad_groupi_n_1037, csa_tree_add_117_21_pad_groupi_n_1038, csa_tree_add_117_21_pad_groupi_n_1039, csa_tree_add_117_21_pad_groupi_n_1040;
  wire csa_tree_add_117_21_pad_groupi_n_1041, csa_tree_add_117_21_pad_groupi_n_1042, csa_tree_add_117_21_pad_groupi_n_1043, csa_tree_add_117_21_pad_groupi_n_1044, csa_tree_add_117_21_pad_groupi_n_1045, csa_tree_add_117_21_pad_groupi_n_1046, csa_tree_add_117_21_pad_groupi_n_1047, csa_tree_add_117_21_pad_groupi_n_1048;
  wire csa_tree_add_117_21_pad_groupi_n_1049, csa_tree_add_117_21_pad_groupi_n_1050, csa_tree_add_117_21_pad_groupi_n_1051, csa_tree_add_117_21_pad_groupi_n_1052, csa_tree_add_117_21_pad_groupi_n_1053, csa_tree_add_117_21_pad_groupi_n_1054, csa_tree_add_117_21_pad_groupi_n_1055, csa_tree_add_117_21_pad_groupi_n_1056;
  wire csa_tree_add_117_21_pad_groupi_n_1057, csa_tree_add_117_21_pad_groupi_n_1058, csa_tree_add_117_21_pad_groupi_n_1059, csa_tree_add_117_21_pad_groupi_n_1060, csa_tree_add_117_21_pad_groupi_n_1061, csa_tree_add_117_21_pad_groupi_n_1062, csa_tree_add_117_21_pad_groupi_n_1063, csa_tree_add_117_21_pad_groupi_n_1064;
  wire csa_tree_add_117_21_pad_groupi_n_1065, csa_tree_add_117_21_pad_groupi_n_1066, csa_tree_add_117_21_pad_groupi_n_1067, csa_tree_add_117_21_pad_groupi_n_1068, csa_tree_add_117_21_pad_groupi_n_1069, csa_tree_add_117_21_pad_groupi_n_1070, csa_tree_add_117_21_pad_groupi_n_1071, csa_tree_add_117_21_pad_groupi_n_1072;
  wire csa_tree_add_117_21_pad_groupi_n_1073, csa_tree_add_117_21_pad_groupi_n_1074, csa_tree_add_117_21_pad_groupi_n_1075, csa_tree_add_117_21_pad_groupi_n_1076, csa_tree_add_117_21_pad_groupi_n_1077, csa_tree_add_117_21_pad_groupi_n_1078, csa_tree_add_117_21_pad_groupi_n_1079, csa_tree_add_117_21_pad_groupi_n_1080;
  wire csa_tree_add_117_21_pad_groupi_n_1081, csa_tree_add_117_21_pad_groupi_n_1082, csa_tree_add_117_21_pad_groupi_n_1083, csa_tree_add_117_21_pad_groupi_n_1084, csa_tree_add_117_21_pad_groupi_n_1085, csa_tree_add_117_21_pad_groupi_n_1086, csa_tree_add_117_21_pad_groupi_n_1087, csa_tree_add_117_21_pad_groupi_n_1088;
  wire csa_tree_add_117_21_pad_groupi_n_1089, csa_tree_add_117_21_pad_groupi_n_1090, csa_tree_add_117_21_pad_groupi_n_1091, csa_tree_add_117_21_pad_groupi_n_1092, csa_tree_add_117_21_pad_groupi_n_1093, csa_tree_add_117_21_pad_groupi_n_1094, csa_tree_add_117_21_pad_groupi_n_1095, csa_tree_add_117_21_pad_groupi_n_1096;
  wire csa_tree_add_117_21_pad_groupi_n_1097, csa_tree_add_117_21_pad_groupi_n_1098, csa_tree_add_117_21_pad_groupi_n_1099, csa_tree_add_117_21_pad_groupi_n_1100, csa_tree_add_117_21_pad_groupi_n_1101, csa_tree_add_117_21_pad_groupi_n_1102, csa_tree_add_117_21_pad_groupi_n_1103, csa_tree_add_117_21_pad_groupi_n_1104;
  wire csa_tree_add_117_21_pad_groupi_n_1105, csa_tree_add_117_21_pad_groupi_n_1106, csa_tree_add_117_21_pad_groupi_n_1107, csa_tree_add_117_21_pad_groupi_n_1108, csa_tree_add_117_21_pad_groupi_n_1109, csa_tree_add_117_21_pad_groupi_n_1110, csa_tree_add_117_21_pad_groupi_n_1111, csa_tree_add_117_21_pad_groupi_n_1112;
  wire csa_tree_add_117_21_pad_groupi_n_1113, csa_tree_add_117_21_pad_groupi_n_1114, csa_tree_add_117_21_pad_groupi_n_1115, csa_tree_add_117_21_pad_groupi_n_1116, csa_tree_add_117_21_pad_groupi_n_1117, csa_tree_add_117_21_pad_groupi_n_1118, csa_tree_add_117_21_pad_groupi_n_1119, csa_tree_add_117_21_pad_groupi_n_1120;
  wire csa_tree_add_117_21_pad_groupi_n_1121, csa_tree_add_117_21_pad_groupi_n_1122, csa_tree_add_117_21_pad_groupi_n_1123, csa_tree_add_117_21_pad_groupi_n_1124, csa_tree_add_117_21_pad_groupi_n_1125, csa_tree_add_117_21_pad_groupi_n_1126, csa_tree_add_117_21_pad_groupi_n_1127, csa_tree_add_117_21_pad_groupi_n_1128;
  wire csa_tree_add_117_21_pad_groupi_n_1129, csa_tree_add_117_21_pad_groupi_n_1130, csa_tree_add_117_21_pad_groupi_n_1131, csa_tree_add_117_21_pad_groupi_n_1132, csa_tree_add_117_21_pad_groupi_n_1133, csa_tree_add_117_21_pad_groupi_n_1134, csa_tree_add_117_21_pad_groupi_n_1135, csa_tree_add_117_21_pad_groupi_n_1136;
  wire csa_tree_add_117_21_pad_groupi_n_1137, csa_tree_add_117_21_pad_groupi_n_1138, csa_tree_add_117_21_pad_groupi_n_1139, csa_tree_add_117_21_pad_groupi_n_1140, csa_tree_add_117_21_pad_groupi_n_1141, csa_tree_add_117_21_pad_groupi_n_1142, csa_tree_add_117_21_pad_groupi_n_1144, csa_tree_add_117_21_pad_groupi_n_1145;
  wire csa_tree_add_117_21_pad_groupi_n_1147, csa_tree_add_117_21_pad_groupi_n_1148, csa_tree_add_117_21_pad_groupi_n_1150, csa_tree_add_117_21_pad_groupi_n_1151, csa_tree_add_117_21_pad_groupi_n_1153, csa_tree_add_117_21_pad_groupi_n_1154, csa_tree_add_117_21_pad_groupi_n_1156, csa_tree_add_117_21_pad_groupi_n_1157;
  wire csa_tree_add_117_21_pad_groupi_n_1159, csa_tree_add_117_21_pad_groupi_n_1160, csa_tree_add_117_21_pad_groupi_n_1162, csa_tree_add_117_21_pad_groupi_n_1163, csa_tree_add_117_21_pad_groupi_n_1165, csa_tree_add_117_21_pad_groupi_n_1166, csa_tree_add_117_21_pad_groupi_n_1167, csa_tree_add_117_21_pad_groupi_n_1168;
  wire csa_tree_add_117_21_pad_groupi_n_1169, csa_tree_add_117_21_pad_groupi_n_1171, csa_tree_add_117_21_pad_groupi_n_1172, csa_tree_add_117_21_pad_groupi_n_1173, csa_tree_add_117_21_pad_groupi_n_1175, csa_tree_add_117_21_pad_groupi_n_1176, csa_tree_add_117_21_pad_groupi_n_1178, csa_tree_add_117_21_pad_groupi_n_1179;
  wire csa_tree_add_117_21_pad_groupi_n_1181, csa_tree_add_118_30_groupi_n_0, csa_tree_add_118_30_groupi_n_1, csa_tree_add_118_30_groupi_n_2, csa_tree_add_118_30_groupi_n_3, csa_tree_add_118_30_groupi_n_4, csa_tree_add_118_30_groupi_n_5, csa_tree_add_118_30_groupi_n_6;
  wire csa_tree_add_118_30_groupi_n_7, csa_tree_add_118_30_groupi_n_8, csa_tree_add_118_30_groupi_n_9, csa_tree_add_118_30_groupi_n_10, csa_tree_add_118_30_groupi_n_11, csa_tree_add_118_30_groupi_n_12, csa_tree_add_118_30_groupi_n_13, csa_tree_add_118_30_groupi_n_14;
  wire csa_tree_add_118_30_groupi_n_15, csa_tree_add_118_30_groupi_n_16, csa_tree_add_118_30_groupi_n_17, csa_tree_add_118_30_groupi_n_18, csa_tree_add_118_30_groupi_n_19, csa_tree_add_118_30_groupi_n_20, csa_tree_add_118_30_groupi_n_21, csa_tree_add_118_30_groupi_n_22;
  wire csa_tree_add_118_30_groupi_n_23, csa_tree_add_118_30_groupi_n_24, csa_tree_add_118_30_groupi_n_25, csa_tree_add_118_30_groupi_n_26, csa_tree_add_118_30_groupi_n_27, csa_tree_add_118_30_groupi_n_28, csa_tree_add_118_30_groupi_n_29, csa_tree_add_118_30_groupi_n_30;
  wire csa_tree_add_118_30_groupi_n_31, csa_tree_add_118_30_groupi_n_32, csa_tree_add_118_30_groupi_n_33, csa_tree_add_118_30_groupi_n_34, csa_tree_add_118_30_groupi_n_35, csa_tree_add_118_30_groupi_n_36, csa_tree_add_118_30_groupi_n_37, csa_tree_add_118_30_groupi_n_38;
  wire csa_tree_add_118_30_groupi_n_39, csa_tree_add_118_30_groupi_n_40, csa_tree_add_118_30_groupi_n_41, csa_tree_add_118_30_groupi_n_42, csa_tree_add_118_30_groupi_n_43, csa_tree_add_118_30_groupi_n_44, csa_tree_add_118_30_groupi_n_45, csa_tree_add_118_30_groupi_n_46;
  wire csa_tree_add_118_30_groupi_n_47, csa_tree_add_118_30_groupi_n_48, csa_tree_add_118_30_groupi_n_49, csa_tree_add_118_30_groupi_n_50, csa_tree_add_118_30_groupi_n_51, csa_tree_add_118_30_groupi_n_52, csa_tree_add_118_30_groupi_n_53, csa_tree_add_118_30_groupi_n_54;
  wire csa_tree_add_118_30_groupi_n_55, csa_tree_add_118_30_groupi_n_56, csa_tree_add_118_30_groupi_n_57, csa_tree_add_118_30_groupi_n_58, csa_tree_add_118_30_groupi_n_59, csa_tree_add_118_30_groupi_n_60, csa_tree_add_118_30_groupi_n_61, csa_tree_add_118_30_groupi_n_62;
  wire csa_tree_add_118_30_groupi_n_63, csa_tree_add_118_30_groupi_n_64, csa_tree_add_118_30_groupi_n_65, csa_tree_add_118_30_groupi_n_66, csa_tree_add_118_30_groupi_n_67, csa_tree_add_118_30_groupi_n_68, csa_tree_add_118_30_groupi_n_69, csa_tree_add_118_30_groupi_n_70;
  wire csa_tree_add_118_30_groupi_n_71, csa_tree_add_118_30_groupi_n_72, csa_tree_add_118_30_groupi_n_73, csa_tree_add_118_30_groupi_n_74, csa_tree_add_118_30_groupi_n_75, csa_tree_add_118_30_groupi_n_76, csa_tree_add_118_30_groupi_n_77, csa_tree_add_118_30_groupi_n_78;
  wire csa_tree_add_118_30_groupi_n_79, csa_tree_add_118_30_groupi_n_80, csa_tree_add_118_30_groupi_n_81, csa_tree_add_118_30_groupi_n_82, csa_tree_add_118_30_groupi_n_83, csa_tree_add_118_30_groupi_n_84, csa_tree_add_118_30_groupi_n_85, csa_tree_add_118_30_groupi_n_86;
  wire csa_tree_add_118_30_groupi_n_87, csa_tree_add_118_30_groupi_n_88, csa_tree_add_118_30_groupi_n_89, csa_tree_add_118_30_groupi_n_90, csa_tree_add_118_30_groupi_n_91, csa_tree_add_118_30_groupi_n_92, csa_tree_add_118_30_groupi_n_93, csa_tree_add_118_30_groupi_n_94;
  wire csa_tree_add_118_30_groupi_n_95, csa_tree_add_118_30_groupi_n_96, csa_tree_add_118_30_groupi_n_97, csa_tree_add_118_30_groupi_n_98, csa_tree_add_118_30_groupi_n_99, csa_tree_add_118_30_groupi_n_100, csa_tree_add_118_30_groupi_n_101, csa_tree_add_118_30_groupi_n_102;
  wire csa_tree_add_118_30_groupi_n_103, csa_tree_add_118_30_groupi_n_104, csa_tree_add_118_30_groupi_n_105, csa_tree_add_118_30_groupi_n_106, csa_tree_add_118_30_groupi_n_107, csa_tree_add_118_30_groupi_n_109, csa_tree_add_118_30_groupi_n_110, csa_tree_add_118_30_groupi_n_111;
  wire csa_tree_add_118_30_groupi_n_112, csa_tree_add_118_30_groupi_n_113, csa_tree_add_118_30_groupi_n_114, csa_tree_add_118_30_groupi_n_115, csa_tree_add_118_30_groupi_n_116, csa_tree_add_118_30_groupi_n_117, csa_tree_add_118_30_groupi_n_118, csa_tree_add_118_30_groupi_n_119;
  wire csa_tree_add_118_30_groupi_n_120, csa_tree_add_118_30_groupi_n_121, csa_tree_add_118_30_groupi_n_122, csa_tree_add_118_30_groupi_n_123, csa_tree_add_118_30_groupi_n_124, csa_tree_add_118_30_groupi_n_125, csa_tree_add_118_30_groupi_n_126, csa_tree_add_118_30_groupi_n_127;
  wire csa_tree_add_118_30_groupi_n_128, csa_tree_add_118_30_groupi_n_129, csa_tree_add_118_30_groupi_n_130, csa_tree_add_118_30_groupi_n_131, csa_tree_add_118_30_groupi_n_132, csa_tree_add_118_30_groupi_n_133, csa_tree_add_118_30_groupi_n_134, csa_tree_add_118_30_groupi_n_135;
  wire csa_tree_add_118_30_groupi_n_136, csa_tree_add_118_30_groupi_n_137, csa_tree_add_118_30_groupi_n_138, csa_tree_add_118_30_groupi_n_139, csa_tree_add_118_30_groupi_n_140, csa_tree_add_118_30_groupi_n_141, csa_tree_add_118_30_groupi_n_142, csa_tree_add_118_30_groupi_n_143;
  wire csa_tree_add_118_30_groupi_n_144, csa_tree_add_118_30_groupi_n_145, csa_tree_add_118_30_groupi_n_146, csa_tree_add_118_30_groupi_n_147, csa_tree_add_118_30_groupi_n_148, csa_tree_add_118_30_groupi_n_149, csa_tree_add_118_30_groupi_n_150, csa_tree_add_118_30_groupi_n_152;
  wire csa_tree_add_118_30_groupi_n_153, csa_tree_add_118_30_groupi_n_154, csa_tree_add_118_30_groupi_n_155, csa_tree_add_118_30_groupi_n_156, csa_tree_add_118_30_groupi_n_157, csa_tree_add_118_30_groupi_n_158, csa_tree_add_118_30_groupi_n_159, csa_tree_add_118_30_groupi_n_160;
  wire csa_tree_add_118_30_groupi_n_161, csa_tree_add_118_30_groupi_n_162, csa_tree_add_118_30_groupi_n_164, csa_tree_add_118_30_groupi_n_165, csa_tree_add_118_30_groupi_n_166, csa_tree_add_118_30_groupi_n_167, csa_tree_add_118_30_groupi_n_168, csa_tree_add_118_30_groupi_n_170;
  wire csa_tree_add_118_30_groupi_n_171, csa_tree_add_118_30_groupi_n_172, csa_tree_add_118_30_groupi_n_173, csa_tree_add_118_30_groupi_n_174, csa_tree_add_118_30_groupi_n_175, csa_tree_add_118_30_groupi_n_176, csa_tree_add_118_30_groupi_n_177, csa_tree_add_118_30_groupi_n_179;
  wire csa_tree_add_118_30_groupi_n_180, csa_tree_add_118_30_groupi_n_181, csa_tree_add_118_30_groupi_n_182, csa_tree_add_118_30_groupi_n_184, csa_tree_add_118_30_groupi_n_185, csa_tree_add_118_30_groupi_n_187, csa_tree_add_118_30_groupi_n_188, csa_tree_add_118_30_groupi_n_190;
  wire csa_tree_add_118_30_groupi_n_191, csa_tree_add_118_30_groupi_n_193, csa_tree_add_118_30_groupi_n_194, csa_tree_add_118_30_groupi_n_196, csa_tree_add_118_30_groupi_n_197, csa_tree_add_118_30_groupi_n_199, csa_tree_add_118_30_groupi_n_200, csa_tree_add_118_30_groupi_n_202;
  wire csa_tree_add_118_30_groupi_n_203, csa_tree_add_118_30_groupi_n_205, csa_tree_add_118_30_groupi_n_206, csa_tree_add_118_30_groupi_n_208, csa_tree_add_118_30_groupi_n_209, csa_tree_add_118_30_groupi_n_211, csa_tree_sub_77_21_n_13, csa_tree_sub_77_21_n_14;
  wire csa_tree_sub_77_21_n_15, csa_tree_sub_77_21_n_17, csa_tree_sub_77_21_n_18, csa_tree_sub_77_21_n_19, csa_tree_sub_77_21_n_20, csa_tree_sub_77_21_n_21, csa_tree_sub_77_21_n_24, csa_tree_sub_77_21_n_25;
  wire csa_tree_sub_77_21_n_26, csa_tree_sub_77_21_n_27, csa_tree_sub_77_21_n_28, csa_tree_sub_77_21_n_29, csa_tree_sub_77_21_n_30, csa_tree_sub_77_21_n_31, csa_tree_sub_77_21_n_32, csa_tree_sub_80_22_n_2;
  wire csa_tree_sub_80_22_n_3, csa_tree_sub_80_22_n_4, csa_tree_sub_80_22_n_6, csa_tree_sub_86_22_n_2, csa_tree_sub_86_22_n_3, csa_tree_sub_86_22_n_4, csa_tree_sub_86_22_n_6, csa_tree_sub_92_22_n_2;
  wire csa_tree_sub_92_22_n_3, csa_tree_sub_92_22_n_4, csa_tree_sub_92_22_n_6, csa_tree_sub_98_22_n_2, csa_tree_sub_98_22_n_3, csa_tree_sub_98_22_n_4, csa_tree_sub_98_22_n_6, csa_tree_sub_104_22_n_2;
  wire csa_tree_sub_104_22_n_3, csa_tree_sub_104_22_n_4, csa_tree_sub_104_22_n_6, mul_84_22_n_0, mul_84_22_n_1, mul_84_22_n_2, mul_84_22_n_3, mul_84_22_n_4;
  wire mul_84_22_n_5, mul_84_22_n_6, mul_84_22_n_7, mul_84_22_n_8, mul_84_22_n_9, mul_84_22_n_10, mul_84_22_n_11, mul_84_22_n_12;
  wire mul_84_22_n_13, mul_84_22_n_14, mul_84_22_n_15, mul_84_22_n_16, mul_84_22_n_17, mul_84_22_n_18, mul_84_22_n_19, mul_84_22_n_20;
  wire mul_84_22_n_21, mul_84_22_n_22, mul_84_22_n_23, mul_84_22_n_24, mul_84_22_n_25, mul_84_22_n_26, mul_84_22_n_27, mul_84_22_n_28;
  wire mul_84_22_n_29, mul_84_22_n_30, mul_84_22_n_31, mul_84_22_n_32, mul_84_22_n_33, mul_84_22_n_34, mul_84_22_n_35, mul_84_22_n_36;
  wire mul_84_22_n_37, mul_84_22_n_38, mul_84_22_n_39, mul_84_22_n_40, mul_84_22_n_41, mul_84_22_n_42, mul_84_22_n_43, mul_84_22_n_44;
  wire mul_84_22_n_45, mul_84_22_n_46, mul_84_22_n_47, mul_84_22_n_48, mul_84_22_n_49, mul_84_22_n_50, mul_84_22_n_51, mul_84_22_n_52;
  wire mul_84_22_n_53, mul_84_22_n_54, mul_84_22_n_55, mul_84_22_n_56, mul_84_22_n_57, mul_84_22_n_58, mul_84_22_n_59, mul_84_22_n_60;
  wire mul_84_22_n_61, mul_84_22_n_62, mul_84_22_n_63, mul_84_22_n_64, mul_84_22_n_65, mul_84_22_n_66, mul_84_22_n_67, mul_84_22_n_68;
  wire mul_84_22_n_69, mul_84_22_n_70, mul_84_22_n_71, mul_84_22_n_72, mul_84_22_n_73, mul_84_22_n_74, mul_84_22_n_75, mul_84_22_n_76;
  wire mul_84_22_n_77, mul_84_22_n_78, mul_84_22_n_79, mul_84_22_n_80, mul_84_22_n_81, mul_84_22_n_82, mul_84_22_n_83, mul_84_22_n_84;
  wire mul_84_22_n_85, mul_84_22_n_86, mul_84_22_n_87, mul_84_22_n_88, mul_84_22_n_89, mul_84_22_n_90, mul_84_22_n_91, mul_84_22_n_92;
  wire mul_84_22_n_93, mul_84_22_n_94, mul_84_22_n_95, mul_84_22_n_96, mul_84_22_n_97, mul_84_22_n_98, mul_84_22_n_99, mul_84_22_n_100;
  wire mul_84_22_n_101, mul_84_22_n_102, mul_84_22_n_103, mul_84_22_n_104, mul_84_22_n_105, mul_84_22_n_106, mul_84_22_n_107, mul_84_22_n_108;
  wire mul_84_22_n_109, mul_84_22_n_110, mul_84_22_n_111, mul_84_22_n_112, mul_84_22_n_113, mul_84_22_n_114, mul_84_22_n_115, mul_84_22_n_116;
  wire mul_84_22_n_117, mul_84_22_n_118, mul_84_22_n_119, mul_84_22_n_120, mul_84_22_n_121, mul_84_22_n_122, mul_84_22_n_123, mul_84_22_n_124;
  wire mul_84_22_n_125, mul_84_22_n_126, mul_84_22_n_127, mul_84_22_n_128, mul_84_22_n_129, mul_84_22_n_130, mul_84_22_n_131, mul_84_22_n_132;
  wire mul_84_22_n_133, mul_84_22_n_134, mul_84_22_n_135, mul_84_22_n_136, mul_84_22_n_137, mul_84_22_n_138, mul_84_22_n_139, mul_84_22_n_140;
  wire mul_84_22_n_141, mul_84_22_n_142, mul_84_22_n_143, mul_84_22_n_144, mul_84_22_n_145, mul_84_22_n_146, mul_84_22_n_147, mul_84_22_n_148;
  wire mul_84_22_n_149, mul_84_22_n_150, mul_84_22_n_151, mul_84_22_n_152, mul_84_22_n_153, mul_84_22_n_154, mul_84_22_n_155, mul_84_22_n_156;
  wire mul_84_22_n_157, mul_84_22_n_158, mul_84_22_n_159, mul_84_22_n_160, mul_84_22_n_161, mul_84_22_n_162, mul_84_22_n_163, mul_84_22_n_164;
  wire mul_84_22_n_165, mul_84_22_n_166, mul_84_22_n_167, mul_84_22_n_168, mul_84_22_n_169, mul_84_22_n_170, mul_84_22_n_171, mul_84_22_n_172;
  wire mul_84_22_n_173, mul_84_22_n_174, mul_84_22_n_175, mul_84_22_n_176, mul_84_22_n_177, mul_84_22_n_178, mul_84_22_n_179, mul_84_22_n_180;
  wire mul_84_22_n_181, mul_84_22_n_182, mul_84_22_n_198, mul_84_22_n_199, mul_84_22_n_200, mul_84_22_n_201, mul_84_22_n_202, mul_84_22_n_203;
  wire mul_84_22_n_204, mul_84_22_n_205, mul_84_22_n_206, mul_84_22_n_207, mul_84_22_n_208, mul_84_22_n_209, mul_84_22_n_210, mul_84_22_n_211;
  wire mul_84_22_n_212, mul_84_22_n_213, mul_84_22_n_214, mul_84_22_n_215, mul_84_22_n_216, mul_84_22_n_217, mul_84_22_n_218, mul_84_22_n_219;
  wire mul_84_22_n_220, mul_84_22_n_221, mul_84_22_n_222, mul_84_22_n_223, mul_84_22_n_224, mul_84_22_n_225, mul_84_22_n_226, mul_84_22_n_227;
  wire mul_84_22_n_228, mul_84_22_n_229, mul_84_22_n_230, mul_84_22_n_231, mul_84_22_n_232, mul_84_22_n_233, mul_84_22_n_234, mul_84_22_n_235;
  wire mul_84_22_n_236, mul_84_22_n_237, mul_84_22_n_238, mul_84_22_n_239, mul_84_22_n_240, mul_84_22_n_241, mul_84_22_n_242, mul_84_22_n_243;
  wire mul_84_22_n_244, mul_84_22_n_245, mul_84_22_n_246, mul_84_22_n_247, mul_84_22_n_248, mul_84_22_n_249, mul_84_22_n_250, mul_84_22_n_251;
  wire mul_84_22_n_252, mul_84_22_n_253, mul_84_22_n_254, mul_84_22_n_255, mul_84_22_n_256, mul_84_22_n_257, mul_84_22_n_258, mul_84_22_n_259;
  wire mul_84_22_n_260, mul_84_22_n_261, mul_84_22_n_262, mul_84_22_n_263, mul_84_22_n_264, mul_84_22_n_265, mul_84_22_n_266, mul_84_22_n_267;
  wire mul_84_22_n_268, mul_84_22_n_269, mul_84_22_n_270, mul_84_22_n_271, mul_84_22_n_272, mul_84_22_n_273, mul_84_22_n_274, mul_84_22_n_275;
  wire mul_84_22_n_276, mul_84_22_n_277, mul_84_22_n_278, mul_84_22_n_279, mul_84_22_n_280, mul_84_22_n_281, mul_84_22_n_282, mul_84_22_n_283;
  wire mul_84_22_n_284, mul_84_22_n_285, mul_84_22_n_286, mul_84_22_n_287, mul_84_22_n_288, mul_84_22_n_289, mul_84_22_n_290, mul_84_22_n_291;
  wire mul_84_22_n_292, mul_84_22_n_293, mul_84_22_n_294, mul_84_22_n_295, mul_84_22_n_296, mul_84_22_n_297, mul_84_22_n_298, mul_84_22_n_299;
  wire mul_84_22_n_300, mul_84_22_n_301, mul_84_22_n_302, mul_84_22_n_303, mul_84_22_n_304, mul_84_22_n_305, mul_84_22_n_306, mul_84_22_n_307;
  wire mul_84_22_n_308, mul_84_22_n_310, mul_84_22_n_311, mul_84_22_n_312, mul_84_22_n_313, mul_84_22_n_314, mul_84_22_n_315, mul_84_22_n_316;
  wire mul_84_22_n_317, mul_84_22_n_318, mul_84_22_n_319, mul_84_22_n_320, mul_84_22_n_321, mul_84_22_n_322, mul_84_22_n_323, mul_84_22_n_324;
  wire mul_84_22_n_325, mul_84_22_n_326, mul_84_22_n_327, mul_84_22_n_328, mul_84_22_n_329, mul_84_22_n_330, mul_84_22_n_331, mul_84_22_n_332;
  wire mul_84_22_n_333, mul_84_22_n_334, mul_84_22_n_335, mul_84_22_n_336, mul_84_22_n_337, mul_84_22_n_338, mul_84_22_n_339, mul_84_22_n_340;
  wire mul_84_22_n_341, mul_84_22_n_342, mul_84_22_n_343, mul_84_22_n_344, mul_84_22_n_345, mul_84_22_n_346, mul_84_22_n_347, mul_84_22_n_348;
  wire mul_84_22_n_349, mul_84_22_n_350, mul_84_22_n_351, mul_84_22_n_352, mul_84_22_n_353, mul_84_22_n_354, mul_84_22_n_355, mul_84_22_n_356;
  wire mul_84_22_n_357, mul_84_22_n_358, mul_84_22_n_359, mul_84_22_n_360, mul_84_22_n_361, mul_84_22_n_362, mul_84_22_n_363, mul_84_22_n_364;
  wire mul_84_22_n_365, mul_84_22_n_366, mul_84_22_n_367, mul_84_22_n_368, mul_84_22_n_369, mul_84_22_n_370, mul_84_22_n_371, mul_84_22_n_372;
  wire mul_84_22_n_373, mul_84_22_n_374, mul_84_22_n_375, mul_84_22_n_376, mul_84_22_n_377, mul_84_22_n_378, mul_84_22_n_379, mul_84_22_n_380;
  wire mul_84_22_n_381, mul_84_22_n_382, mul_84_22_n_383, mul_84_22_n_384, mul_84_22_n_385, mul_84_22_n_386, mul_84_22_n_387, mul_84_22_n_388;
  wire mul_84_22_n_389, mul_84_22_n_390, mul_84_22_n_391, mul_84_22_n_392, mul_84_22_n_393, mul_84_22_n_394, mul_84_22_n_395, mul_84_22_n_396;
  wire mul_84_22_n_397, mul_84_22_n_398, mul_84_22_n_399, mul_84_22_n_400, mul_84_22_n_401, mul_84_22_n_402, mul_84_22_n_403, mul_84_22_n_404;
  wire mul_84_22_n_405, mul_84_22_n_406, mul_84_22_n_407, mul_84_22_n_408, mul_84_22_n_409, mul_84_22_n_410, mul_84_22_n_411, mul_84_22_n_412;
  wire mul_84_22_n_413, mul_84_22_n_414, mul_84_22_n_415, mul_84_22_n_416, mul_84_22_n_417, mul_84_22_n_418, mul_84_22_n_419, mul_84_22_n_420;
  wire mul_84_22_n_421, mul_84_22_n_422, mul_84_22_n_423, mul_84_22_n_424, mul_84_22_n_425, mul_84_22_n_426, mul_84_22_n_427, mul_84_22_n_428;
  wire mul_84_22_n_429, mul_84_22_n_430, mul_84_22_n_431, mul_84_22_n_432, mul_84_22_n_433, mul_84_22_n_434, mul_84_22_n_435, mul_84_22_n_436;
  wire mul_84_22_n_437, mul_84_22_n_438, mul_84_22_n_439, mul_84_22_n_440, mul_84_22_n_441, mul_84_22_n_442, mul_84_22_n_443, mul_84_22_n_444;
  wire mul_84_22_n_445, mul_84_22_n_446, mul_84_22_n_447, mul_84_22_n_448, mul_84_22_n_449, mul_84_22_n_450, mul_84_22_n_451, mul_84_22_n_452;
  wire mul_84_22_n_453, mul_84_22_n_454, mul_84_22_n_455, mul_84_22_n_456, mul_84_22_n_457, mul_84_22_n_458, mul_84_22_n_459, mul_84_22_n_460;
  wire mul_84_22_n_461, mul_84_22_n_462, mul_84_22_n_463, mul_84_22_n_464, mul_84_22_n_465, mul_84_22_n_466, mul_84_22_n_467, mul_84_22_n_468;
  wire mul_84_22_n_469, mul_84_22_n_470, mul_84_22_n_471, mul_84_22_n_472, mul_84_22_n_473, mul_84_22_n_474, mul_84_22_n_475, mul_84_22_n_476;
  wire mul_84_22_n_477, mul_84_22_n_478, mul_84_22_n_479, mul_84_22_n_480, mul_84_22_n_481, mul_84_22_n_482, mul_84_22_n_483, mul_84_22_n_484;
  wire mul_84_22_n_485, mul_84_22_n_486, mul_84_22_n_487, mul_84_22_n_488, mul_84_22_n_489, mul_84_22_n_490, mul_84_22_n_491, mul_84_22_n_492;
  wire mul_84_22_n_493, mul_84_22_n_494, mul_84_22_n_495, mul_84_22_n_496, mul_84_22_n_497, mul_84_22_n_498, mul_84_22_n_499, mul_84_22_n_500;
  wire mul_84_22_n_501, mul_84_22_n_502, mul_84_22_n_503, mul_84_22_n_504, mul_84_22_n_505, mul_84_22_n_506, mul_84_22_n_507, mul_84_22_n_508;
  wire mul_84_22_n_509, mul_84_22_n_510, mul_84_22_n_511, mul_84_22_n_512, mul_84_22_n_513, mul_84_22_n_514, mul_84_22_n_515, mul_84_22_n_516;
  wire mul_84_22_n_517, mul_84_22_n_518, mul_84_22_n_519, mul_84_22_n_520, mul_84_22_n_521, mul_84_22_n_522, mul_84_22_n_523, mul_84_22_n_524;
  wire mul_84_22_n_525, mul_84_22_n_526, mul_84_22_n_527, mul_84_22_n_528, mul_84_22_n_529, mul_84_22_n_530, mul_84_22_n_531, mul_84_22_n_532;
  wire mul_84_22_n_533, mul_84_22_n_534, mul_84_22_n_535, mul_84_22_n_536, mul_84_22_n_537, mul_84_22_n_538, mul_84_22_n_539, mul_84_22_n_540;
  wire mul_84_22_n_541, mul_84_22_n_542, mul_84_22_n_543, mul_84_22_n_544, mul_84_22_n_545, mul_84_22_n_546, mul_84_22_n_547, mul_84_22_n_548;
  wire mul_84_22_n_549, mul_84_22_n_550, mul_84_22_n_551, mul_84_22_n_552, mul_84_22_n_553, mul_84_22_n_554, mul_84_22_n_555, mul_84_22_n_556;
  wire mul_84_22_n_557, mul_84_22_n_558, mul_84_22_n_559, mul_84_22_n_560, mul_84_22_n_561, mul_84_22_n_562, mul_84_22_n_563, mul_84_22_n_564;
  wire mul_84_22_n_565, mul_84_22_n_566, mul_84_22_n_567, mul_84_22_n_568, mul_84_22_n_569, mul_84_22_n_570, mul_84_22_n_571, mul_84_22_n_572;
  wire mul_84_22_n_573, mul_84_22_n_574, mul_84_22_n_575, mul_84_22_n_576, mul_84_22_n_577, mul_84_22_n_578, mul_84_22_n_579, mul_84_22_n_580;
  wire mul_84_22_n_581, mul_84_22_n_582, mul_84_22_n_583, mul_84_22_n_584, mul_84_22_n_585, mul_84_22_n_586, mul_84_22_n_587, mul_84_22_n_588;
  wire mul_84_22_n_589, mul_84_22_n_590, mul_84_22_n_591, mul_84_22_n_592, mul_84_22_n_593, mul_84_22_n_594, mul_84_22_n_595, mul_84_22_n_596;
  wire mul_84_22_n_597, mul_84_22_n_598, mul_84_22_n_599, mul_84_22_n_600, mul_84_22_n_601, mul_84_22_n_602, mul_84_22_n_603, mul_84_22_n_604;
  wire mul_84_22_n_605, mul_84_22_n_606, mul_84_22_n_607, mul_84_22_n_608, mul_84_22_n_609, mul_84_22_n_610, mul_84_22_n_611, mul_84_22_n_612;
  wire mul_84_22_n_613, mul_84_22_n_614, mul_84_22_n_615, mul_84_22_n_616, mul_84_22_n_617, mul_84_22_n_618, mul_84_22_n_619, mul_84_22_n_620;
  wire mul_84_22_n_621, mul_84_22_n_622, mul_84_22_n_623, mul_84_22_n_624, mul_84_22_n_625, mul_84_22_n_626, mul_84_22_n_627, mul_84_22_n_628;
  wire mul_84_22_n_629, mul_84_22_n_630, mul_84_22_n_631, mul_84_22_n_632, mul_84_22_n_633, mul_84_22_n_634, mul_84_22_n_635, mul_84_22_n_636;
  wire mul_84_22_n_637, mul_84_22_n_638, mul_84_22_n_639, mul_84_22_n_640, mul_84_22_n_641, mul_84_22_n_642, mul_84_22_n_643, mul_84_22_n_644;
  wire mul_84_22_n_645, mul_84_22_n_646, mul_84_22_n_647, mul_84_22_n_648, mul_84_22_n_649, mul_84_22_n_650, mul_84_22_n_651, mul_84_22_n_652;
  wire mul_84_22_n_653, mul_84_22_n_654, mul_84_22_n_655, mul_84_22_n_656, mul_84_22_n_657, mul_84_22_n_658, mul_84_22_n_659, mul_84_22_n_660;
  wire mul_84_22_n_661, mul_84_22_n_662, mul_84_22_n_663, mul_84_22_n_664, mul_84_22_n_665, mul_84_22_n_666, mul_84_22_n_667, mul_84_22_n_668;
  wire mul_84_22_n_669, mul_84_22_n_670, mul_84_22_n_671, mul_84_22_n_672, mul_84_22_n_673, mul_84_22_n_674, mul_84_22_n_675, mul_84_22_n_676;
  wire mul_84_22_n_677, mul_84_22_n_678, mul_84_22_n_679, mul_84_22_n_680, mul_84_22_n_681, mul_84_22_n_682, mul_84_22_n_683, mul_84_22_n_684;
  wire mul_84_22_n_685, mul_84_22_n_686, mul_84_22_n_687, mul_84_22_n_688, mul_84_22_n_689, mul_84_22_n_690, mul_84_22_n_691, mul_84_22_n_692;
  wire mul_84_22_n_693, mul_84_22_n_694, mul_84_22_n_695, mul_84_22_n_696, mul_84_22_n_697, mul_84_22_n_698, mul_84_22_n_699, mul_84_22_n_700;
  wire mul_84_22_n_701, mul_84_22_n_702, mul_84_22_n_703, mul_84_22_n_704, mul_84_22_n_705, mul_84_22_n_706, mul_84_22_n_707, mul_84_22_n_708;
  wire mul_84_22_n_709, mul_84_22_n_710, mul_84_22_n_711, mul_84_22_n_712, mul_84_22_n_713, mul_84_22_n_714, mul_84_22_n_715, mul_84_22_n_716;
  wire mul_84_22_n_717, mul_84_22_n_718, mul_84_22_n_719, mul_84_22_n_720, mul_84_22_n_721, mul_84_22_n_722, mul_84_22_n_723, mul_84_22_n_724;
  wire mul_84_22_n_725, mul_84_22_n_726, mul_84_22_n_727, mul_84_22_n_728, mul_84_22_n_729, mul_84_22_n_730, mul_84_22_n_731, mul_84_22_n_732;
  wire mul_84_22_n_733, mul_84_22_n_734, mul_84_22_n_735, mul_84_22_n_736, mul_84_22_n_737, mul_84_22_n_738, mul_84_22_n_739, mul_84_22_n_740;
  wire mul_84_22_n_741, mul_84_22_n_742, mul_84_22_n_743, mul_84_22_n_744, mul_84_22_n_745, mul_84_22_n_746, mul_84_22_n_747, mul_84_22_n_748;
  wire mul_84_22_n_749, mul_84_22_n_750, mul_84_22_n_751, mul_84_22_n_752, mul_84_22_n_753, mul_84_22_n_754, mul_84_22_n_755, mul_84_22_n_756;
  wire mul_84_22_n_757, mul_84_22_n_758, mul_84_22_n_759, mul_84_22_n_760, mul_84_22_n_761, mul_84_22_n_762, mul_84_22_n_763, mul_84_22_n_764;
  wire mul_84_22_n_765, mul_84_22_n_766, mul_84_22_n_767, mul_84_22_n_768, mul_84_22_n_769, mul_84_22_n_770, mul_84_22_n_771, mul_84_22_n_772;
  wire mul_84_22_n_773, mul_84_22_n_774, mul_84_22_n_775, mul_84_22_n_776, mul_84_22_n_777, mul_84_22_n_778, mul_84_22_n_779, mul_84_22_n_780;
  wire mul_84_22_n_781, mul_84_22_n_782, mul_84_22_n_783, mul_84_22_n_784, mul_84_22_n_785, mul_84_22_n_786, mul_84_22_n_787, mul_84_22_n_788;
  wire mul_84_22_n_789, mul_84_22_n_790, mul_84_22_n_791, mul_84_22_n_792, mul_84_22_n_793, mul_84_22_n_794, mul_84_22_n_795, mul_84_22_n_796;
  wire mul_84_22_n_797, mul_84_22_n_798, mul_84_22_n_799, mul_84_22_n_800, mul_84_22_n_801, mul_84_22_n_802, mul_84_22_n_803, mul_84_22_n_804;
  wire mul_84_22_n_805, mul_84_22_n_806, mul_84_22_n_807, mul_84_22_n_808, mul_84_22_n_809, mul_84_22_n_810, mul_84_22_n_811, mul_84_22_n_812;
  wire mul_84_22_n_813, mul_84_22_n_814, mul_84_22_n_815, mul_84_22_n_816, mul_84_22_n_817, mul_84_22_n_818, mul_84_22_n_819, mul_84_22_n_820;
  wire mul_84_22_n_821, mul_84_22_n_822, mul_84_22_n_823, mul_84_22_n_824, mul_84_22_n_825, mul_84_22_n_826, mul_84_22_n_827, mul_84_22_n_828;
  wire mul_84_22_n_829, mul_84_22_n_830, mul_84_22_n_831, mul_84_22_n_832, mul_84_22_n_833, mul_84_22_n_834, mul_84_22_n_835, mul_84_22_n_836;
  wire mul_84_22_n_837, mul_84_22_n_838, mul_84_22_n_839, mul_84_22_n_840, mul_84_22_n_841, mul_84_22_n_842, mul_84_22_n_843, mul_84_22_n_844;
  wire mul_84_22_n_845, mul_84_22_n_846, mul_84_22_n_847, mul_84_22_n_848, mul_84_22_n_849, mul_84_22_n_850, mul_84_22_n_851, mul_84_22_n_852;
  wire mul_84_22_n_853, mul_84_22_n_854, mul_84_22_n_855, mul_84_22_n_856, mul_84_22_n_857, mul_84_22_n_858, mul_84_22_n_859, mul_84_22_n_860;
  wire mul_84_22_n_861, mul_84_22_n_862, mul_84_22_n_863, mul_84_22_n_864, mul_84_22_n_865, mul_84_22_n_866, mul_84_22_n_867, mul_84_22_n_868;
  wire mul_84_22_n_869, mul_84_22_n_870, mul_84_22_n_871, mul_84_22_n_872, mul_84_22_n_873, mul_84_22_n_874, mul_84_22_n_875, mul_84_22_n_876;
  wire mul_84_22_n_877, mul_84_22_n_878, mul_84_22_n_879, mul_84_22_n_880, mul_84_22_n_881, mul_84_22_n_882, mul_84_22_n_883, mul_84_22_n_884;
  wire mul_84_22_n_885, mul_84_22_n_886, mul_84_22_n_887, mul_84_22_n_888, mul_84_22_n_889, mul_84_22_n_890, mul_84_22_n_891, mul_84_22_n_892;
  wire mul_84_22_n_893, mul_84_22_n_894, mul_84_22_n_895, mul_84_22_n_896, mul_84_22_n_897, mul_84_22_n_898, mul_84_22_n_899, mul_84_22_n_900;
  wire mul_84_22_n_901, mul_84_22_n_902, mul_84_22_n_903, mul_84_22_n_904, mul_84_22_n_905, mul_84_22_n_906, mul_84_22_n_907, mul_84_22_n_908;
  wire mul_84_22_n_909, mul_84_22_n_910, mul_84_22_n_911, mul_84_22_n_912, mul_84_22_n_913, mul_84_22_n_914, mul_84_22_n_915, mul_84_22_n_916;
  wire mul_84_22_n_917, mul_84_22_n_918, mul_84_22_n_919, mul_84_22_n_920, mul_84_22_n_921, mul_84_22_n_922, mul_84_22_n_923, mul_84_22_n_924;
  wire mul_84_22_n_925, mul_84_22_n_926, mul_84_22_n_927, mul_84_22_n_928, mul_84_22_n_929, mul_84_22_n_930, mul_84_22_n_931, mul_84_22_n_932;
  wire mul_84_22_n_933, mul_84_22_n_934, mul_84_22_n_935, mul_84_22_n_936, mul_84_22_n_937, mul_84_22_n_938, mul_84_22_n_939, mul_84_22_n_940;
  wire mul_84_22_n_941, mul_84_22_n_942, mul_84_22_n_943, mul_84_22_n_944, mul_84_22_n_945, mul_84_22_n_946, mul_84_22_n_947, mul_84_22_n_948;
  wire mul_84_22_n_949, mul_84_22_n_950, mul_84_22_n_951, mul_84_22_n_952, mul_84_22_n_953, mul_84_22_n_954, mul_84_22_n_955, mul_84_22_n_956;
  wire mul_84_22_n_957, mul_84_22_n_958, mul_84_22_n_959, mul_84_22_n_960, mul_84_22_n_961, mul_84_22_n_962, mul_84_22_n_963, mul_84_22_n_964;
  wire mul_84_22_n_965, mul_84_22_n_966, mul_84_22_n_967, mul_84_22_n_968, mul_84_22_n_969, mul_84_22_n_970, mul_84_22_n_971, mul_84_22_n_972;
  wire mul_84_22_n_973, mul_84_22_n_974, mul_84_22_n_975, mul_84_22_n_976, mul_84_22_n_977, mul_84_22_n_978, mul_84_22_n_979, mul_84_22_n_980;
  wire mul_84_22_n_981, mul_84_22_n_982, mul_84_22_n_983, mul_84_22_n_984, mul_84_22_n_985, mul_84_22_n_986, mul_84_22_n_987, mul_84_22_n_988;
  wire mul_84_22_n_989, mul_84_22_n_990, mul_84_22_n_991, mul_84_22_n_992, mul_84_22_n_993, mul_84_22_n_994, mul_84_22_n_995, mul_84_22_n_996;
  wire mul_84_22_n_997, mul_84_22_n_998, mul_84_22_n_999, mul_84_22_n_1000, mul_84_22_n_1001, mul_84_22_n_1002, mul_84_22_n_1003, mul_84_22_n_1004;
  wire mul_84_22_n_1005, mul_84_22_n_1006, mul_84_22_n_1007, mul_84_22_n_1008, mul_84_22_n_1009, mul_84_22_n_1010, mul_84_22_n_1011, mul_84_22_n_1012;
  wire mul_84_22_n_1013, mul_84_22_n_1014, mul_84_22_n_1015, mul_84_22_n_1016, mul_84_22_n_1017, mul_84_22_n_1018, mul_84_22_n_1019, mul_84_22_n_1020;
  wire mul_84_22_n_1021, mul_84_22_n_1022, mul_84_22_n_1023, mul_84_22_n_1024, mul_84_22_n_1025, mul_84_22_n_1026, mul_84_22_n_1027, mul_84_22_n_1028;
  wire mul_84_22_n_1029, mul_84_22_n_1030, mul_84_22_n_1031, mul_84_22_n_1032, mul_84_22_n_1033, mul_84_22_n_1034, mul_84_22_n_1035, mul_84_22_n_1036;
  wire mul_84_22_n_1037, mul_84_22_n_1038, mul_84_22_n_1039, mul_84_22_n_1040, mul_84_22_n_1041, mul_84_22_n_1042, mul_84_22_n_1043, mul_84_22_n_1044;
  wire mul_84_22_n_1045, mul_84_22_n_1046, mul_84_22_n_1047, mul_84_22_n_1048, mul_84_22_n_1049, mul_84_22_n_1050, mul_84_22_n_1051, mul_84_22_n_1052;
  wire mul_84_22_n_1053, mul_84_22_n_1054, mul_84_22_n_1055, mul_84_22_n_1056, mul_84_22_n_1057, mul_84_22_n_1058, mul_84_22_n_1059, mul_84_22_n_1060;
  wire mul_84_22_n_1061, mul_84_22_n_1062, mul_84_22_n_1063, mul_84_22_n_1064, mul_84_22_n_1065, mul_84_22_n_1066, mul_84_22_n_1067, mul_84_22_n_1068;
  wire mul_84_22_n_1069, mul_84_22_n_1070, mul_84_22_n_1071, mul_84_22_n_1072, mul_84_22_n_1073, mul_84_22_n_1074, mul_84_22_n_1075, mul_84_22_n_1076;
  wire mul_84_22_n_1077, mul_84_22_n_1078, mul_84_22_n_1079, mul_84_22_n_1080, mul_84_22_n_1081, mul_84_22_n_1082, mul_84_22_n_1083, mul_84_22_n_1084;
  wire mul_84_22_n_1085, mul_84_22_n_1086, mul_84_22_n_1087, mul_84_22_n_1088, mul_84_22_n_1089, mul_84_22_n_1090, mul_84_22_n_1091, mul_84_22_n_1092;
  wire mul_84_22_n_1093, mul_84_22_n_1094, mul_84_22_n_1095, mul_84_22_n_1096, mul_84_22_n_1097, mul_84_22_n_1098, mul_84_22_n_1099, mul_84_22_n_1100;
  wire mul_84_22_n_1101, mul_84_22_n_1102, mul_84_22_n_1103, mul_84_22_n_1104, mul_84_22_n_1105, mul_84_22_n_1106, mul_84_22_n_1107, mul_84_22_n_1108;
  wire mul_84_22_n_1109, mul_84_22_n_1110, mul_84_22_n_1111, mul_84_22_n_1112, mul_84_22_n_1113, mul_84_22_n_1114, mul_84_22_n_1115, mul_84_22_n_1116;
  wire mul_84_22_n_1117, mul_84_22_n_1118, mul_84_22_n_1119, mul_84_22_n_1120, mul_84_22_n_1121, mul_84_22_n_1122, mul_84_22_n_1123, mul_84_22_n_1124;
  wire mul_84_22_n_1125, mul_84_22_n_1126, mul_84_22_n_1127, mul_84_22_n_1128, mul_84_22_n_1129, mul_84_22_n_1130, mul_84_22_n_1131, mul_84_22_n_1132;
  wire mul_84_22_n_1133, mul_84_22_n_1134, mul_84_22_n_1135, mul_84_22_n_1136, mul_84_22_n_1137, mul_84_22_n_1138, mul_84_22_n_1139, mul_84_22_n_1140;
  wire mul_84_22_n_1141, mul_84_22_n_1142, mul_84_22_n_1143, mul_84_22_n_1144, mul_84_22_n_1145, mul_84_22_n_1146, mul_84_22_n_1147, mul_84_22_n_1148;
  wire mul_84_22_n_1149, mul_84_22_n_1150, mul_84_22_n_1151, mul_84_22_n_1152, mul_84_22_n_1153, mul_84_22_n_1154, mul_84_22_n_1155, mul_84_22_n_1156;
  wire mul_84_22_n_1157, mul_90_22_n_0, mul_90_22_n_1, mul_90_22_n_2, mul_90_22_n_3, mul_90_22_n_4, mul_90_22_n_5, mul_90_22_n_6;
  wire mul_90_22_n_7, mul_90_22_n_8, mul_90_22_n_9, mul_90_22_n_10, mul_90_22_n_11, mul_90_22_n_12, mul_90_22_n_13, mul_90_22_n_14;
  wire mul_90_22_n_15, mul_90_22_n_16, mul_90_22_n_17, mul_90_22_n_18, mul_90_22_n_19, mul_90_22_n_20, mul_90_22_n_21, mul_90_22_n_22;
  wire mul_90_22_n_23, mul_90_22_n_24, mul_90_22_n_25, mul_90_22_n_26, mul_90_22_n_27, mul_90_22_n_28, mul_90_22_n_29, mul_90_22_n_30;
  wire mul_90_22_n_31, mul_90_22_n_32, mul_90_22_n_33, mul_90_22_n_34, mul_90_22_n_35, mul_90_22_n_36, mul_90_22_n_37, mul_90_22_n_38;
  wire mul_90_22_n_39, mul_90_22_n_40, mul_90_22_n_41, mul_90_22_n_42, mul_90_22_n_43, mul_90_22_n_44, mul_90_22_n_45, mul_90_22_n_46;
  wire mul_90_22_n_47, mul_90_22_n_48, mul_90_22_n_49, mul_90_22_n_50, mul_90_22_n_51, mul_90_22_n_52, mul_90_22_n_53, mul_90_22_n_54;
  wire mul_90_22_n_55, mul_90_22_n_56, mul_90_22_n_57, mul_90_22_n_58, mul_90_22_n_59, mul_90_22_n_60, mul_90_22_n_61, mul_90_22_n_62;
  wire mul_90_22_n_63, mul_90_22_n_64, mul_90_22_n_65, mul_90_22_n_66, mul_90_22_n_67, mul_90_22_n_68, mul_90_22_n_69, mul_90_22_n_70;
  wire mul_90_22_n_71, mul_90_22_n_72, mul_90_22_n_73, mul_90_22_n_74, mul_90_22_n_75, mul_90_22_n_76, mul_90_22_n_77, mul_90_22_n_78;
  wire mul_90_22_n_79, mul_90_22_n_80, mul_90_22_n_81, mul_90_22_n_82, mul_90_22_n_83, mul_90_22_n_84, mul_90_22_n_85, mul_90_22_n_86;
  wire mul_90_22_n_87, mul_90_22_n_88, mul_90_22_n_89, mul_90_22_n_90, mul_90_22_n_91, mul_90_22_n_92, mul_90_22_n_93, mul_90_22_n_94;
  wire mul_90_22_n_95, mul_90_22_n_96, mul_90_22_n_97, mul_90_22_n_98, mul_90_22_n_99, mul_90_22_n_100, mul_90_22_n_101, mul_90_22_n_102;
  wire mul_90_22_n_103, mul_90_22_n_104, mul_90_22_n_105, mul_90_22_n_106, mul_90_22_n_107, mul_90_22_n_108, mul_90_22_n_109, mul_90_22_n_110;
  wire mul_90_22_n_111, mul_90_22_n_112, mul_90_22_n_113, mul_90_22_n_114, mul_90_22_n_115, mul_90_22_n_116, mul_90_22_n_117, mul_90_22_n_118;
  wire mul_90_22_n_119, mul_90_22_n_120, mul_90_22_n_121, mul_90_22_n_122, mul_90_22_n_123, mul_90_22_n_124, mul_90_22_n_125, mul_90_22_n_126;
  wire mul_90_22_n_127, mul_90_22_n_128, mul_90_22_n_129, mul_90_22_n_130, mul_90_22_n_131, mul_90_22_n_132, mul_90_22_n_133, mul_90_22_n_134;
  wire mul_90_22_n_135, mul_90_22_n_136, mul_90_22_n_137, mul_90_22_n_138, mul_90_22_n_139, mul_90_22_n_140, mul_90_22_n_141, mul_90_22_n_142;
  wire mul_90_22_n_143, mul_90_22_n_144, mul_90_22_n_145, mul_90_22_n_146, mul_90_22_n_147, mul_90_22_n_148, mul_90_22_n_149, mul_90_22_n_150;
  wire mul_90_22_n_151, mul_90_22_n_152, mul_90_22_n_153, mul_90_22_n_154, mul_90_22_n_155, mul_90_22_n_156, mul_90_22_n_157, mul_90_22_n_158;
  wire mul_90_22_n_159, mul_90_22_n_160, mul_90_22_n_161, mul_90_22_n_162, mul_90_22_n_163, mul_90_22_n_164, mul_90_22_n_165, mul_90_22_n_166;
  wire mul_90_22_n_167, mul_90_22_n_168, mul_90_22_n_169, mul_90_22_n_170, mul_90_22_n_171, mul_90_22_n_172, mul_90_22_n_173, mul_90_22_n_174;
  wire mul_90_22_n_175, mul_90_22_n_176, mul_90_22_n_177, mul_90_22_n_178, mul_90_22_n_179, mul_90_22_n_180, mul_90_22_n_181, mul_90_22_n_182;
  wire mul_90_22_n_198, mul_90_22_n_199, mul_90_22_n_200, mul_90_22_n_201, mul_90_22_n_202, mul_90_22_n_203, mul_90_22_n_204, mul_90_22_n_205;
  wire mul_90_22_n_206, mul_90_22_n_207, mul_90_22_n_208, mul_90_22_n_209, mul_90_22_n_210, mul_90_22_n_211, mul_90_22_n_212, mul_90_22_n_213;
  wire mul_90_22_n_214, mul_90_22_n_215, mul_90_22_n_216, mul_90_22_n_217, mul_90_22_n_218, mul_90_22_n_219, mul_90_22_n_220, mul_90_22_n_221;
  wire mul_90_22_n_222, mul_90_22_n_223, mul_90_22_n_224, mul_90_22_n_225, mul_90_22_n_226, mul_90_22_n_227, mul_90_22_n_228, mul_90_22_n_229;
  wire mul_90_22_n_230, mul_90_22_n_231, mul_90_22_n_232, mul_90_22_n_233, mul_90_22_n_234, mul_90_22_n_235, mul_90_22_n_236, mul_90_22_n_237;
  wire mul_90_22_n_238, mul_90_22_n_239, mul_90_22_n_240, mul_90_22_n_241, mul_90_22_n_242, mul_90_22_n_243, mul_90_22_n_244, mul_90_22_n_245;
  wire mul_90_22_n_246, mul_90_22_n_247, mul_90_22_n_248, mul_90_22_n_249, mul_90_22_n_250, mul_90_22_n_251, mul_90_22_n_252, mul_90_22_n_253;
  wire mul_90_22_n_254, mul_90_22_n_255, mul_90_22_n_256, mul_90_22_n_257, mul_90_22_n_258, mul_90_22_n_259, mul_90_22_n_260, mul_90_22_n_261;
  wire mul_90_22_n_262, mul_90_22_n_263, mul_90_22_n_264, mul_90_22_n_265, mul_90_22_n_266, mul_90_22_n_267, mul_90_22_n_268, mul_90_22_n_269;
  wire mul_90_22_n_270, mul_90_22_n_271, mul_90_22_n_272, mul_90_22_n_273, mul_90_22_n_274, mul_90_22_n_275, mul_90_22_n_276, mul_90_22_n_277;
  wire mul_90_22_n_278, mul_90_22_n_279, mul_90_22_n_280, mul_90_22_n_281, mul_90_22_n_282, mul_90_22_n_283, mul_90_22_n_284, mul_90_22_n_285;
  wire mul_90_22_n_286, mul_90_22_n_287, mul_90_22_n_288, mul_90_22_n_289, mul_90_22_n_290, mul_90_22_n_291, mul_90_22_n_292, mul_90_22_n_293;
  wire mul_90_22_n_294, mul_90_22_n_295, mul_90_22_n_296, mul_90_22_n_297, mul_90_22_n_298, mul_90_22_n_299, mul_90_22_n_300, mul_90_22_n_301;
  wire mul_90_22_n_302, mul_90_22_n_303, mul_90_22_n_304, mul_90_22_n_305, mul_90_22_n_306, mul_90_22_n_307, mul_90_22_n_308, mul_90_22_n_310;
  wire mul_90_22_n_311, mul_90_22_n_312, mul_90_22_n_313, mul_90_22_n_314, mul_90_22_n_315, mul_90_22_n_316, mul_90_22_n_317, mul_90_22_n_318;
  wire mul_90_22_n_319, mul_90_22_n_320, mul_90_22_n_321, mul_90_22_n_322, mul_90_22_n_323, mul_90_22_n_324, mul_90_22_n_325, mul_90_22_n_326;
  wire mul_90_22_n_327, mul_90_22_n_328, mul_90_22_n_329, mul_90_22_n_330, mul_90_22_n_331, mul_90_22_n_332, mul_90_22_n_333, mul_90_22_n_334;
  wire mul_90_22_n_335, mul_90_22_n_336, mul_90_22_n_337, mul_90_22_n_338, mul_90_22_n_339, mul_90_22_n_340, mul_90_22_n_341, mul_90_22_n_342;
  wire mul_90_22_n_343, mul_90_22_n_344, mul_90_22_n_345, mul_90_22_n_346, mul_90_22_n_347, mul_90_22_n_348, mul_90_22_n_349, mul_90_22_n_350;
  wire mul_90_22_n_351, mul_90_22_n_352, mul_90_22_n_353, mul_90_22_n_354, mul_90_22_n_355, mul_90_22_n_356, mul_90_22_n_357, mul_90_22_n_358;
  wire mul_90_22_n_359, mul_90_22_n_360, mul_90_22_n_361, mul_90_22_n_362, mul_90_22_n_363, mul_90_22_n_364, mul_90_22_n_365, mul_90_22_n_366;
  wire mul_90_22_n_367, mul_90_22_n_368, mul_90_22_n_369, mul_90_22_n_370, mul_90_22_n_371, mul_90_22_n_372, mul_90_22_n_373, mul_90_22_n_374;
  wire mul_90_22_n_375, mul_90_22_n_376, mul_90_22_n_377, mul_90_22_n_378, mul_90_22_n_379, mul_90_22_n_380, mul_90_22_n_381, mul_90_22_n_382;
  wire mul_90_22_n_383, mul_90_22_n_384, mul_90_22_n_385, mul_90_22_n_386, mul_90_22_n_387, mul_90_22_n_388, mul_90_22_n_389, mul_90_22_n_390;
  wire mul_90_22_n_391, mul_90_22_n_392, mul_90_22_n_393, mul_90_22_n_394, mul_90_22_n_395, mul_90_22_n_396, mul_90_22_n_397, mul_90_22_n_398;
  wire mul_90_22_n_399, mul_90_22_n_400, mul_90_22_n_401, mul_90_22_n_402, mul_90_22_n_403, mul_90_22_n_404, mul_90_22_n_405, mul_90_22_n_406;
  wire mul_90_22_n_407, mul_90_22_n_408, mul_90_22_n_409, mul_90_22_n_410, mul_90_22_n_411, mul_90_22_n_412, mul_90_22_n_413, mul_90_22_n_414;
  wire mul_90_22_n_415, mul_90_22_n_416, mul_90_22_n_417, mul_90_22_n_418, mul_90_22_n_419, mul_90_22_n_420, mul_90_22_n_421, mul_90_22_n_422;
  wire mul_90_22_n_423, mul_90_22_n_424, mul_90_22_n_425, mul_90_22_n_426, mul_90_22_n_427, mul_90_22_n_428, mul_90_22_n_429, mul_90_22_n_430;
  wire mul_90_22_n_431, mul_90_22_n_432, mul_90_22_n_433, mul_90_22_n_434, mul_90_22_n_435, mul_90_22_n_436, mul_90_22_n_437, mul_90_22_n_438;
  wire mul_90_22_n_439, mul_90_22_n_440, mul_90_22_n_441, mul_90_22_n_442, mul_90_22_n_443, mul_90_22_n_444, mul_90_22_n_445, mul_90_22_n_446;
  wire mul_90_22_n_447, mul_90_22_n_448, mul_90_22_n_449, mul_90_22_n_450, mul_90_22_n_451, mul_90_22_n_452, mul_90_22_n_453, mul_90_22_n_454;
  wire mul_90_22_n_455, mul_90_22_n_456, mul_90_22_n_457, mul_90_22_n_458, mul_90_22_n_459, mul_90_22_n_460, mul_90_22_n_461, mul_90_22_n_462;
  wire mul_90_22_n_463, mul_90_22_n_464, mul_90_22_n_465, mul_90_22_n_466, mul_90_22_n_467, mul_90_22_n_468, mul_90_22_n_469, mul_90_22_n_470;
  wire mul_90_22_n_471, mul_90_22_n_472, mul_90_22_n_473, mul_90_22_n_474, mul_90_22_n_475, mul_90_22_n_476, mul_90_22_n_477, mul_90_22_n_478;
  wire mul_90_22_n_479, mul_90_22_n_480, mul_90_22_n_481, mul_90_22_n_482, mul_90_22_n_483, mul_90_22_n_484, mul_90_22_n_485, mul_90_22_n_486;
  wire mul_90_22_n_487, mul_90_22_n_488, mul_90_22_n_489, mul_90_22_n_490, mul_90_22_n_491, mul_90_22_n_492, mul_90_22_n_493, mul_90_22_n_494;
  wire mul_90_22_n_495, mul_90_22_n_496, mul_90_22_n_497, mul_90_22_n_498, mul_90_22_n_499, mul_90_22_n_500, mul_90_22_n_501, mul_90_22_n_502;
  wire mul_90_22_n_503, mul_90_22_n_504, mul_90_22_n_505, mul_90_22_n_506, mul_90_22_n_507, mul_90_22_n_508, mul_90_22_n_509, mul_90_22_n_510;
  wire mul_90_22_n_511, mul_90_22_n_512, mul_90_22_n_513, mul_90_22_n_514, mul_90_22_n_515, mul_90_22_n_516, mul_90_22_n_517, mul_90_22_n_518;
  wire mul_90_22_n_519, mul_90_22_n_520, mul_90_22_n_521, mul_90_22_n_522, mul_90_22_n_523, mul_90_22_n_524, mul_90_22_n_525, mul_90_22_n_526;
  wire mul_90_22_n_527, mul_90_22_n_528, mul_90_22_n_529, mul_90_22_n_530, mul_90_22_n_531, mul_90_22_n_532, mul_90_22_n_533, mul_90_22_n_534;
  wire mul_90_22_n_535, mul_90_22_n_536, mul_90_22_n_537, mul_90_22_n_538, mul_90_22_n_539, mul_90_22_n_540, mul_90_22_n_541, mul_90_22_n_542;
  wire mul_90_22_n_543, mul_90_22_n_544, mul_90_22_n_545, mul_90_22_n_546, mul_90_22_n_547, mul_90_22_n_548, mul_90_22_n_549, mul_90_22_n_550;
  wire mul_90_22_n_551, mul_90_22_n_552, mul_90_22_n_553, mul_90_22_n_554, mul_90_22_n_555, mul_90_22_n_556, mul_90_22_n_557, mul_90_22_n_558;
  wire mul_90_22_n_559, mul_90_22_n_560, mul_90_22_n_561, mul_90_22_n_562, mul_90_22_n_563, mul_90_22_n_564, mul_90_22_n_565, mul_90_22_n_566;
  wire mul_90_22_n_567, mul_90_22_n_568, mul_90_22_n_569, mul_90_22_n_570, mul_90_22_n_571, mul_90_22_n_572, mul_90_22_n_573, mul_90_22_n_574;
  wire mul_90_22_n_575, mul_90_22_n_576, mul_90_22_n_577, mul_90_22_n_578, mul_90_22_n_579, mul_90_22_n_580, mul_90_22_n_581, mul_90_22_n_582;
  wire mul_90_22_n_583, mul_90_22_n_584, mul_90_22_n_585, mul_90_22_n_586, mul_90_22_n_587, mul_90_22_n_588, mul_90_22_n_589, mul_90_22_n_590;
  wire mul_90_22_n_591, mul_90_22_n_592, mul_90_22_n_593, mul_90_22_n_594, mul_90_22_n_595, mul_90_22_n_596, mul_90_22_n_597, mul_90_22_n_598;
  wire mul_90_22_n_599, mul_90_22_n_600, mul_90_22_n_601, mul_90_22_n_602, mul_90_22_n_603, mul_90_22_n_604, mul_90_22_n_605, mul_90_22_n_606;
  wire mul_90_22_n_607, mul_90_22_n_608, mul_90_22_n_609, mul_90_22_n_610, mul_90_22_n_611, mul_90_22_n_612, mul_90_22_n_613, mul_90_22_n_614;
  wire mul_90_22_n_615, mul_90_22_n_616, mul_90_22_n_617, mul_90_22_n_618, mul_90_22_n_619, mul_90_22_n_620, mul_90_22_n_621, mul_90_22_n_622;
  wire mul_90_22_n_623, mul_90_22_n_624, mul_90_22_n_625, mul_90_22_n_626, mul_90_22_n_627, mul_90_22_n_628, mul_90_22_n_629, mul_90_22_n_630;
  wire mul_90_22_n_631, mul_90_22_n_632, mul_90_22_n_633, mul_90_22_n_634, mul_90_22_n_635, mul_90_22_n_636, mul_90_22_n_637, mul_90_22_n_638;
  wire mul_90_22_n_639, mul_90_22_n_640, mul_90_22_n_641, mul_90_22_n_642, mul_90_22_n_643, mul_90_22_n_644, mul_90_22_n_645, mul_90_22_n_646;
  wire mul_90_22_n_647, mul_90_22_n_648, mul_90_22_n_649, mul_90_22_n_650, mul_90_22_n_651, mul_90_22_n_652, mul_90_22_n_653, mul_90_22_n_654;
  wire mul_90_22_n_655, mul_90_22_n_656, mul_90_22_n_657, mul_90_22_n_658, mul_90_22_n_659, mul_90_22_n_660, mul_90_22_n_661, mul_90_22_n_662;
  wire mul_90_22_n_663, mul_90_22_n_664, mul_90_22_n_665, mul_90_22_n_666, mul_90_22_n_667, mul_90_22_n_668, mul_90_22_n_669, mul_90_22_n_670;
  wire mul_90_22_n_671, mul_90_22_n_672, mul_90_22_n_673, mul_90_22_n_674, mul_90_22_n_675, mul_90_22_n_676, mul_90_22_n_677, mul_90_22_n_678;
  wire mul_90_22_n_679, mul_90_22_n_680, mul_90_22_n_681, mul_90_22_n_682, mul_90_22_n_683, mul_90_22_n_684, mul_90_22_n_685, mul_90_22_n_686;
  wire mul_90_22_n_687, mul_90_22_n_688, mul_90_22_n_689, mul_90_22_n_690, mul_90_22_n_691, mul_90_22_n_692, mul_90_22_n_693, mul_90_22_n_694;
  wire mul_90_22_n_695, mul_90_22_n_696, mul_90_22_n_697, mul_90_22_n_698, mul_90_22_n_699, mul_90_22_n_700, mul_90_22_n_701, mul_90_22_n_702;
  wire mul_90_22_n_703, mul_90_22_n_704, mul_90_22_n_705, mul_90_22_n_706, mul_90_22_n_707, mul_90_22_n_708, mul_90_22_n_709, mul_90_22_n_710;
  wire mul_90_22_n_711, mul_90_22_n_712, mul_90_22_n_713, mul_90_22_n_714, mul_90_22_n_715, mul_90_22_n_716, mul_90_22_n_717, mul_90_22_n_718;
  wire mul_90_22_n_719, mul_90_22_n_720, mul_90_22_n_721, mul_90_22_n_722, mul_90_22_n_723, mul_90_22_n_724, mul_90_22_n_725, mul_90_22_n_726;
  wire mul_90_22_n_727, mul_90_22_n_728, mul_90_22_n_729, mul_90_22_n_730, mul_90_22_n_731, mul_90_22_n_732, mul_90_22_n_733, mul_90_22_n_734;
  wire mul_90_22_n_735, mul_90_22_n_736, mul_90_22_n_737, mul_90_22_n_738, mul_90_22_n_739, mul_90_22_n_740, mul_90_22_n_741, mul_90_22_n_742;
  wire mul_90_22_n_743, mul_90_22_n_744, mul_90_22_n_745, mul_90_22_n_746, mul_90_22_n_747, mul_90_22_n_748, mul_90_22_n_749, mul_90_22_n_750;
  wire mul_90_22_n_751, mul_90_22_n_752, mul_90_22_n_753, mul_90_22_n_754, mul_90_22_n_755, mul_90_22_n_756, mul_90_22_n_757, mul_90_22_n_758;
  wire mul_90_22_n_759, mul_90_22_n_760, mul_90_22_n_761, mul_90_22_n_762, mul_90_22_n_763, mul_90_22_n_764, mul_90_22_n_765, mul_90_22_n_766;
  wire mul_90_22_n_767, mul_90_22_n_768, mul_90_22_n_769, mul_90_22_n_770, mul_90_22_n_771, mul_90_22_n_772, mul_90_22_n_773, mul_90_22_n_774;
  wire mul_90_22_n_775, mul_90_22_n_776, mul_90_22_n_777, mul_90_22_n_778, mul_90_22_n_779, mul_90_22_n_780, mul_90_22_n_781, mul_90_22_n_782;
  wire mul_90_22_n_783, mul_90_22_n_784, mul_90_22_n_785, mul_90_22_n_786, mul_90_22_n_787, mul_90_22_n_788, mul_90_22_n_789, mul_90_22_n_790;
  wire mul_90_22_n_791, mul_90_22_n_792, mul_90_22_n_793, mul_90_22_n_794, mul_90_22_n_795, mul_90_22_n_796, mul_90_22_n_797, mul_90_22_n_798;
  wire mul_90_22_n_799, mul_90_22_n_800, mul_90_22_n_801, mul_90_22_n_802, mul_90_22_n_803, mul_90_22_n_804, mul_90_22_n_805, mul_90_22_n_806;
  wire mul_90_22_n_807, mul_90_22_n_808, mul_90_22_n_809, mul_90_22_n_810, mul_90_22_n_811, mul_90_22_n_812, mul_90_22_n_813, mul_90_22_n_814;
  wire mul_90_22_n_815, mul_90_22_n_816, mul_90_22_n_817, mul_90_22_n_818, mul_90_22_n_819, mul_90_22_n_820, mul_90_22_n_821, mul_90_22_n_822;
  wire mul_90_22_n_823, mul_90_22_n_824, mul_90_22_n_825, mul_90_22_n_826, mul_90_22_n_827, mul_90_22_n_828, mul_90_22_n_829, mul_90_22_n_830;
  wire mul_90_22_n_831, mul_90_22_n_832, mul_90_22_n_833, mul_90_22_n_834, mul_90_22_n_835, mul_90_22_n_836, mul_90_22_n_837, mul_90_22_n_838;
  wire mul_90_22_n_839, mul_90_22_n_840, mul_90_22_n_841, mul_90_22_n_842, mul_90_22_n_843, mul_90_22_n_844, mul_90_22_n_845, mul_90_22_n_846;
  wire mul_90_22_n_847, mul_90_22_n_848, mul_90_22_n_849, mul_90_22_n_850, mul_90_22_n_851, mul_90_22_n_852, mul_90_22_n_853, mul_90_22_n_854;
  wire mul_90_22_n_855, mul_90_22_n_856, mul_90_22_n_857, mul_90_22_n_858, mul_90_22_n_859, mul_90_22_n_860, mul_90_22_n_861, mul_90_22_n_862;
  wire mul_90_22_n_863, mul_90_22_n_864, mul_90_22_n_865, mul_90_22_n_866, mul_90_22_n_867, mul_90_22_n_868, mul_90_22_n_869, mul_90_22_n_870;
  wire mul_90_22_n_871, mul_90_22_n_872, mul_90_22_n_873, mul_90_22_n_874, mul_90_22_n_875, mul_90_22_n_876, mul_90_22_n_877, mul_90_22_n_878;
  wire mul_90_22_n_879, mul_90_22_n_880, mul_90_22_n_881, mul_90_22_n_882, mul_90_22_n_883, mul_90_22_n_884, mul_90_22_n_885, mul_90_22_n_886;
  wire mul_90_22_n_887, mul_90_22_n_888, mul_90_22_n_889, mul_90_22_n_890, mul_90_22_n_891, mul_90_22_n_892, mul_90_22_n_893, mul_90_22_n_894;
  wire mul_90_22_n_895, mul_90_22_n_896, mul_90_22_n_897, mul_90_22_n_898, mul_90_22_n_899, mul_90_22_n_900, mul_90_22_n_901, mul_90_22_n_902;
  wire mul_90_22_n_903, mul_90_22_n_904, mul_90_22_n_905, mul_90_22_n_906, mul_90_22_n_907, mul_90_22_n_908, mul_90_22_n_909, mul_90_22_n_910;
  wire mul_90_22_n_911, mul_90_22_n_912, mul_90_22_n_913, mul_90_22_n_914, mul_90_22_n_915, mul_90_22_n_916, mul_90_22_n_917, mul_90_22_n_918;
  wire mul_90_22_n_919, mul_90_22_n_920, mul_90_22_n_921, mul_90_22_n_922, mul_90_22_n_923, mul_90_22_n_924, mul_90_22_n_925, mul_90_22_n_926;
  wire mul_90_22_n_927, mul_90_22_n_928, mul_90_22_n_929, mul_90_22_n_930, mul_90_22_n_931, mul_90_22_n_932, mul_90_22_n_933, mul_90_22_n_934;
  wire mul_90_22_n_935, mul_90_22_n_936, mul_90_22_n_937, mul_90_22_n_938, mul_90_22_n_939, mul_90_22_n_940, mul_90_22_n_941, mul_90_22_n_942;
  wire mul_90_22_n_943, mul_90_22_n_944, mul_90_22_n_945, mul_90_22_n_946, mul_90_22_n_947, mul_90_22_n_948, mul_90_22_n_949, mul_90_22_n_950;
  wire mul_90_22_n_951, mul_90_22_n_952, mul_90_22_n_953, mul_90_22_n_954, mul_90_22_n_955, mul_90_22_n_956, mul_90_22_n_957, mul_90_22_n_958;
  wire mul_90_22_n_959, mul_90_22_n_960, mul_90_22_n_961, mul_90_22_n_962, mul_90_22_n_963, mul_90_22_n_964, mul_90_22_n_965, mul_90_22_n_966;
  wire mul_90_22_n_967, mul_90_22_n_968, mul_90_22_n_969, mul_90_22_n_970, mul_90_22_n_971, mul_90_22_n_972, mul_90_22_n_973, mul_90_22_n_974;
  wire mul_90_22_n_975, mul_90_22_n_976, mul_90_22_n_977, mul_90_22_n_978, mul_90_22_n_979, mul_90_22_n_980, mul_90_22_n_981, mul_90_22_n_982;
  wire mul_90_22_n_983, mul_90_22_n_984, mul_90_22_n_985, mul_90_22_n_986, mul_90_22_n_987, mul_90_22_n_988, mul_90_22_n_989, mul_90_22_n_990;
  wire mul_90_22_n_991, mul_90_22_n_992, mul_90_22_n_993, mul_90_22_n_994, mul_90_22_n_995, mul_90_22_n_996, mul_90_22_n_997, mul_90_22_n_998;
  wire mul_90_22_n_999, mul_90_22_n_1000, mul_90_22_n_1001, mul_90_22_n_1002, mul_90_22_n_1003, mul_90_22_n_1004, mul_90_22_n_1005, mul_90_22_n_1006;
  wire mul_90_22_n_1007, mul_90_22_n_1008, mul_90_22_n_1009, mul_90_22_n_1010, mul_90_22_n_1011, mul_90_22_n_1012, mul_90_22_n_1013, mul_90_22_n_1014;
  wire mul_90_22_n_1015, mul_90_22_n_1016, mul_90_22_n_1017, mul_90_22_n_1018, mul_90_22_n_1019, mul_90_22_n_1020, mul_90_22_n_1021, mul_90_22_n_1022;
  wire mul_90_22_n_1023, mul_90_22_n_1024, mul_90_22_n_1025, mul_90_22_n_1026, mul_90_22_n_1027, mul_90_22_n_1028, mul_90_22_n_1029, mul_90_22_n_1030;
  wire mul_90_22_n_1031, mul_90_22_n_1032, mul_90_22_n_1033, mul_90_22_n_1034, mul_90_22_n_1035, mul_90_22_n_1036, mul_90_22_n_1037, mul_90_22_n_1038;
  wire mul_90_22_n_1039, mul_90_22_n_1040, mul_90_22_n_1041, mul_90_22_n_1042, mul_90_22_n_1043, mul_90_22_n_1044, mul_90_22_n_1045, mul_90_22_n_1046;
  wire mul_90_22_n_1047, mul_90_22_n_1048, mul_90_22_n_1049, mul_90_22_n_1050, mul_90_22_n_1051, mul_90_22_n_1052, mul_90_22_n_1053, mul_90_22_n_1054;
  wire mul_90_22_n_1055, mul_90_22_n_1056, mul_90_22_n_1057, mul_90_22_n_1058, mul_90_22_n_1059, mul_90_22_n_1060, mul_90_22_n_1061, mul_90_22_n_1062;
  wire mul_90_22_n_1063, mul_90_22_n_1064, mul_90_22_n_1065, mul_90_22_n_1066, mul_90_22_n_1067, mul_90_22_n_1068, mul_90_22_n_1069, mul_90_22_n_1070;
  wire mul_90_22_n_1071, mul_90_22_n_1072, mul_90_22_n_1073, mul_90_22_n_1074, mul_90_22_n_1075, mul_90_22_n_1076, mul_90_22_n_1077, mul_90_22_n_1078;
  wire mul_90_22_n_1079, mul_90_22_n_1080, mul_90_22_n_1081, mul_90_22_n_1082, mul_90_22_n_1083, mul_90_22_n_1084, mul_90_22_n_1085, mul_90_22_n_1086;
  wire mul_90_22_n_1087, mul_90_22_n_1088, mul_90_22_n_1089, mul_90_22_n_1090, mul_90_22_n_1091, mul_90_22_n_1092, mul_90_22_n_1093, mul_90_22_n_1094;
  wire mul_90_22_n_1095, mul_90_22_n_1096, mul_90_22_n_1097, mul_90_22_n_1098, mul_90_22_n_1099, mul_90_22_n_1100, mul_90_22_n_1101, mul_90_22_n_1102;
  wire mul_90_22_n_1103, mul_90_22_n_1104, mul_90_22_n_1105, mul_90_22_n_1106, mul_90_22_n_1107, mul_90_22_n_1108, mul_90_22_n_1109, mul_90_22_n_1110;
  wire mul_90_22_n_1111, mul_90_22_n_1112, mul_90_22_n_1113, mul_90_22_n_1114, mul_90_22_n_1115, mul_90_22_n_1116, mul_90_22_n_1117, mul_90_22_n_1118;
  wire mul_90_22_n_1119, mul_90_22_n_1120, mul_90_22_n_1121, mul_90_22_n_1122, mul_90_22_n_1123, mul_90_22_n_1124, mul_90_22_n_1125, mul_90_22_n_1126;
  wire mul_90_22_n_1127, mul_90_22_n_1128, mul_90_22_n_1129, mul_90_22_n_1130, mul_90_22_n_1131, mul_90_22_n_1132, mul_90_22_n_1133, mul_90_22_n_1134;
  wire mul_90_22_n_1135, mul_90_22_n_1136, mul_90_22_n_1137, mul_90_22_n_1138, mul_90_22_n_1139, mul_90_22_n_1140, mul_90_22_n_1141, mul_90_22_n_1142;
  wire mul_90_22_n_1143, mul_90_22_n_1144, mul_90_22_n_1145, mul_90_22_n_1146, mul_90_22_n_1147, mul_90_22_n_1148, mul_90_22_n_1149, mul_90_22_n_1150;
  wire mul_90_22_n_1151, mul_90_22_n_1152, mul_90_22_n_1153, mul_90_22_n_1154, mul_90_22_n_1155, mul_90_22_n_1156, mul_90_22_n_1157, mul_102_22_n_0;
  wire mul_102_22_n_1, mul_102_22_n_2, mul_102_22_n_3, mul_102_22_n_4, mul_102_22_n_5, mul_102_22_n_6, mul_102_22_n_7, mul_102_22_n_8;
  wire mul_102_22_n_9, mul_102_22_n_10, mul_102_22_n_11, mul_102_22_n_12, mul_102_22_n_13, mul_102_22_n_14, mul_102_22_n_15, mul_102_22_n_16;
  wire mul_102_22_n_17, mul_102_22_n_18, mul_102_22_n_19, mul_102_22_n_20, mul_102_22_n_21, mul_102_22_n_22, mul_102_22_n_23, mul_102_22_n_24;
  wire mul_102_22_n_25, mul_102_22_n_26, mul_102_22_n_27, mul_102_22_n_28, mul_102_22_n_29, mul_102_22_n_30, mul_102_22_n_31, mul_102_22_n_32;
  wire mul_102_22_n_33, mul_102_22_n_34, mul_102_22_n_35, mul_102_22_n_36, mul_102_22_n_37, mul_102_22_n_38, mul_102_22_n_39, mul_102_22_n_40;
  wire mul_102_22_n_41, mul_102_22_n_42, mul_102_22_n_43, mul_102_22_n_44, mul_102_22_n_45, mul_102_22_n_46, mul_102_22_n_47, mul_102_22_n_48;
  wire mul_102_22_n_49, mul_102_22_n_50, mul_102_22_n_51, mul_102_22_n_52, mul_102_22_n_53, mul_102_22_n_54, mul_102_22_n_55, mul_102_22_n_56;
  wire mul_102_22_n_57, mul_102_22_n_58, mul_102_22_n_59, mul_102_22_n_60, mul_102_22_n_61, mul_102_22_n_62, mul_102_22_n_63, mul_102_22_n_64;
  wire mul_102_22_n_65, mul_102_22_n_66, mul_102_22_n_67, mul_102_22_n_68, mul_102_22_n_69, mul_102_22_n_70, mul_102_22_n_71, mul_102_22_n_72;
  wire mul_102_22_n_73, mul_102_22_n_74, mul_102_22_n_75, mul_102_22_n_76, mul_102_22_n_77, mul_102_22_n_78, mul_102_22_n_79, mul_102_22_n_80;
  wire mul_102_22_n_81, mul_102_22_n_82, mul_102_22_n_83, mul_102_22_n_84, mul_102_22_n_85, mul_102_22_n_86, mul_102_22_n_87, mul_102_22_n_88;
  wire mul_102_22_n_89, mul_102_22_n_90, mul_102_22_n_91, mul_102_22_n_92, mul_102_22_n_93, mul_102_22_n_94, mul_102_22_n_95, mul_102_22_n_96;
  wire mul_102_22_n_97, mul_102_22_n_98, mul_102_22_n_99, mul_102_22_n_100, mul_102_22_n_101, mul_102_22_n_102, mul_102_22_n_103, mul_102_22_n_104;
  wire mul_102_22_n_105, mul_102_22_n_106, mul_102_22_n_107, mul_102_22_n_108, mul_102_22_n_109, mul_102_22_n_110, mul_102_22_n_111, mul_102_22_n_112;
  wire mul_102_22_n_113, mul_102_22_n_114, mul_102_22_n_115, mul_102_22_n_116, mul_102_22_n_117, mul_102_22_n_118, mul_102_22_n_119, mul_102_22_n_120;
  wire mul_102_22_n_121, mul_102_22_n_122, mul_102_22_n_123, mul_102_22_n_124, mul_102_22_n_125, mul_102_22_n_126, mul_102_22_n_127, mul_102_22_n_128;
  wire mul_102_22_n_129, mul_102_22_n_130, mul_102_22_n_131, mul_102_22_n_132, mul_102_22_n_133, mul_102_22_n_134, mul_102_22_n_135, mul_102_22_n_136;
  wire mul_102_22_n_137, mul_102_22_n_138, mul_102_22_n_139, mul_102_22_n_140, mul_102_22_n_141, mul_102_22_n_142, mul_102_22_n_143, mul_102_22_n_144;
  wire mul_102_22_n_145, mul_102_22_n_146, mul_102_22_n_147, mul_102_22_n_148, mul_102_22_n_149, mul_102_22_n_150, mul_102_22_n_151, mul_102_22_n_152;
  wire mul_102_22_n_153, mul_102_22_n_154, mul_102_22_n_155, mul_102_22_n_156, mul_102_22_n_157, mul_102_22_n_158, mul_102_22_n_159, mul_102_22_n_160;
  wire mul_102_22_n_161, mul_102_22_n_162, mul_102_22_n_163, mul_102_22_n_164, mul_102_22_n_165, mul_102_22_n_166, mul_102_22_n_167, mul_102_22_n_168;
  wire mul_102_22_n_169, mul_102_22_n_170, mul_102_22_n_171, mul_102_22_n_172, mul_102_22_n_173, mul_102_22_n_174, mul_102_22_n_175, mul_102_22_n_176;
  wire mul_102_22_n_177, mul_102_22_n_178, mul_102_22_n_179, mul_102_22_n_180, mul_102_22_n_181, mul_102_22_n_182, mul_102_22_n_198, mul_102_22_n_199;
  wire mul_102_22_n_200, mul_102_22_n_201, mul_102_22_n_202, mul_102_22_n_203, mul_102_22_n_204, mul_102_22_n_205, mul_102_22_n_206, mul_102_22_n_207;
  wire mul_102_22_n_208, mul_102_22_n_209, mul_102_22_n_210, mul_102_22_n_211, mul_102_22_n_212, mul_102_22_n_213, mul_102_22_n_214, mul_102_22_n_215;
  wire mul_102_22_n_216, mul_102_22_n_217, mul_102_22_n_218, mul_102_22_n_219, mul_102_22_n_220, mul_102_22_n_221, mul_102_22_n_222, mul_102_22_n_223;
  wire mul_102_22_n_224, mul_102_22_n_225, mul_102_22_n_226, mul_102_22_n_227, mul_102_22_n_228, mul_102_22_n_229, mul_102_22_n_230, mul_102_22_n_231;
  wire mul_102_22_n_232, mul_102_22_n_233, mul_102_22_n_234, mul_102_22_n_235, mul_102_22_n_236, mul_102_22_n_237, mul_102_22_n_238, mul_102_22_n_239;
  wire mul_102_22_n_240, mul_102_22_n_241, mul_102_22_n_242, mul_102_22_n_243, mul_102_22_n_244, mul_102_22_n_245, mul_102_22_n_246, mul_102_22_n_247;
  wire mul_102_22_n_248, mul_102_22_n_249, mul_102_22_n_250, mul_102_22_n_251, mul_102_22_n_252, mul_102_22_n_253, mul_102_22_n_254, mul_102_22_n_255;
  wire mul_102_22_n_256, mul_102_22_n_257, mul_102_22_n_258, mul_102_22_n_259, mul_102_22_n_260, mul_102_22_n_261, mul_102_22_n_262, mul_102_22_n_263;
  wire mul_102_22_n_264, mul_102_22_n_265, mul_102_22_n_266, mul_102_22_n_267, mul_102_22_n_268, mul_102_22_n_269, mul_102_22_n_270, mul_102_22_n_271;
  wire mul_102_22_n_272, mul_102_22_n_273, mul_102_22_n_274, mul_102_22_n_275, mul_102_22_n_276, mul_102_22_n_277, mul_102_22_n_278, mul_102_22_n_279;
  wire mul_102_22_n_280, mul_102_22_n_281, mul_102_22_n_282, mul_102_22_n_283, mul_102_22_n_284, mul_102_22_n_285, mul_102_22_n_286, mul_102_22_n_287;
  wire mul_102_22_n_288, mul_102_22_n_289, mul_102_22_n_290, mul_102_22_n_291, mul_102_22_n_292, mul_102_22_n_293, mul_102_22_n_294, mul_102_22_n_295;
  wire mul_102_22_n_296, mul_102_22_n_297, mul_102_22_n_298, mul_102_22_n_299, mul_102_22_n_300, mul_102_22_n_301, mul_102_22_n_302, mul_102_22_n_303;
  wire mul_102_22_n_304, mul_102_22_n_305, mul_102_22_n_306, mul_102_22_n_307, mul_102_22_n_308, mul_102_22_n_310, mul_102_22_n_311, mul_102_22_n_312;
  wire mul_102_22_n_313, mul_102_22_n_314, mul_102_22_n_315, mul_102_22_n_316, mul_102_22_n_317, mul_102_22_n_318, mul_102_22_n_319, mul_102_22_n_320;
  wire mul_102_22_n_321, mul_102_22_n_322, mul_102_22_n_323, mul_102_22_n_324, mul_102_22_n_325, mul_102_22_n_326, mul_102_22_n_327, mul_102_22_n_328;
  wire mul_102_22_n_329, mul_102_22_n_330, mul_102_22_n_331, mul_102_22_n_332, mul_102_22_n_333, mul_102_22_n_334, mul_102_22_n_335, mul_102_22_n_336;
  wire mul_102_22_n_337, mul_102_22_n_338, mul_102_22_n_339, mul_102_22_n_340, mul_102_22_n_341, mul_102_22_n_342, mul_102_22_n_343, mul_102_22_n_344;
  wire mul_102_22_n_345, mul_102_22_n_346, mul_102_22_n_347, mul_102_22_n_348, mul_102_22_n_349, mul_102_22_n_350, mul_102_22_n_351, mul_102_22_n_352;
  wire mul_102_22_n_353, mul_102_22_n_354, mul_102_22_n_355, mul_102_22_n_356, mul_102_22_n_357, mul_102_22_n_358, mul_102_22_n_359, mul_102_22_n_360;
  wire mul_102_22_n_361, mul_102_22_n_362, mul_102_22_n_363, mul_102_22_n_364, mul_102_22_n_365, mul_102_22_n_366, mul_102_22_n_367, mul_102_22_n_368;
  wire mul_102_22_n_369, mul_102_22_n_370, mul_102_22_n_371, mul_102_22_n_372, mul_102_22_n_373, mul_102_22_n_374, mul_102_22_n_375, mul_102_22_n_376;
  wire mul_102_22_n_377, mul_102_22_n_378, mul_102_22_n_379, mul_102_22_n_380, mul_102_22_n_381, mul_102_22_n_382, mul_102_22_n_383, mul_102_22_n_384;
  wire mul_102_22_n_385, mul_102_22_n_386, mul_102_22_n_387, mul_102_22_n_388, mul_102_22_n_389, mul_102_22_n_390, mul_102_22_n_391, mul_102_22_n_392;
  wire mul_102_22_n_393, mul_102_22_n_394, mul_102_22_n_395, mul_102_22_n_396, mul_102_22_n_397, mul_102_22_n_398, mul_102_22_n_399, mul_102_22_n_400;
  wire mul_102_22_n_401, mul_102_22_n_402, mul_102_22_n_403, mul_102_22_n_404, mul_102_22_n_405, mul_102_22_n_406, mul_102_22_n_407, mul_102_22_n_408;
  wire mul_102_22_n_409, mul_102_22_n_410, mul_102_22_n_411, mul_102_22_n_412, mul_102_22_n_413, mul_102_22_n_414, mul_102_22_n_415, mul_102_22_n_416;
  wire mul_102_22_n_417, mul_102_22_n_418, mul_102_22_n_419, mul_102_22_n_420, mul_102_22_n_421, mul_102_22_n_422, mul_102_22_n_423, mul_102_22_n_424;
  wire mul_102_22_n_425, mul_102_22_n_426, mul_102_22_n_427, mul_102_22_n_428, mul_102_22_n_429, mul_102_22_n_430, mul_102_22_n_431, mul_102_22_n_432;
  wire mul_102_22_n_433, mul_102_22_n_434, mul_102_22_n_435, mul_102_22_n_436, mul_102_22_n_437, mul_102_22_n_438, mul_102_22_n_439, mul_102_22_n_440;
  wire mul_102_22_n_441, mul_102_22_n_442, mul_102_22_n_443, mul_102_22_n_444, mul_102_22_n_445, mul_102_22_n_446, mul_102_22_n_447, mul_102_22_n_448;
  wire mul_102_22_n_449, mul_102_22_n_450, mul_102_22_n_451, mul_102_22_n_452, mul_102_22_n_453, mul_102_22_n_454, mul_102_22_n_455, mul_102_22_n_456;
  wire mul_102_22_n_457, mul_102_22_n_458, mul_102_22_n_459, mul_102_22_n_460, mul_102_22_n_461, mul_102_22_n_462, mul_102_22_n_463, mul_102_22_n_464;
  wire mul_102_22_n_465, mul_102_22_n_466, mul_102_22_n_467, mul_102_22_n_468, mul_102_22_n_469, mul_102_22_n_470, mul_102_22_n_471, mul_102_22_n_472;
  wire mul_102_22_n_473, mul_102_22_n_474, mul_102_22_n_475, mul_102_22_n_476, mul_102_22_n_477, mul_102_22_n_478, mul_102_22_n_479, mul_102_22_n_480;
  wire mul_102_22_n_481, mul_102_22_n_482, mul_102_22_n_483, mul_102_22_n_484, mul_102_22_n_485, mul_102_22_n_486, mul_102_22_n_487, mul_102_22_n_488;
  wire mul_102_22_n_489, mul_102_22_n_490, mul_102_22_n_491, mul_102_22_n_492, mul_102_22_n_493, mul_102_22_n_494, mul_102_22_n_495, mul_102_22_n_496;
  wire mul_102_22_n_497, mul_102_22_n_498, mul_102_22_n_499, mul_102_22_n_500, mul_102_22_n_501, mul_102_22_n_502, mul_102_22_n_503, mul_102_22_n_504;
  wire mul_102_22_n_505, mul_102_22_n_506, mul_102_22_n_507, mul_102_22_n_508, mul_102_22_n_509, mul_102_22_n_510, mul_102_22_n_511, mul_102_22_n_512;
  wire mul_102_22_n_513, mul_102_22_n_514, mul_102_22_n_515, mul_102_22_n_516, mul_102_22_n_517, mul_102_22_n_518, mul_102_22_n_519, mul_102_22_n_520;
  wire mul_102_22_n_521, mul_102_22_n_522, mul_102_22_n_523, mul_102_22_n_524, mul_102_22_n_525, mul_102_22_n_526, mul_102_22_n_527, mul_102_22_n_528;
  wire mul_102_22_n_529, mul_102_22_n_530, mul_102_22_n_531, mul_102_22_n_532, mul_102_22_n_533, mul_102_22_n_534, mul_102_22_n_535, mul_102_22_n_536;
  wire mul_102_22_n_537, mul_102_22_n_538, mul_102_22_n_539, mul_102_22_n_540, mul_102_22_n_541, mul_102_22_n_542, mul_102_22_n_543, mul_102_22_n_544;
  wire mul_102_22_n_545, mul_102_22_n_546, mul_102_22_n_547, mul_102_22_n_548, mul_102_22_n_549, mul_102_22_n_550, mul_102_22_n_551, mul_102_22_n_552;
  wire mul_102_22_n_553, mul_102_22_n_554, mul_102_22_n_555, mul_102_22_n_556, mul_102_22_n_557, mul_102_22_n_558, mul_102_22_n_559, mul_102_22_n_560;
  wire mul_102_22_n_561, mul_102_22_n_562, mul_102_22_n_563, mul_102_22_n_564, mul_102_22_n_565, mul_102_22_n_566, mul_102_22_n_567, mul_102_22_n_568;
  wire mul_102_22_n_569, mul_102_22_n_570, mul_102_22_n_571, mul_102_22_n_572, mul_102_22_n_573, mul_102_22_n_574, mul_102_22_n_575, mul_102_22_n_576;
  wire mul_102_22_n_577, mul_102_22_n_578, mul_102_22_n_579, mul_102_22_n_580, mul_102_22_n_581, mul_102_22_n_582, mul_102_22_n_583, mul_102_22_n_584;
  wire mul_102_22_n_585, mul_102_22_n_586, mul_102_22_n_587, mul_102_22_n_588, mul_102_22_n_589, mul_102_22_n_590, mul_102_22_n_591, mul_102_22_n_592;
  wire mul_102_22_n_593, mul_102_22_n_594, mul_102_22_n_595, mul_102_22_n_596, mul_102_22_n_597, mul_102_22_n_598, mul_102_22_n_599, mul_102_22_n_600;
  wire mul_102_22_n_601, mul_102_22_n_602, mul_102_22_n_603, mul_102_22_n_604, mul_102_22_n_605, mul_102_22_n_606, mul_102_22_n_607, mul_102_22_n_608;
  wire mul_102_22_n_609, mul_102_22_n_610, mul_102_22_n_611, mul_102_22_n_612, mul_102_22_n_613, mul_102_22_n_614, mul_102_22_n_615, mul_102_22_n_616;
  wire mul_102_22_n_617, mul_102_22_n_618, mul_102_22_n_619, mul_102_22_n_620, mul_102_22_n_621, mul_102_22_n_622, mul_102_22_n_623, mul_102_22_n_624;
  wire mul_102_22_n_625, mul_102_22_n_626, mul_102_22_n_627, mul_102_22_n_628, mul_102_22_n_629, mul_102_22_n_630, mul_102_22_n_631, mul_102_22_n_632;
  wire mul_102_22_n_633, mul_102_22_n_634, mul_102_22_n_635, mul_102_22_n_636, mul_102_22_n_637, mul_102_22_n_638, mul_102_22_n_639, mul_102_22_n_640;
  wire mul_102_22_n_641, mul_102_22_n_642, mul_102_22_n_643, mul_102_22_n_644, mul_102_22_n_645, mul_102_22_n_646, mul_102_22_n_647, mul_102_22_n_648;
  wire mul_102_22_n_649, mul_102_22_n_650, mul_102_22_n_651, mul_102_22_n_652, mul_102_22_n_653, mul_102_22_n_654, mul_102_22_n_655, mul_102_22_n_656;
  wire mul_102_22_n_657, mul_102_22_n_658, mul_102_22_n_659, mul_102_22_n_660, mul_102_22_n_661, mul_102_22_n_662, mul_102_22_n_663, mul_102_22_n_664;
  wire mul_102_22_n_665, mul_102_22_n_666, mul_102_22_n_667, mul_102_22_n_668, mul_102_22_n_669, mul_102_22_n_670, mul_102_22_n_671, mul_102_22_n_672;
  wire mul_102_22_n_673, mul_102_22_n_674, mul_102_22_n_675, mul_102_22_n_676, mul_102_22_n_677, mul_102_22_n_678, mul_102_22_n_679, mul_102_22_n_680;
  wire mul_102_22_n_681, mul_102_22_n_682, mul_102_22_n_683, mul_102_22_n_684, mul_102_22_n_685, mul_102_22_n_686, mul_102_22_n_687, mul_102_22_n_688;
  wire mul_102_22_n_689, mul_102_22_n_690, mul_102_22_n_691, mul_102_22_n_692, mul_102_22_n_693, mul_102_22_n_694, mul_102_22_n_695, mul_102_22_n_696;
  wire mul_102_22_n_697, mul_102_22_n_698, mul_102_22_n_699, mul_102_22_n_700, mul_102_22_n_701, mul_102_22_n_702, mul_102_22_n_703, mul_102_22_n_704;
  wire mul_102_22_n_705, mul_102_22_n_706, mul_102_22_n_707, mul_102_22_n_708, mul_102_22_n_709, mul_102_22_n_710, mul_102_22_n_711, mul_102_22_n_712;
  wire mul_102_22_n_713, mul_102_22_n_714, mul_102_22_n_715, mul_102_22_n_716, mul_102_22_n_717, mul_102_22_n_718, mul_102_22_n_719, mul_102_22_n_720;
  wire mul_102_22_n_721, mul_102_22_n_722, mul_102_22_n_723, mul_102_22_n_724, mul_102_22_n_725, mul_102_22_n_726, mul_102_22_n_727, mul_102_22_n_728;
  wire mul_102_22_n_729, mul_102_22_n_730, mul_102_22_n_731, mul_102_22_n_732, mul_102_22_n_733, mul_102_22_n_734, mul_102_22_n_735, mul_102_22_n_736;
  wire mul_102_22_n_737, mul_102_22_n_738, mul_102_22_n_739, mul_102_22_n_740, mul_102_22_n_741, mul_102_22_n_742, mul_102_22_n_743, mul_102_22_n_744;
  wire mul_102_22_n_745, mul_102_22_n_746, mul_102_22_n_747, mul_102_22_n_748, mul_102_22_n_749, mul_102_22_n_750, mul_102_22_n_751, mul_102_22_n_752;
  wire mul_102_22_n_753, mul_102_22_n_754, mul_102_22_n_755, mul_102_22_n_756, mul_102_22_n_757, mul_102_22_n_758, mul_102_22_n_759, mul_102_22_n_760;
  wire mul_102_22_n_761, mul_102_22_n_762, mul_102_22_n_763, mul_102_22_n_764, mul_102_22_n_765, mul_102_22_n_766, mul_102_22_n_767, mul_102_22_n_768;
  wire mul_102_22_n_769, mul_102_22_n_770, mul_102_22_n_771, mul_102_22_n_772, mul_102_22_n_773, mul_102_22_n_774, mul_102_22_n_775, mul_102_22_n_776;
  wire mul_102_22_n_777, mul_102_22_n_778, mul_102_22_n_779, mul_102_22_n_780, mul_102_22_n_781, mul_102_22_n_782, mul_102_22_n_783, mul_102_22_n_784;
  wire mul_102_22_n_785, mul_102_22_n_786, mul_102_22_n_787, mul_102_22_n_788, mul_102_22_n_789, mul_102_22_n_790, mul_102_22_n_791, mul_102_22_n_792;
  wire mul_102_22_n_793, mul_102_22_n_794, mul_102_22_n_795, mul_102_22_n_796, mul_102_22_n_797, mul_102_22_n_798, mul_102_22_n_799, mul_102_22_n_800;
  wire mul_102_22_n_801, mul_102_22_n_802, mul_102_22_n_803, mul_102_22_n_804, mul_102_22_n_805, mul_102_22_n_806, mul_102_22_n_807, mul_102_22_n_808;
  wire mul_102_22_n_809, mul_102_22_n_810, mul_102_22_n_811, mul_102_22_n_812, mul_102_22_n_813, mul_102_22_n_814, mul_102_22_n_815, mul_102_22_n_816;
  wire mul_102_22_n_817, mul_102_22_n_818, mul_102_22_n_819, mul_102_22_n_820, mul_102_22_n_821, mul_102_22_n_822, mul_102_22_n_823, mul_102_22_n_824;
  wire mul_102_22_n_825, mul_102_22_n_826, mul_102_22_n_827, mul_102_22_n_828, mul_102_22_n_829, mul_102_22_n_830, mul_102_22_n_831, mul_102_22_n_832;
  wire mul_102_22_n_833, mul_102_22_n_834, mul_102_22_n_835, mul_102_22_n_836, mul_102_22_n_837, mul_102_22_n_838, mul_102_22_n_839, mul_102_22_n_840;
  wire mul_102_22_n_841, mul_102_22_n_842, mul_102_22_n_843, mul_102_22_n_844, mul_102_22_n_845, mul_102_22_n_846, mul_102_22_n_847, mul_102_22_n_848;
  wire mul_102_22_n_849, mul_102_22_n_850, mul_102_22_n_851, mul_102_22_n_852, mul_102_22_n_853, mul_102_22_n_854, mul_102_22_n_855, mul_102_22_n_856;
  wire mul_102_22_n_857, mul_102_22_n_858, mul_102_22_n_859, mul_102_22_n_860, mul_102_22_n_861, mul_102_22_n_862, mul_102_22_n_863, mul_102_22_n_864;
  wire mul_102_22_n_865, mul_102_22_n_866, mul_102_22_n_867, mul_102_22_n_868, mul_102_22_n_869, mul_102_22_n_870, mul_102_22_n_871, mul_102_22_n_872;
  wire mul_102_22_n_873, mul_102_22_n_874, mul_102_22_n_875, mul_102_22_n_876, mul_102_22_n_877, mul_102_22_n_878, mul_102_22_n_879, mul_102_22_n_880;
  wire mul_102_22_n_881, mul_102_22_n_882, mul_102_22_n_883, mul_102_22_n_884, mul_102_22_n_885, mul_102_22_n_886, mul_102_22_n_887, mul_102_22_n_888;
  wire mul_102_22_n_889, mul_102_22_n_890, mul_102_22_n_891, mul_102_22_n_892, mul_102_22_n_893, mul_102_22_n_894, mul_102_22_n_895, mul_102_22_n_896;
  wire mul_102_22_n_897, mul_102_22_n_898, mul_102_22_n_899, mul_102_22_n_900, mul_102_22_n_901, mul_102_22_n_902, mul_102_22_n_903, mul_102_22_n_904;
  wire mul_102_22_n_905, mul_102_22_n_906, mul_102_22_n_907, mul_102_22_n_908, mul_102_22_n_909, mul_102_22_n_910, mul_102_22_n_911, mul_102_22_n_912;
  wire mul_102_22_n_913, mul_102_22_n_914, mul_102_22_n_915, mul_102_22_n_916, mul_102_22_n_917, mul_102_22_n_918, mul_102_22_n_919, mul_102_22_n_920;
  wire mul_102_22_n_921, mul_102_22_n_922, mul_102_22_n_923, mul_102_22_n_924, mul_102_22_n_925, mul_102_22_n_926, mul_102_22_n_927, mul_102_22_n_928;
  wire mul_102_22_n_929, mul_102_22_n_930, mul_102_22_n_931, mul_102_22_n_932, mul_102_22_n_933, mul_102_22_n_934, mul_102_22_n_935, mul_102_22_n_936;
  wire mul_102_22_n_937, mul_102_22_n_938, mul_102_22_n_939, mul_102_22_n_940, mul_102_22_n_941, mul_102_22_n_942, mul_102_22_n_943, mul_102_22_n_944;
  wire mul_102_22_n_945, mul_102_22_n_946, mul_102_22_n_947, mul_102_22_n_948, mul_102_22_n_949, mul_102_22_n_950, mul_102_22_n_951, mul_102_22_n_952;
  wire mul_102_22_n_953, mul_102_22_n_954, mul_102_22_n_955, mul_102_22_n_956, mul_102_22_n_957, mul_102_22_n_958, mul_102_22_n_959, mul_102_22_n_960;
  wire mul_102_22_n_961, mul_102_22_n_962, mul_102_22_n_963, mul_102_22_n_964, mul_102_22_n_965, mul_102_22_n_966, mul_102_22_n_967, mul_102_22_n_968;
  wire mul_102_22_n_969, mul_102_22_n_970, mul_102_22_n_971, mul_102_22_n_972, mul_102_22_n_973, mul_102_22_n_974, mul_102_22_n_975, mul_102_22_n_976;
  wire mul_102_22_n_977, mul_102_22_n_978, mul_102_22_n_979, mul_102_22_n_980, mul_102_22_n_981, mul_102_22_n_982, mul_102_22_n_983, mul_102_22_n_984;
  wire mul_102_22_n_985, mul_102_22_n_986, mul_102_22_n_987, mul_102_22_n_988, mul_102_22_n_989, mul_102_22_n_990, mul_102_22_n_991, mul_102_22_n_992;
  wire mul_102_22_n_993, mul_102_22_n_994, mul_102_22_n_995, mul_102_22_n_996, mul_102_22_n_997, mul_102_22_n_998, mul_102_22_n_999, mul_102_22_n_1000;
  wire mul_102_22_n_1001, mul_102_22_n_1002, mul_102_22_n_1003, mul_102_22_n_1004, mul_102_22_n_1005, mul_102_22_n_1006, mul_102_22_n_1007, mul_102_22_n_1008;
  wire mul_102_22_n_1009, mul_102_22_n_1010, mul_102_22_n_1011, mul_102_22_n_1012, mul_102_22_n_1013, mul_102_22_n_1014, mul_102_22_n_1015, mul_102_22_n_1016;
  wire mul_102_22_n_1017, mul_102_22_n_1018, mul_102_22_n_1019, mul_102_22_n_1020, mul_102_22_n_1021, mul_102_22_n_1022, mul_102_22_n_1023, mul_102_22_n_1024;
  wire mul_102_22_n_1025, mul_102_22_n_1026, mul_102_22_n_1027, mul_102_22_n_1028, mul_102_22_n_1029, mul_102_22_n_1030, mul_102_22_n_1031, mul_102_22_n_1032;
  wire mul_102_22_n_1033, mul_102_22_n_1034, mul_102_22_n_1035, mul_102_22_n_1036, mul_102_22_n_1037, mul_102_22_n_1038, mul_102_22_n_1039, mul_102_22_n_1040;
  wire mul_102_22_n_1041, mul_102_22_n_1042, mul_102_22_n_1043, mul_102_22_n_1044, mul_102_22_n_1045, mul_102_22_n_1046, mul_102_22_n_1047, mul_102_22_n_1048;
  wire mul_102_22_n_1049, mul_102_22_n_1050, mul_102_22_n_1051, mul_102_22_n_1052, mul_102_22_n_1053, mul_102_22_n_1054, mul_102_22_n_1055, mul_102_22_n_1056;
  wire mul_102_22_n_1057, mul_102_22_n_1058, mul_102_22_n_1059, mul_102_22_n_1060, mul_102_22_n_1061, mul_102_22_n_1062, mul_102_22_n_1063, mul_102_22_n_1064;
  wire mul_102_22_n_1065, mul_102_22_n_1066, mul_102_22_n_1067, mul_102_22_n_1068, mul_102_22_n_1069, mul_102_22_n_1070, mul_102_22_n_1071, mul_102_22_n_1072;
  wire mul_102_22_n_1073, mul_102_22_n_1074, mul_102_22_n_1075, mul_102_22_n_1076, mul_102_22_n_1077, mul_102_22_n_1078, mul_102_22_n_1079, mul_102_22_n_1080;
  wire mul_102_22_n_1081, mul_102_22_n_1082, mul_102_22_n_1083, mul_102_22_n_1084, mul_102_22_n_1085, mul_102_22_n_1086, mul_102_22_n_1087, mul_102_22_n_1088;
  wire mul_102_22_n_1089, mul_102_22_n_1090, mul_102_22_n_1091, mul_102_22_n_1092, mul_102_22_n_1093, mul_102_22_n_1094, mul_102_22_n_1095, mul_102_22_n_1096;
  wire mul_102_22_n_1097, mul_102_22_n_1098, mul_102_22_n_1099, mul_102_22_n_1100, mul_102_22_n_1101, mul_102_22_n_1102, mul_102_22_n_1103, mul_102_22_n_1104;
  wire mul_102_22_n_1105, mul_102_22_n_1106, mul_102_22_n_1107, mul_102_22_n_1108, mul_102_22_n_1109, mul_102_22_n_1110, mul_102_22_n_1111, mul_102_22_n_1112;
  wire mul_102_22_n_1113, mul_102_22_n_1114, mul_102_22_n_1115, mul_102_22_n_1116, mul_102_22_n_1117, mul_102_22_n_1118, mul_102_22_n_1119, mul_102_22_n_1120;
  wire mul_102_22_n_1121, mul_102_22_n_1122, mul_102_22_n_1123, mul_102_22_n_1124, mul_102_22_n_1125, mul_102_22_n_1126, mul_102_22_n_1127, mul_102_22_n_1128;
  wire mul_102_22_n_1129, mul_102_22_n_1130, mul_102_22_n_1131, mul_102_22_n_1132, mul_102_22_n_1133, mul_102_22_n_1134, mul_102_22_n_1135, mul_102_22_n_1136;
  wire mul_102_22_n_1137, mul_102_22_n_1138, mul_102_22_n_1139, mul_102_22_n_1140, mul_102_22_n_1141, mul_102_22_n_1142, mul_102_22_n_1143, mul_102_22_n_1144;
  wire mul_102_22_n_1145, mul_102_22_n_1146, mul_102_22_n_1147, mul_102_22_n_1148, mul_102_22_n_1149, mul_102_22_n_1150, mul_102_22_n_1151, mul_102_22_n_1152;
  wire mul_102_22_n_1153, mul_102_22_n_1154, mul_102_22_n_1155, mul_102_22_n_1156, mul_102_22_n_1157, mul_108_22_n_0, mul_108_22_n_1, mul_108_22_n_2;
  wire mul_108_22_n_3, mul_108_22_n_4, mul_108_22_n_5, mul_108_22_n_6, mul_108_22_n_7, mul_108_22_n_8, mul_108_22_n_9, mul_108_22_n_10;
  wire mul_108_22_n_11, mul_108_22_n_12, mul_108_22_n_13, mul_108_22_n_14, mul_108_22_n_15, mul_108_22_n_16, mul_108_22_n_17, mul_108_22_n_18;
  wire mul_108_22_n_19, mul_108_22_n_20, mul_108_22_n_21, mul_108_22_n_22, mul_108_22_n_23, mul_108_22_n_24, mul_108_22_n_25, mul_108_22_n_26;
  wire mul_108_22_n_27, mul_108_22_n_28, mul_108_22_n_29, mul_108_22_n_30, mul_108_22_n_31, mul_108_22_n_32, mul_108_22_n_33, mul_108_22_n_34;
  wire mul_108_22_n_35, mul_108_22_n_36, mul_108_22_n_37, mul_108_22_n_38, mul_108_22_n_39, mul_108_22_n_40, mul_108_22_n_41, mul_108_22_n_42;
  wire mul_108_22_n_43, mul_108_22_n_44, mul_108_22_n_45, mul_108_22_n_46, mul_108_22_n_47, mul_108_22_n_48, mul_108_22_n_49, mul_108_22_n_50;
  wire mul_108_22_n_51, mul_108_22_n_52, mul_108_22_n_53, mul_108_22_n_54, mul_108_22_n_55, mul_108_22_n_56, mul_108_22_n_57, mul_108_22_n_58;
  wire mul_108_22_n_59, mul_108_22_n_60, mul_108_22_n_61, mul_108_22_n_62, mul_108_22_n_63, mul_108_22_n_64, mul_108_22_n_65, mul_108_22_n_66;
  wire mul_108_22_n_67, mul_108_22_n_68, mul_108_22_n_69, mul_108_22_n_70, mul_108_22_n_71, mul_108_22_n_72, mul_108_22_n_73, mul_108_22_n_74;
  wire mul_108_22_n_75, mul_108_22_n_76, mul_108_22_n_77, mul_108_22_n_78, mul_108_22_n_79, mul_108_22_n_80, mul_108_22_n_81, mul_108_22_n_82;
  wire mul_108_22_n_83, mul_108_22_n_84, mul_108_22_n_85, mul_108_22_n_86, mul_108_22_n_87, mul_108_22_n_88, mul_108_22_n_89, mul_108_22_n_90;
  wire mul_108_22_n_91, mul_108_22_n_92, mul_108_22_n_93, mul_108_22_n_94, mul_108_22_n_95, mul_108_22_n_96, mul_108_22_n_97, mul_108_22_n_98;
  wire mul_108_22_n_99, mul_108_22_n_100, mul_108_22_n_101, mul_108_22_n_102, mul_108_22_n_103, mul_108_22_n_104, mul_108_22_n_105, mul_108_22_n_106;
  wire mul_108_22_n_107, mul_108_22_n_108, mul_108_22_n_109, mul_108_22_n_110, mul_108_22_n_111, mul_108_22_n_112, mul_108_22_n_113, mul_108_22_n_114;
  wire mul_108_22_n_115, mul_108_22_n_116, mul_108_22_n_117, mul_108_22_n_118, mul_108_22_n_119, mul_108_22_n_120, mul_108_22_n_121, mul_108_22_n_122;
  wire mul_108_22_n_123, mul_108_22_n_124, mul_108_22_n_125, mul_108_22_n_126, mul_108_22_n_127, mul_108_22_n_128, mul_108_22_n_129, mul_108_22_n_130;
  wire mul_108_22_n_131, mul_108_22_n_132, mul_108_22_n_133, mul_108_22_n_134, mul_108_22_n_135, mul_108_22_n_136, mul_108_22_n_137, mul_108_22_n_138;
  wire mul_108_22_n_139, mul_108_22_n_140, mul_108_22_n_141, mul_108_22_n_142, mul_108_22_n_143, mul_108_22_n_144, mul_108_22_n_145, mul_108_22_n_146;
  wire mul_108_22_n_147, mul_108_22_n_148, mul_108_22_n_149, mul_108_22_n_150, mul_108_22_n_151, mul_108_22_n_152, mul_108_22_n_153, mul_108_22_n_154;
  wire mul_108_22_n_155, mul_108_22_n_156, mul_108_22_n_157, mul_108_22_n_158, mul_108_22_n_159, mul_108_22_n_160, mul_108_22_n_161, mul_108_22_n_162;
  wire mul_108_22_n_163, mul_108_22_n_164, mul_108_22_n_165, mul_108_22_n_166, mul_108_22_n_167, mul_108_22_n_168, mul_108_22_n_169, mul_108_22_n_170;
  wire mul_108_22_n_171, mul_108_22_n_172, mul_108_22_n_173, mul_108_22_n_174, mul_108_22_n_175, mul_108_22_n_176, mul_108_22_n_177, mul_108_22_n_178;
  wire mul_108_22_n_179, mul_108_22_n_180, mul_108_22_n_181, mul_108_22_n_182, mul_108_22_n_198, mul_108_22_n_199, mul_108_22_n_200, mul_108_22_n_201;
  wire mul_108_22_n_202, mul_108_22_n_203, mul_108_22_n_204, mul_108_22_n_205, mul_108_22_n_206, mul_108_22_n_207, mul_108_22_n_208, mul_108_22_n_209;
  wire mul_108_22_n_210, mul_108_22_n_211, mul_108_22_n_212, mul_108_22_n_213, mul_108_22_n_214, mul_108_22_n_215, mul_108_22_n_216, mul_108_22_n_217;
  wire mul_108_22_n_218, mul_108_22_n_219, mul_108_22_n_220, mul_108_22_n_221, mul_108_22_n_222, mul_108_22_n_223, mul_108_22_n_224, mul_108_22_n_225;
  wire mul_108_22_n_226, mul_108_22_n_227, mul_108_22_n_228, mul_108_22_n_229, mul_108_22_n_230, mul_108_22_n_231, mul_108_22_n_232, mul_108_22_n_233;
  wire mul_108_22_n_234, mul_108_22_n_235, mul_108_22_n_236, mul_108_22_n_237, mul_108_22_n_238, mul_108_22_n_239, mul_108_22_n_240, mul_108_22_n_241;
  wire mul_108_22_n_242, mul_108_22_n_243, mul_108_22_n_244, mul_108_22_n_245, mul_108_22_n_246, mul_108_22_n_247, mul_108_22_n_248, mul_108_22_n_249;
  wire mul_108_22_n_250, mul_108_22_n_251, mul_108_22_n_252, mul_108_22_n_253, mul_108_22_n_254, mul_108_22_n_255, mul_108_22_n_256, mul_108_22_n_257;
  wire mul_108_22_n_258, mul_108_22_n_259, mul_108_22_n_260, mul_108_22_n_261, mul_108_22_n_262, mul_108_22_n_263, mul_108_22_n_264, mul_108_22_n_265;
  wire mul_108_22_n_266, mul_108_22_n_267, mul_108_22_n_268, mul_108_22_n_269, mul_108_22_n_270, mul_108_22_n_271, mul_108_22_n_272, mul_108_22_n_273;
  wire mul_108_22_n_274, mul_108_22_n_275, mul_108_22_n_276, mul_108_22_n_277, mul_108_22_n_278, mul_108_22_n_279, mul_108_22_n_280, mul_108_22_n_281;
  wire mul_108_22_n_282, mul_108_22_n_283, mul_108_22_n_284, mul_108_22_n_285, mul_108_22_n_286, mul_108_22_n_287, mul_108_22_n_288, mul_108_22_n_289;
  wire mul_108_22_n_290, mul_108_22_n_291, mul_108_22_n_292, mul_108_22_n_293, mul_108_22_n_294, mul_108_22_n_295, mul_108_22_n_296, mul_108_22_n_297;
  wire mul_108_22_n_298, mul_108_22_n_299, mul_108_22_n_300, mul_108_22_n_301, mul_108_22_n_302, mul_108_22_n_303, mul_108_22_n_304, mul_108_22_n_305;
  wire mul_108_22_n_306, mul_108_22_n_307, mul_108_22_n_308, mul_108_22_n_310, mul_108_22_n_311, mul_108_22_n_312, mul_108_22_n_313, mul_108_22_n_314;
  wire mul_108_22_n_315, mul_108_22_n_316, mul_108_22_n_317, mul_108_22_n_318, mul_108_22_n_319, mul_108_22_n_320, mul_108_22_n_321, mul_108_22_n_322;
  wire mul_108_22_n_323, mul_108_22_n_324, mul_108_22_n_325, mul_108_22_n_326, mul_108_22_n_327, mul_108_22_n_328, mul_108_22_n_329, mul_108_22_n_330;
  wire mul_108_22_n_331, mul_108_22_n_332, mul_108_22_n_333, mul_108_22_n_334, mul_108_22_n_335, mul_108_22_n_336, mul_108_22_n_337, mul_108_22_n_338;
  wire mul_108_22_n_339, mul_108_22_n_340, mul_108_22_n_341, mul_108_22_n_342, mul_108_22_n_343, mul_108_22_n_344, mul_108_22_n_345, mul_108_22_n_346;
  wire mul_108_22_n_347, mul_108_22_n_348, mul_108_22_n_349, mul_108_22_n_350, mul_108_22_n_351, mul_108_22_n_352, mul_108_22_n_353, mul_108_22_n_354;
  wire mul_108_22_n_355, mul_108_22_n_356, mul_108_22_n_357, mul_108_22_n_358, mul_108_22_n_359, mul_108_22_n_360, mul_108_22_n_361, mul_108_22_n_362;
  wire mul_108_22_n_363, mul_108_22_n_364, mul_108_22_n_365, mul_108_22_n_366, mul_108_22_n_367, mul_108_22_n_368, mul_108_22_n_369, mul_108_22_n_370;
  wire mul_108_22_n_371, mul_108_22_n_372, mul_108_22_n_373, mul_108_22_n_374, mul_108_22_n_375, mul_108_22_n_376, mul_108_22_n_377, mul_108_22_n_378;
  wire mul_108_22_n_379, mul_108_22_n_380, mul_108_22_n_381, mul_108_22_n_382, mul_108_22_n_383, mul_108_22_n_384, mul_108_22_n_385, mul_108_22_n_386;
  wire mul_108_22_n_387, mul_108_22_n_388, mul_108_22_n_389, mul_108_22_n_390, mul_108_22_n_391, mul_108_22_n_392, mul_108_22_n_393, mul_108_22_n_394;
  wire mul_108_22_n_395, mul_108_22_n_396, mul_108_22_n_397, mul_108_22_n_398, mul_108_22_n_399, mul_108_22_n_400, mul_108_22_n_401, mul_108_22_n_402;
  wire mul_108_22_n_403, mul_108_22_n_404, mul_108_22_n_405, mul_108_22_n_406, mul_108_22_n_407, mul_108_22_n_408, mul_108_22_n_409, mul_108_22_n_410;
  wire mul_108_22_n_411, mul_108_22_n_412, mul_108_22_n_413, mul_108_22_n_414, mul_108_22_n_415, mul_108_22_n_416, mul_108_22_n_417, mul_108_22_n_418;
  wire mul_108_22_n_419, mul_108_22_n_420, mul_108_22_n_421, mul_108_22_n_422, mul_108_22_n_423, mul_108_22_n_424, mul_108_22_n_425, mul_108_22_n_426;
  wire mul_108_22_n_427, mul_108_22_n_428, mul_108_22_n_429, mul_108_22_n_430, mul_108_22_n_431, mul_108_22_n_432, mul_108_22_n_433, mul_108_22_n_434;
  wire mul_108_22_n_435, mul_108_22_n_436, mul_108_22_n_437, mul_108_22_n_438, mul_108_22_n_439, mul_108_22_n_440, mul_108_22_n_441, mul_108_22_n_442;
  wire mul_108_22_n_443, mul_108_22_n_444, mul_108_22_n_445, mul_108_22_n_446, mul_108_22_n_447, mul_108_22_n_448, mul_108_22_n_449, mul_108_22_n_450;
  wire mul_108_22_n_451, mul_108_22_n_452, mul_108_22_n_453, mul_108_22_n_454, mul_108_22_n_455, mul_108_22_n_456, mul_108_22_n_457, mul_108_22_n_458;
  wire mul_108_22_n_459, mul_108_22_n_460, mul_108_22_n_461, mul_108_22_n_462, mul_108_22_n_463, mul_108_22_n_464, mul_108_22_n_465, mul_108_22_n_466;
  wire mul_108_22_n_467, mul_108_22_n_468, mul_108_22_n_469, mul_108_22_n_470, mul_108_22_n_471, mul_108_22_n_472, mul_108_22_n_473, mul_108_22_n_474;
  wire mul_108_22_n_475, mul_108_22_n_476, mul_108_22_n_477, mul_108_22_n_478, mul_108_22_n_479, mul_108_22_n_480, mul_108_22_n_481, mul_108_22_n_482;
  wire mul_108_22_n_483, mul_108_22_n_484, mul_108_22_n_485, mul_108_22_n_486, mul_108_22_n_487, mul_108_22_n_488, mul_108_22_n_489, mul_108_22_n_490;
  wire mul_108_22_n_491, mul_108_22_n_492, mul_108_22_n_493, mul_108_22_n_494, mul_108_22_n_495, mul_108_22_n_496, mul_108_22_n_497, mul_108_22_n_498;
  wire mul_108_22_n_499, mul_108_22_n_500, mul_108_22_n_501, mul_108_22_n_502, mul_108_22_n_503, mul_108_22_n_504, mul_108_22_n_505, mul_108_22_n_506;
  wire mul_108_22_n_507, mul_108_22_n_508, mul_108_22_n_509, mul_108_22_n_510, mul_108_22_n_511, mul_108_22_n_512, mul_108_22_n_513, mul_108_22_n_514;
  wire mul_108_22_n_515, mul_108_22_n_516, mul_108_22_n_517, mul_108_22_n_518, mul_108_22_n_519, mul_108_22_n_520, mul_108_22_n_521, mul_108_22_n_522;
  wire mul_108_22_n_523, mul_108_22_n_524, mul_108_22_n_525, mul_108_22_n_526, mul_108_22_n_527, mul_108_22_n_528, mul_108_22_n_529, mul_108_22_n_530;
  wire mul_108_22_n_531, mul_108_22_n_532, mul_108_22_n_533, mul_108_22_n_534, mul_108_22_n_535, mul_108_22_n_536, mul_108_22_n_537, mul_108_22_n_538;
  wire mul_108_22_n_539, mul_108_22_n_540, mul_108_22_n_541, mul_108_22_n_542, mul_108_22_n_543, mul_108_22_n_544, mul_108_22_n_545, mul_108_22_n_546;
  wire mul_108_22_n_547, mul_108_22_n_548, mul_108_22_n_549, mul_108_22_n_550, mul_108_22_n_551, mul_108_22_n_552, mul_108_22_n_553, mul_108_22_n_554;
  wire mul_108_22_n_555, mul_108_22_n_556, mul_108_22_n_557, mul_108_22_n_558, mul_108_22_n_559, mul_108_22_n_560, mul_108_22_n_561, mul_108_22_n_562;
  wire mul_108_22_n_563, mul_108_22_n_564, mul_108_22_n_565, mul_108_22_n_566, mul_108_22_n_567, mul_108_22_n_568, mul_108_22_n_569, mul_108_22_n_570;
  wire mul_108_22_n_571, mul_108_22_n_572, mul_108_22_n_573, mul_108_22_n_574, mul_108_22_n_575, mul_108_22_n_576, mul_108_22_n_577, mul_108_22_n_578;
  wire mul_108_22_n_579, mul_108_22_n_580, mul_108_22_n_581, mul_108_22_n_582, mul_108_22_n_583, mul_108_22_n_584, mul_108_22_n_585, mul_108_22_n_586;
  wire mul_108_22_n_587, mul_108_22_n_588, mul_108_22_n_589, mul_108_22_n_590, mul_108_22_n_591, mul_108_22_n_592, mul_108_22_n_593, mul_108_22_n_594;
  wire mul_108_22_n_595, mul_108_22_n_596, mul_108_22_n_597, mul_108_22_n_598, mul_108_22_n_599, mul_108_22_n_600, mul_108_22_n_601, mul_108_22_n_602;
  wire mul_108_22_n_603, mul_108_22_n_604, mul_108_22_n_605, mul_108_22_n_606, mul_108_22_n_607, mul_108_22_n_608, mul_108_22_n_609, mul_108_22_n_610;
  wire mul_108_22_n_611, mul_108_22_n_612, mul_108_22_n_613, mul_108_22_n_614, mul_108_22_n_615, mul_108_22_n_616, mul_108_22_n_617, mul_108_22_n_618;
  wire mul_108_22_n_619, mul_108_22_n_620, mul_108_22_n_621, mul_108_22_n_622, mul_108_22_n_623, mul_108_22_n_624, mul_108_22_n_625, mul_108_22_n_626;
  wire mul_108_22_n_627, mul_108_22_n_628, mul_108_22_n_629, mul_108_22_n_630, mul_108_22_n_631, mul_108_22_n_632, mul_108_22_n_633, mul_108_22_n_634;
  wire mul_108_22_n_635, mul_108_22_n_636, mul_108_22_n_637, mul_108_22_n_638, mul_108_22_n_639, mul_108_22_n_640, mul_108_22_n_641, mul_108_22_n_642;
  wire mul_108_22_n_643, mul_108_22_n_644, mul_108_22_n_645, mul_108_22_n_646, mul_108_22_n_647, mul_108_22_n_648, mul_108_22_n_649, mul_108_22_n_650;
  wire mul_108_22_n_651, mul_108_22_n_652, mul_108_22_n_653, mul_108_22_n_654, mul_108_22_n_655, mul_108_22_n_656, mul_108_22_n_657, mul_108_22_n_658;
  wire mul_108_22_n_659, mul_108_22_n_660, mul_108_22_n_661, mul_108_22_n_662, mul_108_22_n_663, mul_108_22_n_664, mul_108_22_n_665, mul_108_22_n_666;
  wire mul_108_22_n_667, mul_108_22_n_668, mul_108_22_n_669, mul_108_22_n_670, mul_108_22_n_671, mul_108_22_n_672, mul_108_22_n_673, mul_108_22_n_674;
  wire mul_108_22_n_675, mul_108_22_n_676, mul_108_22_n_677, mul_108_22_n_678, mul_108_22_n_679, mul_108_22_n_680, mul_108_22_n_681, mul_108_22_n_682;
  wire mul_108_22_n_683, mul_108_22_n_684, mul_108_22_n_685, mul_108_22_n_686, mul_108_22_n_687, mul_108_22_n_688, mul_108_22_n_689, mul_108_22_n_690;
  wire mul_108_22_n_691, mul_108_22_n_692, mul_108_22_n_693, mul_108_22_n_694, mul_108_22_n_695, mul_108_22_n_696, mul_108_22_n_697, mul_108_22_n_698;
  wire mul_108_22_n_699, mul_108_22_n_700, mul_108_22_n_701, mul_108_22_n_702, mul_108_22_n_703, mul_108_22_n_704, mul_108_22_n_705, mul_108_22_n_706;
  wire mul_108_22_n_707, mul_108_22_n_708, mul_108_22_n_709, mul_108_22_n_710, mul_108_22_n_711, mul_108_22_n_712, mul_108_22_n_713, mul_108_22_n_714;
  wire mul_108_22_n_715, mul_108_22_n_716, mul_108_22_n_717, mul_108_22_n_718, mul_108_22_n_719, mul_108_22_n_720, mul_108_22_n_721, mul_108_22_n_722;
  wire mul_108_22_n_723, mul_108_22_n_724, mul_108_22_n_725, mul_108_22_n_726, mul_108_22_n_727, mul_108_22_n_728, mul_108_22_n_729, mul_108_22_n_730;
  wire mul_108_22_n_731, mul_108_22_n_732, mul_108_22_n_733, mul_108_22_n_734, mul_108_22_n_735, mul_108_22_n_736, mul_108_22_n_737, mul_108_22_n_738;
  wire mul_108_22_n_739, mul_108_22_n_740, mul_108_22_n_741, mul_108_22_n_742, mul_108_22_n_743, mul_108_22_n_744, mul_108_22_n_745, mul_108_22_n_746;
  wire mul_108_22_n_747, mul_108_22_n_748, mul_108_22_n_749, mul_108_22_n_750, mul_108_22_n_751, mul_108_22_n_752, mul_108_22_n_753, mul_108_22_n_754;
  wire mul_108_22_n_755, mul_108_22_n_756, mul_108_22_n_757, mul_108_22_n_758, mul_108_22_n_759, mul_108_22_n_760, mul_108_22_n_761, mul_108_22_n_762;
  wire mul_108_22_n_763, mul_108_22_n_764, mul_108_22_n_765, mul_108_22_n_766, mul_108_22_n_767, mul_108_22_n_768, mul_108_22_n_769, mul_108_22_n_770;
  wire mul_108_22_n_771, mul_108_22_n_772, mul_108_22_n_773, mul_108_22_n_774, mul_108_22_n_775, mul_108_22_n_776, mul_108_22_n_777, mul_108_22_n_778;
  wire mul_108_22_n_779, mul_108_22_n_780, mul_108_22_n_781, mul_108_22_n_782, mul_108_22_n_783, mul_108_22_n_784, mul_108_22_n_785, mul_108_22_n_786;
  wire mul_108_22_n_787, mul_108_22_n_788, mul_108_22_n_789, mul_108_22_n_790, mul_108_22_n_791, mul_108_22_n_792, mul_108_22_n_793, mul_108_22_n_794;
  wire mul_108_22_n_795, mul_108_22_n_796, mul_108_22_n_797, mul_108_22_n_798, mul_108_22_n_799, mul_108_22_n_800, mul_108_22_n_801, mul_108_22_n_802;
  wire mul_108_22_n_803, mul_108_22_n_804, mul_108_22_n_805, mul_108_22_n_806, mul_108_22_n_807, mul_108_22_n_808, mul_108_22_n_809, mul_108_22_n_810;
  wire mul_108_22_n_811, mul_108_22_n_812, mul_108_22_n_813, mul_108_22_n_814, mul_108_22_n_815, mul_108_22_n_816, mul_108_22_n_817, mul_108_22_n_818;
  wire mul_108_22_n_819, mul_108_22_n_820, mul_108_22_n_821, mul_108_22_n_822, mul_108_22_n_823, mul_108_22_n_824, mul_108_22_n_825, mul_108_22_n_826;
  wire mul_108_22_n_827, mul_108_22_n_828, mul_108_22_n_829, mul_108_22_n_830, mul_108_22_n_831, mul_108_22_n_832, mul_108_22_n_833, mul_108_22_n_834;
  wire mul_108_22_n_835, mul_108_22_n_836, mul_108_22_n_837, mul_108_22_n_838, mul_108_22_n_839, mul_108_22_n_840, mul_108_22_n_841, mul_108_22_n_842;
  wire mul_108_22_n_843, mul_108_22_n_844, mul_108_22_n_845, mul_108_22_n_846, mul_108_22_n_847, mul_108_22_n_848, mul_108_22_n_849, mul_108_22_n_850;
  wire mul_108_22_n_851, mul_108_22_n_852, mul_108_22_n_853, mul_108_22_n_854, mul_108_22_n_855, mul_108_22_n_856, mul_108_22_n_857, mul_108_22_n_858;
  wire mul_108_22_n_859, mul_108_22_n_860, mul_108_22_n_861, mul_108_22_n_862, mul_108_22_n_863, mul_108_22_n_864, mul_108_22_n_865, mul_108_22_n_866;
  wire mul_108_22_n_867, mul_108_22_n_868, mul_108_22_n_869, mul_108_22_n_870, mul_108_22_n_871, mul_108_22_n_872, mul_108_22_n_873, mul_108_22_n_874;
  wire mul_108_22_n_875, mul_108_22_n_876, mul_108_22_n_877, mul_108_22_n_878, mul_108_22_n_879, mul_108_22_n_880, mul_108_22_n_881, mul_108_22_n_882;
  wire mul_108_22_n_883, mul_108_22_n_884, mul_108_22_n_885, mul_108_22_n_886, mul_108_22_n_887, mul_108_22_n_888, mul_108_22_n_889, mul_108_22_n_890;
  wire mul_108_22_n_891, mul_108_22_n_892, mul_108_22_n_893, mul_108_22_n_894, mul_108_22_n_895, mul_108_22_n_896, mul_108_22_n_897, mul_108_22_n_898;
  wire mul_108_22_n_899, mul_108_22_n_900, mul_108_22_n_901, mul_108_22_n_902, mul_108_22_n_903, mul_108_22_n_904, mul_108_22_n_905, mul_108_22_n_906;
  wire mul_108_22_n_907, mul_108_22_n_908, mul_108_22_n_909, mul_108_22_n_910, mul_108_22_n_911, mul_108_22_n_912, mul_108_22_n_913, mul_108_22_n_914;
  wire mul_108_22_n_915, mul_108_22_n_916, mul_108_22_n_917, mul_108_22_n_918, mul_108_22_n_919, mul_108_22_n_920, mul_108_22_n_921, mul_108_22_n_922;
  wire mul_108_22_n_923, mul_108_22_n_924, mul_108_22_n_925, mul_108_22_n_926, mul_108_22_n_927, mul_108_22_n_928, mul_108_22_n_929, mul_108_22_n_930;
  wire mul_108_22_n_931, mul_108_22_n_932, mul_108_22_n_933, mul_108_22_n_934, mul_108_22_n_935, mul_108_22_n_936, mul_108_22_n_937, mul_108_22_n_938;
  wire mul_108_22_n_939, mul_108_22_n_940, mul_108_22_n_941, mul_108_22_n_942, mul_108_22_n_943, mul_108_22_n_944, mul_108_22_n_945, mul_108_22_n_946;
  wire mul_108_22_n_947, mul_108_22_n_948, mul_108_22_n_949, mul_108_22_n_950, mul_108_22_n_951, mul_108_22_n_952, mul_108_22_n_953, mul_108_22_n_954;
  wire mul_108_22_n_955, mul_108_22_n_956, mul_108_22_n_957, mul_108_22_n_958, mul_108_22_n_959, mul_108_22_n_960, mul_108_22_n_961, mul_108_22_n_962;
  wire mul_108_22_n_963, mul_108_22_n_964, mul_108_22_n_965, mul_108_22_n_966, mul_108_22_n_967, mul_108_22_n_968, mul_108_22_n_969, mul_108_22_n_970;
  wire mul_108_22_n_971, mul_108_22_n_972, mul_108_22_n_973, mul_108_22_n_974, mul_108_22_n_975, mul_108_22_n_976, mul_108_22_n_977, mul_108_22_n_978;
  wire mul_108_22_n_979, mul_108_22_n_980, mul_108_22_n_981, mul_108_22_n_982, mul_108_22_n_983, mul_108_22_n_984, mul_108_22_n_985, mul_108_22_n_986;
  wire mul_108_22_n_987, mul_108_22_n_988, mul_108_22_n_989, mul_108_22_n_990, mul_108_22_n_991, mul_108_22_n_992, mul_108_22_n_993, mul_108_22_n_994;
  wire mul_108_22_n_995, mul_108_22_n_996, mul_108_22_n_997, mul_108_22_n_998, mul_108_22_n_999, mul_108_22_n_1000, mul_108_22_n_1001, mul_108_22_n_1002;
  wire mul_108_22_n_1003, mul_108_22_n_1004, mul_108_22_n_1005, mul_108_22_n_1006, mul_108_22_n_1007, mul_108_22_n_1008, mul_108_22_n_1009, mul_108_22_n_1010;
  wire mul_108_22_n_1011, mul_108_22_n_1012, mul_108_22_n_1013, mul_108_22_n_1014, mul_108_22_n_1015, mul_108_22_n_1016, mul_108_22_n_1017, mul_108_22_n_1018;
  wire mul_108_22_n_1019, mul_108_22_n_1020, mul_108_22_n_1021, mul_108_22_n_1022, mul_108_22_n_1023, mul_108_22_n_1024, mul_108_22_n_1025, mul_108_22_n_1026;
  wire mul_108_22_n_1027, mul_108_22_n_1028, mul_108_22_n_1029, mul_108_22_n_1030, mul_108_22_n_1031, mul_108_22_n_1032, mul_108_22_n_1033, mul_108_22_n_1034;
  wire mul_108_22_n_1035, mul_108_22_n_1036, mul_108_22_n_1037, mul_108_22_n_1038, mul_108_22_n_1039, mul_108_22_n_1040, mul_108_22_n_1041, mul_108_22_n_1042;
  wire mul_108_22_n_1043, mul_108_22_n_1044, mul_108_22_n_1045, mul_108_22_n_1046, mul_108_22_n_1047, mul_108_22_n_1048, mul_108_22_n_1049, mul_108_22_n_1050;
  wire mul_108_22_n_1051, mul_108_22_n_1052, mul_108_22_n_1053, mul_108_22_n_1054, mul_108_22_n_1055, mul_108_22_n_1056, mul_108_22_n_1057, mul_108_22_n_1058;
  wire mul_108_22_n_1059, mul_108_22_n_1060, mul_108_22_n_1061, mul_108_22_n_1062, mul_108_22_n_1063, mul_108_22_n_1064, mul_108_22_n_1065, mul_108_22_n_1066;
  wire mul_108_22_n_1067, mul_108_22_n_1068, mul_108_22_n_1069, mul_108_22_n_1070, mul_108_22_n_1071, mul_108_22_n_1072, mul_108_22_n_1073, mul_108_22_n_1074;
  wire mul_108_22_n_1075, mul_108_22_n_1076, mul_108_22_n_1077, mul_108_22_n_1078, mul_108_22_n_1079, mul_108_22_n_1080, mul_108_22_n_1081, mul_108_22_n_1082;
  wire mul_108_22_n_1083, mul_108_22_n_1084, mul_108_22_n_1085, mul_108_22_n_1086, mul_108_22_n_1087, mul_108_22_n_1088, mul_108_22_n_1089, mul_108_22_n_1090;
  wire mul_108_22_n_1091, mul_108_22_n_1092, mul_108_22_n_1093, mul_108_22_n_1094, mul_108_22_n_1095, mul_108_22_n_1096, mul_108_22_n_1097, mul_108_22_n_1098;
  wire mul_108_22_n_1099, mul_108_22_n_1100, mul_108_22_n_1101, mul_108_22_n_1102, mul_108_22_n_1103, mul_108_22_n_1104, mul_108_22_n_1105, mul_108_22_n_1106;
  wire mul_108_22_n_1107, mul_108_22_n_1108, mul_108_22_n_1109, mul_108_22_n_1110, mul_108_22_n_1111, mul_108_22_n_1112, mul_108_22_n_1113, mul_108_22_n_1114;
  wire mul_108_22_n_1115, mul_108_22_n_1116, mul_108_22_n_1117, mul_108_22_n_1118, mul_108_22_n_1119, mul_108_22_n_1120, mul_108_22_n_1121, mul_108_22_n_1122;
  wire mul_108_22_n_1123, mul_108_22_n_1124, mul_108_22_n_1125, mul_108_22_n_1126, mul_108_22_n_1127, mul_108_22_n_1128, mul_108_22_n_1129, mul_108_22_n_1130;
  wire mul_108_22_n_1131, mul_108_22_n_1132, mul_108_22_n_1133, mul_108_22_n_1134, mul_108_22_n_1135, mul_108_22_n_1136, mul_108_22_n_1137, mul_108_22_n_1138;
  wire mul_108_22_n_1139, mul_108_22_n_1140, mul_108_22_n_1141, mul_108_22_n_1142, mul_108_22_n_1143, mul_108_22_n_1144, mul_108_22_n_1145, mul_108_22_n_1146;
  wire mul_108_22_n_1147, mul_108_22_n_1148, mul_108_22_n_1149, mul_108_22_n_1150, mul_108_22_n_1151, mul_108_22_n_1152, mul_108_22_n_1153, mul_108_22_n_1154;
  wire mul_108_22_n_1155, mul_108_22_n_1156, mul_108_22_n_1157, mul_113_23_n_0, mul_113_23_n_1, mul_113_23_n_2, mul_113_23_n_3, mul_113_23_n_4;
  wire mul_113_23_n_5, mul_113_23_n_6, mul_113_23_n_7, mul_113_23_n_8, mul_113_23_n_9, mul_113_23_n_10, mul_113_23_n_11, mul_113_23_n_12;
  wire mul_113_23_n_13, mul_113_23_n_14, mul_113_23_n_15, mul_113_23_n_16, mul_113_23_n_17, mul_113_23_n_18, mul_113_23_n_19, mul_113_23_n_20;
  wire mul_113_23_n_21, mul_113_23_n_22, mul_113_23_n_23, mul_113_23_n_24, mul_113_23_n_25, mul_113_23_n_26, mul_113_23_n_27, mul_113_23_n_28;
  wire mul_113_23_n_29, mul_113_23_n_30, mul_113_23_n_31, mul_113_23_n_32, mul_113_23_n_33, mul_113_23_n_34, mul_113_23_n_35, mul_113_23_n_36;
  wire mul_113_23_n_37, mul_113_23_n_38, mul_113_23_n_39, mul_113_23_n_40, mul_113_23_n_41, mul_113_23_n_42, mul_113_23_n_43, mul_113_23_n_44;
  wire mul_113_23_n_45, mul_113_23_n_46, mul_113_23_n_47, mul_113_23_n_48, mul_113_23_n_49, mul_113_23_n_50, mul_113_23_n_51, mul_113_23_n_52;
  wire mul_113_23_n_53, mul_113_23_n_54, mul_113_23_n_55, mul_113_23_n_56, mul_113_23_n_57, mul_113_23_n_58, mul_113_23_n_59, mul_113_23_n_60;
  wire mul_113_23_n_61, mul_113_23_n_62, mul_113_23_n_63, mul_113_23_n_64, mul_113_23_n_65, mul_113_23_n_66, mul_113_23_n_67, mul_113_23_n_68;
  wire mul_113_23_n_69, mul_113_23_n_70, mul_113_23_n_71, mul_113_23_n_72, mul_113_23_n_73, mul_113_23_n_74, mul_113_23_n_75, mul_113_23_n_76;
  wire mul_113_23_n_77, mul_113_23_n_78, mul_113_23_n_79, mul_113_23_n_80, mul_113_23_n_81, mul_113_23_n_82, mul_113_23_n_83, mul_113_23_n_84;
  wire mul_113_23_n_85, mul_113_23_n_86, mul_113_23_n_87, mul_113_23_n_88, mul_113_23_n_89, mul_113_23_n_90, mul_113_23_n_91, mul_113_23_n_92;
  wire mul_113_23_n_93, mul_113_23_n_94, mul_113_23_n_95, mul_113_23_n_96, mul_113_23_n_97, mul_113_23_n_110, mul_113_23_n_111, mul_113_23_n_112;
  wire mul_113_23_n_113, mul_113_23_n_114, mul_113_23_n_115, mul_113_23_n_116, mul_113_23_n_117, mul_113_23_n_118, mul_113_23_n_119, mul_113_23_n_120;
  wire mul_113_23_n_121, mul_113_23_n_122, mul_113_23_n_123, mul_113_23_n_124, mul_113_23_n_125, mul_113_23_n_126, mul_113_23_n_127, mul_113_23_n_128;
  wire mul_113_23_n_129, mul_113_23_n_130, mul_113_23_n_131, mul_113_23_n_132, mul_113_23_n_133, mul_113_23_n_134, mul_113_23_n_135, mul_113_23_n_137;
  wire mul_113_23_n_138, mul_113_23_n_139, mul_113_23_n_140, mul_113_23_n_141, mul_113_23_n_142, mul_113_23_n_143, mul_113_23_n_144, mul_113_23_n_145;
  wire mul_113_23_n_146, mul_113_23_n_147, mul_113_23_n_148, mul_113_23_n_149, mul_113_23_n_150, mul_113_23_n_151, mul_113_23_n_152, mul_113_23_n_153;
  wire mul_113_23_n_154, mul_113_23_n_155, mul_113_23_n_156, mul_113_23_n_157, mul_113_23_n_158, mul_113_23_n_159, mul_113_23_n_160, mul_113_23_n_161;
  wire mul_113_23_n_162, mul_113_23_n_163, mul_113_23_n_164, mul_113_23_n_165, mul_113_23_n_166, mul_113_23_n_167, mul_113_23_n_168, mul_113_23_n_169;
  wire mul_113_23_n_170, mul_113_23_n_171, mul_113_23_n_172, mul_113_23_n_173, mul_113_23_n_174, mul_113_23_n_175, mul_113_23_n_176, mul_113_23_n_177;
  wire mul_113_23_n_178, mul_113_23_n_179, mul_113_23_n_180, mul_113_23_n_181, mul_113_23_n_182, mul_113_23_n_183, mul_113_23_n_184, mul_113_23_n_185;
  wire mul_113_23_n_186, mul_113_23_n_187, mul_113_23_n_188, mul_113_23_n_189, mul_113_23_n_190, mul_113_23_n_191, mul_113_23_n_192, mul_113_23_n_193;
  wire mul_113_23_n_194, mul_113_23_n_195, mul_113_23_n_196, mul_113_23_n_197, mul_113_23_n_198, mul_113_23_n_199, mul_113_23_n_200, mul_113_23_n_201;
  wire mul_113_23_n_202, mul_113_23_n_203, mul_113_23_n_204, mul_113_23_n_205, mul_113_23_n_206, mul_113_23_n_207, mul_113_23_n_208, mul_113_23_n_209;
  wire mul_113_23_n_210, mul_113_23_n_211, mul_113_23_n_212, mul_113_23_n_213, mul_113_23_n_214, mul_113_23_n_215, mul_113_23_n_216, mul_113_23_n_217;
  wire mul_113_23_n_218, mul_113_23_n_219, mul_113_23_n_220, mul_113_23_n_221, mul_113_23_n_222, mul_113_23_n_223, mul_113_23_n_224, mul_113_23_n_225;
  wire mul_113_23_n_226, mul_113_23_n_227, mul_113_23_n_228, mul_113_23_n_229, mul_113_23_n_230, mul_113_23_n_231, mul_113_23_n_232, mul_113_23_n_233;
  wire mul_113_23_n_234, mul_113_23_n_235, mul_113_23_n_236, mul_113_23_n_237, mul_113_23_n_238, mul_113_23_n_239, mul_113_23_n_240, mul_113_23_n_241;
  wire mul_113_23_n_242, mul_113_23_n_243, mul_113_23_n_244, mul_113_23_n_245, mul_113_23_n_246, mul_113_23_n_247, mul_113_23_n_248, mul_113_23_n_249;
  wire mul_113_23_n_250, mul_113_23_n_251, mul_113_23_n_252, mul_113_23_n_253, mul_113_23_n_254, mul_113_23_n_255, mul_113_23_n_256, mul_113_23_n_257;
  wire mul_113_23_n_258, mul_113_23_n_259, mul_113_23_n_260, mul_113_23_n_261, mul_113_23_n_262, mul_113_23_n_263, mul_113_23_n_264, mul_113_23_n_265;
  wire mul_113_23_n_266, mul_113_23_n_267, mul_113_23_n_268, mul_113_23_n_269, mul_113_23_n_270, mul_113_23_n_271, mul_113_23_n_272, mul_113_23_n_273;
  wire mul_113_23_n_274, mul_113_23_n_275, mul_113_23_n_276, mul_113_23_n_277, mul_113_23_n_278, mul_113_23_n_279, mul_113_23_n_280, mul_113_23_n_281;
  wire mul_113_23_n_282, mul_113_23_n_283, mul_113_23_n_284, mul_113_23_n_285, mul_113_23_n_286, mul_113_23_n_287, mul_113_23_n_288, mul_113_23_n_289;
  wire mul_113_23_n_290, mul_113_23_n_291, mul_113_23_n_292, mul_113_23_n_293, mul_113_23_n_294, mul_113_23_n_295, mul_113_23_n_296, mul_113_23_n_297;
  wire mul_113_23_n_298, mul_113_23_n_299, mul_113_23_n_300, mul_113_23_n_301, mul_113_23_n_302, mul_113_23_n_303, mul_113_23_n_304, mul_113_23_n_305;
  wire mul_113_23_n_306, mul_113_23_n_307, mul_113_23_n_308, mul_113_23_n_309, mul_113_23_n_310, mul_113_23_n_311, mul_113_23_n_312, mul_113_23_n_313;
  wire mul_113_23_n_314, mul_113_23_n_315, mul_113_23_n_316, mul_113_23_n_317, mul_113_23_n_318, mul_113_23_n_319, mul_113_23_n_320, mul_113_23_n_321;
  wire mul_113_23_n_322, mul_113_23_n_323, mul_113_23_n_324, mul_113_23_n_325, mul_113_23_n_326, mul_113_23_n_327, mul_113_23_n_328, mul_113_23_n_329;
  wire mul_113_23_n_330, mul_113_23_n_331, mul_113_23_n_332, mul_113_23_n_333, mul_113_23_n_334, mul_113_23_n_335, mul_113_23_n_336, mul_113_23_n_337;
  wire mul_113_23_n_338, mul_113_23_n_339, mul_113_23_n_340, mul_113_23_n_341, mul_113_23_n_342, mul_113_23_n_343, mul_113_23_n_344, mul_113_23_n_345;
  wire mul_113_23_n_346, mul_113_23_n_347, mul_113_23_n_348, mul_113_23_n_349, mul_113_23_n_350, mul_113_23_n_351, mul_113_23_n_352, mul_113_23_n_353;
  wire mul_113_23_n_354, mul_113_23_n_355, mul_113_23_n_356, mul_113_23_n_357, mul_113_23_n_358, mul_113_23_n_359, mul_113_23_n_360, mul_113_23_n_361;
  wire mul_113_23_n_362, mul_113_23_n_363, mul_113_23_n_364, mul_113_23_n_365, mul_113_23_n_366, mul_113_23_n_367, mul_113_23_n_368, mul_113_23_n_369;
  wire mul_113_23_n_370, mul_113_23_n_371, mul_113_23_n_372, mul_113_23_n_373, mul_113_23_n_374, mul_113_23_n_375, mul_113_23_n_376, mul_113_23_n_377;
  wire mul_113_23_n_378, mul_113_23_n_379, mul_113_23_n_380, mul_113_23_n_381, mul_113_23_n_382, mul_113_23_n_383, mul_113_23_n_384, mul_113_23_n_385;
  wire mul_113_23_n_386, mul_113_23_n_387, mul_113_23_n_388, mul_113_23_n_389, mul_113_23_n_390, mul_113_23_n_391, mul_113_23_n_392, mul_113_23_n_393;
  wire mul_113_23_n_394, mul_113_23_n_395, mul_113_23_n_396, mul_113_23_n_397, mul_113_23_n_398, mul_113_23_n_399, mul_113_23_n_400, mul_113_23_n_401;
  wire mul_113_23_n_402, mul_113_23_n_403, mul_113_23_n_404, mul_113_23_n_405, mul_113_23_n_406, mul_113_23_n_407, mul_113_23_n_408, mul_113_23_n_409;
  wire mul_113_23_n_410, mul_113_23_n_411, mul_113_23_n_412, mul_113_23_n_413, mul_113_23_n_414, mul_113_23_n_415, mul_113_23_n_416, mul_113_23_n_417;
  wire mul_113_23_n_418, mul_113_23_n_419, mul_113_23_n_420, mul_113_23_n_421, mul_113_23_n_422, mul_113_23_n_423, mul_113_23_n_424, mul_113_23_n_425;
  wire mul_113_23_n_426, mul_113_23_n_427, mul_113_23_n_428, mul_113_23_n_429, mul_113_23_n_430, mul_113_23_n_431, mul_113_23_n_432, mul_113_23_n_433;
  wire mul_113_23_n_434, mul_113_23_n_435, mul_113_23_n_436, mul_113_23_n_437, mul_113_23_n_438, mul_113_23_n_439, mul_113_23_n_440, mul_113_23_n_441;
  wire mul_113_23_n_442, mul_113_23_n_443, mul_113_23_n_444, mul_113_23_n_445, mul_113_23_n_446, mul_113_23_n_447, mul_113_23_n_448, mul_113_23_n_449;
  wire mul_113_23_n_450, mul_113_23_n_451, mul_113_23_n_452, mul_113_23_n_453, mul_113_23_n_454, mul_113_23_n_455, mul_113_23_n_456, mul_113_23_n_457;
  wire mul_113_23_n_458, mul_113_23_n_459, mul_113_23_n_460, mul_113_23_n_461, mul_113_23_n_462, mul_113_23_n_463, mul_113_23_n_464, mul_113_23_n_465;
  wire mul_113_23_n_466, mul_113_23_n_467, mul_113_23_n_468, mul_113_23_n_469, mul_113_23_n_470, mul_113_23_n_471, mul_113_23_n_472, mul_113_23_n_473;
  wire mul_113_23_n_474, mul_113_23_n_475, mul_113_23_n_476, mul_113_23_n_477, mul_113_23_n_478, mul_113_23_n_479, mul_113_23_n_480, mul_113_23_n_481;
  wire mul_113_23_n_482, mul_113_23_n_483, mul_113_23_n_484, mul_113_23_n_485, mul_113_23_n_486, mul_113_23_n_487, mul_113_23_n_488, mul_113_23_n_489;
  wire mul_113_23_n_490, mul_113_23_n_491, mul_113_23_n_492, mul_113_23_n_493, mul_113_23_n_494, mul_113_23_n_495, mul_113_23_n_496, mul_113_23_n_497;
  wire mul_113_23_n_498, mul_113_23_n_499, mul_113_23_n_500, mul_113_23_n_501, mul_113_23_n_502, mul_113_23_n_503, mul_113_23_n_504, mul_113_23_n_505;
  wire mul_113_23_n_506, mul_113_23_n_507, mul_113_23_n_508, mul_113_23_n_509, mul_113_23_n_510, mul_113_23_n_511, mul_113_23_n_512, mul_113_23_n_513;
  wire mul_113_23_n_514, mul_113_23_n_515, mul_113_23_n_516, mul_113_23_n_517, mul_113_23_n_518, mul_113_23_n_519, mul_113_23_n_520, mul_113_23_n_521;
  wire mul_113_23_n_522, mul_113_23_n_523, mul_113_23_n_524, mul_113_23_n_525, mul_113_23_n_526, mul_113_23_n_527, mul_113_23_n_528, mul_113_23_n_529;
  wire mul_113_23_n_530, mul_113_23_n_531, mul_113_23_n_532, mul_113_23_n_533, mul_113_23_n_534, mul_113_23_n_535, mul_113_23_n_536, mul_113_23_n_537;
  wire mul_113_23_n_538, mul_113_23_n_539, mul_113_23_n_540, mul_113_23_n_541, mul_113_23_n_542, mul_113_23_n_543, mul_113_23_n_544, mul_113_23_n_545;
  wire mul_113_23_n_546, mul_113_23_n_547, mul_113_23_n_548, mul_113_23_n_549, mul_113_23_n_550, mul_113_23_n_551, mul_113_23_n_552, mul_113_23_n_553;
  wire mul_113_23_n_554, mul_113_23_n_555, mul_113_23_n_556, mul_113_23_n_557, mul_113_23_n_558, mul_113_23_n_559, mul_113_23_n_560, mul_113_23_n_561;
  wire mul_113_23_n_562, mul_113_23_n_563, mul_113_23_n_564, mul_113_23_n_565, mul_113_23_n_566, mul_113_23_n_567, mul_113_23_n_568, mul_113_23_n_569;
  wire mul_113_23_n_570, mul_113_23_n_571, mul_113_23_n_572, mul_113_23_n_573, mul_113_23_n_574, mul_113_23_n_575, mul_113_23_n_576, mul_113_23_n_577;
  wire mul_113_23_n_578, mul_113_23_n_579, mul_113_23_n_580, mul_113_23_n_581, mul_113_23_n_582, mul_113_23_n_583, mul_113_23_n_584, mul_113_23_n_585;
  wire mul_113_23_n_586, mul_113_23_n_587, mul_113_23_n_588, mul_113_23_n_589, mul_113_23_n_590, mul_113_23_n_591, mul_113_23_n_592, mul_113_23_n_593;
  wire mul_113_23_n_594, mul_113_23_n_595, mul_113_23_n_596, mul_113_23_n_597, mul_113_23_n_598, mul_113_23_n_599, mul_113_23_n_600, mul_113_23_n_601;
  wire mul_113_23_n_602, mul_113_23_n_603, mul_113_23_n_604, mul_113_23_n_605, mul_113_23_n_606, mul_113_23_n_607, mul_113_23_n_608, mul_113_23_n_609;
  wire mul_113_23_n_610, mul_113_23_n_611, mul_113_23_n_612, mul_113_23_n_613, mul_113_23_n_614, mul_113_23_n_615, mul_113_23_n_616, mul_113_23_n_617;
  wire mul_113_23_n_618, mul_113_23_n_619, mul_113_23_n_620, mul_113_23_n_621, mul_113_23_n_622, mul_113_23_n_623, mul_113_23_n_624, mul_113_23_n_625;
  wire mul_113_23_n_627, mul_113_23_n_628, mul_113_23_n_629, mul_113_23_n_630, mul_113_23_n_631, mul_113_23_n_632, mul_113_23_n_633, mul_113_23_n_634;
  wire mul_113_23_n_635, mul_113_23_n_636, mul_113_23_n_637, mul_113_23_n_638, mul_113_23_n_639, mul_113_23_n_640, mul_113_23_n_641, mul_113_23_n_642;
  wire mul_113_23_n_643, mul_113_23_n_644, mul_113_23_n_645, mul_113_23_n_646, mul_113_23_n_647, mul_113_23_n_648, mul_113_23_n_649, mul_113_23_n_650;
  wire mul_113_23_n_651, mul_113_23_n_652, mul_113_23_n_653, mul_113_23_n_654, mul_113_23_n_655, mul_113_23_n_656, mul_113_23_n_657, mul_113_23_n_658;
  wire mul_113_23_n_659, mul_113_23_n_660, mul_113_23_n_661, mul_113_23_n_662, mul_113_23_n_664, n_0, n_1, n_2;
  wire n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10;
  wire n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18;
  wire n_19, n_20, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
  wire n_317, n_318, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339;
  wire n_340, n_341, n_342, n_343, n_344, n_456, n_457, n_458;
  wire n_459, n_460, n_462, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_550, n_551, n_552, n_554, n_556;
  wire n_557, n_558, n_559, n_560, n_561, n_580, n_581, n_582;
  wire n_584, n_586, n_587, n_588, n_589, n_590, n_591, n_626;
  wire n_627, n_628, n_630, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_672, n_673, n_674, n_676, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_718, n_719, n_720, n_722, n_724;
  wire n_725, n_726, n_727, n_728, n_729, sub_112_23_n_1, sub_112_23_n_2, sub_112_23_n_3;
  wire sub_112_23_n_4, sub_112_23_n_5, sub_112_23_n_6, sub_112_23_n_7, sub_112_23_n_8, sub_112_23_n_9, sub_112_23_n_10, sub_112_23_n_11;
  wire sub_112_23_n_12, sub_112_23_n_13, sub_112_23_n_14, sub_112_23_n_15, sub_112_23_n_17, sub_112_23_n_18, sub_112_23_n_20, sub_112_23_n_21;
  wire sub_112_23_n_22, sub_112_23_n_23;
  and g336__2398(n_20 ,in5 ,n_127);
  and g337__5107(n_19 ,in5 ,n_141);
  and g338__6260(n_18 ,in5 ,n_139);
  and g339__4319(n_17 ,in5 ,n_135);
  and g340__8428(n_126 ,in5 ,n_142);
  and g341__5526(n_118 ,in5 ,n_134);
  and g342__6783(n_16 ,in5 ,n_138);
  and g343__3680(n_117 ,in5 ,n_133);
  and g344__1617(n_15 ,in5 ,n_130);
  and g345__2802(n_14 ,in5 ,n_140);
  and g346__1705(n_13 ,in5 ,n_137);
  and g347__5122(n_12 ,in5 ,n_131);
  and g348__8246(n_11 ,in5 ,n_132);
  and g349__7098(n_10 ,in5 ,n_136);
  and g350__6131(n_9 ,in5 ,n_129);
  and g351__1881(n_8 ,in5 ,n_128);
  buf drc_bufs(n_113 ,n_9);
  buf drc_bufs352(n_112 ,n_8);
  buf drc_bufs353(n_114 ,n_15);
  buf drc_bufs354(n_120 ,n_10);
  buf drc_bufs355(n_116 ,n_11);
  buf drc_bufs356(n_115 ,n_12);
  buf drc_bufs357(n_121 ,n_13);
  buf drc_bufs358(n_124 ,n_14);
  buf drc_bufs359(n_111 ,n_20);
  buf drc_bufs360(n_122 ,n_16);
  buf drc_bufs361(n_119 ,n_17);
  buf drc_bufs362(n_123 ,n_18);
  buf drc_bufs363(n_125 ,n_19);
  and g364__5115(n_7 ,in28 ,n_303);
  and g365__7482(n_301 ,in28 ,n_317);
  and g366__4733(n_299 ,in28 ,n_315);
  and g367__6161(n_295 ,in28 ,n_311);
  and g368__9315(n_302 ,in28 ,n_318);
  and g369__9945(n_6 ,in28 ,n_310);
  and g370__2883(n_298 ,in28 ,n_314);
  and g371__2346(n_5 ,in28 ,n_309);
  and g372__1666(n_4 ,in28 ,n_306);
  and g373__7410(n_300 ,in28 ,n_316);
  and g374__6417(n_3 ,in28 ,n_313);
  and g375__5477(n_2 ,in28 ,n_307);
  and g376__2398(n_1 ,in28 ,n_308);
  and g377__5107(n_296 ,in28 ,n_312);
  and g378__6260(n_0 ,in28 ,n_305);
  and g379__4319(n_288 ,in28 ,n_304);
  buf drc_bufs380(n_294 ,n_6);
  buf drc_bufs381(n_289 ,n_0);
  buf drc_bufs382(n_293 ,n_5);
  buf drc_bufs383(n_291 ,n_2);
  buf drc_bufs384(n_297 ,n_3);
  buf drc_bufs385(n_287 ,n_7);
  buf drc_bufs386(n_292 ,n_1);
  buf drc_bufs387(n_290 ,n_4);
  xnor add_115_23_pad_g341__8428(n_317 ,add_115_23_pad_n_94 ,n_339);
  xnor add_115_23_pad_g343__5526(n_316 ,add_115_23_pad_n_92 ,n_339);
  or add_115_23_pad_g344__6783(add_115_23_pad_n_94 ,add_115_23_pad_n_10 ,add_115_23_pad_n_92);
  and add_115_23_pad_g345__3680(n_315 ,add_115_23_pad_n_92 ,add_115_23_pad_n_91);
  or add_115_23_pad_g346__1617(add_115_23_pad_n_92 ,add_115_23_pad_n_16 ,add_115_23_pad_n_89);
  or add_115_23_pad_g347__2802(add_115_23_pad_n_91 ,n_338 ,add_115_23_pad_n_90);
  not add_115_23_pad_g348(add_115_23_pad_n_90 ,add_115_23_pad_n_89);
  and add_115_23_pad_g349__1705(add_115_23_pad_n_89 ,add_115_23_pad_n_33 ,add_115_23_pad_n_88);
  or add_115_23_pad_g351__5122(add_115_23_pad_n_88 ,add_115_23_pad_n_31 ,add_115_23_pad_n_87);
  and add_115_23_pad_g353__8246(add_115_23_pad_n_87 ,add_115_23_pad_n_37 ,add_115_23_pad_n_86);
  or add_115_23_pad_g355__7098(add_115_23_pad_n_86 ,add_115_23_pad_n_35 ,add_115_23_pad_n_85);
  and add_115_23_pad_g357__6131(add_115_23_pad_n_85 ,add_115_23_pad_n_41 ,add_115_23_pad_n_84);
  or add_115_23_pad_g359__1881(add_115_23_pad_n_84 ,add_115_23_pad_n_36 ,add_115_23_pad_n_83);
  and add_115_23_pad_g361__5115(add_115_23_pad_n_83 ,add_115_23_pad_n_34 ,add_115_23_pad_n_82);
  or add_115_23_pad_g363__7482(add_115_23_pad_n_82 ,add_115_23_pad_n_39 ,add_115_23_pad_n_81);
  and add_115_23_pad_g365__4733(add_115_23_pad_n_81 ,add_115_23_pad_n_28 ,add_115_23_pad_n_80);
  or add_115_23_pad_g367__6161(add_115_23_pad_n_80 ,add_115_23_pad_n_47 ,add_115_23_pad_n_79);
  and add_115_23_pad_g369__9315(add_115_23_pad_n_79 ,add_115_23_pad_n_32 ,add_115_23_pad_n_78);
  or add_115_23_pad_g371__9945(add_115_23_pad_n_78 ,add_115_23_pad_n_38 ,add_115_23_pad_n_77);
  and add_115_23_pad_g373__2883(add_115_23_pad_n_77 ,add_115_23_pad_n_46 ,add_115_23_pad_n_75);
  xnor add_115_23_pad_g374__2346(n_308 ,add_115_23_pad_n_73 ,add_115_23_pad_n_57);
  or add_115_23_pad_g375__1666(add_115_23_pad_n_75 ,add_115_23_pad_n_43 ,add_115_23_pad_n_74);
  not add_115_23_pad_g376(add_115_23_pad_n_74 ,add_115_23_pad_n_73);
  or add_115_23_pad_g377__7410(add_115_23_pad_n_73 ,add_115_23_pad_n_45 ,add_115_23_pad_n_71);
  xnor add_115_23_pad_g378__6417(n_307 ,add_115_23_pad_n_70 ,add_115_23_pad_n_56);
  and add_115_23_pad_g379__5477(add_115_23_pad_n_71 ,add_115_23_pad_n_26 ,add_115_23_pad_n_70);
  or add_115_23_pad_g380__2398(add_115_23_pad_n_70 ,add_115_23_pad_n_29 ,add_115_23_pad_n_68);
  xnor add_115_23_pad_g381__5107(n_306 ,add_115_23_pad_n_67 ,add_115_23_pad_n_58);
  and add_115_23_pad_g382__6260(add_115_23_pad_n_68 ,add_115_23_pad_n_30 ,add_115_23_pad_n_67);
  or add_115_23_pad_g383__4319(add_115_23_pad_n_67 ,add_115_23_pad_n_27 ,add_115_23_pad_n_65);
  xnor add_115_23_pad_g384__8428(n_305 ,add_115_23_pad_n_63 ,add_115_23_pad_n_59);
  and add_115_23_pad_g385__5526(add_115_23_pad_n_65 ,add_115_23_pad_n_42 ,add_115_23_pad_n_63);
  xor add_115_23_pad_g386__6783(n_304 ,add_115_23_pad_n_49 ,add_115_23_pad_n_60);
  or add_115_23_pad_g387__3680(add_115_23_pad_n_63 ,add_115_23_pad_n_44 ,add_115_23_pad_n_62);
  nor add_115_23_pad_g388__1617(add_115_23_pad_n_62 ,add_115_23_pad_n_49 ,add_115_23_pad_n_48);
  and add_115_23_pad_g389__2802(n_303 ,add_115_23_pad_n_49 ,add_115_23_pad_n_40);
  xnor add_115_23_pad_g390__1705(add_115_23_pad_n_60 ,n_327 ,in30[1]);
  xnor add_115_23_pad_g391__5122(add_115_23_pad_n_59 ,n_328 ,in30[2]);
  xnor add_115_23_pad_g392__8246(add_115_23_pad_n_58 ,n_329 ,in30[3]);
  xnor add_115_23_pad_g393__7098(add_115_23_pad_n_57 ,n_331 ,in30[5]);
  xnor add_115_23_pad_g394__6131(add_115_23_pad_n_56 ,n_330 ,in30[4]);
  xnor add_115_23_pad_g395__1881(add_115_23_pad_n_55 ,n_336 ,in30[10]);
  xnor add_115_23_pad_g396__5115(add_115_23_pad_n_54 ,n_335 ,in30[9]);
  xnor add_115_23_pad_g397__7482(add_115_23_pad_n_53 ,n_334 ,in30[8]);
  xnor add_115_23_pad_g398__4733(add_115_23_pad_n_52 ,n_333 ,in30[7]);
  xnor add_115_23_pad_g399__6161(add_115_23_pad_n_51 ,n_332 ,in30[6]);
  xnor add_115_23_pad_g400__9315(add_115_23_pad_n_50 ,n_337 ,in30[11]);
  nor add_115_23_pad_g401__9945(add_115_23_pad_n_48 ,in30[1] ,n_327);
  nor add_115_23_pad_g402__2883(add_115_23_pad_n_47 ,in30[7] ,n_333);
  or add_115_23_pad_g403__2346(add_115_23_pad_n_46 ,add_115_23_pad_n_24 ,add_115_23_pad_n_23);
  and add_115_23_pad_g404__1666(add_115_23_pad_n_45 ,in30[4] ,n_330);
  and add_115_23_pad_g405__7410(add_115_23_pad_n_44 ,in30[1] ,n_327);
  nor add_115_23_pad_g406__6417(add_115_23_pad_n_43 ,in30[5] ,n_331);
  or add_115_23_pad_g407__5477(add_115_23_pad_n_42 ,in30[2] ,n_328);
  or add_115_23_pad_g408__2398(add_115_23_pad_n_41 ,add_115_23_pad_n_12 ,add_115_23_pad_n_19);
  or add_115_23_pad_g409__5107(add_115_23_pad_n_40 ,in30[0] ,n_326);
  nor add_115_23_pad_g410__6260(add_115_23_pad_n_39 ,in30[8] ,n_334);
  nor add_115_23_pad_g411__4319(add_115_23_pad_n_38 ,in30[6] ,n_332);
  or add_115_23_pad_g412__8428(add_115_23_pad_n_49 ,add_115_23_pad_n_14 ,add_115_23_pad_n_15);
  or add_115_23_pad_g413__5526(add_115_23_pad_n_37 ,add_115_23_pad_n_18 ,add_115_23_pad_n_9);
  nor add_115_23_pad_g414__6783(add_115_23_pad_n_36 ,in30[9] ,n_335);
  nor add_115_23_pad_g415__3680(add_115_23_pad_n_35 ,in30[10] ,n_336);
  or add_115_23_pad_g416__1617(add_115_23_pad_n_34 ,add_115_23_pad_n_21 ,add_115_23_pad_n_22);
  or add_115_23_pad_g417__2802(add_115_23_pad_n_33 ,add_115_23_pad_n_17 ,add_115_23_pad_n_13);
  or add_115_23_pad_g418__1705(add_115_23_pad_n_32 ,add_115_23_pad_n_25 ,add_115_23_pad_n_8);
  nor add_115_23_pad_g419__5122(add_115_23_pad_n_31 ,in30[11] ,n_337);
  or add_115_23_pad_g420__8246(add_115_23_pad_n_30 ,in30[3] ,n_329);
  and add_115_23_pad_g421__7098(add_115_23_pad_n_29 ,in30[3] ,n_329);
  or add_115_23_pad_g422__6131(add_115_23_pad_n_28 ,add_115_23_pad_n_11 ,add_115_23_pad_n_20);
  and add_115_23_pad_g423__1881(add_115_23_pad_n_27 ,in30[2] ,n_328);
  or add_115_23_pad_g424__5115(add_115_23_pad_n_26 ,in30[4] ,n_330);
  not add_115_23_pad_g425(add_115_23_pad_n_25 ,in30[6]);
  not add_115_23_pad_g426(add_115_23_pad_n_24 ,in30[5]);
  not add_115_23_pad_g427(add_115_23_pad_n_23 ,n_331);
  not add_115_23_pad_g428(add_115_23_pad_n_22 ,n_334);
  not add_115_23_pad_g429(add_115_23_pad_n_21 ,in30[8]);
  not add_115_23_pad_g430(add_115_23_pad_n_20 ,n_333);
  not add_115_23_pad_g431(add_115_23_pad_n_19 ,n_335);
  not add_115_23_pad_g432(add_115_23_pad_n_18 ,in30[10]);
  not add_115_23_pad_g433(add_115_23_pad_n_17 ,in30[11]);
  not add_115_23_pad_g434(add_115_23_pad_n_16 ,n_338);
  not add_115_23_pad_g435(add_115_23_pad_n_15 ,n_326);
  not add_115_23_pad_g436(add_115_23_pad_n_14 ,in30[0]);
  not add_115_23_pad_g437(add_115_23_pad_n_13 ,n_337);
  not add_115_23_pad_g438(add_115_23_pad_n_12 ,in30[9]);
  not add_115_23_pad_g439(add_115_23_pad_n_11 ,in30[7]);
  not add_115_23_pad_g440(add_115_23_pad_n_10 ,n_339);
  not add_115_23_pad_g441(add_115_23_pad_n_9 ,n_336);
  not add_115_23_pad_g442(add_115_23_pad_n_8 ,n_332);
  buf add_115_23_pad_drc_bufs(n_318 ,add_115_23_pad_n_96);
  xor add_115_23_pad_g2__7482(n_314 ,add_115_23_pad_n_87 ,add_115_23_pad_n_50);
  xor add_115_23_pad_g444__4733(n_313 ,add_115_23_pad_n_85 ,add_115_23_pad_n_55);
  xor add_115_23_pad_g445__6161(n_312 ,add_115_23_pad_n_83 ,add_115_23_pad_n_54);
  xor add_115_23_pad_g446__9315(n_311 ,add_115_23_pad_n_81 ,add_115_23_pad_n_53);
  xor add_115_23_pad_g447__9945(n_310 ,add_115_23_pad_n_79 ,add_115_23_pad_n_52);
  xor add_115_23_pad_g448__2883(n_309 ,add_115_23_pad_n_77 ,add_115_23_pad_n_51);
  xnor csa_tree_add_83_21_pad_groupi_g4151__2346(n_206 ,csa_tree_add_83_21_pad_groupi_n_1336 ,csa_tree_add_83_21_pad_groupi_n_1558);
  or csa_tree_add_83_21_pad_groupi_g4152__1666(csa_tree_add_83_21_pad_groupi_n_1558 ,csa_tree_add_83_21_pad_groupi_n_1393 ,csa_tree_add_83_21_pad_groupi_n_1556);
  xnor csa_tree_add_83_21_pad_groupi_g4153__7410(n_205 ,csa_tree_add_83_21_pad_groupi_n_1555 ,csa_tree_add_83_21_pad_groupi_n_1404);
  and csa_tree_add_83_21_pad_groupi_g4154__6417(csa_tree_add_83_21_pad_groupi_n_1556 ,csa_tree_add_83_21_pad_groupi_n_1389 ,csa_tree_add_83_21_pad_groupi_n_1555);
  or csa_tree_add_83_21_pad_groupi_g4155__5477(csa_tree_add_83_21_pad_groupi_n_1555 ,csa_tree_add_83_21_pad_groupi_n_1407 ,csa_tree_add_83_21_pad_groupi_n_1553);
  xnor csa_tree_add_83_21_pad_groupi_g4156__2398(n_204 ,csa_tree_add_83_21_pad_groupi_n_1552 ,csa_tree_add_83_21_pad_groupi_n_1434);
  and csa_tree_add_83_21_pad_groupi_g4157__5107(csa_tree_add_83_21_pad_groupi_n_1553 ,csa_tree_add_83_21_pad_groupi_n_1410 ,csa_tree_add_83_21_pad_groupi_n_1552);
  or csa_tree_add_83_21_pad_groupi_g4158__6260(csa_tree_add_83_21_pad_groupi_n_1552 ,csa_tree_add_83_21_pad_groupi_n_1453 ,csa_tree_add_83_21_pad_groupi_n_1550);
  xnor csa_tree_add_83_21_pad_groupi_g4159__4319(n_203 ,csa_tree_add_83_21_pad_groupi_n_1549 ,csa_tree_add_83_21_pad_groupi_n_1462);
  and csa_tree_add_83_21_pad_groupi_g4160__8428(csa_tree_add_83_21_pad_groupi_n_1550 ,csa_tree_add_83_21_pad_groupi_n_1459 ,csa_tree_add_83_21_pad_groupi_n_1549);
  or csa_tree_add_83_21_pad_groupi_g4161__5526(csa_tree_add_83_21_pad_groupi_n_1549 ,csa_tree_add_83_21_pad_groupi_n_1463 ,csa_tree_add_83_21_pad_groupi_n_1547);
  xnor csa_tree_add_83_21_pad_groupi_g4162__6783(n_202 ,csa_tree_add_83_21_pad_groupi_n_1546 ,csa_tree_add_83_21_pad_groupi_n_1483);
  nor csa_tree_add_83_21_pad_groupi_g4163__3680(csa_tree_add_83_21_pad_groupi_n_1547 ,csa_tree_add_83_21_pad_groupi_n_1546 ,csa_tree_add_83_21_pad_groupi_n_1464);
  and csa_tree_add_83_21_pad_groupi_g4164__1617(csa_tree_add_83_21_pad_groupi_n_1546 ,csa_tree_add_83_21_pad_groupi_n_1500 ,csa_tree_add_83_21_pad_groupi_n_1544);
  xnor csa_tree_add_83_21_pad_groupi_g4165__2802(n_201 ,csa_tree_add_83_21_pad_groupi_n_1542 ,csa_tree_add_83_21_pad_groupi_n_1501);
  or csa_tree_add_83_21_pad_groupi_g4166__1705(csa_tree_add_83_21_pad_groupi_n_1544 ,csa_tree_add_83_21_pad_groupi_n_1494 ,csa_tree_add_83_21_pad_groupi_n_1543);
  not csa_tree_add_83_21_pad_groupi_g4167(csa_tree_add_83_21_pad_groupi_n_1543 ,csa_tree_add_83_21_pad_groupi_n_1542);
  or csa_tree_add_83_21_pad_groupi_g4168__5122(csa_tree_add_83_21_pad_groupi_n_1542 ,csa_tree_add_83_21_pad_groupi_n_1499 ,csa_tree_add_83_21_pad_groupi_n_1540);
  xnor csa_tree_add_83_21_pad_groupi_g4169__8246(n_200 ,csa_tree_add_83_21_pad_groupi_n_1539 ,csa_tree_add_83_21_pad_groupi_n_1503);
  nor csa_tree_add_83_21_pad_groupi_g4170__7098(csa_tree_add_83_21_pad_groupi_n_1540 ,csa_tree_add_83_21_pad_groupi_n_1496 ,csa_tree_add_83_21_pad_groupi_n_1539);
  and csa_tree_add_83_21_pad_groupi_g4171__6131(csa_tree_add_83_21_pad_groupi_n_1539 ,csa_tree_add_83_21_pad_groupi_n_1538 ,csa_tree_add_83_21_pad_groupi_n_1510);
  or csa_tree_add_83_21_pad_groupi_g4173__1881(csa_tree_add_83_21_pad_groupi_n_1538 ,csa_tree_add_83_21_pad_groupi_n_1513 ,csa_tree_add_83_21_pad_groupi_n_1537);
  and csa_tree_add_83_21_pad_groupi_g4175__5115(csa_tree_add_83_21_pad_groupi_n_1537 ,csa_tree_add_83_21_pad_groupi_n_1512 ,csa_tree_add_83_21_pad_groupi_n_1535);
  xnor csa_tree_add_83_21_pad_groupi_g4176__7482(n_198 ,csa_tree_add_83_21_pad_groupi_n_1534 ,csa_tree_add_83_21_pad_groupi_n_1519);
  or csa_tree_add_83_21_pad_groupi_g4177__4733(csa_tree_add_83_21_pad_groupi_n_1535 ,csa_tree_add_83_21_pad_groupi_n_1514 ,csa_tree_add_83_21_pad_groupi_n_1534);
  and csa_tree_add_83_21_pad_groupi_g4178__6161(csa_tree_add_83_21_pad_groupi_n_1534 ,csa_tree_add_83_21_pad_groupi_n_1533 ,csa_tree_add_83_21_pad_groupi_n_1511);
  or csa_tree_add_83_21_pad_groupi_g4180__9315(csa_tree_add_83_21_pad_groupi_n_1533 ,csa_tree_add_83_21_pad_groupi_n_1505 ,csa_tree_add_83_21_pad_groupi_n_1532);
  and csa_tree_add_83_21_pad_groupi_g4182__9945(csa_tree_add_83_21_pad_groupi_n_1532 ,csa_tree_add_83_21_pad_groupi_n_1506 ,csa_tree_add_83_21_pad_groupi_n_1530);
  xnor csa_tree_add_83_21_pad_groupi_g4183__2883(n_196 ,csa_tree_add_83_21_pad_groupi_n_1529 ,csa_tree_add_83_21_pad_groupi_n_1517);
  or csa_tree_add_83_21_pad_groupi_g4184__2346(csa_tree_add_83_21_pad_groupi_n_1530 ,csa_tree_add_83_21_pad_groupi_n_1507 ,csa_tree_add_83_21_pad_groupi_n_1529);
  and csa_tree_add_83_21_pad_groupi_g4185__1666(csa_tree_add_83_21_pad_groupi_n_1529 ,csa_tree_add_83_21_pad_groupi_n_1508 ,csa_tree_add_83_21_pad_groupi_n_1527);
  xnor csa_tree_add_83_21_pad_groupi_g4186__7410(n_195 ,csa_tree_add_83_21_pad_groupi_n_1526 ,csa_tree_add_83_21_pad_groupi_n_1516);
  or csa_tree_add_83_21_pad_groupi_g4187__6417(csa_tree_add_83_21_pad_groupi_n_1527 ,csa_tree_add_83_21_pad_groupi_n_1526 ,csa_tree_add_83_21_pad_groupi_n_1509);
  and csa_tree_add_83_21_pad_groupi_g4188__5477(csa_tree_add_83_21_pad_groupi_n_1526 ,csa_tree_add_83_21_pad_groupi_n_1471 ,csa_tree_add_83_21_pad_groupi_n_1525);
  or csa_tree_add_83_21_pad_groupi_g4190__2398(csa_tree_add_83_21_pad_groupi_n_1525 ,csa_tree_add_83_21_pad_groupi_n_1470 ,csa_tree_add_83_21_pad_groupi_n_1524);
  and csa_tree_add_83_21_pad_groupi_g4192__5107(csa_tree_add_83_21_pad_groupi_n_1524 ,csa_tree_add_83_21_pad_groupi_n_1498 ,csa_tree_add_83_21_pad_groupi_n_1523);
  or csa_tree_add_83_21_pad_groupi_g4194__6260(csa_tree_add_83_21_pad_groupi_n_1523 ,csa_tree_add_83_21_pad_groupi_n_1497 ,csa_tree_add_83_21_pad_groupi_n_1522);
  and csa_tree_add_83_21_pad_groupi_g4196__4319(csa_tree_add_83_21_pad_groupi_n_1522 ,csa_tree_add_83_21_pad_groupi_n_1452 ,csa_tree_add_83_21_pad_groupi_n_1521);
  or csa_tree_add_83_21_pad_groupi_g4198__8428(csa_tree_add_83_21_pad_groupi_n_1521 ,csa_tree_add_83_21_pad_groupi_n_1451 ,csa_tree_add_83_21_pad_groupi_n_1515);
  xnor csa_tree_add_83_21_pad_groupi_g4199__5526(csa_tree_add_83_21_pad_groupi_n_1520 ,csa_tree_add_83_21_pad_groupi_n_1475 ,csa_tree_add_83_21_pad_groupi_n_1491);
  xnor csa_tree_add_83_21_pad_groupi_g4200__6783(csa_tree_add_83_21_pad_groupi_n_1519 ,csa_tree_add_83_21_pad_groupi_n_1473 ,csa_tree_add_83_21_pad_groupi_n_1489);
  xnor csa_tree_add_83_21_pad_groupi_g4201__3680(csa_tree_add_83_21_pad_groupi_n_1518 ,csa_tree_add_83_21_pad_groupi_n_1480 ,csa_tree_add_83_21_pad_groupi_n_1487);
  xnor csa_tree_add_83_21_pad_groupi_g4202__1617(csa_tree_add_83_21_pad_groupi_n_1517 ,csa_tree_add_83_21_pad_groupi_n_1477 ,csa_tree_add_83_21_pad_groupi_n_1493);
  xnor csa_tree_add_83_21_pad_groupi_g4203__2802(csa_tree_add_83_21_pad_groupi_n_1516 ,csa_tree_add_83_21_pad_groupi_n_1448 ,csa_tree_add_83_21_pad_groupi_n_1485);
  nor csa_tree_add_83_21_pad_groupi_g4205__1705(csa_tree_add_83_21_pad_groupi_n_1514 ,csa_tree_add_83_21_pad_groupi_n_1472 ,csa_tree_add_83_21_pad_groupi_n_1489);
  nor csa_tree_add_83_21_pad_groupi_g4206__5122(csa_tree_add_83_21_pad_groupi_n_1513 ,csa_tree_add_83_21_pad_groupi_n_1475 ,csa_tree_add_83_21_pad_groupi_n_1491);
  or csa_tree_add_83_21_pad_groupi_g4207__8246(csa_tree_add_83_21_pad_groupi_n_1512 ,csa_tree_add_83_21_pad_groupi_n_1473 ,csa_tree_add_83_21_pad_groupi_n_1488);
  or csa_tree_add_83_21_pad_groupi_g4208__7098(csa_tree_add_83_21_pad_groupi_n_1511 ,csa_tree_add_83_21_pad_groupi_n_1479 ,csa_tree_add_83_21_pad_groupi_n_1486);
  or csa_tree_add_83_21_pad_groupi_g4209__6131(csa_tree_add_83_21_pad_groupi_n_1510 ,csa_tree_add_83_21_pad_groupi_n_1474 ,csa_tree_add_83_21_pad_groupi_n_1490);
  nor csa_tree_add_83_21_pad_groupi_g4210__1881(csa_tree_add_83_21_pad_groupi_n_1509 ,csa_tree_add_83_21_pad_groupi_n_1447 ,csa_tree_add_83_21_pad_groupi_n_1485);
  and csa_tree_add_83_21_pad_groupi_g4211__5115(csa_tree_add_83_21_pad_groupi_n_1515 ,csa_tree_add_83_21_pad_groupi_n_1450 ,csa_tree_add_83_21_pad_groupi_n_1495);
  or csa_tree_add_83_21_pad_groupi_g4212__7482(csa_tree_add_83_21_pad_groupi_n_1508 ,csa_tree_add_83_21_pad_groupi_n_1448 ,csa_tree_add_83_21_pad_groupi_n_1484);
  nor csa_tree_add_83_21_pad_groupi_g4213__4733(csa_tree_add_83_21_pad_groupi_n_1507 ,csa_tree_add_83_21_pad_groupi_n_1476 ,csa_tree_add_83_21_pad_groupi_n_1493);
  or csa_tree_add_83_21_pad_groupi_g4214__6161(csa_tree_add_83_21_pad_groupi_n_1506 ,csa_tree_add_83_21_pad_groupi_n_1477 ,csa_tree_add_83_21_pad_groupi_n_1492);
  nor csa_tree_add_83_21_pad_groupi_g4215__9315(csa_tree_add_83_21_pad_groupi_n_1505 ,csa_tree_add_83_21_pad_groupi_n_1480 ,csa_tree_add_83_21_pad_groupi_n_1487);
  xnor csa_tree_add_83_21_pad_groupi_g4216__9945(n_191 ,csa_tree_add_83_21_pad_groupi_n_1481 ,csa_tree_add_83_21_pad_groupi_n_1460);
  xnor csa_tree_add_83_21_pad_groupi_g4217__2883(csa_tree_add_83_21_pad_groupi_n_1503 ,csa_tree_add_83_21_pad_groupi_n_1478 ,csa_tree_add_83_21_pad_groupi_n_1467);
  xnor csa_tree_add_83_21_pad_groupi_g4218__2346(csa_tree_add_83_21_pad_groupi_n_1502 ,csa_tree_add_83_21_pad_groupi_n_1412 ,csa_tree_add_83_21_pad_groupi_n_1466);
  xnor csa_tree_add_83_21_pad_groupi_g4219__1666(csa_tree_add_83_21_pad_groupi_n_1501 ,csa_tree_add_83_21_pad_groupi_n_1442 ,csa_tree_add_83_21_pad_groupi_n_1469);
  or csa_tree_add_83_21_pad_groupi_g4220__7410(csa_tree_add_83_21_pad_groupi_n_1500 ,csa_tree_add_83_21_pad_groupi_n_1441 ,csa_tree_add_83_21_pad_groupi_n_6);
  nor csa_tree_add_83_21_pad_groupi_g4221__6417(csa_tree_add_83_21_pad_groupi_n_1499 ,csa_tree_add_83_21_pad_groupi_n_1478 ,csa_tree_add_83_21_pad_groupi_n_1468);
  or csa_tree_add_83_21_pad_groupi_g4222__5477(csa_tree_add_83_21_pad_groupi_n_1498 ,csa_tree_add_83_21_pad_groupi_n_1411 ,csa_tree_add_83_21_pad_groupi_n_1465);
  nor csa_tree_add_83_21_pad_groupi_g4223__2398(csa_tree_add_83_21_pad_groupi_n_1497 ,csa_tree_add_83_21_pad_groupi_n_1412 ,csa_tree_add_83_21_pad_groupi_n_1466);
  and csa_tree_add_83_21_pad_groupi_g4224__5107(csa_tree_add_83_21_pad_groupi_n_1496 ,csa_tree_add_83_21_pad_groupi_n_1478 ,csa_tree_add_83_21_pad_groupi_n_1468);
  or csa_tree_add_83_21_pad_groupi_g4225__6260(csa_tree_add_83_21_pad_groupi_n_1495 ,csa_tree_add_83_21_pad_groupi_n_1449 ,csa_tree_add_83_21_pad_groupi_n_1481);
  nor csa_tree_add_83_21_pad_groupi_g4226__4319(csa_tree_add_83_21_pad_groupi_n_1494 ,csa_tree_add_83_21_pad_groupi_n_1442 ,csa_tree_add_83_21_pad_groupi_n_1469);
  not csa_tree_add_83_21_pad_groupi_g4227(csa_tree_add_83_21_pad_groupi_n_1493 ,csa_tree_add_83_21_pad_groupi_n_1492);
  not csa_tree_add_83_21_pad_groupi_g4228(csa_tree_add_83_21_pad_groupi_n_1491 ,csa_tree_add_83_21_pad_groupi_n_1490);
  not csa_tree_add_83_21_pad_groupi_g4229(csa_tree_add_83_21_pad_groupi_n_1489 ,csa_tree_add_83_21_pad_groupi_n_1488);
  not csa_tree_add_83_21_pad_groupi_g4230(csa_tree_add_83_21_pad_groupi_n_1487 ,csa_tree_add_83_21_pad_groupi_n_1486);
  not csa_tree_add_83_21_pad_groupi_g4231(csa_tree_add_83_21_pad_groupi_n_1485 ,csa_tree_add_83_21_pad_groupi_n_1484);
  xnor csa_tree_add_83_21_pad_groupi_g4232__8428(csa_tree_add_83_21_pad_groupi_n_1483 ,csa_tree_add_83_21_pad_groupi_n_1440 ,csa_tree_add_83_21_pad_groupi_n_1445);
  xnor csa_tree_add_83_21_pad_groupi_g4233__5526(csa_tree_add_83_21_pad_groupi_n_1482 ,csa_tree_add_83_21_pad_groupi_n_1419 ,csa_tree_add_83_21_pad_groupi_n_1444);
  xnor csa_tree_add_83_21_pad_groupi_g4234__6783(csa_tree_add_83_21_pad_groupi_n_1492 ,csa_tree_add_83_21_pad_groupi_n_1387 ,csa_tree_add_83_21_pad_groupi_n_1438);
  xnor csa_tree_add_83_21_pad_groupi_g4235__3680(csa_tree_add_83_21_pad_groupi_n_1490 ,csa_tree_add_83_21_pad_groupi_n_1400 ,csa_tree_add_83_21_pad_groupi_n_1433);
  xnor csa_tree_add_83_21_pad_groupi_g4236__1617(csa_tree_add_83_21_pad_groupi_n_1488 ,csa_tree_add_83_21_pad_groupi_n_1401 ,csa_tree_add_83_21_pad_groupi_n_1436);
  xnor csa_tree_add_83_21_pad_groupi_g4237__2802(csa_tree_add_83_21_pad_groupi_n_1486 ,csa_tree_add_83_21_pad_groupi_n_1402 ,csa_tree_add_83_21_pad_groupi_n_1437);
  xnor csa_tree_add_83_21_pad_groupi_g4238__1705(csa_tree_add_83_21_pad_groupi_n_1484 ,csa_tree_add_83_21_pad_groupi_n_1403 ,csa_tree_add_83_21_pad_groupi_n_1435);
  not csa_tree_add_83_21_pad_groupi_g4239(csa_tree_add_83_21_pad_groupi_n_1479 ,csa_tree_add_83_21_pad_groupi_n_1480);
  not csa_tree_add_83_21_pad_groupi_g4240(csa_tree_add_83_21_pad_groupi_n_1477 ,csa_tree_add_83_21_pad_groupi_n_1476);
  not csa_tree_add_83_21_pad_groupi_g4241(csa_tree_add_83_21_pad_groupi_n_1474 ,csa_tree_add_83_21_pad_groupi_n_1475);
  not csa_tree_add_83_21_pad_groupi_g4242(csa_tree_add_83_21_pad_groupi_n_1473 ,csa_tree_add_83_21_pad_groupi_n_1472);
  or csa_tree_add_83_21_pad_groupi_g4243__5122(csa_tree_add_83_21_pad_groupi_n_1471 ,csa_tree_add_83_21_pad_groupi_n_1418 ,csa_tree_add_83_21_pad_groupi_n_1443);
  nor csa_tree_add_83_21_pad_groupi_g4244__8246(csa_tree_add_83_21_pad_groupi_n_1470 ,csa_tree_add_83_21_pad_groupi_n_1419 ,csa_tree_add_83_21_pad_groupi_n_1444);
  and csa_tree_add_83_21_pad_groupi_g4245__7098(csa_tree_add_83_21_pad_groupi_n_1481 ,csa_tree_add_83_21_pad_groupi_n_1371 ,csa_tree_add_83_21_pad_groupi_n_1439);
  or csa_tree_add_83_21_pad_groupi_g4246__6131(csa_tree_add_83_21_pad_groupi_n_1480 ,csa_tree_add_83_21_pad_groupi_n_1424 ,csa_tree_add_83_21_pad_groupi_n_1456);
  and csa_tree_add_83_21_pad_groupi_g4247__1881(csa_tree_add_83_21_pad_groupi_n_1478 ,csa_tree_add_83_21_pad_groupi_n_1431 ,csa_tree_add_83_21_pad_groupi_n_1454);
  or csa_tree_add_83_21_pad_groupi_g4248__5115(csa_tree_add_83_21_pad_groupi_n_1476 ,csa_tree_add_83_21_pad_groupi_n_1422 ,csa_tree_add_83_21_pad_groupi_n_1455);
  or csa_tree_add_83_21_pad_groupi_g4249__7482(csa_tree_add_83_21_pad_groupi_n_1475 ,csa_tree_add_83_21_pad_groupi_n_1429 ,csa_tree_add_83_21_pad_groupi_n_1458);
  or csa_tree_add_83_21_pad_groupi_g4250__4733(csa_tree_add_83_21_pad_groupi_n_1472 ,csa_tree_add_83_21_pad_groupi_n_1426 ,csa_tree_add_83_21_pad_groupi_n_1457);
  not csa_tree_add_83_21_pad_groupi_g4251(csa_tree_add_83_21_pad_groupi_n_1469 ,csa_tree_add_83_21_pad_groupi_n_6);
  not csa_tree_add_83_21_pad_groupi_g4252(csa_tree_add_83_21_pad_groupi_n_1468 ,csa_tree_add_83_21_pad_groupi_n_1467);
  not csa_tree_add_83_21_pad_groupi_g4253(csa_tree_add_83_21_pad_groupi_n_1466 ,csa_tree_add_83_21_pad_groupi_n_1465);
  and csa_tree_add_83_21_pad_groupi_g4254__6161(csa_tree_add_83_21_pad_groupi_n_1464 ,csa_tree_add_83_21_pad_groupi_n_1440 ,csa_tree_add_83_21_pad_groupi_n_1446);
  nor csa_tree_add_83_21_pad_groupi_g4255__9315(csa_tree_add_83_21_pad_groupi_n_1463 ,csa_tree_add_83_21_pad_groupi_n_1440 ,csa_tree_add_83_21_pad_groupi_n_1446);
  xnor csa_tree_add_83_21_pad_groupi_g4256__9945(csa_tree_add_83_21_pad_groupi_n_1462 ,csa_tree_add_83_21_pad_groupi_n_1432 ,csa_tree_add_83_21_pad_groupi_n_1413);
  xnor csa_tree_add_83_21_pad_groupi_g4257__2883(csa_tree_add_83_21_pad_groupi_n_1461 ,csa_tree_add_83_21_pad_groupi_n_1397 ,csa_tree_add_83_21_pad_groupi_n_1417);
  xnor csa_tree_add_83_21_pad_groupi_g4258__2346(csa_tree_add_83_21_pad_groupi_n_1460 ,csa_tree_add_83_21_pad_groupi_n_1367 ,csa_tree_add_83_21_pad_groupi_n_1415);
  xnor csa_tree_add_83_21_pad_groupi_g4260__1666(csa_tree_add_83_21_pad_groupi_n_1467 ,csa_tree_add_83_21_pad_groupi_n_1384 ,csa_tree_add_83_21_pad_groupi_n_1405);
  xnor csa_tree_add_83_21_pad_groupi_g4261__7410(csa_tree_add_83_21_pad_groupi_n_1465 ,csa_tree_add_83_21_pad_groupi_n_1295 ,csa_tree_add_83_21_pad_groupi_n_5);
  or csa_tree_add_83_21_pad_groupi_g4262__6417(csa_tree_add_83_21_pad_groupi_n_1459 ,csa_tree_add_83_21_pad_groupi_n_1432 ,csa_tree_add_83_21_pad_groupi_n_1413);
  and csa_tree_add_83_21_pad_groupi_g4263__5477(csa_tree_add_83_21_pad_groupi_n_1458 ,csa_tree_add_83_21_pad_groupi_n_1401 ,csa_tree_add_83_21_pad_groupi_n_1427);
  and csa_tree_add_83_21_pad_groupi_g4264__2398(csa_tree_add_83_21_pad_groupi_n_1457 ,csa_tree_add_83_21_pad_groupi_n_1402 ,csa_tree_add_83_21_pad_groupi_n_1425);
  and csa_tree_add_83_21_pad_groupi_g4265__5107(csa_tree_add_83_21_pad_groupi_n_1456 ,csa_tree_add_83_21_pad_groupi_n_1387 ,csa_tree_add_83_21_pad_groupi_n_1423);
  and csa_tree_add_83_21_pad_groupi_g4266__6260(csa_tree_add_83_21_pad_groupi_n_1455 ,csa_tree_add_83_21_pad_groupi_n_1403 ,csa_tree_add_83_21_pad_groupi_n_1421);
  or csa_tree_add_83_21_pad_groupi_g4267__4319(csa_tree_add_83_21_pad_groupi_n_1454 ,csa_tree_add_83_21_pad_groupi_n_1430 ,csa_tree_add_83_21_pad_groupi_n_1386);
  and csa_tree_add_83_21_pad_groupi_g4268__8428(csa_tree_add_83_21_pad_groupi_n_1453 ,csa_tree_add_83_21_pad_groupi_n_1432 ,csa_tree_add_83_21_pad_groupi_n_1413);
  or csa_tree_add_83_21_pad_groupi_g4269__5526(csa_tree_add_83_21_pad_groupi_n_1452 ,csa_tree_add_83_21_pad_groupi_n_1396 ,csa_tree_add_83_21_pad_groupi_n_1416);
  nor csa_tree_add_83_21_pad_groupi_g4270__6783(csa_tree_add_83_21_pad_groupi_n_1451 ,csa_tree_add_83_21_pad_groupi_n_1397 ,csa_tree_add_83_21_pad_groupi_n_1417);
  or csa_tree_add_83_21_pad_groupi_g4271__3680(csa_tree_add_83_21_pad_groupi_n_1450 ,csa_tree_add_83_21_pad_groupi_n_1367 ,csa_tree_add_83_21_pad_groupi_n_1414);
  nor csa_tree_add_83_21_pad_groupi_g4272__1617(csa_tree_add_83_21_pad_groupi_n_1449 ,csa_tree_add_83_21_pad_groupi_n_1366 ,csa_tree_add_83_21_pad_groupi_n_1415);
  not csa_tree_add_83_21_pad_groupi_g4273(csa_tree_add_83_21_pad_groupi_n_1448 ,csa_tree_add_83_21_pad_groupi_n_1447);
  not csa_tree_add_83_21_pad_groupi_g4274(csa_tree_add_83_21_pad_groupi_n_1446 ,csa_tree_add_83_21_pad_groupi_n_1445);
  not csa_tree_add_83_21_pad_groupi_g4275(csa_tree_add_83_21_pad_groupi_n_1444 ,csa_tree_add_83_21_pad_groupi_n_1443);
  not csa_tree_add_83_21_pad_groupi_g4276(csa_tree_add_83_21_pad_groupi_n_1441 ,csa_tree_add_83_21_pad_groupi_n_1442);
  or csa_tree_add_83_21_pad_groupi_g4277__2802(csa_tree_add_83_21_pad_groupi_n_1439 ,csa_tree_add_83_21_pad_groupi_n_1372 ,csa_tree_add_83_21_pad_groupi_n_1428);
  xnor csa_tree_add_83_21_pad_groupi_g4278__1705(csa_tree_add_83_21_pad_groupi_n_1438 ,csa_tree_add_83_21_pad_groupi_n_1291 ,csa_tree_add_83_21_pad_groupi_n_1379);
  xnor csa_tree_add_83_21_pad_groupi_g4279__5122(csa_tree_add_83_21_pad_groupi_n_1437 ,csa_tree_add_83_21_pad_groupi_n_1293 ,csa_tree_add_83_21_pad_groupi_n_1381);
  xnor csa_tree_add_83_21_pad_groupi_g4280__8246(csa_tree_add_83_21_pad_groupi_n_1436 ,csa_tree_add_83_21_pad_groupi_n_1301 ,csa_tree_add_83_21_pad_groupi_n_1376);
  xnor csa_tree_add_83_21_pad_groupi_g4281__7098(csa_tree_add_83_21_pad_groupi_n_1435 ,csa_tree_add_83_21_pad_groupi_n_1303 ,csa_tree_add_83_21_pad_groupi_n_1383);
  xnor csa_tree_add_83_21_pad_groupi_g4282__6131(csa_tree_add_83_21_pad_groupi_n_1434 ,csa_tree_add_83_21_pad_groupi_n_1377 ,csa_tree_add_83_21_pad_groupi_n_1398);
  xnor csa_tree_add_83_21_pad_groupi_g4283__1881(csa_tree_add_83_21_pad_groupi_n_1433 ,csa_tree_add_83_21_pad_groupi_n_1298 ,csa_tree_add_83_21_pad_groupi_n_1386);
  or csa_tree_add_83_21_pad_groupi_g4284__5115(csa_tree_add_83_21_pad_groupi_n_1447 ,csa_tree_add_83_21_pad_groupi_n_1340 ,csa_tree_add_83_21_pad_groupi_n_1420);
  xnor csa_tree_add_83_21_pad_groupi_g4285__7482(csa_tree_add_83_21_pad_groupi_n_1445 ,csa_tree_add_83_21_pad_groupi_n_1334 ,csa_tree_add_83_21_pad_groupi_n_1370);
  xnor csa_tree_add_83_21_pad_groupi_g4286__4733(csa_tree_add_83_21_pad_groupi_n_1443 ,csa_tree_add_83_21_pad_groupi_n_1385 ,csa_tree_add_83_21_pad_groupi_n_1369);
  or csa_tree_add_83_21_pad_groupi_g4287__6161(csa_tree_add_83_21_pad_groupi_n_1442 ,csa_tree_add_83_21_pad_groupi_n_1374 ,csa_tree_add_83_21_pad_groupi_n_1409);
  and csa_tree_add_83_21_pad_groupi_g4288__9315(csa_tree_add_83_21_pad_groupi_n_1440 ,csa_tree_add_83_21_pad_groupi_n_1395 ,csa_tree_add_83_21_pad_groupi_n_1408);
  or csa_tree_add_83_21_pad_groupi_g4289__9945(csa_tree_add_83_21_pad_groupi_n_1431 ,csa_tree_add_83_21_pad_groupi_n_1297 ,csa_tree_add_83_21_pad_groupi_n_1399);
  nor csa_tree_add_83_21_pad_groupi_g4290__2883(csa_tree_add_83_21_pad_groupi_n_1430 ,csa_tree_add_83_21_pad_groupi_n_1298 ,csa_tree_add_83_21_pad_groupi_n_1400);
  nor csa_tree_add_83_21_pad_groupi_g4291__2346(csa_tree_add_83_21_pad_groupi_n_1429 ,csa_tree_add_83_21_pad_groupi_n_1300 ,csa_tree_add_83_21_pad_groupi_n_1376);
  nor csa_tree_add_83_21_pad_groupi_g4292__1666(csa_tree_add_83_21_pad_groupi_n_1428 ,csa_tree_add_83_21_pad_groupi_n_1363 ,csa_tree_add_83_21_pad_groupi_n_1394);
  or csa_tree_add_83_21_pad_groupi_g4293__7410(csa_tree_add_83_21_pad_groupi_n_1427 ,csa_tree_add_83_21_pad_groupi_n_1301 ,csa_tree_add_83_21_pad_groupi_n_1375);
  nor csa_tree_add_83_21_pad_groupi_g4294__6417(csa_tree_add_83_21_pad_groupi_n_1426 ,csa_tree_add_83_21_pad_groupi_n_1292 ,csa_tree_add_83_21_pad_groupi_n_1381);
  or csa_tree_add_83_21_pad_groupi_g4295__5477(csa_tree_add_83_21_pad_groupi_n_1425 ,csa_tree_add_83_21_pad_groupi_n_1293 ,csa_tree_add_83_21_pad_groupi_n_1380);
  nor csa_tree_add_83_21_pad_groupi_g4296__2398(csa_tree_add_83_21_pad_groupi_n_1424 ,csa_tree_add_83_21_pad_groupi_n_1290 ,csa_tree_add_83_21_pad_groupi_n_1379);
  or csa_tree_add_83_21_pad_groupi_g4297__5107(csa_tree_add_83_21_pad_groupi_n_1423 ,csa_tree_add_83_21_pad_groupi_n_1291 ,csa_tree_add_83_21_pad_groupi_n_1378);
  nor csa_tree_add_83_21_pad_groupi_g4298__6260(csa_tree_add_83_21_pad_groupi_n_1422 ,csa_tree_add_83_21_pad_groupi_n_1302 ,csa_tree_add_83_21_pad_groupi_n_1383);
  or csa_tree_add_83_21_pad_groupi_g4299__4319(csa_tree_add_83_21_pad_groupi_n_1421 ,csa_tree_add_83_21_pad_groupi_n_1303 ,csa_tree_add_83_21_pad_groupi_n_1382);
  nor csa_tree_add_83_21_pad_groupi_g4300__8428(csa_tree_add_83_21_pad_groupi_n_1420 ,csa_tree_add_83_21_pad_groupi_n_1355 ,csa_tree_add_83_21_pad_groupi_n_1385);
  or csa_tree_add_83_21_pad_groupi_g4301__5526(csa_tree_add_83_21_pad_groupi_n_1432 ,csa_tree_add_83_21_pad_groupi_n_1365 ,csa_tree_add_83_21_pad_groupi_n_1391);
  not csa_tree_add_83_21_pad_groupi_g4302(csa_tree_add_83_21_pad_groupi_n_1419 ,csa_tree_add_83_21_pad_groupi_n_1418);
  not csa_tree_add_83_21_pad_groupi_g4303(csa_tree_add_83_21_pad_groupi_n_1417 ,csa_tree_add_83_21_pad_groupi_n_1416);
  not csa_tree_add_83_21_pad_groupi_g4304(csa_tree_add_83_21_pad_groupi_n_1415 ,csa_tree_add_83_21_pad_groupi_n_1414);
  not csa_tree_add_83_21_pad_groupi_g4305(csa_tree_add_83_21_pad_groupi_n_1412 ,csa_tree_add_83_21_pad_groupi_n_1411);
  or csa_tree_add_83_21_pad_groupi_g4306__6783(csa_tree_add_83_21_pad_groupi_n_1410 ,csa_tree_add_83_21_pad_groupi_n_1377 ,csa_tree_add_83_21_pad_groupi_n_1398);
  nor csa_tree_add_83_21_pad_groupi_g4307__3680(csa_tree_add_83_21_pad_groupi_n_1409 ,csa_tree_add_83_21_pad_groupi_n_1384 ,csa_tree_add_83_21_pad_groupi_n_1392);
  or csa_tree_add_83_21_pad_groupi_g4308__1617(csa_tree_add_83_21_pad_groupi_n_1408 ,csa_tree_add_83_21_pad_groupi_n_1368 ,csa_tree_add_83_21_pad_groupi_n_1373);
  and csa_tree_add_83_21_pad_groupi_g4309__2802(csa_tree_add_83_21_pad_groupi_n_1407 ,csa_tree_add_83_21_pad_groupi_n_1377 ,csa_tree_add_83_21_pad_groupi_n_1398);
  xnor csa_tree_add_83_21_pad_groupi_g4310__1705(csa_tree_add_83_21_pad_groupi_n_1406 ,csa_tree_add_83_21_pad_groupi_n_1280 ,csa_tree_add_83_21_pad_groupi_n_1346);
  xnor csa_tree_add_83_21_pad_groupi_g4312__5122(csa_tree_add_83_21_pad_groupi_n_1405 ,csa_tree_add_83_21_pad_groupi_n_1304 ,csa_tree_add_83_21_pad_groupi_n_1348);
  xnor csa_tree_add_83_21_pad_groupi_g4313__8246(csa_tree_add_83_21_pad_groupi_n_1404 ,csa_tree_add_83_21_pad_groupi_n_1309 ,csa_tree_add_83_21_pad_groupi_n_1345);
  and csa_tree_add_83_21_pad_groupi_g4314__7098(csa_tree_add_83_21_pad_groupi_n_1418 ,csa_tree_add_83_21_pad_groupi_n_1354 ,csa_tree_add_83_21_pad_groupi_n_1390);
  xnor csa_tree_add_83_21_pad_groupi_g4315__6131(csa_tree_add_83_21_pad_groupi_n_1416 ,csa_tree_add_83_21_pad_groupi_n_1311 ,csa_tree_add_83_21_pad_groupi_n_1337);
  xnor csa_tree_add_83_21_pad_groupi_g4316__1881(csa_tree_add_83_21_pad_groupi_n_1414 ,csa_tree_add_83_21_pad_groupi_n_1320 ,csa_tree_add_83_21_pad_groupi_n_1335);
  xnor csa_tree_add_83_21_pad_groupi_g4317__5115(csa_tree_add_83_21_pad_groupi_n_1413 ,csa_tree_add_83_21_pad_groupi_n_1333 ,csa_tree_add_83_21_pad_groupi_n_1338);
  and csa_tree_add_83_21_pad_groupi_g4318__7482(csa_tree_add_83_21_pad_groupi_n_1411 ,csa_tree_add_83_21_pad_groupi_n_1356 ,csa_tree_add_83_21_pad_groupi_n_1388);
  not csa_tree_add_83_21_pad_groupi_g4319(csa_tree_add_83_21_pad_groupi_n_1400 ,csa_tree_add_83_21_pad_groupi_n_1399);
  not csa_tree_add_83_21_pad_groupi_g4320(csa_tree_add_83_21_pad_groupi_n_1396 ,csa_tree_add_83_21_pad_groupi_n_1397);
  or csa_tree_add_83_21_pad_groupi_g4321__4733(csa_tree_add_83_21_pad_groupi_n_1395 ,csa_tree_add_83_21_pad_groupi_n_1280 ,csa_tree_add_83_21_pad_groupi_n_1347);
  nor csa_tree_add_83_21_pad_groupi_g4322__6161(csa_tree_add_83_21_pad_groupi_n_1394 ,csa_tree_add_83_21_pad_groupi_n_1362 ,csa_tree_add_83_21_pad_groupi_n_1361);
  and csa_tree_add_83_21_pad_groupi_g4323__9315(csa_tree_add_83_21_pad_groupi_n_1393 ,csa_tree_add_83_21_pad_groupi_n_1309 ,csa_tree_add_83_21_pad_groupi_n_1345);
  and csa_tree_add_83_21_pad_groupi_g4324__9945(csa_tree_add_83_21_pad_groupi_n_1392 ,csa_tree_add_83_21_pad_groupi_n_1304 ,csa_tree_add_83_21_pad_groupi_n_1349);
  and csa_tree_add_83_21_pad_groupi_g4325__2883(csa_tree_add_83_21_pad_groupi_n_1391 ,csa_tree_add_83_21_pad_groupi_n_1334 ,csa_tree_add_83_21_pad_groupi_n_1360);
  or csa_tree_add_83_21_pad_groupi_g4326__2346(csa_tree_add_83_21_pad_groupi_n_1390 ,csa_tree_add_83_21_pad_groupi_n_1353 ,csa_tree_add_83_21_pad_groupi_n_1350);
  or csa_tree_add_83_21_pad_groupi_g4327__1666(csa_tree_add_83_21_pad_groupi_n_1389 ,csa_tree_add_83_21_pad_groupi_n_1309 ,csa_tree_add_83_21_pad_groupi_n_1345);
  or csa_tree_add_83_21_pad_groupi_g4328__7410(csa_tree_add_83_21_pad_groupi_n_1388 ,csa_tree_add_83_21_pad_groupi_n_1305 ,csa_tree_add_83_21_pad_groupi_n_1342);
  or csa_tree_add_83_21_pad_groupi_g4329__6417(csa_tree_add_83_21_pad_groupi_n_1403 ,csa_tree_add_83_21_pad_groupi_n_1246 ,csa_tree_add_83_21_pad_groupi_n_1359);
  or csa_tree_add_83_21_pad_groupi_g4330__5477(csa_tree_add_83_21_pad_groupi_n_1402 ,csa_tree_add_83_21_pad_groupi_n_1230 ,csa_tree_add_83_21_pad_groupi_n_1343);
  or csa_tree_add_83_21_pad_groupi_g4331__2398(csa_tree_add_83_21_pad_groupi_n_1401 ,csa_tree_add_83_21_pad_groupi_n_1232 ,csa_tree_add_83_21_pad_groupi_n_1339);
  and csa_tree_add_83_21_pad_groupi_g4332__5107(csa_tree_add_83_21_pad_groupi_n_1399 ,csa_tree_add_83_21_pad_groupi_n_1254 ,csa_tree_add_83_21_pad_groupi_n_1364);
  or csa_tree_add_83_21_pad_groupi_g4333__6260(csa_tree_add_83_21_pad_groupi_n_1398 ,csa_tree_add_83_21_pad_groupi_n_1329 ,csa_tree_add_83_21_pad_groupi_n_1357);
  or csa_tree_add_83_21_pad_groupi_g4334__4319(csa_tree_add_83_21_pad_groupi_n_1397 ,csa_tree_add_83_21_pad_groupi_n_1323 ,csa_tree_add_83_21_pad_groupi_n_1358);
  not csa_tree_add_83_21_pad_groupi_g4335(csa_tree_add_83_21_pad_groupi_n_1383 ,csa_tree_add_83_21_pad_groupi_n_1382);
  not csa_tree_add_83_21_pad_groupi_g4336(csa_tree_add_83_21_pad_groupi_n_1381 ,csa_tree_add_83_21_pad_groupi_n_1380);
  not csa_tree_add_83_21_pad_groupi_g4337(csa_tree_add_83_21_pad_groupi_n_1379 ,csa_tree_add_83_21_pad_groupi_n_1378);
  not csa_tree_add_83_21_pad_groupi_g4338(csa_tree_add_83_21_pad_groupi_n_1376 ,csa_tree_add_83_21_pad_groupi_n_1375);
  nor csa_tree_add_83_21_pad_groupi_g4339__8428(csa_tree_add_83_21_pad_groupi_n_1374 ,csa_tree_add_83_21_pad_groupi_n_1304 ,csa_tree_add_83_21_pad_groupi_n_1349);
  and csa_tree_add_83_21_pad_groupi_g4340__5526(csa_tree_add_83_21_pad_groupi_n_1373 ,csa_tree_add_83_21_pad_groupi_n_1280 ,csa_tree_add_83_21_pad_groupi_n_1347);
  nor csa_tree_add_83_21_pad_groupi_g4341__6783(csa_tree_add_83_21_pad_groupi_n_1372 ,csa_tree_add_83_21_pad_groupi_n_1306 ,csa_tree_add_83_21_pad_groupi_n_1352);
  or csa_tree_add_83_21_pad_groupi_g4342__3680(csa_tree_add_83_21_pad_groupi_n_1371 ,csa_tree_add_83_21_pad_groupi_n_1307 ,csa_tree_add_83_21_pad_groupi_n_1351);
  xnor csa_tree_add_83_21_pad_groupi_g4343__1617(csa_tree_add_83_21_pad_groupi_n_1370 ,csa_tree_add_83_21_pad_groupi_n_1261 ,csa_tree_add_83_21_pad_groupi_n_1310);
  xnor csa_tree_add_83_21_pad_groupi_g4344__2802(csa_tree_add_83_21_pad_groupi_n_1369 ,csa_tree_add_83_21_pad_groupi_n_1299 ,csa_tree_add_83_21_pad_groupi_n_1330);
  or csa_tree_add_83_21_pad_groupi_g4345__1705(csa_tree_add_83_21_pad_groupi_n_1387 ,csa_tree_add_83_21_pad_groupi_n_1227 ,csa_tree_add_83_21_pad_groupi_n_1341);
  xnor csa_tree_add_83_21_pad_groupi_g4346__5122(csa_tree_add_83_21_pad_groupi_n_1386 ,csa_tree_add_83_21_pad_groupi_n_1317 ,csa_tree_add_83_21_pad_groupi_n_1273);
  xnor csa_tree_add_83_21_pad_groupi_g4347__8246(csa_tree_add_83_21_pad_groupi_n_1385 ,csa_tree_add_83_21_pad_groupi_n_1316 ,csa_tree_add_83_21_pad_groupi_n_1268);
  and csa_tree_add_83_21_pad_groupi_g4348__7098(csa_tree_add_83_21_pad_groupi_n_1384 ,csa_tree_add_83_21_pad_groupi_n_1225 ,csa_tree_add_83_21_pad_groupi_n_1344);
  xnor csa_tree_add_83_21_pad_groupi_g4349__6131(csa_tree_add_83_21_pad_groupi_n_1382 ,csa_tree_add_83_21_pad_groupi_n_1313 ,csa_tree_add_83_21_pad_groupi_n_1266);
  xnor csa_tree_add_83_21_pad_groupi_g4350__1881(csa_tree_add_83_21_pad_groupi_n_1380 ,csa_tree_add_83_21_pad_groupi_n_1315 ,csa_tree_add_83_21_pad_groupi_n_1270);
  xnor csa_tree_add_83_21_pad_groupi_g4351__5115(csa_tree_add_83_21_pad_groupi_n_1378 ,csa_tree_add_83_21_pad_groupi_n_1314 ,csa_tree_add_83_21_pad_groupi_n_1267);
  xnor csa_tree_add_83_21_pad_groupi_g4352__7482(csa_tree_add_83_21_pad_groupi_n_1377 ,csa_tree_add_83_21_pad_groupi_n_1262 ,csa_tree_add_83_21_pad_groupi_n_1308);
  xnor csa_tree_add_83_21_pad_groupi_g4353__4733(csa_tree_add_83_21_pad_groupi_n_1375 ,csa_tree_add_83_21_pad_groupi_n_1318 ,csa_tree_add_83_21_pad_groupi_n_1271);
  not csa_tree_add_83_21_pad_groupi_g4355(csa_tree_add_83_21_pad_groupi_n_1367 ,csa_tree_add_83_21_pad_groupi_n_1366);
  and csa_tree_add_83_21_pad_groupi_g4356__6161(csa_tree_add_83_21_pad_groupi_n_1365 ,csa_tree_add_83_21_pad_groupi_n_1261 ,csa_tree_add_83_21_pad_groupi_n_1310);
  or csa_tree_add_83_21_pad_groupi_g4357__9315(csa_tree_add_83_21_pad_groupi_n_1364 ,csa_tree_add_83_21_pad_groupi_n_1224 ,csa_tree_add_83_21_pad_groupi_n_1319);
  and csa_tree_add_83_21_pad_groupi_g4358__9945(csa_tree_add_83_21_pad_groupi_n_1363 ,csa_tree_add_83_21_pad_groupi_n_1265 ,csa_tree_add_83_21_pad_groupi_n_1321);
  nor csa_tree_add_83_21_pad_groupi_g4359__2883(csa_tree_add_83_21_pad_groupi_n_1362 ,csa_tree_add_83_21_pad_groupi_n_1265 ,csa_tree_add_83_21_pad_groupi_n_1321);
  nor csa_tree_add_83_21_pad_groupi_g4360__2346(csa_tree_add_83_21_pad_groupi_n_1361 ,csa_tree_add_83_21_pad_groupi_n_1285 ,csa_tree_add_83_21_pad_groupi_n_1326);
  or csa_tree_add_83_21_pad_groupi_g4361__1666(csa_tree_add_83_21_pad_groupi_n_1360 ,csa_tree_add_83_21_pad_groupi_n_1261 ,csa_tree_add_83_21_pad_groupi_n_1310);
  nor csa_tree_add_83_21_pad_groupi_g4362__7410(csa_tree_add_83_21_pad_groupi_n_1359 ,csa_tree_add_83_21_pad_groupi_n_1245 ,csa_tree_add_83_21_pad_groupi_n_1316);
  nor csa_tree_add_83_21_pad_groupi_g4363__6417(csa_tree_add_83_21_pad_groupi_n_1358 ,csa_tree_add_83_21_pad_groupi_n_1328 ,csa_tree_add_83_21_pad_groupi_n_1320);
  nor csa_tree_add_83_21_pad_groupi_g4364__5477(csa_tree_add_83_21_pad_groupi_n_1357 ,csa_tree_add_83_21_pad_groupi_n_1333 ,csa_tree_add_83_21_pad_groupi_n_1322);
  or csa_tree_add_83_21_pad_groupi_g4365__2398(csa_tree_add_83_21_pad_groupi_n_1356 ,csa_tree_add_83_21_pad_groupi_n_1278 ,csa_tree_add_83_21_pad_groupi_n_1312);
  nor csa_tree_add_83_21_pad_groupi_g4366__5107(csa_tree_add_83_21_pad_groupi_n_1355 ,csa_tree_add_83_21_pad_groupi_n_1299 ,csa_tree_add_83_21_pad_groupi_n_1330);
  or csa_tree_add_83_21_pad_groupi_g4367__6260(csa_tree_add_83_21_pad_groupi_n_1354 ,csa_tree_add_83_21_pad_groupi_n_1294 ,csa_tree_add_83_21_pad_groupi_n_1332);
  nor csa_tree_add_83_21_pad_groupi_g4368__4319(csa_tree_add_83_21_pad_groupi_n_1353 ,csa_tree_add_83_21_pad_groupi_n_1295 ,csa_tree_add_83_21_pad_groupi_n_1331);
  and csa_tree_add_83_21_pad_groupi_g4369__8428(csa_tree_add_83_21_pad_groupi_n_1368 ,csa_tree_add_83_21_pad_groupi_n_1243 ,csa_tree_add_83_21_pad_groupi_n_1324);
  or csa_tree_add_83_21_pad_groupi_g4370__5526(csa_tree_add_83_21_pad_groupi_n_1366 ,csa_tree_add_83_21_pad_groupi_n_1185 ,csa_tree_add_83_21_pad_groupi_n_1327);
  not csa_tree_add_83_21_pad_groupi_g4371(csa_tree_add_83_21_pad_groupi_n_1352 ,csa_tree_add_83_21_pad_groupi_n_1351);
  not csa_tree_add_83_21_pad_groupi_g4373(csa_tree_add_83_21_pad_groupi_n_1349 ,csa_tree_add_83_21_pad_groupi_n_1348);
  not csa_tree_add_83_21_pad_groupi_g4374(csa_tree_add_83_21_pad_groupi_n_1347 ,csa_tree_add_83_21_pad_groupi_n_1346);
  or csa_tree_add_83_21_pad_groupi_g4375__6783(csa_tree_add_83_21_pad_groupi_n_1344 ,csa_tree_add_83_21_pad_groupi_n_1223 ,csa_tree_add_83_21_pad_groupi_n_1317);
  and csa_tree_add_83_21_pad_groupi_g4376__3680(csa_tree_add_83_21_pad_groupi_n_1343 ,csa_tree_add_83_21_pad_groupi_n_1228 ,csa_tree_add_83_21_pad_groupi_n_1314);
  and csa_tree_add_83_21_pad_groupi_g4377__1617(csa_tree_add_83_21_pad_groupi_n_1342 ,csa_tree_add_83_21_pad_groupi_n_1278 ,csa_tree_add_83_21_pad_groupi_n_1312);
  and csa_tree_add_83_21_pad_groupi_g4378__2802(csa_tree_add_83_21_pad_groupi_n_1341 ,csa_tree_add_83_21_pad_groupi_n_1226 ,csa_tree_add_83_21_pad_groupi_n_1313);
  and csa_tree_add_83_21_pad_groupi_g4379__1705(csa_tree_add_83_21_pad_groupi_n_1340 ,csa_tree_add_83_21_pad_groupi_n_1299 ,csa_tree_add_83_21_pad_groupi_n_1330);
  and csa_tree_add_83_21_pad_groupi_g4380__5122(csa_tree_add_83_21_pad_groupi_n_1339 ,csa_tree_add_83_21_pad_groupi_n_1231 ,csa_tree_add_83_21_pad_groupi_n_1315);
  xnor csa_tree_add_83_21_pad_groupi_g4381__8246(csa_tree_add_83_21_pad_groupi_n_1338 ,csa_tree_add_83_21_pad_groupi_n_1201 ,csa_tree_add_83_21_pad_groupi_n_1279);
  xnor csa_tree_add_83_21_pad_groupi_g4382__7098(csa_tree_add_83_21_pad_groupi_n_1351 ,csa_tree_add_83_21_pad_groupi_n_1281 ,csa_tree_add_83_21_pad_groupi_n_1211);
  xor csa_tree_add_83_21_pad_groupi_g4383__6131(csa_tree_add_83_21_pad_groupi_n_1337 ,csa_tree_add_83_21_pad_groupi_n_1278 ,csa_tree_add_83_21_pad_groupi_n_1305);
  xnor csa_tree_add_83_21_pad_groupi_g4384__1881(csa_tree_add_83_21_pad_groupi_n_1336 ,csa_tree_add_83_21_pad_groupi_n_1075 ,csa_tree_add_83_21_pad_groupi_n_1274);
  xnor csa_tree_add_83_21_pad_groupi_g4385__5115(csa_tree_add_83_21_pad_groupi_n_1335 ,csa_tree_add_83_21_pad_groupi_n_1235 ,csa_tree_add_83_21_pad_groupi_n_1296);
  xnor csa_tree_add_83_21_pad_groupi_g4386__7482(csa_tree_add_83_21_pad_groupi_n_1350 ,csa_tree_add_83_21_pad_groupi_n_1264 ,csa_tree_add_83_21_pad_groupi_n_1272);
  xnor csa_tree_add_83_21_pad_groupi_g4387__4733(csa_tree_add_83_21_pad_groupi_n_1348 ,csa_tree_add_83_21_pad_groupi_n_1282 ,csa_tree_add_83_21_pad_groupi_n_1269);
  xnor csa_tree_add_83_21_pad_groupi_g4388__6161(csa_tree_add_83_21_pad_groupi_n_1346 ,csa_tree_add_83_21_pad_groupi_n_1263 ,csa_tree_add_83_21_pad_groupi_n_1275);
  or csa_tree_add_83_21_pad_groupi_g4389__9315(csa_tree_add_83_21_pad_groupi_n_1345 ,csa_tree_add_83_21_pad_groupi_n_1277 ,csa_tree_add_83_21_pad_groupi_n_1325);
  not csa_tree_add_83_21_pad_groupi_g4390(csa_tree_add_83_21_pad_groupi_n_1332 ,csa_tree_add_83_21_pad_groupi_n_1331);
  nor csa_tree_add_83_21_pad_groupi_g4391__9945(csa_tree_add_83_21_pad_groupi_n_1329 ,csa_tree_add_83_21_pad_groupi_n_1202 ,csa_tree_add_83_21_pad_groupi_n_1279);
  nor csa_tree_add_83_21_pad_groupi_g4392__2883(csa_tree_add_83_21_pad_groupi_n_1328 ,csa_tree_add_83_21_pad_groupi_n_1235 ,csa_tree_add_83_21_pad_groupi_n_1296);
  nor csa_tree_add_83_21_pad_groupi_g4393__2346(csa_tree_add_83_21_pad_groupi_n_1327 ,csa_tree_add_83_21_pad_groupi_n_1184 ,csa_tree_add_83_21_pad_groupi_n_1281);
  nor csa_tree_add_83_21_pad_groupi_g4394__1666(csa_tree_add_83_21_pad_groupi_n_1326 ,csa_tree_add_83_21_pad_groupi_n_1287 ,csa_tree_add_83_21_pad_groupi_n_1288);
  nor csa_tree_add_83_21_pad_groupi_g4395__7410(csa_tree_add_83_21_pad_groupi_n_1325 ,csa_tree_add_83_21_pad_groupi_n_1276 ,csa_tree_add_83_21_pad_groupi_n_1262);
  or csa_tree_add_83_21_pad_groupi_g4396__6417(csa_tree_add_83_21_pad_groupi_n_1324 ,csa_tree_add_83_21_pad_groupi_n_1252 ,csa_tree_add_83_21_pad_groupi_n_1283);
  and csa_tree_add_83_21_pad_groupi_g4397__5477(csa_tree_add_83_21_pad_groupi_n_1323 ,csa_tree_add_83_21_pad_groupi_n_1235 ,csa_tree_add_83_21_pad_groupi_n_1296);
  and csa_tree_add_83_21_pad_groupi_g4398__2398(csa_tree_add_83_21_pad_groupi_n_1322 ,csa_tree_add_83_21_pad_groupi_n_1202 ,csa_tree_add_83_21_pad_groupi_n_1279);
  or csa_tree_add_83_21_pad_groupi_g4399__5107(csa_tree_add_83_21_pad_groupi_n_1334 ,csa_tree_add_83_21_pad_groupi_n_1240 ,csa_tree_add_83_21_pad_groupi_n_1284);
  and csa_tree_add_83_21_pad_groupi_g4400__6260(csa_tree_add_83_21_pad_groupi_n_1333 ,csa_tree_add_83_21_pad_groupi_n_1156 ,csa_tree_add_83_21_pad_groupi_n_1286);
  xnor csa_tree_add_83_21_pad_groupi_g4401__4319(csa_tree_add_83_21_pad_groupi_n_1331 ,csa_tree_add_83_21_pad_groupi_n_1039 ,csa_tree_add_83_21_pad_groupi_n_1216);
  or csa_tree_add_83_21_pad_groupi_g4402__8428(csa_tree_add_83_21_pad_groupi_n_1330 ,csa_tree_add_83_21_pad_groupi_n_1242 ,csa_tree_add_83_21_pad_groupi_n_1289);
  not csa_tree_add_83_21_pad_groupi_g4403(csa_tree_add_83_21_pad_groupi_n_1319 ,csa_tree_add_83_21_pad_groupi_n_1318);
  not csa_tree_add_83_21_pad_groupi_g4404(csa_tree_add_83_21_pad_groupi_n_1312 ,csa_tree_add_83_21_pad_groupi_n_1311);
  xnor csa_tree_add_83_21_pad_groupi_g4405__5526(csa_tree_add_83_21_pad_groupi_n_1321 ,csa_tree_add_83_21_pad_groupi_n_1176 ,csa_tree_add_83_21_pad_groupi_n_1210);
  xnor csa_tree_add_83_21_pad_groupi_g4406__6783(csa_tree_add_83_21_pad_groupi_n_1308 ,csa_tree_add_83_21_pad_groupi_n_1132 ,csa_tree_add_83_21_pad_groupi_n_1233);
  xnor csa_tree_add_83_21_pad_groupi_g4407__3680(csa_tree_add_83_21_pad_groupi_n_1320 ,csa_tree_add_83_21_pad_groupi_n_1084 ,csa_tree_add_83_21_pad_groupi_n_1220);
  xnor csa_tree_add_83_21_pad_groupi_g4408__1617(csa_tree_add_83_21_pad_groupi_n_1318 ,csa_tree_add_83_21_pad_groupi_n_1138 ,csa_tree_add_83_21_pad_groupi_n_1221);
  xnor csa_tree_add_83_21_pad_groupi_g4409__2802(csa_tree_add_83_21_pad_groupi_n_1317 ,csa_tree_add_83_21_pad_groupi_n_1092 ,csa_tree_add_83_21_pad_groupi_n_1213);
  xnor csa_tree_add_83_21_pad_groupi_g4410__1705(csa_tree_add_83_21_pad_groupi_n_1316 ,csa_tree_add_83_21_pad_groupi_n_1088 ,csa_tree_add_83_21_pad_groupi_n_1214);
  xnor csa_tree_add_83_21_pad_groupi_g4411__5122(csa_tree_add_83_21_pad_groupi_n_1315 ,csa_tree_add_83_21_pad_groupi_n_1141 ,csa_tree_add_83_21_pad_groupi_n_1218);
  xnor csa_tree_add_83_21_pad_groupi_g4412__8246(csa_tree_add_83_21_pad_groupi_n_1314 ,csa_tree_add_83_21_pad_groupi_n_1102 ,csa_tree_add_83_21_pad_groupi_n_1217);
  xnor csa_tree_add_83_21_pad_groupi_g4413__7098(csa_tree_add_83_21_pad_groupi_n_1313 ,csa_tree_add_83_21_pad_groupi_n_1107 ,csa_tree_add_83_21_pad_groupi_n_1222);
  xnor csa_tree_add_83_21_pad_groupi_g4414__6131(csa_tree_add_83_21_pad_groupi_n_1311 ,csa_tree_add_83_21_pad_groupi_n_1209 ,csa_tree_add_83_21_pad_groupi_n_1215);
  xnor csa_tree_add_83_21_pad_groupi_g4415__1881(csa_tree_add_83_21_pad_groupi_n_1310 ,csa_tree_add_83_21_pad_groupi_n_1236 ,csa_tree_add_83_21_pad_groupi_n_1212);
  xnor csa_tree_add_83_21_pad_groupi_g4416__5115(csa_tree_add_83_21_pad_groupi_n_1309 ,csa_tree_add_83_21_pad_groupi_n_1175 ,csa_tree_add_83_21_pad_groupi_n_1219);
  not csa_tree_add_83_21_pad_groupi_g4417(csa_tree_add_83_21_pad_groupi_n_1307 ,csa_tree_add_83_21_pad_groupi_n_1306);
  not csa_tree_add_83_21_pad_groupi_g4418(csa_tree_add_83_21_pad_groupi_n_1302 ,csa_tree_add_83_21_pad_groupi_n_1303);
  not csa_tree_add_83_21_pad_groupi_g4419(csa_tree_add_83_21_pad_groupi_n_1300 ,csa_tree_add_83_21_pad_groupi_n_1301);
  not csa_tree_add_83_21_pad_groupi_g4420(csa_tree_add_83_21_pad_groupi_n_1297 ,csa_tree_add_83_21_pad_groupi_n_1298);
  not csa_tree_add_83_21_pad_groupi_g4421(csa_tree_add_83_21_pad_groupi_n_1295 ,csa_tree_add_83_21_pad_groupi_n_1294);
  not csa_tree_add_83_21_pad_groupi_g4422(csa_tree_add_83_21_pad_groupi_n_1292 ,csa_tree_add_83_21_pad_groupi_n_1293);
  not csa_tree_add_83_21_pad_groupi_g4423(csa_tree_add_83_21_pad_groupi_n_1290 ,csa_tree_add_83_21_pad_groupi_n_1291);
  nor csa_tree_add_83_21_pad_groupi_g4424__7482(csa_tree_add_83_21_pad_groupi_n_1289 ,csa_tree_add_83_21_pad_groupi_n_1247 ,csa_tree_add_83_21_pad_groupi_n_1264);
  nor csa_tree_add_83_21_pad_groupi_g4425__4733(csa_tree_add_83_21_pad_groupi_n_1288 ,csa_tree_add_83_21_pad_groupi_n_1048 ,csa_tree_add_83_21_pad_groupi_n_1238);
  nor csa_tree_add_83_21_pad_groupi_g4426__6161(csa_tree_add_83_21_pad_groupi_n_1287 ,csa_tree_add_83_21_pad_groupi_n_1178 ,csa_tree_add_83_21_pad_groupi_n_1251);
  or csa_tree_add_83_21_pad_groupi_g4427__9315(csa_tree_add_83_21_pad_groupi_n_1286 ,csa_tree_add_83_21_pad_groupi_n_1150 ,csa_tree_add_83_21_pad_groupi_n_1237);
  nor csa_tree_add_83_21_pad_groupi_g4428__9945(csa_tree_add_83_21_pad_groupi_n_1285 ,csa_tree_add_83_21_pad_groupi_n_1047 ,csa_tree_add_83_21_pad_groupi_n_1239);
  and csa_tree_add_83_21_pad_groupi_g4429__2883(csa_tree_add_83_21_pad_groupi_n_1284 ,csa_tree_add_83_21_pad_groupi_n_1241 ,csa_tree_add_83_21_pad_groupi_n_1263);
  or csa_tree_add_83_21_pad_groupi_g4430__2346(csa_tree_add_83_21_pad_groupi_n_1306 ,csa_tree_add_83_21_pad_groupi_n_1183 ,csa_tree_add_83_21_pad_groupi_n_1253);
  and csa_tree_add_83_21_pad_groupi_g4431__1666(csa_tree_add_83_21_pad_groupi_n_1305 ,csa_tree_add_83_21_pad_groupi_n_1192 ,csa_tree_add_83_21_pad_groupi_n_1257);
  and csa_tree_add_83_21_pad_groupi_g4432__7410(csa_tree_add_83_21_pad_groupi_n_1304 ,csa_tree_add_83_21_pad_groupi_n_1155 ,csa_tree_add_83_21_pad_groupi_n_1260);
  or csa_tree_add_83_21_pad_groupi_g4433__6417(csa_tree_add_83_21_pad_groupi_n_1303 ,csa_tree_add_83_21_pad_groupi_n_1154 ,csa_tree_add_83_21_pad_groupi_n_1248);
  or csa_tree_add_83_21_pad_groupi_g4434__5477(csa_tree_add_83_21_pad_groupi_n_1301 ,csa_tree_add_83_21_pad_groupi_n_1187 ,csa_tree_add_83_21_pad_groupi_n_1255);
  or csa_tree_add_83_21_pad_groupi_g4435__2398(csa_tree_add_83_21_pad_groupi_n_1299 ,csa_tree_add_83_21_pad_groupi_n_1147 ,csa_tree_add_83_21_pad_groupi_n_1244);
  or csa_tree_add_83_21_pad_groupi_g4436__5107(csa_tree_add_83_21_pad_groupi_n_1298 ,csa_tree_add_83_21_pad_groupi_n_1198 ,csa_tree_add_83_21_pad_groupi_n_1258);
  or csa_tree_add_83_21_pad_groupi_g4437__6260(csa_tree_add_83_21_pad_groupi_n_1296 ,csa_tree_add_83_21_pad_groupi_n_1188 ,csa_tree_add_83_21_pad_groupi_n_1256);
  and csa_tree_add_83_21_pad_groupi_g4438__4319(csa_tree_add_83_21_pad_groupi_n_1294 ,csa_tree_add_83_21_pad_groupi_n_1197 ,csa_tree_add_83_21_pad_groupi_n_1259);
  or csa_tree_add_83_21_pad_groupi_g4439__8428(csa_tree_add_83_21_pad_groupi_n_1293 ,csa_tree_add_83_21_pad_groupi_n_1179 ,csa_tree_add_83_21_pad_groupi_n_1250);
  or csa_tree_add_83_21_pad_groupi_g4440__5526(csa_tree_add_83_21_pad_groupi_n_1291 ,csa_tree_add_83_21_pad_groupi_n_1200 ,csa_tree_add_83_21_pad_groupi_n_1249);
  not csa_tree_add_83_21_pad_groupi_g4441(csa_tree_add_83_21_pad_groupi_n_1283 ,csa_tree_add_83_21_pad_groupi_n_1282);
  nor csa_tree_add_83_21_pad_groupi_g4442__6783(csa_tree_add_83_21_pad_groupi_n_1277 ,csa_tree_add_83_21_pad_groupi_n_1132 ,csa_tree_add_83_21_pad_groupi_n_1234);
  and csa_tree_add_83_21_pad_groupi_g4443__3680(csa_tree_add_83_21_pad_groupi_n_1276 ,csa_tree_add_83_21_pad_groupi_n_1132 ,csa_tree_add_83_21_pad_groupi_n_1234);
  xnor csa_tree_add_83_21_pad_groupi_g4444__1617(csa_tree_add_83_21_pad_groupi_n_1275 ,csa_tree_add_83_21_pad_groupi_n_1207 ,csa_tree_add_83_21_pad_groupi_n_1098);
  nor csa_tree_add_83_21_pad_groupi_g4445__2802(csa_tree_add_83_21_pad_groupi_n_1274 ,csa_tree_add_83_21_pad_groupi_n_1157 ,csa_tree_add_83_21_pad_groupi_n_1229);
  xnor csa_tree_add_83_21_pad_groupi_g4446__1705(csa_tree_add_83_21_pad_groupi_n_1273 ,csa_tree_add_83_21_pad_groupi_n_1163 ,csa_tree_add_83_21_pad_groupi_n_1166);
  xnor csa_tree_add_83_21_pad_groupi_g4447__5122(csa_tree_add_83_21_pad_groupi_n_1272 ,csa_tree_add_83_21_pad_groupi_n_1099 ,csa_tree_add_83_21_pad_groupi_n_1169);
  xnor csa_tree_add_83_21_pad_groupi_g4448__8246(csa_tree_add_83_21_pad_groupi_n_1271 ,csa_tree_add_83_21_pad_groupi_n_1204 ,csa_tree_add_83_21_pad_groupi_n_1160);
  xnor csa_tree_add_83_21_pad_groupi_g4449__7098(csa_tree_add_83_21_pad_groupi_n_1270 ,csa_tree_add_83_21_pad_groupi_n_1208 ,csa_tree_add_83_21_pad_groupi_n_1174);
  xnor csa_tree_add_83_21_pad_groupi_g4450__6131(csa_tree_add_83_21_pad_groupi_n_1269 ,csa_tree_add_83_21_pad_groupi_n_1206 ,csa_tree_add_83_21_pad_groupi_n_1171);
  xnor csa_tree_add_83_21_pad_groupi_g4451__1881(csa_tree_add_83_21_pad_groupi_n_1268 ,csa_tree_add_83_21_pad_groupi_n_1164 ,csa_tree_add_83_21_pad_groupi_n_1167);
  xnor csa_tree_add_83_21_pad_groupi_g4452__5115(csa_tree_add_83_21_pad_groupi_n_1267 ,csa_tree_add_83_21_pad_groupi_n_1173 ,csa_tree_add_83_21_pad_groupi_n_1172);
  xnor csa_tree_add_83_21_pad_groupi_g4453__7482(csa_tree_add_83_21_pad_groupi_n_1266 ,csa_tree_add_83_21_pad_groupi_n_1161 ,csa_tree_add_83_21_pad_groupi_n_1168);
  xnor csa_tree_add_83_21_pad_groupi_g4454__4733(csa_tree_add_83_21_pad_groupi_n_1282 ,csa_tree_add_83_21_pad_groupi_n_1106 ,csa_tree_add_83_21_pad_groupi_n_1143);
  xnor csa_tree_add_83_21_pad_groupi_g4455__6161(csa_tree_add_83_21_pad_groupi_n_1281 ,csa_tree_add_83_21_pad_groupi_n_1080 ,csa_tree_add_83_21_pad_groupi_n_1145);
  xnor csa_tree_add_83_21_pad_groupi_g4456__9315(csa_tree_add_83_21_pad_groupi_n_1280 ,csa_tree_add_83_21_pad_groupi_n_1103 ,csa_tree_add_83_21_pad_groupi_n_1146);
  xnor csa_tree_add_83_21_pad_groupi_g4457__9945(csa_tree_add_83_21_pad_groupi_n_1279 ,csa_tree_add_83_21_pad_groupi_n_1101 ,csa_tree_add_83_21_pad_groupi_n_1142);
  xnor csa_tree_add_83_21_pad_groupi_g4458__2883(csa_tree_add_83_21_pad_groupi_n_1278 ,csa_tree_add_83_21_pad_groupi_n_1105 ,csa_tree_add_83_21_pad_groupi_n_1144);
  or csa_tree_add_83_21_pad_groupi_g4459__2346(csa_tree_add_83_21_pad_groupi_n_1260 ,csa_tree_add_83_21_pad_groupi_n_1104 ,csa_tree_add_83_21_pad_groupi_n_1151);
  or csa_tree_add_83_21_pad_groupi_g4460__1666(csa_tree_add_83_21_pad_groupi_n_1259 ,csa_tree_add_83_21_pad_groupi_n_1209 ,csa_tree_add_83_21_pad_groupi_n_1193);
  nor csa_tree_add_83_21_pad_groupi_g4461__7410(csa_tree_add_83_21_pad_groupi_n_1258 ,csa_tree_add_83_21_pad_groupi_n_1074 ,csa_tree_add_83_21_pad_groupi_n_1195);
  or csa_tree_add_83_21_pad_groupi_g4462__6417(csa_tree_add_83_21_pad_groupi_n_1257 ,csa_tree_add_83_21_pad_groupi_n_1072 ,csa_tree_add_83_21_pad_groupi_n_1190);
  nor csa_tree_add_83_21_pad_groupi_g4463__5477(csa_tree_add_83_21_pad_groupi_n_1256 ,csa_tree_add_83_21_pad_groupi_n_1067 ,csa_tree_add_83_21_pad_groupi_n_1186);
  and csa_tree_add_83_21_pad_groupi_g4464__2398(csa_tree_add_83_21_pad_groupi_n_1255 ,csa_tree_add_83_21_pad_groupi_n_1141 ,csa_tree_add_83_21_pad_groupi_n_1189);
  or csa_tree_add_83_21_pad_groupi_g4465__5107(csa_tree_add_83_21_pad_groupi_n_1254 ,csa_tree_add_83_21_pad_groupi_n_1203 ,csa_tree_add_83_21_pad_groupi_n_1159);
  and csa_tree_add_83_21_pad_groupi_g4466__6260(csa_tree_add_83_21_pad_groupi_n_1253 ,csa_tree_add_83_21_pad_groupi_n_1181 ,csa_tree_add_83_21_pad_groupi_n_1176);
  nor csa_tree_add_83_21_pad_groupi_g4467__4319(csa_tree_add_83_21_pad_groupi_n_1252 ,csa_tree_add_83_21_pad_groupi_n_1206 ,csa_tree_add_83_21_pad_groupi_n_1171);
  nor csa_tree_add_83_21_pad_groupi_g4468__8428(csa_tree_add_83_21_pad_groupi_n_1251 ,csa_tree_add_83_21_pad_groupi_n_1177 ,csa_tree_add_83_21_pad_groupi_n_1191);
  and csa_tree_add_83_21_pad_groupi_g4469__5526(csa_tree_add_83_21_pad_groupi_n_1250 ,csa_tree_add_83_21_pad_groupi_n_1102 ,csa_tree_add_83_21_pad_groupi_n_1194);
  and csa_tree_add_83_21_pad_groupi_g4470__6783(csa_tree_add_83_21_pad_groupi_n_1249 ,csa_tree_add_83_21_pad_groupi_n_1107 ,csa_tree_add_83_21_pad_groupi_n_1158);
  nor csa_tree_add_83_21_pad_groupi_g4471__3680(csa_tree_add_83_21_pad_groupi_n_1248 ,csa_tree_add_83_21_pad_groupi_n_1042 ,csa_tree_add_83_21_pad_groupi_n_1153);
  nor csa_tree_add_83_21_pad_groupi_g4472__1617(csa_tree_add_83_21_pad_groupi_n_1247 ,csa_tree_add_83_21_pad_groupi_n_1099 ,csa_tree_add_83_21_pad_groupi_n_1169);
  and csa_tree_add_83_21_pad_groupi_g4473__2802(csa_tree_add_83_21_pad_groupi_n_1246 ,csa_tree_add_83_21_pad_groupi_n_1164 ,csa_tree_add_83_21_pad_groupi_n_1167);
  nor csa_tree_add_83_21_pad_groupi_g4474__1705(csa_tree_add_83_21_pad_groupi_n_1245 ,csa_tree_add_83_21_pad_groupi_n_1164 ,csa_tree_add_83_21_pad_groupi_n_1167);
  nor csa_tree_add_83_21_pad_groupi_g4475__5122(csa_tree_add_83_21_pad_groupi_n_1244 ,csa_tree_add_83_21_pad_groupi_n_1039 ,csa_tree_add_83_21_pad_groupi_n_1148);
  or csa_tree_add_83_21_pad_groupi_g4476__8246(csa_tree_add_83_21_pad_groupi_n_1243 ,csa_tree_add_83_21_pad_groupi_n_1205 ,csa_tree_add_83_21_pad_groupi_n_1170);
  and csa_tree_add_83_21_pad_groupi_g4477__7098(csa_tree_add_83_21_pad_groupi_n_1242 ,csa_tree_add_83_21_pad_groupi_n_1099 ,csa_tree_add_83_21_pad_groupi_n_1169);
  or csa_tree_add_83_21_pad_groupi_g4478__6131(csa_tree_add_83_21_pad_groupi_n_1241 ,csa_tree_add_83_21_pad_groupi_n_1207 ,csa_tree_add_83_21_pad_groupi_n_1098);
  and csa_tree_add_83_21_pad_groupi_g4479__1881(csa_tree_add_83_21_pad_groupi_n_1240 ,csa_tree_add_83_21_pad_groupi_n_1207 ,csa_tree_add_83_21_pad_groupi_n_1098);
  or csa_tree_add_83_21_pad_groupi_g4480__5115(csa_tree_add_83_21_pad_groupi_n_1265 ,csa_tree_add_83_21_pad_groupi_n_1051 ,csa_tree_add_83_21_pad_groupi_n_1180);
  and csa_tree_add_83_21_pad_groupi_g4481__7482(csa_tree_add_83_21_pad_groupi_n_1264 ,csa_tree_add_83_21_pad_groupi_n_1115 ,csa_tree_add_83_21_pad_groupi_n_1199);
  or csa_tree_add_83_21_pad_groupi_g4482__4733(csa_tree_add_83_21_pad_groupi_n_1263 ,csa_tree_add_83_21_pad_groupi_n_1123 ,csa_tree_add_83_21_pad_groupi_n_1182);
  and csa_tree_add_83_21_pad_groupi_g4483__6161(csa_tree_add_83_21_pad_groupi_n_1262 ,csa_tree_add_83_21_pad_groupi_n_1114 ,csa_tree_add_83_21_pad_groupi_n_1149);
  or csa_tree_add_83_21_pad_groupi_g4484__9315(csa_tree_add_83_21_pad_groupi_n_1261 ,csa_tree_add_83_21_pad_groupi_n_1124 ,csa_tree_add_83_21_pad_groupi_n_1196);
  not csa_tree_add_83_21_pad_groupi_g4485(csa_tree_add_83_21_pad_groupi_n_1239 ,csa_tree_add_83_21_pad_groupi_n_1238);
  not csa_tree_add_83_21_pad_groupi_g4486(csa_tree_add_83_21_pad_groupi_n_1237 ,csa_tree_add_83_21_pad_groupi_n_1236);
  not csa_tree_add_83_21_pad_groupi_g4487(csa_tree_add_83_21_pad_groupi_n_1234 ,csa_tree_add_83_21_pad_groupi_n_1233);
  and csa_tree_add_83_21_pad_groupi_g4488__9945(csa_tree_add_83_21_pad_groupi_n_1232 ,csa_tree_add_83_21_pad_groupi_n_1208 ,csa_tree_add_83_21_pad_groupi_n_1174);
  or csa_tree_add_83_21_pad_groupi_g4489__2883(csa_tree_add_83_21_pad_groupi_n_1231 ,csa_tree_add_83_21_pad_groupi_n_1208 ,csa_tree_add_83_21_pad_groupi_n_1174);
  and csa_tree_add_83_21_pad_groupi_g4490__2346(csa_tree_add_83_21_pad_groupi_n_1230 ,csa_tree_add_83_21_pad_groupi_n_1173 ,csa_tree_add_83_21_pad_groupi_n_1172);
  nor csa_tree_add_83_21_pad_groupi_g4491__1666(csa_tree_add_83_21_pad_groupi_n_1229 ,csa_tree_add_83_21_pad_groupi_n_1152 ,csa_tree_add_83_21_pad_groupi_n_1175);
  or csa_tree_add_83_21_pad_groupi_g4492__7410(csa_tree_add_83_21_pad_groupi_n_1228 ,csa_tree_add_83_21_pad_groupi_n_1173 ,csa_tree_add_83_21_pad_groupi_n_1172);
  and csa_tree_add_83_21_pad_groupi_g4493__6417(csa_tree_add_83_21_pad_groupi_n_1227 ,csa_tree_add_83_21_pad_groupi_n_1161 ,csa_tree_add_83_21_pad_groupi_n_1168);
  or csa_tree_add_83_21_pad_groupi_g4494__5477(csa_tree_add_83_21_pad_groupi_n_1226 ,csa_tree_add_83_21_pad_groupi_n_1161 ,csa_tree_add_83_21_pad_groupi_n_1168);
  or csa_tree_add_83_21_pad_groupi_g4495__2398(csa_tree_add_83_21_pad_groupi_n_1225 ,csa_tree_add_83_21_pad_groupi_n_1162 ,csa_tree_add_83_21_pad_groupi_n_1165);
  nor csa_tree_add_83_21_pad_groupi_g4496__5107(csa_tree_add_83_21_pad_groupi_n_1224 ,csa_tree_add_83_21_pad_groupi_n_1204 ,csa_tree_add_83_21_pad_groupi_n_1160);
  nor csa_tree_add_83_21_pad_groupi_g4497__6260(csa_tree_add_83_21_pad_groupi_n_1223 ,csa_tree_add_83_21_pad_groupi_n_1163 ,csa_tree_add_83_21_pad_groupi_n_1166);
  xnor csa_tree_add_83_21_pad_groupi_g4498__4319(csa_tree_add_83_21_pad_groupi_n_1222 ,csa_tree_add_83_21_pad_groupi_n_1035 ,csa_tree_add_83_21_pad_groupi_n_1094);
  xnor csa_tree_add_83_21_pad_groupi_g4499__8428(csa_tree_add_83_21_pad_groupi_n_1221 ,csa_tree_add_83_21_pad_groupi_n_1100 ,csa_tree_add_83_21_pad_groupi_n_1074);
  xnor csa_tree_add_83_21_pad_groupi_g4500__5526(csa_tree_add_83_21_pad_groupi_n_1220 ,csa_tree_add_83_21_pad_groupi_n_1072 ,csa_tree_add_83_21_pad_groupi_n_1090);
  xnor csa_tree_add_83_21_pad_groupi_g4501__6783(csa_tree_add_83_21_pad_groupi_n_1219 ,csa_tree_add_83_21_pad_groupi_n_1016 ,csa_tree_add_83_21_pad_groupi_n_1097);
  xnor csa_tree_add_83_21_pad_groupi_g4502__3680(csa_tree_add_83_21_pad_groupi_n_1218 ,csa_tree_add_83_21_pad_groupi_n_1056 ,csa_tree_add_83_21_pad_groupi_n_3);
  xnor csa_tree_add_83_21_pad_groupi_g4503__1617(csa_tree_add_83_21_pad_groupi_n_1238 ,csa_tree_add_83_21_pad_groupi_n_1140 ,csa_tree_add_83_21_pad_groupi_n_1076);
  xnor csa_tree_add_83_21_pad_groupi_g4504__2802(csa_tree_add_83_21_pad_groupi_n_1217 ,csa_tree_add_83_21_pad_groupi_n_1055 ,csa_tree_add_83_21_pad_groupi_n_1095);
  xnor csa_tree_add_83_21_pad_groupi_g4505__1705(csa_tree_add_83_21_pad_groupi_n_1216 ,csa_tree_add_83_21_pad_groupi_n_1036 ,csa_tree_add_83_21_pad_groupi_n_1087);
  xnor csa_tree_add_83_21_pad_groupi_g4506__5122(csa_tree_add_83_21_pad_groupi_n_1215 ,csa_tree_add_83_21_pad_groupi_n_1137 ,csa_tree_add_83_21_pad_groupi_n_1086);
  xnor csa_tree_add_83_21_pad_groupi_g4507__8246(csa_tree_add_83_21_pad_groupi_n_1214 ,csa_tree_add_83_21_pad_groupi_n_1042 ,csa_tree_add_83_21_pad_groupi_n_1093);
  xnor csa_tree_add_83_21_pad_groupi_g4508__7098(csa_tree_add_83_21_pad_groupi_n_1213 ,csa_tree_add_83_21_pad_groupi_n_1034 ,csa_tree_add_83_21_pad_groupi_n_1104);
  xnor csa_tree_add_83_21_pad_groupi_g4509__6131(csa_tree_add_83_21_pad_groupi_n_1212 ,csa_tree_add_83_21_pad_groupi_n_1131 ,csa_tree_add_83_21_pad_groupi_n_1082);
  xnor csa_tree_add_83_21_pad_groupi_g4510__1881(csa_tree_add_83_21_pad_groupi_n_1211 ,csa_tree_add_83_21_pad_groupi_n_1134 ,csa_tree_add_83_21_pad_groupi_n_1135);
  xnor csa_tree_add_83_21_pad_groupi_g4511__5115(csa_tree_add_83_21_pad_groupi_n_1210 ,csa_tree_add_83_21_pad_groupi_n_1062 ,csa_tree_add_83_21_pad_groupi_n_1133);
  xnor csa_tree_add_83_21_pad_groupi_g4512__7482(csa_tree_add_83_21_pad_groupi_n_1236 ,csa_tree_add_83_21_pad_groupi_n_1043 ,csa_tree_add_83_21_pad_groupi_n_1078);
  xnor csa_tree_add_83_21_pad_groupi_g4513__4733(csa_tree_add_83_21_pad_groupi_n_1235 ,csa_tree_add_83_21_pad_groupi_n_1070 ,csa_tree_add_83_21_pad_groupi_n_1079);
  xnor csa_tree_add_83_21_pad_groupi_g4514__6161(csa_tree_add_83_21_pad_groupi_n_1233 ,csa_tree_add_83_21_pad_groupi_n_976 ,csa_tree_add_83_21_pad_groupi_n_1077);
  not csa_tree_add_83_21_pad_groupi_g4515(csa_tree_add_83_21_pad_groupi_n_1206 ,csa_tree_add_83_21_pad_groupi_n_1205);
  not csa_tree_add_83_21_pad_groupi_g4516(csa_tree_add_83_21_pad_groupi_n_1204 ,csa_tree_add_83_21_pad_groupi_n_1203);
  not csa_tree_add_83_21_pad_groupi_g4517(csa_tree_add_83_21_pad_groupi_n_1202 ,csa_tree_add_83_21_pad_groupi_n_1201);
  and csa_tree_add_83_21_pad_groupi_g4518__9315(csa_tree_add_83_21_pad_groupi_n_1200 ,csa_tree_add_83_21_pad_groupi_n_1035 ,csa_tree_add_83_21_pad_groupi_n_1094);
  or csa_tree_add_83_21_pad_groupi_g4519__9945(csa_tree_add_83_21_pad_groupi_n_1199 ,csa_tree_add_83_21_pad_groupi_n_1105 ,csa_tree_add_83_21_pad_groupi_n_1128);
  nor csa_tree_add_83_21_pad_groupi_g4520__2883(csa_tree_add_83_21_pad_groupi_n_1198 ,csa_tree_add_83_21_pad_groupi_n_1100 ,csa_tree_add_83_21_pad_groupi_n_1139);
  or csa_tree_add_83_21_pad_groupi_g4521__2346(csa_tree_add_83_21_pad_groupi_n_1197 ,csa_tree_add_83_21_pad_groupi_n_1136 ,csa_tree_add_83_21_pad_groupi_n_1086);
  and csa_tree_add_83_21_pad_groupi_g4522__1666(csa_tree_add_83_21_pad_groupi_n_1196 ,csa_tree_add_83_21_pad_groupi_n_1118 ,csa_tree_add_83_21_pad_groupi_n_1103);
  and csa_tree_add_83_21_pad_groupi_g4523__7410(csa_tree_add_83_21_pad_groupi_n_1195 ,csa_tree_add_83_21_pad_groupi_n_1100 ,csa_tree_add_83_21_pad_groupi_n_1139);
  or csa_tree_add_83_21_pad_groupi_g4524__6417(csa_tree_add_83_21_pad_groupi_n_1194 ,csa_tree_add_83_21_pad_groupi_n_1055 ,csa_tree_add_83_21_pad_groupi_n_1095);
  nor csa_tree_add_83_21_pad_groupi_g4525__5477(csa_tree_add_83_21_pad_groupi_n_1193 ,csa_tree_add_83_21_pad_groupi_n_1137 ,csa_tree_add_83_21_pad_groupi_n_1085);
  or csa_tree_add_83_21_pad_groupi_g4526__2398(csa_tree_add_83_21_pad_groupi_n_1192 ,csa_tree_add_83_21_pad_groupi_n_1083 ,csa_tree_add_83_21_pad_groupi_n_1089);
  nor csa_tree_add_83_21_pad_groupi_g4527__5107(csa_tree_add_83_21_pad_groupi_n_1191 ,csa_tree_add_83_21_pad_groupi_n_1022 ,csa_tree_add_83_21_pad_groupi_n_1109);
  nor csa_tree_add_83_21_pad_groupi_g4528__6260(csa_tree_add_83_21_pad_groupi_n_1190 ,csa_tree_add_83_21_pad_groupi_n_1084 ,csa_tree_add_83_21_pad_groupi_n_1090);
  or csa_tree_add_83_21_pad_groupi_g4529__4319(csa_tree_add_83_21_pad_groupi_n_1189 ,csa_tree_add_83_21_pad_groupi_n_1056 ,csa_tree_add_83_21_pad_groupi_n_3);
  nor csa_tree_add_83_21_pad_groupi_g4530__8428(csa_tree_add_83_21_pad_groupi_n_1188 ,csa_tree_add_83_21_pad_groupi_n_1019 ,csa_tree_add_83_21_pad_groupi_n_1080);
  and csa_tree_add_83_21_pad_groupi_g4531__5526(csa_tree_add_83_21_pad_groupi_n_1187 ,csa_tree_add_83_21_pad_groupi_n_1056 ,csa_tree_add_83_21_pad_groupi_n_3);
  and csa_tree_add_83_21_pad_groupi_g4532__6783(csa_tree_add_83_21_pad_groupi_n_1186 ,csa_tree_add_83_21_pad_groupi_n_1019 ,csa_tree_add_83_21_pad_groupi_n_1080);
  and csa_tree_add_83_21_pad_groupi_g4533__3680(csa_tree_add_83_21_pad_groupi_n_1185 ,csa_tree_add_83_21_pad_groupi_n_1134 ,csa_tree_add_83_21_pad_groupi_n_1135);
  nor csa_tree_add_83_21_pad_groupi_g4534__1617(csa_tree_add_83_21_pad_groupi_n_1184 ,csa_tree_add_83_21_pad_groupi_n_1134 ,csa_tree_add_83_21_pad_groupi_n_1135);
  and csa_tree_add_83_21_pad_groupi_g4535__2802(csa_tree_add_83_21_pad_groupi_n_1183 ,csa_tree_add_83_21_pad_groupi_n_1062 ,csa_tree_add_83_21_pad_groupi_n_1133);
  and csa_tree_add_83_21_pad_groupi_g4536__1705(csa_tree_add_83_21_pad_groupi_n_1182 ,csa_tree_add_83_21_pad_groupi_n_1120 ,csa_tree_add_83_21_pad_groupi_n_1106);
  or csa_tree_add_83_21_pad_groupi_g4537__5122(csa_tree_add_83_21_pad_groupi_n_1181 ,csa_tree_add_83_21_pad_groupi_n_1062 ,csa_tree_add_83_21_pad_groupi_n_1133);
  and csa_tree_add_83_21_pad_groupi_g4538__8246(csa_tree_add_83_21_pad_groupi_n_1180 ,csa_tree_add_83_21_pad_groupi_n_1050 ,csa_tree_add_83_21_pad_groupi_n_1140);
  and csa_tree_add_83_21_pad_groupi_g4539__7098(csa_tree_add_83_21_pad_groupi_n_1179 ,csa_tree_add_83_21_pad_groupi_n_1055 ,csa_tree_add_83_21_pad_groupi_n_1095);
  nor csa_tree_add_83_21_pad_groupi_g4540__6131(csa_tree_add_83_21_pad_groupi_n_1178 ,csa_tree_add_83_21_pad_groupi_n_1023 ,csa_tree_add_83_21_pad_groupi_n_1108);
  nor csa_tree_add_83_21_pad_groupi_g4541__1881(csa_tree_add_83_21_pad_groupi_n_1177 ,csa_tree_add_83_21_pad_groupi_n_1031 ,csa_tree_add_83_21_pad_groupi_n_1119);
  and csa_tree_add_83_21_pad_groupi_g4542__5115(csa_tree_add_83_21_pad_groupi_n_1209 ,csa_tree_add_83_21_pad_groupi_n_1054 ,csa_tree_add_83_21_pad_groupi_n_1127);
  or csa_tree_add_83_21_pad_groupi_g4543__7482(csa_tree_add_83_21_pad_groupi_n_1208 ,csa_tree_add_83_21_pad_groupi_n_901 ,csa_tree_add_83_21_pad_groupi_n_1122);
  or csa_tree_add_83_21_pad_groupi_g4544__4733(csa_tree_add_83_21_pad_groupi_n_1207 ,csa_tree_add_83_21_pad_groupi_n_914 ,csa_tree_add_83_21_pad_groupi_n_1125);
  and csa_tree_add_83_21_pad_groupi_g4545__6161(csa_tree_add_83_21_pad_groupi_n_1205 ,csa_tree_add_83_21_pad_groupi_n_884 ,csa_tree_add_83_21_pad_groupi_n_1116);
  and csa_tree_add_83_21_pad_groupi_g4546__9315(csa_tree_add_83_21_pad_groupi_n_1203 ,csa_tree_add_83_21_pad_groupi_n_921 ,csa_tree_add_83_21_pad_groupi_n_1126);
  or csa_tree_add_83_21_pad_groupi_g4547__9945(csa_tree_add_83_21_pad_groupi_n_1201 ,csa_tree_add_83_21_pad_groupi_n_1049 ,csa_tree_add_83_21_pad_groupi_n_1117);
  not csa_tree_add_83_21_pad_groupi_g4548(csa_tree_add_83_21_pad_groupi_n_1170 ,csa_tree_add_83_21_pad_groupi_n_1171);
  not csa_tree_add_83_21_pad_groupi_g4549(csa_tree_add_83_21_pad_groupi_n_1166 ,csa_tree_add_83_21_pad_groupi_n_1165);
  not csa_tree_add_83_21_pad_groupi_g4550(csa_tree_add_83_21_pad_groupi_n_1163 ,csa_tree_add_83_21_pad_groupi_n_1162);
  not csa_tree_add_83_21_pad_groupi_g4551(csa_tree_add_83_21_pad_groupi_n_1160 ,csa_tree_add_83_21_pad_groupi_n_1159);
  or csa_tree_add_83_21_pad_groupi_g4552__2883(csa_tree_add_83_21_pad_groupi_n_1158 ,csa_tree_add_83_21_pad_groupi_n_1035 ,csa_tree_add_83_21_pad_groupi_n_1094);
  and csa_tree_add_83_21_pad_groupi_g4553__2346(csa_tree_add_83_21_pad_groupi_n_1157 ,csa_tree_add_83_21_pad_groupi_n_1015 ,csa_tree_add_83_21_pad_groupi_n_1097);
  or csa_tree_add_83_21_pad_groupi_g4554__1666(csa_tree_add_83_21_pad_groupi_n_1156 ,csa_tree_add_83_21_pad_groupi_n_1130 ,csa_tree_add_83_21_pad_groupi_n_1081);
  or csa_tree_add_83_21_pad_groupi_g4555__7410(csa_tree_add_83_21_pad_groupi_n_1155 ,csa_tree_add_83_21_pad_groupi_n_1033 ,csa_tree_add_83_21_pad_groupi_n_1091);
  and csa_tree_add_83_21_pad_groupi_g4556__6417(csa_tree_add_83_21_pad_groupi_n_1154 ,csa_tree_add_83_21_pad_groupi_n_1093 ,csa_tree_add_83_21_pad_groupi_n_1088);
  nor csa_tree_add_83_21_pad_groupi_g4557__5477(csa_tree_add_83_21_pad_groupi_n_1153 ,csa_tree_add_83_21_pad_groupi_n_1093 ,csa_tree_add_83_21_pad_groupi_n_1088);
  and csa_tree_add_83_21_pad_groupi_g4558__2398(csa_tree_add_83_21_pad_groupi_n_1152 ,csa_tree_add_83_21_pad_groupi_n_1016 ,csa_tree_add_83_21_pad_groupi_n_1096);
  nor csa_tree_add_83_21_pad_groupi_g4559__5107(csa_tree_add_83_21_pad_groupi_n_1151 ,csa_tree_add_83_21_pad_groupi_n_1034 ,csa_tree_add_83_21_pad_groupi_n_1092);
  nor csa_tree_add_83_21_pad_groupi_g4560__6260(csa_tree_add_83_21_pad_groupi_n_1150 ,csa_tree_add_83_21_pad_groupi_n_1131 ,csa_tree_add_83_21_pad_groupi_n_1082);
  or csa_tree_add_83_21_pad_groupi_g4561__4319(csa_tree_add_83_21_pad_groupi_n_1149 ,csa_tree_add_83_21_pad_groupi_n_1110 ,csa_tree_add_83_21_pad_groupi_n_1101);
  and csa_tree_add_83_21_pad_groupi_g4562__8428(csa_tree_add_83_21_pad_groupi_n_1148 ,csa_tree_add_83_21_pad_groupi_n_1037 ,csa_tree_add_83_21_pad_groupi_n_1087);
  nor csa_tree_add_83_21_pad_groupi_g4563__5526(csa_tree_add_83_21_pad_groupi_n_1147 ,csa_tree_add_83_21_pad_groupi_n_1037 ,csa_tree_add_83_21_pad_groupi_n_1087);
  xnor csa_tree_add_83_21_pad_groupi_g4564__6783(csa_tree_add_83_21_pad_groupi_n_1146 ,csa_tree_add_83_21_pad_groupi_n_1010 ,csa_tree_add_83_21_pad_groupi_n_1064);
  xnor csa_tree_add_83_21_pad_groupi_g4565__3680(csa_tree_add_83_21_pad_groupi_n_1145 ,csa_tree_add_83_21_pad_groupi_n_1067 ,csa_tree_add_83_21_pad_groupi_n_1019);
  xnor csa_tree_add_83_21_pad_groupi_g4566__1617(csa_tree_add_83_21_pad_groupi_n_1144 ,csa_tree_add_83_21_pad_groupi_n_1058 ,csa_tree_add_83_21_pad_groupi_n_1061);
  xnor csa_tree_add_83_21_pad_groupi_g4567__2802(csa_tree_add_83_21_pad_groupi_n_1143 ,csa_tree_add_83_21_pad_groupi_n_1011 ,csa_tree_add_83_21_pad_groupi_n_1059);
  xnor csa_tree_add_83_21_pad_groupi_g4568__1705(csa_tree_add_83_21_pad_groupi_n_1142 ,csa_tree_add_83_21_pad_groupi_n_1018 ,csa_tree_add_83_21_pad_groupi_n_1066);
  xnor csa_tree_add_83_21_pad_groupi_g4569__5122(csa_tree_add_83_21_pad_groupi_n_1176 ,csa_tree_add_83_21_pad_groupi_n_1020 ,csa_tree_add_83_21_pad_groupi_n_1025);
  and csa_tree_add_83_21_pad_groupi_g4570__8246(csa_tree_add_83_21_pad_groupi_n_1175 ,csa_tree_add_83_21_pad_groupi_n_1030 ,csa_tree_add_83_21_pad_groupi_n_1111);
  xnor csa_tree_add_83_21_pad_groupi_g4571__7098(csa_tree_add_83_21_pad_groupi_n_1174 ,csa_tree_add_83_21_pad_groupi_n_1068 ,csa_tree_add_83_21_pad_groupi_n_950);
  or csa_tree_add_83_21_pad_groupi_g4572__6131(csa_tree_add_83_21_pad_groupi_n_1173 ,csa_tree_add_83_21_pad_groupi_n_908 ,csa_tree_add_83_21_pad_groupi_n_1121);
  xnor csa_tree_add_83_21_pad_groupi_g4573__1881(csa_tree_add_83_21_pad_groupi_n_1172 ,csa_tree_add_83_21_pad_groupi_n_1045 ,csa_tree_add_83_21_pad_groupi_n_944);
  xnor csa_tree_add_83_21_pad_groupi_g4574__5115(csa_tree_add_83_21_pad_groupi_n_1171 ,csa_tree_add_83_21_pad_groupi_n_1073 ,csa_tree_add_83_21_pad_groupi_n_941);
  xnor csa_tree_add_83_21_pad_groupi_g4575__7482(csa_tree_add_83_21_pad_groupi_n_1169 ,csa_tree_add_83_21_pad_groupi_n_1041 ,csa_tree_add_83_21_pad_groupi_n_974);
  xnor csa_tree_add_83_21_pad_groupi_g4576__4733(csa_tree_add_83_21_pad_groupi_n_1168 ,csa_tree_add_83_21_pad_groupi_n_1044 ,csa_tree_add_83_21_pad_groupi_n_939);
  xnor csa_tree_add_83_21_pad_groupi_g4577__6161(csa_tree_add_83_21_pad_groupi_n_1167 ,csa_tree_add_83_21_pad_groupi_n_1040 ,csa_tree_add_83_21_pad_groupi_n_969);
  xnor csa_tree_add_83_21_pad_groupi_g4578__9315(csa_tree_add_83_21_pad_groupi_n_1165 ,csa_tree_add_83_21_pad_groupi_n_1038 ,csa_tree_add_83_21_pad_groupi_n_970);
  or csa_tree_add_83_21_pad_groupi_g4579__9945(csa_tree_add_83_21_pad_groupi_n_1164 ,csa_tree_add_83_21_pad_groupi_n_858 ,csa_tree_add_83_21_pad_groupi_n_1113);
  and csa_tree_add_83_21_pad_groupi_g4580__2883(csa_tree_add_83_21_pad_groupi_n_1162 ,csa_tree_add_83_21_pad_groupi_n_857 ,csa_tree_add_83_21_pad_groupi_n_1112);
  or csa_tree_add_83_21_pad_groupi_g4581__2346(csa_tree_add_83_21_pad_groupi_n_1161 ,csa_tree_add_83_21_pad_groupi_n_873 ,csa_tree_add_83_21_pad_groupi_n_1129);
  xnor csa_tree_add_83_21_pad_groupi_g4582__1666(csa_tree_add_83_21_pad_groupi_n_1159 ,csa_tree_add_83_21_pad_groupi_n_1046 ,csa_tree_add_83_21_pad_groupi_n_955);
  not csa_tree_add_83_21_pad_groupi_g4583(csa_tree_add_83_21_pad_groupi_n_1139 ,csa_tree_add_83_21_pad_groupi_n_1138);
  not csa_tree_add_83_21_pad_groupi_g4584(csa_tree_add_83_21_pad_groupi_n_1136 ,csa_tree_add_83_21_pad_groupi_n_1137);
  not csa_tree_add_83_21_pad_groupi_g4585(csa_tree_add_83_21_pad_groupi_n_1130 ,csa_tree_add_83_21_pad_groupi_n_1131);
  and csa_tree_add_83_21_pad_groupi_g4586__7410(csa_tree_add_83_21_pad_groupi_n_1129 ,csa_tree_add_83_21_pad_groupi_n_871 ,csa_tree_add_83_21_pad_groupi_n_1040);
  nor csa_tree_add_83_21_pad_groupi_g4587__6417(csa_tree_add_83_21_pad_groupi_n_1128 ,csa_tree_add_83_21_pad_groupi_n_1058 ,csa_tree_add_83_21_pad_groupi_n_1061);
  or csa_tree_add_83_21_pad_groupi_g4588__5477(csa_tree_add_83_21_pad_groupi_n_1127 ,csa_tree_add_83_21_pad_groupi_n_1053 ,csa_tree_add_83_21_pad_groupi_n_1071);
  or csa_tree_add_83_21_pad_groupi_g4589__2398(csa_tree_add_83_21_pad_groupi_n_1126 ,csa_tree_add_83_21_pad_groupi_n_918 ,csa_tree_add_83_21_pad_groupi_n_1069);
  and csa_tree_add_83_21_pad_groupi_g4590__5107(csa_tree_add_83_21_pad_groupi_n_1125 ,csa_tree_add_83_21_pad_groupi_n_932 ,csa_tree_add_83_21_pad_groupi_n_1073);
  nor csa_tree_add_83_21_pad_groupi_g4591__6260(csa_tree_add_83_21_pad_groupi_n_1124 ,csa_tree_add_83_21_pad_groupi_n_1010 ,csa_tree_add_83_21_pad_groupi_n_1063);
  and csa_tree_add_83_21_pad_groupi_g4592__4319(csa_tree_add_83_21_pad_groupi_n_1123 ,csa_tree_add_83_21_pad_groupi_n_1011 ,csa_tree_add_83_21_pad_groupi_n_1059);
  and csa_tree_add_83_21_pad_groupi_g4593__8428(csa_tree_add_83_21_pad_groupi_n_1122 ,csa_tree_add_83_21_pad_groupi_n_880 ,csa_tree_add_83_21_pad_groupi_n_1045);
  and csa_tree_add_83_21_pad_groupi_g4594__5526(csa_tree_add_83_21_pad_groupi_n_1121 ,csa_tree_add_83_21_pad_groupi_n_867 ,csa_tree_add_83_21_pad_groupi_n_1044);
  or csa_tree_add_83_21_pad_groupi_g4595__6783(csa_tree_add_83_21_pad_groupi_n_1120 ,csa_tree_add_83_21_pad_groupi_n_1011 ,csa_tree_add_83_21_pad_groupi_n_1059);
  nor csa_tree_add_83_21_pad_groupi_g4596__3680(csa_tree_add_83_21_pad_groupi_n_1119 ,csa_tree_add_83_21_pad_groupi_n_1026 ,csa_tree_add_83_21_pad_groupi_n_980);
  or csa_tree_add_83_21_pad_groupi_g4597__1617(csa_tree_add_83_21_pad_groupi_n_1118 ,csa_tree_add_83_21_pad_groupi_n_1009 ,csa_tree_add_83_21_pad_groupi_n_1064);
  and csa_tree_add_83_21_pad_groupi_g4598__2802(csa_tree_add_83_21_pad_groupi_n_1117 ,csa_tree_add_83_21_pad_groupi_n_1029 ,csa_tree_add_83_21_pad_groupi_n_1043);
  or csa_tree_add_83_21_pad_groupi_g4599__1705(csa_tree_add_83_21_pad_groupi_n_1116 ,csa_tree_add_83_21_pad_groupi_n_882 ,csa_tree_add_83_21_pad_groupi_n_1038);
  or csa_tree_add_83_21_pad_groupi_g4600__5122(csa_tree_add_83_21_pad_groupi_n_1115 ,csa_tree_add_83_21_pad_groupi_n_1057 ,csa_tree_add_83_21_pad_groupi_n_1060);
  or csa_tree_add_83_21_pad_groupi_g4601__8246(csa_tree_add_83_21_pad_groupi_n_1114 ,csa_tree_add_83_21_pad_groupi_n_1017 ,csa_tree_add_83_21_pad_groupi_n_1065);
  and csa_tree_add_83_21_pad_groupi_g4602__7098(csa_tree_add_83_21_pad_groupi_n_1113 ,csa_tree_add_83_21_pad_groupi_n_860 ,csa_tree_add_83_21_pad_groupi_n_1041);
  or csa_tree_add_83_21_pad_groupi_g4603__6131(csa_tree_add_83_21_pad_groupi_n_1112 ,csa_tree_add_83_21_pad_groupi_n_854 ,csa_tree_add_83_21_pad_groupi_n_1046);
  or csa_tree_add_83_21_pad_groupi_g4604__1881(csa_tree_add_83_21_pad_groupi_n_1111 ,csa_tree_add_83_21_pad_groupi_n_1028 ,csa_tree_add_83_21_pad_groupi_n_976);
  nor csa_tree_add_83_21_pad_groupi_g4605__5115(csa_tree_add_83_21_pad_groupi_n_1110 ,csa_tree_add_83_21_pad_groupi_n_1018 ,csa_tree_add_83_21_pad_groupi_n_1066);
  xnor csa_tree_add_83_21_pad_groupi_g4606__7482(csa_tree_add_83_21_pad_groupi_n_1141 ,csa_tree_add_83_21_pad_groupi_n_842 ,csa_tree_add_83_21_pad_groupi_n_951);
  xnor csa_tree_add_83_21_pad_groupi_g4607__4733(csa_tree_add_83_21_pad_groupi_n_1140 ,csa_tree_add_83_21_pad_groupi_n_803 ,csa_tree_add_83_21_pad_groupi_n_964);
  xnor csa_tree_add_83_21_pad_groupi_g4608__6161(csa_tree_add_83_21_pad_groupi_n_1138 ,csa_tree_add_83_21_pad_groupi_n_773 ,csa_tree_add_83_21_pad_groupi_n_962);
  xnor csa_tree_add_83_21_pad_groupi_g4609__9315(csa_tree_add_83_21_pad_groupi_n_1137 ,csa_tree_add_83_21_pad_groupi_n_783 ,csa_tree_add_83_21_pad_groupi_n_960);
  xnor csa_tree_add_83_21_pad_groupi_g4610__9945(csa_tree_add_83_21_pad_groupi_n_1135 ,csa_tree_add_83_21_pad_groupi_n_840 ,csa_tree_add_83_21_pad_groupi_n_965);
  or csa_tree_add_83_21_pad_groupi_g4611__2883(csa_tree_add_83_21_pad_groupi_n_1134 ,csa_tree_add_83_21_pad_groupi_n_1000 ,csa_tree_add_83_21_pad_groupi_n_1052);
  xnor csa_tree_add_83_21_pad_groupi_g4612__2346(csa_tree_add_83_21_pad_groupi_n_1133 ,csa_tree_add_83_21_pad_groupi_n_778 ,csa_tree_add_83_21_pad_groupi_n_949);
  and csa_tree_add_83_21_pad_groupi_g4613__1666(csa_tree_add_83_21_pad_groupi_n_1132 ,csa_tree_add_83_21_pad_groupi_n_888 ,csa_tree_add_83_21_pad_groupi_n_1032);
  or csa_tree_add_83_21_pad_groupi_g4614__7410(csa_tree_add_83_21_pad_groupi_n_1131 ,csa_tree_add_83_21_pad_groupi_n_868 ,csa_tree_add_83_21_pad_groupi_n_1027);
  not csa_tree_add_83_21_pad_groupi_g4615(csa_tree_add_83_21_pad_groupi_n_1109 ,csa_tree_add_83_21_pad_groupi_n_1108);
  not csa_tree_add_83_21_pad_groupi_g4616(csa_tree_add_83_21_pad_groupi_n_1097 ,csa_tree_add_83_21_pad_groupi_n_1096);
  not csa_tree_add_83_21_pad_groupi_g4617(csa_tree_add_83_21_pad_groupi_n_1091 ,csa_tree_add_83_21_pad_groupi_n_1092);
  not csa_tree_add_83_21_pad_groupi_g4618(csa_tree_add_83_21_pad_groupi_n_1090 ,csa_tree_add_83_21_pad_groupi_n_1089);
  not csa_tree_add_83_21_pad_groupi_g4619(csa_tree_add_83_21_pad_groupi_n_1085 ,csa_tree_add_83_21_pad_groupi_n_1086);
  not csa_tree_add_83_21_pad_groupi_g4620(csa_tree_add_83_21_pad_groupi_n_1083 ,csa_tree_add_83_21_pad_groupi_n_1084);
  not csa_tree_add_83_21_pad_groupi_g4621(csa_tree_add_83_21_pad_groupi_n_1081 ,csa_tree_add_83_21_pad_groupi_n_1082);
  xnor csa_tree_add_83_21_pad_groupi_g4622__6417(csa_tree_add_83_21_pad_groupi_n_1079 ,csa_tree_add_83_21_pad_groupi_n_975 ,csa_tree_add_83_21_pad_groupi_n_934);
  xnor csa_tree_add_83_21_pad_groupi_g4623__5477(csa_tree_add_83_21_pad_groupi_n_1108 ,csa_tree_add_83_21_pad_groupi_n_892 ,csa_tree_add_83_21_pad_groupi_n_961);
  xnor csa_tree_add_83_21_pad_groupi_g4624__2398(csa_tree_add_83_21_pad_groupi_n_1078 ,csa_tree_add_83_21_pad_groupi_n_797 ,csa_tree_add_83_21_pad_groupi_n_4);
  xnor csa_tree_add_83_21_pad_groupi_g4625__5107(csa_tree_add_83_21_pad_groupi_n_1077 ,csa_tree_add_83_21_pad_groupi_n_746 ,csa_tree_add_83_21_pad_groupi_n_1014);
  xnor csa_tree_add_83_21_pad_groupi_g4626__6260(csa_tree_add_83_21_pad_groupi_n_1076 ,csa_tree_add_83_21_pad_groupi_n_1012 ,csa_tree_add_83_21_pad_groupi_n_933);
  xnor csa_tree_add_83_21_pad_groupi_g4628__4319(csa_tree_add_83_21_pad_groupi_n_1107 ,csa_tree_add_83_21_pad_groupi_n_768 ,csa_tree_add_83_21_pad_groupi_n_942);
  xnor csa_tree_add_83_21_pad_groupi_g4629__8428(csa_tree_add_83_21_pad_groupi_n_1106 ,csa_tree_add_83_21_pad_groupi_n_764 ,csa_tree_add_83_21_pad_groupi_n_968);
  xnor csa_tree_add_83_21_pad_groupi_g4630__5526(csa_tree_add_83_21_pad_groupi_n_1105 ,csa_tree_add_83_21_pad_groupi_n_740 ,csa_tree_add_83_21_pad_groupi_n_963);
  xnor csa_tree_add_83_21_pad_groupi_g4631__6783(csa_tree_add_83_21_pad_groupi_n_1104 ,csa_tree_add_83_21_pad_groupi_n_782 ,csa_tree_add_83_21_pad_groupi_n_967);
  xnor csa_tree_add_83_21_pad_groupi_g4632__3680(csa_tree_add_83_21_pad_groupi_n_1103 ,csa_tree_add_83_21_pad_groupi_n_1021 ,csa_tree_add_83_21_pad_groupi_n_957);
  xnor csa_tree_add_83_21_pad_groupi_g4633__1617(csa_tree_add_83_21_pad_groupi_n_1102 ,csa_tree_add_83_21_pad_groupi_n_769 ,csa_tree_add_83_21_pad_groupi_n_945);
  xnor csa_tree_add_83_21_pad_groupi_g4634__2802(csa_tree_add_83_21_pad_groupi_n_1101 ,csa_tree_add_83_21_pad_groupi_n_977 ,csa_tree_add_83_21_pad_groupi_n_966);
  xnor csa_tree_add_83_21_pad_groupi_g4635__1705(csa_tree_add_83_21_pad_groupi_n_1100 ,csa_tree_add_83_21_pad_groupi_n_838 ,csa_tree_add_83_21_pad_groupi_n_946);
  xnor csa_tree_add_83_21_pad_groupi_g4637__5122(csa_tree_add_83_21_pad_groupi_n_1099 ,csa_tree_add_83_21_pad_groupi_n_750 ,csa_tree_add_83_21_pad_groupi_n_952);
  xnor csa_tree_add_83_21_pad_groupi_g4638__8246(csa_tree_add_83_21_pad_groupi_n_1098 ,csa_tree_add_83_21_pad_groupi_n_743 ,csa_tree_add_83_21_pad_groupi_n_972);
  xnor csa_tree_add_83_21_pad_groupi_g4639__7098(csa_tree_add_83_21_pad_groupi_n_1096 ,csa_tree_add_83_21_pad_groupi_n_971 ,csa_tree_add_83_21_pad_groupi_n_578);
  xnor csa_tree_add_83_21_pad_groupi_g4640__6131(csa_tree_add_83_21_pad_groupi_n_1095 ,csa_tree_add_83_21_pad_groupi_n_770 ,csa_tree_add_83_21_pad_groupi_n_947);
  xnor csa_tree_add_83_21_pad_groupi_g4641__1881(csa_tree_add_83_21_pad_groupi_n_1094 ,csa_tree_add_83_21_pad_groupi_n_830 ,csa_tree_add_83_21_pad_groupi_n_943);
  xnor csa_tree_add_83_21_pad_groupi_g4642__5115(csa_tree_add_83_21_pad_groupi_n_1093 ,csa_tree_add_83_21_pad_groupi_n_780 ,csa_tree_add_83_21_pad_groupi_n_938);
  xnor csa_tree_add_83_21_pad_groupi_g4643__7482(csa_tree_add_83_21_pad_groupi_n_1092 ,csa_tree_add_83_21_pad_groupi_n_775 ,csa_tree_add_83_21_pad_groupi_n_937);
  xnor csa_tree_add_83_21_pad_groupi_g4644__4733(csa_tree_add_83_21_pad_groupi_n_1089 ,csa_tree_add_83_21_pad_groupi_n_827 ,csa_tree_add_83_21_pad_groupi_n_973);
  xnor csa_tree_add_83_21_pad_groupi_g4645__6161(csa_tree_add_83_21_pad_groupi_n_1088 ,csa_tree_add_83_21_pad_groupi_n_777 ,csa_tree_add_83_21_pad_groupi_n_940);
  xnor csa_tree_add_83_21_pad_groupi_g4646__9315(csa_tree_add_83_21_pad_groupi_n_1087 ,csa_tree_add_83_21_pad_groupi_n_774 ,csa_tree_add_83_21_pad_groupi_n_954);
  xnor csa_tree_add_83_21_pad_groupi_g4647__9945(csa_tree_add_83_21_pad_groupi_n_1086 ,csa_tree_add_83_21_pad_groupi_n_893 ,csa_tree_add_83_21_pad_groupi_n_959);
  xnor csa_tree_add_83_21_pad_groupi_g4648__2883(csa_tree_add_83_21_pad_groupi_n_1084 ,csa_tree_add_83_21_pad_groupi_n_785 ,csa_tree_add_83_21_pad_groupi_n_956);
  xnor csa_tree_add_83_21_pad_groupi_g4649__2346(csa_tree_add_83_21_pad_groupi_n_1082 ,csa_tree_add_83_21_pad_groupi_n_839 ,csa_tree_add_83_21_pad_groupi_n_958);
  xnor csa_tree_add_83_21_pad_groupi_g4650__1666(csa_tree_add_83_21_pad_groupi_n_1080 ,csa_tree_add_83_21_pad_groupi_n_936 ,csa_tree_add_83_21_pad_groupi_n_953);
  not csa_tree_add_83_21_pad_groupi_g4651(csa_tree_add_83_21_pad_groupi_n_1071 ,csa_tree_add_83_21_pad_groupi_n_1070);
  not csa_tree_add_83_21_pad_groupi_g4652(csa_tree_add_83_21_pad_groupi_n_1069 ,csa_tree_add_83_21_pad_groupi_n_1068);
  not csa_tree_add_83_21_pad_groupi_g4653(csa_tree_add_83_21_pad_groupi_n_1065 ,csa_tree_add_83_21_pad_groupi_n_1066);
  not csa_tree_add_83_21_pad_groupi_g4654(csa_tree_add_83_21_pad_groupi_n_1063 ,csa_tree_add_83_21_pad_groupi_n_1064);
  not csa_tree_add_83_21_pad_groupi_g4655(csa_tree_add_83_21_pad_groupi_n_1060 ,csa_tree_add_83_21_pad_groupi_n_1061);
  not csa_tree_add_83_21_pad_groupi_g4656(csa_tree_add_83_21_pad_groupi_n_1057 ,csa_tree_add_83_21_pad_groupi_n_1058);
  or csa_tree_add_83_21_pad_groupi_g4657__7410(csa_tree_add_83_21_pad_groupi_n_1054 ,csa_tree_add_83_21_pad_groupi_n_276 ,csa_tree_add_83_21_pad_groupi_n_975);
  and csa_tree_add_83_21_pad_groupi_g4658__6417(csa_tree_add_83_21_pad_groupi_n_1053 ,csa_tree_add_83_21_pad_groupi_n_934 ,csa_tree_add_83_21_pad_groupi_n_975);
  and csa_tree_add_83_21_pad_groupi_g4659__5477(csa_tree_add_83_21_pad_groupi_n_1052 ,csa_tree_add_83_21_pad_groupi_n_998 ,csa_tree_add_83_21_pad_groupi_n_1020);
  and csa_tree_add_83_21_pad_groupi_g4660__2398(csa_tree_add_83_21_pad_groupi_n_1051 ,csa_tree_add_83_21_pad_groupi_n_933 ,csa_tree_add_83_21_pad_groupi_n_1012);
  or csa_tree_add_83_21_pad_groupi_g4661__5107(csa_tree_add_83_21_pad_groupi_n_1050 ,csa_tree_add_83_21_pad_groupi_n_933 ,csa_tree_add_83_21_pad_groupi_n_1012);
  and csa_tree_add_83_21_pad_groupi_g4662__6260(csa_tree_add_83_21_pad_groupi_n_1049 ,csa_tree_add_83_21_pad_groupi_n_797 ,csa_tree_add_83_21_pad_groupi_n_4);
  and csa_tree_add_83_21_pad_groupi_g4663__4319(csa_tree_add_83_21_pad_groupi_n_1074 ,csa_tree_add_83_21_pad_groupi_n_913 ,csa_tree_add_83_21_pad_groupi_n_1007);
  or csa_tree_add_83_21_pad_groupi_g4664__8428(csa_tree_add_83_21_pad_groupi_n_1073 ,csa_tree_add_83_21_pad_groupi_n_910 ,csa_tree_add_83_21_pad_groupi_n_999);
  and csa_tree_add_83_21_pad_groupi_g4665__5526(csa_tree_add_83_21_pad_groupi_n_1072 ,csa_tree_add_83_21_pad_groupi_n_915 ,csa_tree_add_83_21_pad_groupi_n_996);
  or csa_tree_add_83_21_pad_groupi_g4666__6783(csa_tree_add_83_21_pad_groupi_n_1070 ,csa_tree_add_83_21_pad_groupi_n_890 ,csa_tree_add_83_21_pad_groupi_n_1005);
  or csa_tree_add_83_21_pad_groupi_g4667__3680(csa_tree_add_83_21_pad_groupi_n_1068 ,csa_tree_add_83_21_pad_groupi_n_905 ,csa_tree_add_83_21_pad_groupi_n_1003);
  and csa_tree_add_83_21_pad_groupi_g4668__1617(csa_tree_add_83_21_pad_groupi_n_1067 ,csa_tree_add_83_21_pad_groupi_n_912 ,csa_tree_add_83_21_pad_groupi_n_1002);
  or csa_tree_add_83_21_pad_groupi_g4669__2802(csa_tree_add_83_21_pad_groupi_n_1066 ,csa_tree_add_83_21_pad_groupi_n_903 ,csa_tree_add_83_21_pad_groupi_n_1004);
  or csa_tree_add_83_21_pad_groupi_g4670__1705(csa_tree_add_83_21_pad_groupi_n_1064 ,csa_tree_add_83_21_pad_groupi_n_925 ,csa_tree_add_83_21_pad_groupi_n_1006);
  or csa_tree_add_83_21_pad_groupi_g4671__5122(csa_tree_add_83_21_pad_groupi_n_1062 ,csa_tree_add_83_21_pad_groupi_n_874 ,csa_tree_add_83_21_pad_groupi_n_987);
  or csa_tree_add_83_21_pad_groupi_g4672__8246(csa_tree_add_83_21_pad_groupi_n_1061 ,csa_tree_add_83_21_pad_groupi_n_929 ,csa_tree_add_83_21_pad_groupi_n_979);
  or csa_tree_add_83_21_pad_groupi_g4673__7098(csa_tree_add_83_21_pad_groupi_n_1059 ,csa_tree_add_83_21_pad_groupi_n_889 ,csa_tree_add_83_21_pad_groupi_n_995);
  or csa_tree_add_83_21_pad_groupi_g4674__6131(csa_tree_add_83_21_pad_groupi_n_1058 ,csa_tree_add_83_21_pad_groupi_n_911 ,csa_tree_add_83_21_pad_groupi_n_1008);
  or csa_tree_add_83_21_pad_groupi_g4675__1881(csa_tree_add_83_21_pad_groupi_n_1056 ,csa_tree_add_83_21_pad_groupi_n_869 ,csa_tree_add_83_21_pad_groupi_n_1001);
  or csa_tree_add_83_21_pad_groupi_g4676__5115(csa_tree_add_83_21_pad_groupi_n_1055 ,csa_tree_add_83_21_pad_groupi_n_886 ,csa_tree_add_83_21_pad_groupi_n_993);
  not csa_tree_add_83_21_pad_groupi_g4677(csa_tree_add_83_21_pad_groupi_n_1048 ,csa_tree_add_83_21_pad_groupi_n_1047);
  not csa_tree_add_83_21_pad_groupi_g4678(csa_tree_add_83_21_pad_groupi_n_1037 ,csa_tree_add_83_21_pad_groupi_n_1036);
  not csa_tree_add_83_21_pad_groupi_g4679(csa_tree_add_83_21_pad_groupi_n_1033 ,csa_tree_add_83_21_pad_groupi_n_1034);
  or csa_tree_add_83_21_pad_groupi_g4680__7482(csa_tree_add_83_21_pad_groupi_n_1032 ,csa_tree_add_83_21_pad_groupi_n_876 ,csa_tree_add_83_21_pad_groupi_n_977);
  nor csa_tree_add_83_21_pad_groupi_g4681__4733(csa_tree_add_83_21_pad_groupi_n_1031 ,csa_tree_add_83_21_pad_groupi_n_646 ,csa_tree_add_83_21_pad_groupi_n_1024);
  or csa_tree_add_83_21_pad_groupi_g4682__6161(csa_tree_add_83_21_pad_groupi_n_1030 ,csa_tree_add_83_21_pad_groupi_n_745 ,csa_tree_add_83_21_pad_groupi_n_1014);
  or csa_tree_add_83_21_pad_groupi_g4683__9315(csa_tree_add_83_21_pad_groupi_n_1029 ,csa_tree_add_83_21_pad_groupi_n_797 ,csa_tree_add_83_21_pad_groupi_n_4);
  nor csa_tree_add_83_21_pad_groupi_g4684__9945(csa_tree_add_83_21_pad_groupi_n_1028 ,csa_tree_add_83_21_pad_groupi_n_746 ,csa_tree_add_83_21_pad_groupi_n_1013);
  and csa_tree_add_83_21_pad_groupi_g4685__2883(csa_tree_add_83_21_pad_groupi_n_1027 ,csa_tree_add_83_21_pad_groupi_n_865 ,csa_tree_add_83_21_pad_groupi_n_1021);
  and csa_tree_add_83_21_pad_groupi_g4686__2346(csa_tree_add_83_21_pad_groupi_n_1026 ,csa_tree_add_83_21_pad_groupi_n_646 ,csa_tree_add_83_21_pad_groupi_n_1024);
  and csa_tree_add_83_21_pad_groupi_g4687__1666(csa_tree_add_83_21_pad_groupi_n_1047 ,csa_tree_add_83_21_pad_groupi_n_895 ,csa_tree_add_83_21_pad_groupi_n_994);
  xnor csa_tree_add_83_21_pad_groupi_g4688__7410(csa_tree_add_83_21_pad_groupi_n_1025 ,csa_tree_add_83_21_pad_groupi_n_935 ,csa_tree_add_83_21_pad_groupi_n_820);
  and csa_tree_add_83_21_pad_groupi_g4689__6417(csa_tree_add_83_21_pad_groupi_n_1046 ,csa_tree_add_83_21_pad_groupi_n_853 ,csa_tree_add_83_21_pad_groupi_n_982);
  or csa_tree_add_83_21_pad_groupi_g4690__5477(csa_tree_add_83_21_pad_groupi_n_1045 ,csa_tree_add_83_21_pad_groupi_n_906 ,csa_tree_add_83_21_pad_groupi_n_997);
  or csa_tree_add_83_21_pad_groupi_g4691__2398(csa_tree_add_83_21_pad_groupi_n_1044 ,csa_tree_add_83_21_pad_groupi_n_887 ,csa_tree_add_83_21_pad_groupi_n_992);
  or csa_tree_add_83_21_pad_groupi_g4692__5107(csa_tree_add_83_21_pad_groupi_n_1043 ,csa_tree_add_83_21_pad_groupi_n_926 ,csa_tree_add_83_21_pad_groupi_n_991);
  and csa_tree_add_83_21_pad_groupi_g4693__6260(csa_tree_add_83_21_pad_groupi_n_1042 ,csa_tree_add_83_21_pad_groupi_n_864 ,csa_tree_add_83_21_pad_groupi_n_985);
  or csa_tree_add_83_21_pad_groupi_g4694__4319(csa_tree_add_83_21_pad_groupi_n_1041 ,csa_tree_add_83_21_pad_groupi_n_879 ,csa_tree_add_83_21_pad_groupi_n_984);
  or csa_tree_add_83_21_pad_groupi_g4695__8428(csa_tree_add_83_21_pad_groupi_n_1040 ,csa_tree_add_83_21_pad_groupi_n_870 ,csa_tree_add_83_21_pad_groupi_n_988);
  and csa_tree_add_83_21_pad_groupi_g4696__5526(csa_tree_add_83_21_pad_groupi_n_1039 ,csa_tree_add_83_21_pad_groupi_n_852 ,csa_tree_add_83_21_pad_groupi_n_981);
  and csa_tree_add_83_21_pad_groupi_g4697__6783(csa_tree_add_83_21_pad_groupi_n_1038 ,csa_tree_add_83_21_pad_groupi_n_878 ,csa_tree_add_83_21_pad_groupi_n_989);
  or csa_tree_add_83_21_pad_groupi_g4698__3680(csa_tree_add_83_21_pad_groupi_n_1036 ,csa_tree_add_83_21_pad_groupi_n_897 ,csa_tree_add_83_21_pad_groupi_n_983);
  or csa_tree_add_83_21_pad_groupi_g4699__1617(csa_tree_add_83_21_pad_groupi_n_1035 ,csa_tree_add_83_21_pad_groupi_n_907 ,csa_tree_add_83_21_pad_groupi_n_990);
  or csa_tree_add_83_21_pad_groupi_g4700__2802(csa_tree_add_83_21_pad_groupi_n_1034 ,csa_tree_add_83_21_pad_groupi_n_866 ,csa_tree_add_83_21_pad_groupi_n_986);
  not csa_tree_add_83_21_pad_groupi_g4701(csa_tree_add_83_21_pad_groupi_n_1023 ,csa_tree_add_83_21_pad_groupi_n_1022);
  not csa_tree_add_83_21_pad_groupi_g4702(csa_tree_add_83_21_pad_groupi_n_1018 ,csa_tree_add_83_21_pad_groupi_n_1017);
  not csa_tree_add_83_21_pad_groupi_g4703(csa_tree_add_83_21_pad_groupi_n_1016 ,csa_tree_add_83_21_pad_groupi_n_1015);
  not csa_tree_add_83_21_pad_groupi_g4704(csa_tree_add_83_21_pad_groupi_n_1014 ,csa_tree_add_83_21_pad_groupi_n_1013);
  not csa_tree_add_83_21_pad_groupi_g4705(csa_tree_add_83_21_pad_groupi_n_1010 ,csa_tree_add_83_21_pad_groupi_n_1009);
  nor csa_tree_add_83_21_pad_groupi_g4706__1705(csa_tree_add_83_21_pad_groupi_n_1008 ,csa_tree_add_83_21_pad_groupi_n_841 ,csa_tree_add_83_21_pad_groupi_n_930);
  or csa_tree_add_83_21_pad_groupi_g4707__5122(csa_tree_add_83_21_pad_groupi_n_1007 ,csa_tree_add_83_21_pad_groupi_n_843 ,csa_tree_add_83_21_pad_groupi_n_917);
  nor csa_tree_add_83_21_pad_groupi_g4708__8246(csa_tree_add_83_21_pad_groupi_n_1006 ,csa_tree_add_83_21_pad_groupi_n_824 ,csa_tree_add_83_21_pad_groupi_n_872);
  and csa_tree_add_83_21_pad_groupi_g4709__7098(csa_tree_add_83_21_pad_groupi_n_1005 ,csa_tree_add_83_21_pad_groupi_n_840 ,csa_tree_add_83_21_pad_groupi_n_922);
  and csa_tree_add_83_21_pad_groupi_g4710__6131(csa_tree_add_83_21_pad_groupi_n_1004 ,csa_tree_add_83_21_pad_groupi_n_839 ,csa_tree_add_83_21_pad_groupi_n_909);
  and csa_tree_add_83_21_pad_groupi_g4711__1881(csa_tree_add_83_21_pad_groupi_n_1003 ,csa_tree_add_83_21_pad_groupi_n_770 ,csa_tree_add_83_21_pad_groupi_n_916);
  or csa_tree_add_83_21_pad_groupi_g4712__5115(csa_tree_add_83_21_pad_groupi_n_1002 ,csa_tree_add_83_21_pad_groupi_n_779 ,csa_tree_add_83_21_pad_groupi_n_902);
  and csa_tree_add_83_21_pad_groupi_g4713__7482(csa_tree_add_83_21_pad_groupi_n_1001 ,csa_tree_add_83_21_pad_groupi_n_769 ,csa_tree_add_83_21_pad_groupi_n_904);
  and csa_tree_add_83_21_pad_groupi_g4714__4733(csa_tree_add_83_21_pad_groupi_n_1000 ,csa_tree_add_83_21_pad_groupi_n_820 ,csa_tree_add_83_21_pad_groupi_n_935);
  nor csa_tree_add_83_21_pad_groupi_g4715__6161(csa_tree_add_83_21_pad_groupi_n_999 ,csa_tree_add_83_21_pad_groupi_n_834 ,csa_tree_add_83_21_pad_groupi_n_896);
  or csa_tree_add_83_21_pad_groupi_g4716__9315(csa_tree_add_83_21_pad_groupi_n_998 ,csa_tree_add_83_21_pad_groupi_n_820 ,csa_tree_add_83_21_pad_groupi_n_935);
  and csa_tree_add_83_21_pad_groupi_g4717__9945(csa_tree_add_83_21_pad_groupi_n_997 ,csa_tree_add_83_21_pad_groupi_n_830 ,csa_tree_add_83_21_pad_groupi_n_856);
  or csa_tree_add_83_21_pad_groupi_g4718__2883(csa_tree_add_83_21_pad_groupi_n_996 ,csa_tree_add_83_21_pad_groupi_n_936 ,csa_tree_add_83_21_pad_groupi_n_919);
  and csa_tree_add_83_21_pad_groupi_g4719__2346(csa_tree_add_83_21_pad_groupi_n_995 ,csa_tree_add_83_21_pad_groupi_n_775 ,csa_tree_add_83_21_pad_groupi_n_891);
  or csa_tree_add_83_21_pad_groupi_g4720__1666(csa_tree_add_83_21_pad_groupi_n_994 ,csa_tree_add_83_21_pad_groupi_n_892 ,csa_tree_add_83_21_pad_groupi_n_894);
  and csa_tree_add_83_21_pad_groupi_g4721__7410(csa_tree_add_83_21_pad_groupi_n_993 ,csa_tree_add_83_21_pad_groupi_n_768 ,csa_tree_add_83_21_pad_groupi_n_924);
  and csa_tree_add_83_21_pad_groupi_g4722__6417(csa_tree_add_83_21_pad_groupi_n_992 ,csa_tree_add_83_21_pad_groupi_n_780 ,csa_tree_add_83_21_pad_groupi_n_885);
  nor csa_tree_add_83_21_pad_groupi_g4723__5477(csa_tree_add_83_21_pad_groupi_n_991 ,csa_tree_add_83_21_pad_groupi_n_837 ,csa_tree_add_83_21_pad_groupi_n_877);
  and csa_tree_add_83_21_pad_groupi_g4724__2398(csa_tree_add_83_21_pad_groupi_n_990 ,csa_tree_add_83_21_pad_groupi_n_777 ,csa_tree_add_83_21_pad_groupi_n_928);
  or csa_tree_add_83_21_pad_groupi_g4725__5107(csa_tree_add_83_21_pad_groupi_n_989 ,csa_tree_add_83_21_pad_groupi_n_838 ,csa_tree_add_83_21_pad_groupi_n_875);
  nor csa_tree_add_83_21_pad_groupi_g4726__6260(csa_tree_add_83_21_pad_groupi_n_988 ,csa_tree_add_83_21_pad_groupi_n_774 ,csa_tree_add_83_21_pad_groupi_n_855);
  nor csa_tree_add_83_21_pad_groupi_g4727__4319(csa_tree_add_83_21_pad_groupi_n_987 ,csa_tree_add_83_21_pad_groupi_n_776 ,csa_tree_add_83_21_pad_groupi_n_883);
  and csa_tree_add_83_21_pad_groupi_g4728__8428(csa_tree_add_83_21_pad_groupi_n_986 ,csa_tree_add_83_21_pad_groupi_n_773 ,csa_tree_add_83_21_pad_groupi_n_863);
  or csa_tree_add_83_21_pad_groupi_g4729__5526(csa_tree_add_83_21_pad_groupi_n_985 ,csa_tree_add_83_21_pad_groupi_n_823 ,csa_tree_add_83_21_pad_groupi_n_862);
  nor csa_tree_add_83_21_pad_groupi_g4730__6783(csa_tree_add_83_21_pad_groupi_n_984 ,csa_tree_add_83_21_pad_groupi_n_772 ,csa_tree_add_83_21_pad_groupi_n_859);
  nor csa_tree_add_83_21_pad_groupi_g4731__3680(csa_tree_add_83_21_pad_groupi_n_983 ,csa_tree_add_83_21_pad_groupi_n_771 ,csa_tree_add_83_21_pad_groupi_n_900);
  or csa_tree_add_83_21_pad_groupi_g4732__1617(csa_tree_add_83_21_pad_groupi_n_982 ,csa_tree_add_83_21_pad_groupi_n_835 ,csa_tree_add_83_21_pad_groupi_n_851);
  or csa_tree_add_83_21_pad_groupi_g4733__2802(csa_tree_add_83_21_pad_groupi_n_981 ,csa_tree_add_83_21_pad_groupi_n_893 ,csa_tree_add_83_21_pad_groupi_n_920);
  xnor csa_tree_add_83_21_pad_groupi_g4734__1705(csa_tree_add_83_21_pad_groupi_n_980 ,csa_tree_add_83_21_pad_groupi_n_846 ,csa_tree_add_83_21_pad_groupi_n_848);
  and csa_tree_add_83_21_pad_groupi_g4735__5122(csa_tree_add_83_21_pad_groupi_n_979 ,csa_tree_add_83_21_pad_groupi_n_827 ,csa_tree_add_83_21_pad_groupi_n_927);
  or csa_tree_add_83_21_pad_groupi_g4736__8246(csa_tree_add_83_21_pad_groupi_n_1024 ,csa_tree_add_83_21_pad_groupi_n_19 ,csa_tree_add_83_21_pad_groupi_n_898);
  xnor csa_tree_add_83_21_pad_groupi_g4737__7098(csa_tree_add_83_21_pad_groupi_n_1022 ,csa_tree_add_83_21_pad_groupi_n_706 ,csa_tree_add_83_21_pad_groupi_n_844);
  xnor csa_tree_add_83_21_pad_groupi_g4739__6131(csa_tree_add_83_21_pad_groupi_n_1021 ,csa_tree_add_83_21_pad_groupi_n_711 ,in8[9]);
  xnor csa_tree_add_83_21_pad_groupi_g4740__1881(csa_tree_add_83_21_pad_groupi_n_1020 ,csa_tree_add_83_21_pad_groupi_n_645 ,csa_tree_add_83_21_pad_groupi_n_832);
  and csa_tree_add_83_21_pad_groupi_g4741__5115(csa_tree_add_83_21_pad_groupi_n_1019 ,csa_tree_add_83_21_pad_groupi_n_899 ,csa_tree_add_83_21_pad_groupi_n_359);
  and csa_tree_add_83_21_pad_groupi_g4742__7482(csa_tree_add_83_21_pad_groupi_n_1017 ,csa_tree_add_83_21_pad_groupi_n_656 ,csa_tree_add_83_21_pad_groupi_n_923);
  or csa_tree_add_83_21_pad_groupi_g4743__4733(csa_tree_add_83_21_pad_groupi_n_1015 ,csa_tree_add_83_21_pad_groupi_n_682 ,csa_tree_add_83_21_pad_groupi_n_881);
  or csa_tree_add_83_21_pad_groupi_g4744__6161(csa_tree_add_83_21_pad_groupi_n_1013 ,csa_tree_add_83_21_pad_groupi_n_666 ,csa_tree_add_83_21_pad_groupi_n_861);
  xnor csa_tree_add_83_21_pad_groupi_g4745__9315(csa_tree_add_83_21_pad_groupi_n_1012 ,csa_tree_add_83_21_pad_groupi_n_704 ,csa_tree_add_83_21_pad_groupi_n_767);
  xnor csa_tree_add_83_21_pad_groupi_g4746__9945(csa_tree_add_83_21_pad_groupi_n_1011 ,csa_tree_add_83_21_pad_groupi_n_831 ,csa_tree_add_83_21_pad_groupi_n_1);
  or csa_tree_add_83_21_pad_groupi_g4747__2883(csa_tree_add_83_21_pad_groupi_n_1009 ,csa_tree_add_83_21_pad_groupi_n_702 ,csa_tree_add_83_21_pad_groupi_n_931);
  xnor csa_tree_add_83_21_pad_groupi_g4748__2346(csa_tree_add_83_21_pad_groupi_n_974 ,csa_tree_add_83_21_pad_groupi_n_726 ,csa_tree_add_83_21_pad_groupi_n_821);
  xnor csa_tree_add_83_21_pad_groupi_g4749__1666(csa_tree_add_83_21_pad_groupi_n_973 ,csa_tree_add_83_21_pad_groupi_n_802 ,csa_tree_add_83_21_pad_groupi_n_795);
  xnor csa_tree_add_83_21_pad_groupi_g4750__7410(csa_tree_add_83_21_pad_groupi_n_972 ,csa_tree_add_83_21_pad_groupi_n_837 ,csa_tree_add_83_21_pad_groupi_n_766);
  xnor csa_tree_add_83_21_pad_groupi_g4751__6417(csa_tree_add_83_21_pad_groupi_n_971 ,csa_tree_add_83_21_pad_groupi_n_829 ,in8[12]);
  xnor csa_tree_add_83_21_pad_groupi_g4752__5477(csa_tree_add_83_21_pad_groupi_n_970 ,csa_tree_add_83_21_pad_groupi_n_739 ,csa_tree_add_83_21_pad_groupi_n_728);
  xnor csa_tree_add_83_21_pad_groupi_g4753__2398(csa_tree_add_83_21_pad_groupi_n_969 ,csa_tree_add_83_21_pad_groupi_n_758 ,csa_tree_add_83_21_pad_groupi_n_757);
  xor csa_tree_add_83_21_pad_groupi_g4754__5107(csa_tree_add_83_21_pad_groupi_n_968 ,csa_tree_add_83_21_pad_groupi_n_824 ,csa_tree_add_83_21_pad_groupi_n_809);
  xor csa_tree_add_83_21_pad_groupi_g4755__6260(csa_tree_add_83_21_pad_groupi_n_967 ,csa_tree_add_83_21_pad_groupi_n_834 ,in8[8]);
  xnor csa_tree_add_83_21_pad_groupi_g4756__4319(csa_tree_add_83_21_pad_groupi_n_966 ,csa_tree_add_83_21_pad_groupi_n_733 ,csa_tree_add_83_21_pad_groupi_n_755);
  xnor csa_tree_add_83_21_pad_groupi_g4757__8428(csa_tree_add_83_21_pad_groupi_n_965 ,csa_tree_add_83_21_pad_groupi_n_800 ,csa_tree_add_83_21_pad_groupi_n_799);
  xor csa_tree_add_83_21_pad_groupi_g4758__5526(csa_tree_add_83_21_pad_groupi_n_964 ,csa_tree_add_83_21_pad_groupi_n_776 ,csa_tree_add_83_21_pad_groupi_n_721);
  xor csa_tree_add_83_21_pad_groupi_g4759__6783(csa_tree_add_83_21_pad_groupi_n_963 ,csa_tree_add_83_21_pad_groupi_n_772 ,in8[1]);
  xnor csa_tree_add_83_21_pad_groupi_g4760__3680(csa_tree_add_83_21_pad_groupi_n_962 ,csa_tree_add_83_21_pad_groupi_n_765 ,csa_tree_add_83_21_pad_groupi_n_751);
  xnor csa_tree_add_83_21_pad_groupi_g4761__1617(csa_tree_add_83_21_pad_groupi_n_961 ,csa_tree_add_83_21_pad_groupi_n_735 ,csa_tree_add_83_21_pad_groupi_n_792);
  xor csa_tree_add_83_21_pad_groupi_g4762__2802(csa_tree_add_83_21_pad_groupi_n_960 ,csa_tree_add_83_21_pad_groupi_n_771 ,csa_tree_add_83_21_pad_groupi_n_729);
  xnor csa_tree_add_83_21_pad_groupi_g4763__1705(csa_tree_add_83_21_pad_groupi_n_959 ,csa_tree_add_83_21_pad_groupi_n_725 ,csa_tree_add_83_21_pad_groupi_n_723);
  xnor csa_tree_add_83_21_pad_groupi_g4764__5122(csa_tree_add_83_21_pad_groupi_n_958 ,csa_tree_add_83_21_pad_groupi_n_814 ,csa_tree_add_83_21_pad_groupi_n_796);
  xnor csa_tree_add_83_21_pad_groupi_g4765__8246(csa_tree_add_83_21_pad_groupi_n_957 ,csa_tree_add_83_21_pad_groupi_n_784 ,csa_tree_add_83_21_pad_groupi_n_747);
  xor csa_tree_add_83_21_pad_groupi_g4766__7098(csa_tree_add_83_21_pad_groupi_n_956 ,csa_tree_add_83_21_pad_groupi_n_841 ,csa_tree_add_83_21_pad_groupi_n_748);
  xnor csa_tree_add_83_21_pad_groupi_g4767__6131(csa_tree_add_83_21_pad_groupi_n_955 ,csa_tree_add_83_21_pad_groupi_n_760 ,csa_tree_add_83_21_pad_groupi_n_737);
  xnor csa_tree_add_83_21_pad_groupi_g4768__1881(csa_tree_add_83_21_pad_groupi_n_954 ,csa_tree_add_83_21_pad_groupi_n_756 ,in8[2]);
  xnor csa_tree_add_83_21_pad_groupi_g4769__5115(csa_tree_add_83_21_pad_groupi_n_953 ,csa_tree_add_83_21_pad_groupi_n_763 ,csa_tree_add_83_21_pad_groupi_n_817);
  xor csa_tree_add_83_21_pad_groupi_g4770__7482(csa_tree_add_83_21_pad_groupi_n_952 ,csa_tree_add_83_21_pad_groupi_n_823 ,csa_tree_add_83_21_pad_groupi_n_742);
  xnor csa_tree_add_83_21_pad_groupi_g4771__4733(csa_tree_add_83_21_pad_groupi_n_951 ,csa_tree_add_83_21_pad_groupi_n_806 ,csa_tree_add_83_21_pad_groupi_n_753);
  xnor csa_tree_add_83_21_pad_groupi_g4772__6161(csa_tree_add_83_21_pad_groupi_n_950 ,csa_tree_add_83_21_pad_groupi_n_790 ,csa_tree_add_83_21_pad_groupi_n_819);
  xnor csa_tree_add_83_21_pad_groupi_g4773__9315(csa_tree_add_83_21_pad_groupi_n_949 ,csa_tree_add_83_21_pad_groupi_n_813 ,csa_tree_add_83_21_pad_groupi_n_716);
  xnor csa_tree_add_83_21_pad_groupi_g4774__9945(csa_tree_add_83_21_pad_groupi_n_948 ,csa_tree_add_83_21_pad_groupi_n_731 ,in8[6]);
  xnor csa_tree_add_83_21_pad_groupi_g4775__2883(csa_tree_add_83_21_pad_groupi_n_947 ,csa_tree_add_83_21_pad_groupi_n_787 ,in8[5]);
  xnor csa_tree_add_83_21_pad_groupi_g4776__2346(csa_tree_add_83_21_pad_groupi_n_946 ,csa_tree_add_83_21_pad_groupi_n_713 ,in8[7]);
  xnor csa_tree_add_83_21_pad_groupi_g4777__1666(csa_tree_add_83_21_pad_groupi_n_945 ,csa_tree_add_83_21_pad_groupi_n_808 ,csa_tree_add_83_21_pad_groupi_n_788);
  xnor csa_tree_add_83_21_pad_groupi_g4778__7410(csa_tree_add_83_21_pad_groupi_n_944 ,csa_tree_add_83_21_pad_groupi_n_761 ,csa_tree_add_83_21_pad_groupi_n_786);
  xnor csa_tree_add_83_21_pad_groupi_g4779__6417(csa_tree_add_83_21_pad_groupi_n_943 ,csa_tree_add_83_21_pad_groupi_n_798 ,in8[4]);
  xnor csa_tree_add_83_21_pad_groupi_g4780__5477(csa_tree_add_83_21_pad_groupi_n_942 ,csa_tree_add_83_21_pad_groupi_n_719 ,csa_tree_add_83_21_pad_groupi_n_720);
  xnor csa_tree_add_83_21_pad_groupi_g4781__2398(csa_tree_add_83_21_pad_groupi_n_941 ,csa_tree_add_83_21_pad_groupi_n_815 ,csa_tree_add_83_21_pad_groupi_n_717);
  xnor csa_tree_add_83_21_pad_groupi_g4782__5107(csa_tree_add_83_21_pad_groupi_n_940 ,csa_tree_add_83_21_pad_groupi_n_807 ,csa_tree_add_83_21_pad_groupi_n_714);
  xnor csa_tree_add_83_21_pad_groupi_g4783__6260(csa_tree_add_83_21_pad_groupi_n_939 ,csa_tree_add_83_21_pad_groupi_n_810 ,csa_tree_add_83_21_pad_groupi_n_811);
  xnor csa_tree_add_83_21_pad_groupi_g4784__4319(csa_tree_add_83_21_pad_groupi_n_938 ,csa_tree_add_83_21_pad_groupi_n_804 ,in8[3]);
  xnor csa_tree_add_83_21_pad_groupi_g4785__8428(csa_tree_add_83_21_pad_groupi_n_937 ,csa_tree_add_83_21_pad_groupi_n_718 ,csa_tree_add_83_21_pad_groupi_n_793);
  xnor csa_tree_add_83_21_pad_groupi_g4786__5526(csa_tree_add_83_21_pad_groupi_n_977 ,csa_tree_add_83_21_pad_groupi_n_822 ,csa_tree_add_83_21_pad_groupi_n_709);
  xnor csa_tree_add_83_21_pad_groupi_g4787__6783(csa_tree_add_83_21_pad_groupi_n_976 ,csa_tree_add_83_21_pad_groupi_n_828 ,csa_tree_add_83_21_pad_groupi_n_710);
  xnor csa_tree_add_83_21_pad_groupi_g4788__3680(csa_tree_add_83_21_pad_groupi_n_975 ,csa_tree_add_83_21_pad_groupi_n_825 ,in8[0]);
  or csa_tree_add_83_21_pad_groupi_g4791__1617(csa_tree_add_83_21_pad_groupi_n_932 ,csa_tree_add_83_21_pad_groupi_n_815 ,csa_tree_add_83_21_pad_groupi_n_717);
  nor csa_tree_add_83_21_pad_groupi_g4792__2802(csa_tree_add_83_21_pad_groupi_n_931 ,csa_tree_add_83_21_pad_groupi_n_673 ,csa_tree_add_83_21_pad_groupi_n_831);
  nor csa_tree_add_83_21_pad_groupi_g4793__1705(csa_tree_add_83_21_pad_groupi_n_930 ,csa_tree_add_83_21_pad_groupi_n_748 ,csa_tree_add_83_21_pad_groupi_n_785);
  nor csa_tree_add_83_21_pad_groupi_g4794__5122(csa_tree_add_83_21_pad_groupi_n_929 ,csa_tree_add_83_21_pad_groupi_n_802 ,csa_tree_add_83_21_pad_groupi_n_794);
  or csa_tree_add_83_21_pad_groupi_g4795__8246(csa_tree_add_83_21_pad_groupi_n_928 ,csa_tree_add_83_21_pad_groupi_n_807 ,csa_tree_add_83_21_pad_groupi_n_714);
  or csa_tree_add_83_21_pad_groupi_g4796__7098(csa_tree_add_83_21_pad_groupi_n_927 ,csa_tree_add_83_21_pad_groupi_n_801 ,csa_tree_add_83_21_pad_groupi_n_795);
  nor csa_tree_add_83_21_pad_groupi_g4797__6131(csa_tree_add_83_21_pad_groupi_n_926 ,csa_tree_add_83_21_pad_groupi_n_766 ,csa_tree_add_83_21_pad_groupi_n_744);
  and csa_tree_add_83_21_pad_groupi_g4798__1881(csa_tree_add_83_21_pad_groupi_n_925 ,csa_tree_add_83_21_pad_groupi_n_764 ,csa_tree_add_83_21_pad_groupi_n_809);
  or csa_tree_add_83_21_pad_groupi_g4799__5115(csa_tree_add_83_21_pad_groupi_n_924 ,csa_tree_add_83_21_pad_groupi_n_719 ,csa_tree_add_83_21_pad_groupi_n_720);
  or csa_tree_add_83_21_pad_groupi_g4800__7482(csa_tree_add_83_21_pad_groupi_n_923 ,csa_tree_add_83_21_pad_groupi_n_593 ,csa_tree_add_83_21_pad_groupi_n_836);
  or csa_tree_add_83_21_pad_groupi_g4801__4733(csa_tree_add_83_21_pad_groupi_n_922 ,csa_tree_add_83_21_pad_groupi_n_800 ,csa_tree_add_83_21_pad_groupi_n_799);
  or csa_tree_add_83_21_pad_groupi_g4802__6161(csa_tree_add_83_21_pad_groupi_n_921 ,csa_tree_add_83_21_pad_groupi_n_789 ,csa_tree_add_83_21_pad_groupi_n_818);
  nor csa_tree_add_83_21_pad_groupi_g4803__9315(csa_tree_add_83_21_pad_groupi_n_920 ,csa_tree_add_83_21_pad_groupi_n_725 ,csa_tree_add_83_21_pad_groupi_n_723);
  nor csa_tree_add_83_21_pad_groupi_g4804__9945(csa_tree_add_83_21_pad_groupi_n_919 ,csa_tree_add_83_21_pad_groupi_n_763 ,csa_tree_add_83_21_pad_groupi_n_817);
  nor csa_tree_add_83_21_pad_groupi_g4805__2883(csa_tree_add_83_21_pad_groupi_n_918 ,csa_tree_add_83_21_pad_groupi_n_790 ,csa_tree_add_83_21_pad_groupi_n_819);
  nor csa_tree_add_83_21_pad_groupi_g4806__2346(csa_tree_add_83_21_pad_groupi_n_917 ,csa_tree_add_83_21_pad_groupi_n_806 ,csa_tree_add_83_21_pad_groupi_n_753);
  or csa_tree_add_83_21_pad_groupi_g4807__1666(csa_tree_add_83_21_pad_groupi_n_916 ,in8[5] ,csa_tree_add_83_21_pad_groupi_n_787);
  or csa_tree_add_83_21_pad_groupi_g4808__7410(csa_tree_add_83_21_pad_groupi_n_915 ,csa_tree_add_83_21_pad_groupi_n_762 ,csa_tree_add_83_21_pad_groupi_n_816);
  and csa_tree_add_83_21_pad_groupi_g4809__6417(csa_tree_add_83_21_pad_groupi_n_914 ,csa_tree_add_83_21_pad_groupi_n_815 ,csa_tree_add_83_21_pad_groupi_n_717);
  or csa_tree_add_83_21_pad_groupi_g4810__5477(csa_tree_add_83_21_pad_groupi_n_913 ,csa_tree_add_83_21_pad_groupi_n_805 ,csa_tree_add_83_21_pad_groupi_n_752);
  or csa_tree_add_83_21_pad_groupi_g4811__2398(csa_tree_add_83_21_pad_groupi_n_912 ,csa_tree_add_83_21_pad_groupi_n_812 ,csa_tree_add_83_21_pad_groupi_n_715);
  and csa_tree_add_83_21_pad_groupi_g4812__5107(csa_tree_add_83_21_pad_groupi_n_911 ,csa_tree_add_83_21_pad_groupi_n_748 ,csa_tree_add_83_21_pad_groupi_n_785);
  nor csa_tree_add_83_21_pad_groupi_g4813__6260(csa_tree_add_83_21_pad_groupi_n_910 ,csa_tree_add_83_21_pad_groupi_n_372 ,csa_tree_add_83_21_pad_groupi_n_782);
  or csa_tree_add_83_21_pad_groupi_g4814__4319(csa_tree_add_83_21_pad_groupi_n_909 ,csa_tree_add_83_21_pad_groupi_n_814 ,csa_tree_add_83_21_pad_groupi_n_796);
  and csa_tree_add_83_21_pad_groupi_g4815__8428(csa_tree_add_83_21_pad_groupi_n_908 ,csa_tree_add_83_21_pad_groupi_n_810 ,csa_tree_add_83_21_pad_groupi_n_811);
  and csa_tree_add_83_21_pad_groupi_g4816__5526(csa_tree_add_83_21_pad_groupi_n_907 ,csa_tree_add_83_21_pad_groupi_n_807 ,csa_tree_add_83_21_pad_groupi_n_714);
  and csa_tree_add_83_21_pad_groupi_g4817__6783(csa_tree_add_83_21_pad_groupi_n_906 ,in8[4] ,csa_tree_add_83_21_pad_groupi_n_798);
  and csa_tree_add_83_21_pad_groupi_g4818__3680(csa_tree_add_83_21_pad_groupi_n_905 ,in8[5] ,csa_tree_add_83_21_pad_groupi_n_787);
  or csa_tree_add_83_21_pad_groupi_g4819__1617(csa_tree_add_83_21_pad_groupi_n_904 ,csa_tree_add_83_21_pad_groupi_n_808 ,csa_tree_add_83_21_pad_groupi_n_788);
  and csa_tree_add_83_21_pad_groupi_g4820__2802(csa_tree_add_83_21_pad_groupi_n_903 ,csa_tree_add_83_21_pad_groupi_n_814 ,csa_tree_add_83_21_pad_groupi_n_796);
  nor csa_tree_add_83_21_pad_groupi_g4821__1705(csa_tree_add_83_21_pad_groupi_n_902 ,csa_tree_add_83_21_pad_groupi_n_813 ,csa_tree_add_83_21_pad_groupi_n_716);
  and csa_tree_add_83_21_pad_groupi_g4822__5122(csa_tree_add_83_21_pad_groupi_n_901 ,csa_tree_add_83_21_pad_groupi_n_761 ,csa_tree_add_83_21_pad_groupi_n_786);
  nor csa_tree_add_83_21_pad_groupi_g4823__8246(csa_tree_add_83_21_pad_groupi_n_900 ,csa_tree_add_83_21_pad_groupi_n_783 ,csa_tree_add_83_21_pad_groupi_n_729);
  or csa_tree_add_83_21_pad_groupi_g4824__7098(csa_tree_add_83_21_pad_groupi_n_899 ,csa_tree_add_83_21_pad_groupi_n_708 ,csa_tree_add_83_21_pad_groupi_n_845);
  or csa_tree_add_83_21_pad_groupi_g4825__6131(csa_tree_add_83_21_pad_groupi_n_898 ,csa_tree_add_83_21_pad_groupi_n_112 ,csa_tree_add_83_21_pad_groupi_n_781);
  and csa_tree_add_83_21_pad_groupi_g4826__1881(csa_tree_add_83_21_pad_groupi_n_897 ,csa_tree_add_83_21_pad_groupi_n_783 ,csa_tree_add_83_21_pad_groupi_n_729);
  and csa_tree_add_83_21_pad_groupi_g4827__5115(csa_tree_add_83_21_pad_groupi_n_896 ,csa_tree_add_83_21_pad_groupi_n_372 ,csa_tree_add_83_21_pad_groupi_n_782);
  or csa_tree_add_83_21_pad_groupi_g4828__7482(csa_tree_add_83_21_pad_groupi_n_895 ,csa_tree_add_83_21_pad_groupi_n_734 ,csa_tree_add_83_21_pad_groupi_n_791);
  nor csa_tree_add_83_21_pad_groupi_g4829__4733(csa_tree_add_83_21_pad_groupi_n_894 ,csa_tree_add_83_21_pad_groupi_n_735 ,csa_tree_add_83_21_pad_groupi_n_792);
  or csa_tree_add_83_21_pad_groupi_g4830__6161(csa_tree_add_83_21_pad_groupi_n_936 ,csa_tree_add_83_21_pad_groupi_n_645 ,csa_tree_add_83_21_pad_groupi_n_833);
  and csa_tree_add_83_21_pad_groupi_g4831__9315(csa_tree_add_83_21_pad_groupi_n_935 ,csa_tree_add_83_21_pad_groupi_n_705 ,csa_tree_add_83_21_pad_groupi_n_767);
  and csa_tree_add_83_21_pad_groupi_g4832__9945(csa_tree_add_83_21_pad_groupi_n_934 ,csa_tree_add_83_21_pad_groupi_n_708 ,csa_tree_add_83_21_pad_groupi_n_845);
  and csa_tree_add_83_21_pad_groupi_g4833__2883(csa_tree_add_83_21_pad_groupi_n_933 ,csa_tree_add_83_21_pad_groupi_n_707 ,csa_tree_add_83_21_pad_groupi_n_844);
  or csa_tree_add_83_21_pad_groupi_g4834__2346(csa_tree_add_83_21_pad_groupi_n_891 ,csa_tree_add_83_21_pad_groupi_n_718 ,csa_tree_add_83_21_pad_groupi_n_793);
  and csa_tree_add_83_21_pad_groupi_g4835__1666(csa_tree_add_83_21_pad_groupi_n_890 ,csa_tree_add_83_21_pad_groupi_n_800 ,csa_tree_add_83_21_pad_groupi_n_799);
  and csa_tree_add_83_21_pad_groupi_g4836__7410(csa_tree_add_83_21_pad_groupi_n_889 ,csa_tree_add_83_21_pad_groupi_n_718 ,csa_tree_add_83_21_pad_groupi_n_793);
  or csa_tree_add_83_21_pad_groupi_g4837__6417(csa_tree_add_83_21_pad_groupi_n_888 ,csa_tree_add_83_21_pad_groupi_n_732 ,csa_tree_add_83_21_pad_groupi_n_754);
  and csa_tree_add_83_21_pad_groupi_g4838__5477(csa_tree_add_83_21_pad_groupi_n_887 ,in8[3] ,csa_tree_add_83_21_pad_groupi_n_804);
  and csa_tree_add_83_21_pad_groupi_g4839__2398(csa_tree_add_83_21_pad_groupi_n_886 ,csa_tree_add_83_21_pad_groupi_n_719 ,csa_tree_add_83_21_pad_groupi_n_720);
  or csa_tree_add_83_21_pad_groupi_g4840__5107(csa_tree_add_83_21_pad_groupi_n_885 ,in8[3] ,csa_tree_add_83_21_pad_groupi_n_804);
  or csa_tree_add_83_21_pad_groupi_g4841__6260(csa_tree_add_83_21_pad_groupi_n_884 ,csa_tree_add_83_21_pad_groupi_n_738 ,csa_tree_add_83_21_pad_groupi_n_727);
  nor csa_tree_add_83_21_pad_groupi_g4842__4319(csa_tree_add_83_21_pad_groupi_n_883 ,csa_tree_add_83_21_pad_groupi_n_803 ,csa_tree_add_83_21_pad_groupi_n_721);
  nor csa_tree_add_83_21_pad_groupi_g4843__8428(csa_tree_add_83_21_pad_groupi_n_882 ,csa_tree_add_83_21_pad_groupi_n_739 ,csa_tree_add_83_21_pad_groupi_n_728);
  nor csa_tree_add_83_21_pad_groupi_g4844__5526(csa_tree_add_83_21_pad_groupi_n_881 ,csa_tree_add_83_21_pad_groupi_n_700 ,csa_tree_add_83_21_pad_groupi_n_828);
  or csa_tree_add_83_21_pad_groupi_g4845__6783(csa_tree_add_83_21_pad_groupi_n_880 ,csa_tree_add_83_21_pad_groupi_n_761 ,csa_tree_add_83_21_pad_groupi_n_786);
  nor csa_tree_add_83_21_pad_groupi_g4846__3680(csa_tree_add_83_21_pad_groupi_n_879 ,csa_tree_add_83_21_pad_groupi_n_371 ,csa_tree_add_83_21_pad_groupi_n_740);
  or csa_tree_add_83_21_pad_groupi_g4847__1617(csa_tree_add_83_21_pad_groupi_n_878 ,csa_tree_add_83_21_pad_groupi_n_387 ,csa_tree_add_83_21_pad_groupi_n_712);
  and csa_tree_add_83_21_pad_groupi_g4848__2802(csa_tree_add_83_21_pad_groupi_n_877 ,csa_tree_add_83_21_pad_groupi_n_766 ,csa_tree_add_83_21_pad_groupi_n_744);
  nor csa_tree_add_83_21_pad_groupi_g4849__1705(csa_tree_add_83_21_pad_groupi_n_876 ,csa_tree_add_83_21_pad_groupi_n_733 ,csa_tree_add_83_21_pad_groupi_n_755);
  nor csa_tree_add_83_21_pad_groupi_g4850__5122(csa_tree_add_83_21_pad_groupi_n_875 ,in8[7] ,csa_tree_add_83_21_pad_groupi_n_713);
  and csa_tree_add_83_21_pad_groupi_g4851__8246(csa_tree_add_83_21_pad_groupi_n_874 ,csa_tree_add_83_21_pad_groupi_n_803 ,csa_tree_add_83_21_pad_groupi_n_721);
  and csa_tree_add_83_21_pad_groupi_g4852__7098(csa_tree_add_83_21_pad_groupi_n_873 ,csa_tree_add_83_21_pad_groupi_n_758 ,csa_tree_add_83_21_pad_groupi_n_757);
  nor csa_tree_add_83_21_pad_groupi_g4853__6131(csa_tree_add_83_21_pad_groupi_n_872 ,csa_tree_add_83_21_pad_groupi_n_764 ,csa_tree_add_83_21_pad_groupi_n_809);
  or csa_tree_add_83_21_pad_groupi_g4854__1881(csa_tree_add_83_21_pad_groupi_n_871 ,csa_tree_add_83_21_pad_groupi_n_758 ,csa_tree_add_83_21_pad_groupi_n_757);
  and csa_tree_add_83_21_pad_groupi_g4855__5115(csa_tree_add_83_21_pad_groupi_n_870 ,in8[2] ,csa_tree_add_83_21_pad_groupi_n_756);
  and csa_tree_add_83_21_pad_groupi_g4856__7482(csa_tree_add_83_21_pad_groupi_n_869 ,csa_tree_add_83_21_pad_groupi_n_808 ,csa_tree_add_83_21_pad_groupi_n_788);
  and csa_tree_add_83_21_pad_groupi_g4857__4733(csa_tree_add_83_21_pad_groupi_n_868 ,csa_tree_add_83_21_pad_groupi_n_784 ,csa_tree_add_83_21_pad_groupi_n_747);
  or csa_tree_add_83_21_pad_groupi_g4858__6161(csa_tree_add_83_21_pad_groupi_n_867 ,csa_tree_add_83_21_pad_groupi_n_810 ,csa_tree_add_83_21_pad_groupi_n_811);
  and csa_tree_add_83_21_pad_groupi_g4859__9315(csa_tree_add_83_21_pad_groupi_n_866 ,csa_tree_add_83_21_pad_groupi_n_765 ,csa_tree_add_83_21_pad_groupi_n_751);
  or csa_tree_add_83_21_pad_groupi_g4860__9945(csa_tree_add_83_21_pad_groupi_n_865 ,csa_tree_add_83_21_pad_groupi_n_784 ,csa_tree_add_83_21_pad_groupi_n_747);
  or csa_tree_add_83_21_pad_groupi_g4861__2883(csa_tree_add_83_21_pad_groupi_n_864 ,csa_tree_add_83_21_pad_groupi_n_749 ,csa_tree_add_83_21_pad_groupi_n_741);
  or csa_tree_add_83_21_pad_groupi_g4862__2346(csa_tree_add_83_21_pad_groupi_n_863 ,csa_tree_add_83_21_pad_groupi_n_765 ,csa_tree_add_83_21_pad_groupi_n_751);
  nor csa_tree_add_83_21_pad_groupi_g4863__1666(csa_tree_add_83_21_pad_groupi_n_862 ,csa_tree_add_83_21_pad_groupi_n_750 ,csa_tree_add_83_21_pad_groupi_n_742);
  nor csa_tree_add_83_21_pad_groupi_g4864__7410(csa_tree_add_83_21_pad_groupi_n_861 ,csa_tree_add_83_21_pad_groupi_n_600 ,csa_tree_add_83_21_pad_groupi_n_822);
  or csa_tree_add_83_21_pad_groupi_g4865__6417(csa_tree_add_83_21_pad_groupi_n_860 ,csa_tree_add_83_21_pad_groupi_n_726 ,csa_tree_add_83_21_pad_groupi_n_821);
  and csa_tree_add_83_21_pad_groupi_g4866__5477(csa_tree_add_83_21_pad_groupi_n_859 ,csa_tree_add_83_21_pad_groupi_n_371 ,csa_tree_add_83_21_pad_groupi_n_740);
  and csa_tree_add_83_21_pad_groupi_g4867__2398(csa_tree_add_83_21_pad_groupi_n_858 ,csa_tree_add_83_21_pad_groupi_n_726 ,csa_tree_add_83_21_pad_groupi_n_821);
  or csa_tree_add_83_21_pad_groupi_g4868__5107(csa_tree_add_83_21_pad_groupi_n_857 ,csa_tree_add_83_21_pad_groupi_n_759 ,csa_tree_add_83_21_pad_groupi_n_736);
  or csa_tree_add_83_21_pad_groupi_g4869__6260(csa_tree_add_83_21_pad_groupi_n_856 ,in8[4] ,csa_tree_add_83_21_pad_groupi_n_798);
  nor csa_tree_add_83_21_pad_groupi_g4870__4319(csa_tree_add_83_21_pad_groupi_n_855 ,in8[2] ,csa_tree_add_83_21_pad_groupi_n_756);
  nor csa_tree_add_83_21_pad_groupi_g4871__8428(csa_tree_add_83_21_pad_groupi_n_854 ,csa_tree_add_83_21_pad_groupi_n_760 ,csa_tree_add_83_21_pad_groupi_n_737);
  or csa_tree_add_83_21_pad_groupi_g4872__5526(csa_tree_add_83_21_pad_groupi_n_853 ,csa_tree_add_83_21_pad_groupi_n_370 ,csa_tree_add_83_21_pad_groupi_n_730);
  or csa_tree_add_83_21_pad_groupi_g4873__6783(csa_tree_add_83_21_pad_groupi_n_852 ,csa_tree_add_83_21_pad_groupi_n_724 ,csa_tree_add_83_21_pad_groupi_n_722);
  nor csa_tree_add_83_21_pad_groupi_g4874__3680(csa_tree_add_83_21_pad_groupi_n_851 ,in8[6] ,csa_tree_add_83_21_pad_groupi_n_731);
  or csa_tree_add_83_21_pad_groupi_g4876__1617(csa_tree_add_83_21_pad_groupi_n_893 ,csa_tree_add_83_21_pad_groupi_n_374 ,csa_tree_add_83_21_pad_groupi_n_826);
  or csa_tree_add_83_21_pad_groupi_g4877__2802(csa_tree_add_83_21_pad_groupi_n_892 ,csa_tree_add_83_21_pad_groupi_n_847 ,csa_tree_add_83_21_pad_groupi_n_849);
  not csa_tree_add_83_21_pad_groupi_g4878(csa_tree_add_83_21_pad_groupi_n_849 ,csa_tree_add_83_21_pad_groupi_n_848);
  not csa_tree_add_83_21_pad_groupi_g4879(csa_tree_add_83_21_pad_groupi_n_847 ,csa_tree_add_83_21_pad_groupi_n_846);
  not csa_tree_add_83_21_pad_groupi_g4880(csa_tree_add_83_21_pad_groupi_n_843 ,csa_tree_add_83_21_pad_groupi_n_842);
  not csa_tree_add_83_21_pad_groupi_g4883(csa_tree_add_83_21_pad_groupi_n_833 ,csa_tree_add_83_21_pad_groupi_n_832);
  not csa_tree_add_83_21_pad_groupi_g4884(csa_tree_add_83_21_pad_groupi_n_826 ,csa_tree_add_83_21_pad_groupi_n_825);
  not csa_tree_add_83_21_pad_groupi_g4885(csa_tree_add_83_21_pad_groupi_n_818 ,csa_tree_add_83_21_pad_groupi_n_819);
  not csa_tree_add_83_21_pad_groupi_g4886(csa_tree_add_83_21_pad_groupi_n_816 ,csa_tree_add_83_21_pad_groupi_n_817);
  not csa_tree_add_83_21_pad_groupi_g4887(csa_tree_add_83_21_pad_groupi_n_812 ,csa_tree_add_83_21_pad_groupi_n_813);
  not csa_tree_add_83_21_pad_groupi_g4888(csa_tree_add_83_21_pad_groupi_n_805 ,csa_tree_add_83_21_pad_groupi_n_806);
  not csa_tree_add_83_21_pad_groupi_g4889(csa_tree_add_83_21_pad_groupi_n_801 ,csa_tree_add_83_21_pad_groupi_n_802);
  not csa_tree_add_83_21_pad_groupi_g4890(csa_tree_add_83_21_pad_groupi_n_794 ,csa_tree_add_83_21_pad_groupi_n_795);
  not csa_tree_add_83_21_pad_groupi_g4891(csa_tree_add_83_21_pad_groupi_n_791 ,csa_tree_add_83_21_pad_groupi_n_792);
  not csa_tree_add_83_21_pad_groupi_g4892(csa_tree_add_83_21_pad_groupi_n_789 ,csa_tree_add_83_21_pad_groupi_n_790);
  and csa_tree_add_83_21_pad_groupi_g4893__1705(csa_tree_add_83_21_pad_groupi_n_781 ,csa_tree_add_83_21_pad_groupi_n_459 ,csa_tree_add_83_21_pad_groupi_n_612);
  or csa_tree_add_83_21_pad_groupi_g4894__5122(csa_tree_add_83_21_pad_groupi_n_848 ,csa_tree_add_83_21_pad_groupi_n_466 ,csa_tree_add_83_21_pad_groupi_n_621);
  or csa_tree_add_83_21_pad_groupi_g4895__8246(csa_tree_add_83_21_pad_groupi_n_846 ,csa_tree_add_83_21_pad_groupi_n_576 ,csa_tree_add_83_21_pad_groupi_n_703);
  and csa_tree_add_83_21_pad_groupi_g4896__7098(csa_tree_add_83_21_pad_groupi_n_845 ,csa_tree_add_83_21_pad_groupi_n_531 ,csa_tree_add_83_21_pad_groupi_n_685);
  or csa_tree_add_83_21_pad_groupi_g4897__6131(csa_tree_add_83_21_pad_groupi_n_844 ,csa_tree_add_83_21_pad_groupi_n_526 ,csa_tree_add_83_21_pad_groupi_n_652);
  or csa_tree_add_83_21_pad_groupi_g4898__1881(csa_tree_add_83_21_pad_groupi_n_842 ,csa_tree_add_83_21_pad_groupi_n_533 ,csa_tree_add_83_21_pad_groupi_n_618);
  and csa_tree_add_83_21_pad_groupi_g4899__5115(csa_tree_add_83_21_pad_groupi_n_841 ,csa_tree_add_83_21_pad_groupi_n_472 ,csa_tree_add_83_21_pad_groupi_n_642);
  or csa_tree_add_83_21_pad_groupi_g4900__7482(csa_tree_add_83_21_pad_groupi_n_840 ,csa_tree_add_83_21_pad_groupi_n_557 ,csa_tree_add_83_21_pad_groupi_n_598);
  or csa_tree_add_83_21_pad_groupi_g4901__4733(csa_tree_add_83_21_pad_groupi_n_839 ,csa_tree_add_83_21_pad_groupi_n_574 ,csa_tree_add_83_21_pad_groupi_n_588);
  and csa_tree_add_83_21_pad_groupi_g4903__6161(csa_tree_add_83_21_pad_groupi_n_837 ,csa_tree_add_83_21_pad_groupi_n_483 ,csa_tree_add_83_21_pad_groupi_n_587);
  and csa_tree_add_83_21_pad_groupi_g4906__9315(csa_tree_add_83_21_pad_groupi_n_834 ,csa_tree_add_83_21_pad_groupi_n_460 ,csa_tree_add_83_21_pad_groupi_n_586);
  or csa_tree_add_83_21_pad_groupi_g4907__9945(csa_tree_add_83_21_pad_groupi_n_832 ,csa_tree_add_83_21_pad_groupi_n_548 ,csa_tree_add_83_21_pad_groupi_n_699);
  or csa_tree_add_83_21_pad_groupi_g4912__2883(csa_tree_add_83_21_pad_groupi_n_827 ,csa_tree_add_83_21_pad_groupi_n_487 ,csa_tree_add_83_21_pad_groupi_n_647);
  or csa_tree_add_83_21_pad_groupi_g4913__2346(csa_tree_add_83_21_pad_groupi_n_825 ,csa_tree_add_83_21_pad_groupi_n_462 ,csa_tree_add_83_21_pad_groupi_n_662);
  and csa_tree_add_83_21_pad_groupi_g4914__1666(csa_tree_add_83_21_pad_groupi_n_824 ,csa_tree_add_83_21_pad_groupi_n_485 ,csa_tree_add_83_21_pad_groupi_n_683);
  and csa_tree_add_83_21_pad_groupi_g4915__7410(csa_tree_add_83_21_pad_groupi_n_823 ,csa_tree_add_83_21_pad_groupi_n_518 ,csa_tree_add_83_21_pad_groupi_n_595);
  or csa_tree_add_83_21_pad_groupi_g4917__6417(csa_tree_add_83_21_pad_groupi_n_821 ,csa_tree_add_83_21_pad_groupi_n_551 ,csa_tree_add_83_21_pad_groupi_n_665);
  or csa_tree_add_83_21_pad_groupi_g4918__5477(csa_tree_add_83_21_pad_groupi_n_820 ,csa_tree_add_83_21_pad_groupi_n_556 ,csa_tree_add_83_21_pad_groupi_n_677);
  or csa_tree_add_83_21_pad_groupi_g4919__2398(csa_tree_add_83_21_pad_groupi_n_819 ,csa_tree_add_83_21_pad_groupi_n_516 ,csa_tree_add_83_21_pad_groupi_n_681);
  or csa_tree_add_83_21_pad_groupi_g4920__5107(csa_tree_add_83_21_pad_groupi_n_817 ,csa_tree_add_83_21_pad_groupi_n_527 ,csa_tree_add_83_21_pad_groupi_n_674);
  or csa_tree_add_83_21_pad_groupi_g4921__6260(csa_tree_add_83_21_pad_groupi_n_815 ,csa_tree_add_83_21_pad_groupi_n_491 ,csa_tree_add_83_21_pad_groupi_n_649);
  or csa_tree_add_83_21_pad_groupi_g4922__4319(csa_tree_add_83_21_pad_groupi_n_814 ,csa_tree_add_83_21_pad_groupi_n_475 ,csa_tree_add_83_21_pad_groupi_n_633);
  or csa_tree_add_83_21_pad_groupi_g4923__8428(csa_tree_add_83_21_pad_groupi_n_813 ,csa_tree_add_83_21_pad_groupi_n_525 ,csa_tree_add_83_21_pad_groupi_n_695);
  or csa_tree_add_83_21_pad_groupi_g4924__5526(csa_tree_add_83_21_pad_groupi_n_811 ,csa_tree_add_83_21_pad_groupi_n_476 ,csa_tree_add_83_21_pad_groupi_n_599);
  or csa_tree_add_83_21_pad_groupi_g4925__6783(csa_tree_add_83_21_pad_groupi_n_810 ,csa_tree_add_83_21_pad_groupi_n_470 ,csa_tree_add_83_21_pad_groupi_n_627);
  or csa_tree_add_83_21_pad_groupi_g4926__3680(csa_tree_add_83_21_pad_groupi_n_809 ,csa_tree_add_83_21_pad_groupi_n_528 ,csa_tree_add_83_21_pad_groupi_n_651);
  or csa_tree_add_83_21_pad_groupi_g4927__1617(csa_tree_add_83_21_pad_groupi_n_808 ,csa_tree_add_83_21_pad_groupi_n_541 ,csa_tree_add_83_21_pad_groupi_n_635);
  or csa_tree_add_83_21_pad_groupi_g4928__2802(csa_tree_add_83_21_pad_groupi_n_807 ,csa_tree_add_83_21_pad_groupi_n_512 ,csa_tree_add_83_21_pad_groupi_n_625);
  or csa_tree_add_83_21_pad_groupi_g4929__1705(csa_tree_add_83_21_pad_groupi_n_806 ,csa_tree_add_83_21_pad_groupi_n_523 ,csa_tree_add_83_21_pad_groupi_n_623);
  or csa_tree_add_83_21_pad_groupi_g4930__5122(csa_tree_add_83_21_pad_groupi_n_804 ,csa_tree_add_83_21_pad_groupi_n_461 ,csa_tree_add_83_21_pad_groupi_n_694);
  or csa_tree_add_83_21_pad_groupi_g4931__8246(csa_tree_add_83_21_pad_groupi_n_803 ,csa_tree_add_83_21_pad_groupi_n_529 ,csa_tree_add_83_21_pad_groupi_n_653);
  or csa_tree_add_83_21_pad_groupi_g4933__7098(csa_tree_add_83_21_pad_groupi_n_800 ,csa_tree_add_83_21_pad_groupi_n_477 ,csa_tree_add_83_21_pad_groupi_n_658);
  or csa_tree_add_83_21_pad_groupi_g4934__6131(csa_tree_add_83_21_pad_groupi_n_799 ,csa_tree_add_83_21_pad_groupi_n_467 ,csa_tree_add_83_21_pad_groupi_n_680);
  or csa_tree_add_83_21_pad_groupi_g4935__1881(csa_tree_add_83_21_pad_groupi_n_798 ,csa_tree_add_83_21_pad_groupi_n_468 ,csa_tree_add_83_21_pad_groupi_n_607);
  or csa_tree_add_83_21_pad_groupi_g4936__5115(csa_tree_add_83_21_pad_groupi_n_797 ,csa_tree_add_83_21_pad_groupi_n_394 ,csa_tree_add_83_21_pad_groupi_n_663);
  or csa_tree_add_83_21_pad_groupi_g4937__7482(csa_tree_add_83_21_pad_groupi_n_796 ,csa_tree_add_83_21_pad_groupi_n_555 ,csa_tree_add_83_21_pad_groupi_n_669);
  or csa_tree_add_83_21_pad_groupi_g4938__4733(csa_tree_add_83_21_pad_groupi_n_795 ,csa_tree_add_83_21_pad_groupi_n_547 ,csa_tree_add_83_21_pad_groupi_n_696);
  or csa_tree_add_83_21_pad_groupi_g4939__6161(csa_tree_add_83_21_pad_groupi_n_793 ,csa_tree_add_83_21_pad_groupi_n_540 ,csa_tree_add_83_21_pad_groupi_n_697);
  or csa_tree_add_83_21_pad_groupi_g4940__9315(csa_tree_add_83_21_pad_groupi_n_792 ,csa_tree_add_83_21_pad_groupi_n_456 ,csa_tree_add_83_21_pad_groupi_n_638);
  or csa_tree_add_83_21_pad_groupi_g4941__9945(csa_tree_add_83_21_pad_groupi_n_790 ,csa_tree_add_83_21_pad_groupi_n_524 ,csa_tree_add_83_21_pad_groupi_n_661);
  or csa_tree_add_83_21_pad_groupi_g4942__2883(csa_tree_add_83_21_pad_groupi_n_788 ,csa_tree_add_83_21_pad_groupi_n_537 ,csa_tree_add_83_21_pad_groupi_n_616);
  or csa_tree_add_83_21_pad_groupi_g4943__2346(csa_tree_add_83_21_pad_groupi_n_787 ,csa_tree_add_83_21_pad_groupi_n_469 ,csa_tree_add_83_21_pad_groupi_n_672);
  or csa_tree_add_83_21_pad_groupi_g4944__1666(csa_tree_add_83_21_pad_groupi_n_786 ,csa_tree_add_83_21_pad_groupi_n_473 ,csa_tree_add_83_21_pad_groupi_n_589);
  or csa_tree_add_83_21_pad_groupi_g4945__7410(csa_tree_add_83_21_pad_groupi_n_785 ,csa_tree_add_83_21_pad_groupi_n_484 ,csa_tree_add_83_21_pad_groupi_n_698);
  or csa_tree_add_83_21_pad_groupi_g4946__6417(csa_tree_add_83_21_pad_groupi_n_784 ,csa_tree_add_83_21_pad_groupi_n_488 ,csa_tree_add_83_21_pad_groupi_n_608);
  or csa_tree_add_83_21_pad_groupi_g4947__5477(csa_tree_add_83_21_pad_groupi_n_783 ,csa_tree_add_83_21_pad_groupi_n_546 ,csa_tree_add_83_21_pad_groupi_n_648);
  not csa_tree_add_83_21_pad_groupi_g4949(csa_tree_add_83_21_pad_groupi_n_779 ,csa_tree_add_83_21_pad_groupi_n_778);
  not csa_tree_add_83_21_pad_groupi_g4950(csa_tree_add_83_21_pad_groupi_n_762 ,csa_tree_add_83_21_pad_groupi_n_763);
  not csa_tree_add_83_21_pad_groupi_g4951(csa_tree_add_83_21_pad_groupi_n_759 ,csa_tree_add_83_21_pad_groupi_n_760);
  not csa_tree_add_83_21_pad_groupi_g4952(csa_tree_add_83_21_pad_groupi_n_754 ,csa_tree_add_83_21_pad_groupi_n_755);
  not csa_tree_add_83_21_pad_groupi_g4953(csa_tree_add_83_21_pad_groupi_n_752 ,csa_tree_add_83_21_pad_groupi_n_753);
  not csa_tree_add_83_21_pad_groupi_g4954(csa_tree_add_83_21_pad_groupi_n_749 ,csa_tree_add_83_21_pad_groupi_n_750);
  not csa_tree_add_83_21_pad_groupi_g4955(csa_tree_add_83_21_pad_groupi_n_745 ,csa_tree_add_83_21_pad_groupi_n_746);
  not csa_tree_add_83_21_pad_groupi_g4956(csa_tree_add_83_21_pad_groupi_n_744 ,csa_tree_add_83_21_pad_groupi_n_743);
  not csa_tree_add_83_21_pad_groupi_g4957(csa_tree_add_83_21_pad_groupi_n_741 ,csa_tree_add_83_21_pad_groupi_n_742);
  not csa_tree_add_83_21_pad_groupi_g4958(csa_tree_add_83_21_pad_groupi_n_738 ,csa_tree_add_83_21_pad_groupi_n_739);
  not csa_tree_add_83_21_pad_groupi_g4959(csa_tree_add_83_21_pad_groupi_n_736 ,csa_tree_add_83_21_pad_groupi_n_737);
  not csa_tree_add_83_21_pad_groupi_g4960(csa_tree_add_83_21_pad_groupi_n_734 ,csa_tree_add_83_21_pad_groupi_n_735);
  not csa_tree_add_83_21_pad_groupi_g4961(csa_tree_add_83_21_pad_groupi_n_732 ,csa_tree_add_83_21_pad_groupi_n_733);
  not csa_tree_add_83_21_pad_groupi_g4962(csa_tree_add_83_21_pad_groupi_n_730 ,csa_tree_add_83_21_pad_groupi_n_731);
  not csa_tree_add_83_21_pad_groupi_g4963(csa_tree_add_83_21_pad_groupi_n_727 ,csa_tree_add_83_21_pad_groupi_n_728);
  not csa_tree_add_83_21_pad_groupi_g4964(csa_tree_add_83_21_pad_groupi_n_724 ,csa_tree_add_83_21_pad_groupi_n_725);
  not csa_tree_add_83_21_pad_groupi_g4965(csa_tree_add_83_21_pad_groupi_n_722 ,csa_tree_add_83_21_pad_groupi_n_723);
  not csa_tree_add_83_21_pad_groupi_g4966(csa_tree_add_83_21_pad_groupi_n_715 ,csa_tree_add_83_21_pad_groupi_n_716);
  not csa_tree_add_83_21_pad_groupi_g4967(csa_tree_add_83_21_pad_groupi_n_712 ,csa_tree_add_83_21_pad_groupi_n_713);
  xnor csa_tree_add_83_21_pad_groupi_g4968__2398(csa_tree_add_83_21_pad_groupi_n_711 ,csa_tree_add_83_21_pad_groupi_n_583 ,in8[10]);
  xnor csa_tree_add_83_21_pad_groupi_g4970__5107(csa_tree_add_83_21_pad_groupi_n_710 ,csa_tree_add_83_21_pad_groupi_n_282 ,in8[12]);
  xnor csa_tree_add_83_21_pad_groupi_g4972__6260(csa_tree_add_83_21_pad_groupi_n_709 ,csa_tree_add_83_21_pad_groupi_n_582 ,in8[12]);
  or csa_tree_add_83_21_pad_groupi_g4975__4319(csa_tree_add_83_21_pad_groupi_n_778 ,csa_tree_add_83_21_pad_groupi_n_539 ,csa_tree_add_83_21_pad_groupi_n_626);
  or csa_tree_add_83_21_pad_groupi_g4976__8428(csa_tree_add_83_21_pad_groupi_n_777 ,csa_tree_add_83_21_pad_groupi_n_550 ,csa_tree_add_83_21_pad_groupi_n_624);
  and csa_tree_add_83_21_pad_groupi_g4977__5526(csa_tree_add_83_21_pad_groupi_n_776 ,csa_tree_add_83_21_pad_groupi_n_464 ,csa_tree_add_83_21_pad_groupi_n_655);
  or csa_tree_add_83_21_pad_groupi_g4978__6783(csa_tree_add_83_21_pad_groupi_n_775 ,csa_tree_add_83_21_pad_groupi_n_482 ,csa_tree_add_83_21_pad_groupi_n_637);
  or csa_tree_add_83_21_pad_groupi_g4980__3680(csa_tree_add_83_21_pad_groupi_n_773 ,csa_tree_add_83_21_pad_groupi_n_519 ,csa_tree_add_83_21_pad_groupi_n_605);
  and csa_tree_add_83_21_pad_groupi_g4981__1617(csa_tree_add_83_21_pad_groupi_n_772 ,csa_tree_add_83_21_pad_groupi_n_457 ,csa_tree_add_83_21_pad_groupi_n_594);
  and csa_tree_add_83_21_pad_groupi_g4982__2802(csa_tree_add_83_21_pad_groupi_n_771 ,csa_tree_add_83_21_pad_groupi_n_492 ,csa_tree_add_83_21_pad_groupi_n_606);
  or csa_tree_add_83_21_pad_groupi_g4984__1705(csa_tree_add_83_21_pad_groupi_n_769 ,csa_tree_add_83_21_pad_groupi_n_490 ,csa_tree_add_83_21_pad_groupi_n_689);
  or csa_tree_add_83_21_pad_groupi_g4985__5122(csa_tree_add_83_21_pad_groupi_n_768 ,csa_tree_add_83_21_pad_groupi_n_545 ,csa_tree_add_83_21_pad_groupi_n_640);
  or csa_tree_add_83_21_pad_groupi_g4986__8246(csa_tree_add_83_21_pad_groupi_n_767 ,csa_tree_add_83_21_pad_groupi_n_552 ,csa_tree_add_83_21_pad_groupi_n_659);
  or csa_tree_add_83_21_pad_groupi_g4988__7098(csa_tree_add_83_21_pad_groupi_n_765 ,csa_tree_add_83_21_pad_groupi_n_517 ,csa_tree_add_83_21_pad_groupi_n_688);
  or csa_tree_add_83_21_pad_groupi_g4989__6131(csa_tree_add_83_21_pad_groupi_n_764 ,csa_tree_add_83_21_pad_groupi_n_554 ,csa_tree_add_83_21_pad_groupi_n_654);
  or csa_tree_add_83_21_pad_groupi_g4990__1881(csa_tree_add_83_21_pad_groupi_n_763 ,csa_tree_add_83_21_pad_groupi_n_480 ,csa_tree_add_83_21_pad_groupi_n_602);
  or csa_tree_add_83_21_pad_groupi_g4991__5115(csa_tree_add_83_21_pad_groupi_n_761 ,csa_tree_add_83_21_pad_groupi_n_577 ,csa_tree_add_83_21_pad_groupi_n_693);
  or csa_tree_add_83_21_pad_groupi_g4992__7482(csa_tree_add_83_21_pad_groupi_n_760 ,csa_tree_add_83_21_pad_groupi_n_478 ,csa_tree_add_83_21_pad_groupi_n_591);
  or csa_tree_add_83_21_pad_groupi_g4993__4733(csa_tree_add_83_21_pad_groupi_n_758 ,csa_tree_add_83_21_pad_groupi_n_514 ,csa_tree_add_83_21_pad_groupi_n_604);
  or csa_tree_add_83_21_pad_groupi_g4994__6161(csa_tree_add_83_21_pad_groupi_n_757 ,csa_tree_add_83_21_pad_groupi_n_532 ,csa_tree_add_83_21_pad_groupi_n_617);
  or csa_tree_add_83_21_pad_groupi_g4995__9315(csa_tree_add_83_21_pad_groupi_n_756 ,csa_tree_add_83_21_pad_groupi_n_455 ,csa_tree_add_83_21_pad_groupi_n_670);
  or csa_tree_add_83_21_pad_groupi_g4996__9945(csa_tree_add_83_21_pad_groupi_n_755 ,csa_tree_add_83_21_pad_groupi_n_544 ,csa_tree_add_83_21_pad_groupi_n_660);
  or csa_tree_add_83_21_pad_groupi_g4997__2883(csa_tree_add_83_21_pad_groupi_n_753 ,csa_tree_add_83_21_pad_groupi_n_486 ,csa_tree_add_83_21_pad_groupi_n_679);
  or csa_tree_add_83_21_pad_groupi_g4998__2346(csa_tree_add_83_21_pad_groupi_n_751 ,csa_tree_add_83_21_pad_groupi_n_575 ,csa_tree_add_83_21_pad_groupi_n_619);
  or csa_tree_add_83_21_pad_groupi_g4999__1666(csa_tree_add_83_21_pad_groupi_n_750 ,csa_tree_add_83_21_pad_groupi_n_522 ,csa_tree_add_83_21_pad_groupi_n_671);
  or csa_tree_add_83_21_pad_groupi_g5000__7410(csa_tree_add_83_21_pad_groupi_n_748 ,csa_tree_add_83_21_pad_groupi_n_515 ,csa_tree_add_83_21_pad_groupi_n_631);
  or csa_tree_add_83_21_pad_groupi_g5001__6417(csa_tree_add_83_21_pad_groupi_n_747 ,csa_tree_add_83_21_pad_groupi_n_573 ,csa_tree_add_83_21_pad_groupi_n_620);
  or csa_tree_add_83_21_pad_groupi_g5002__5477(csa_tree_add_83_21_pad_groupi_n_746 ,csa_tree_add_83_21_pad_groupi_n_534 ,csa_tree_add_83_21_pad_groupi_n_643);
  or csa_tree_add_83_21_pad_groupi_g5003__2398(csa_tree_add_83_21_pad_groupi_n_743 ,csa_tree_add_83_21_pad_groupi_n_481 ,csa_tree_add_83_21_pad_groupi_n_629);
  or csa_tree_add_83_21_pad_groupi_g5004__5107(csa_tree_add_83_21_pad_groupi_n_742 ,csa_tree_add_83_21_pad_groupi_n_536 ,csa_tree_add_83_21_pad_groupi_n_650);
  or csa_tree_add_83_21_pad_groupi_g5006__6260(csa_tree_add_83_21_pad_groupi_n_739 ,csa_tree_add_83_21_pad_groupi_n_564 ,csa_tree_add_83_21_pad_groupi_n_628);
  or csa_tree_add_83_21_pad_groupi_g5007__4319(csa_tree_add_83_21_pad_groupi_n_737 ,csa_tree_add_83_21_pad_groupi_n_513 ,csa_tree_add_83_21_pad_groupi_n_603);
  or csa_tree_add_83_21_pad_groupi_g5008__8428(csa_tree_add_83_21_pad_groupi_n_735 ,csa_tree_add_83_21_pad_groupi_n_553 ,csa_tree_add_83_21_pad_groupi_n_691);
  or csa_tree_add_83_21_pad_groupi_g5009__5526(csa_tree_add_83_21_pad_groupi_n_733 ,csa_tree_add_83_21_pad_groupi_n_530 ,csa_tree_add_83_21_pad_groupi_n_622);
  or csa_tree_add_83_21_pad_groupi_g5010__6783(csa_tree_add_83_21_pad_groupi_n_731 ,csa_tree_add_83_21_pad_groupi_n_463 ,csa_tree_add_83_21_pad_groupi_n_590);
  or csa_tree_add_83_21_pad_groupi_g5011__3680(csa_tree_add_83_21_pad_groupi_n_729 ,csa_tree_add_83_21_pad_groupi_n_471 ,csa_tree_add_83_21_pad_groupi_n_610);
  or csa_tree_add_83_21_pad_groupi_g5012__1617(csa_tree_add_83_21_pad_groupi_n_728 ,csa_tree_add_83_21_pad_groupi_n_520 ,csa_tree_add_83_21_pad_groupi_n_639);
  or csa_tree_add_83_21_pad_groupi_g5013__2802(csa_tree_add_83_21_pad_groupi_n_726 ,csa_tree_add_83_21_pad_groupi_n_535 ,csa_tree_add_83_21_pad_groupi_n_690);
  or csa_tree_add_83_21_pad_groupi_g5014__1705(csa_tree_add_83_21_pad_groupi_n_725 ,csa_tree_add_83_21_pad_groupi_n_538 ,csa_tree_add_83_21_pad_groupi_n_675);
  or csa_tree_add_83_21_pad_groupi_g5015__5122(csa_tree_add_83_21_pad_groupi_n_723 ,csa_tree_add_83_21_pad_groupi_n_543 ,csa_tree_add_83_21_pad_groupi_n_676);
  or csa_tree_add_83_21_pad_groupi_g5016__8246(csa_tree_add_83_21_pad_groupi_n_721 ,csa_tree_add_83_21_pad_groupi_n_542 ,csa_tree_add_83_21_pad_groupi_n_634);
  or csa_tree_add_83_21_pad_groupi_g5017__7098(csa_tree_add_83_21_pad_groupi_n_720 ,csa_tree_add_83_21_pad_groupi_n_479 ,csa_tree_add_83_21_pad_groupi_n_644);
  or csa_tree_add_83_21_pad_groupi_g5018__6131(csa_tree_add_83_21_pad_groupi_n_719 ,csa_tree_add_83_21_pad_groupi_n_521 ,csa_tree_add_83_21_pad_groupi_n_611);
  or csa_tree_add_83_21_pad_groupi_g5019__1881(csa_tree_add_83_21_pad_groupi_n_718 ,csa_tree_add_83_21_pad_groupi_n_489 ,csa_tree_add_83_21_pad_groupi_n_609);
  or csa_tree_add_83_21_pad_groupi_g5020__5115(csa_tree_add_83_21_pad_groupi_n_717 ,csa_tree_add_83_21_pad_groupi_n_549 ,csa_tree_add_83_21_pad_groupi_n_692);
  or csa_tree_add_83_21_pad_groupi_g5021__7482(csa_tree_add_83_21_pad_groupi_n_716 ,csa_tree_add_83_21_pad_groupi_n_465 ,csa_tree_add_83_21_pad_groupi_n_613);
  or csa_tree_add_83_21_pad_groupi_g5022__4733(csa_tree_add_83_21_pad_groupi_n_714 ,csa_tree_add_83_21_pad_groupi_n_474 ,csa_tree_add_83_21_pad_groupi_n_657);
  or csa_tree_add_83_21_pad_groupi_g5023__6161(csa_tree_add_83_21_pad_groupi_n_713 ,csa_tree_add_83_21_pad_groupi_n_458 ,csa_tree_add_83_21_pad_groupi_n_667);
  not csa_tree_add_83_21_pad_groupi_g5024(csa_tree_add_83_21_pad_groupi_n_707 ,csa_tree_add_83_21_pad_groupi_n_706);
  not csa_tree_add_83_21_pad_groupi_g5025(csa_tree_add_83_21_pad_groupi_n_705 ,csa_tree_add_83_21_pad_groupi_n_704);
  nor csa_tree_add_83_21_pad_groupi_g5026__9315(csa_tree_add_83_21_pad_groupi_n_703 ,csa_tree_add_83_21_pad_groupi_n_113 ,csa_tree_add_83_21_pad_groupi_n_218);
  nor csa_tree_add_83_21_pad_groupi_g5027__9945(csa_tree_add_83_21_pad_groupi_n_702 ,in8[9] ,csa_tree_add_83_21_pad_groupi_n_358);
  nor csa_tree_add_83_21_pad_groupi_g5029__2883(csa_tree_add_83_21_pad_groupi_n_700 ,in8[12] ,csa_tree_add_83_21_pad_groupi_n_579);
  nor csa_tree_add_83_21_pad_groupi_g5030__2346(csa_tree_add_83_21_pad_groupi_n_699 ,csa_tree_add_83_21_pad_groupi_n_115 ,csa_tree_add_83_21_pad_groupi_n_189);
  and csa_tree_add_83_21_pad_groupi_g5031__1666(csa_tree_add_83_21_pad_groupi_n_698 ,in9[5] ,csa_tree_add_83_21_pad_groupi_n_172);
  nor csa_tree_add_83_21_pad_groupi_g5032__7410(csa_tree_add_83_21_pad_groupi_n_697 ,csa_tree_add_83_21_pad_groupi_n_119 ,csa_tree_add_83_21_pad_groupi_n_38);
  nor csa_tree_add_83_21_pad_groupi_g5033__6417(csa_tree_add_83_21_pad_groupi_n_696 ,csa_tree_add_83_21_pad_groupi_n_93 ,csa_tree_add_83_21_pad_groupi_n_66);
  and csa_tree_add_83_21_pad_groupi_g5034__5477(csa_tree_add_83_21_pad_groupi_n_695 ,in9[2] ,csa_tree_add_83_21_pad_groupi_n_133);
  and csa_tree_add_83_21_pad_groupi_g5035__2398(csa_tree_add_83_21_pad_groupi_n_694 ,in9[10] ,csa_tree_add_83_21_pad_groupi_n_433);
  and csa_tree_add_83_21_pad_groupi_g5036__5107(csa_tree_add_83_21_pad_groupi_n_693 ,in9[8] ,csa_tree_add_83_21_pad_groupi_n_287);
  and csa_tree_add_83_21_pad_groupi_g5037__6260(csa_tree_add_83_21_pad_groupi_n_692 ,in9[14] ,csa_tree_add_83_21_pad_groupi_n_169);
  and csa_tree_add_83_21_pad_groupi_g5038__4319(csa_tree_add_83_21_pad_groupi_n_691 ,in9[1] ,csa_tree_add_83_21_pad_groupi_n_168);
  and csa_tree_add_83_21_pad_groupi_g5039__8428(csa_tree_add_83_21_pad_groupi_n_690 ,in9[5] ,csa_tree_add_83_21_pad_groupi_n_142);
  and csa_tree_add_83_21_pad_groupi_g5040__5526(csa_tree_add_83_21_pad_groupi_n_689 ,in9[7] ,csa_tree_add_83_21_pad_groupi_n_126);
  and csa_tree_add_83_21_pad_groupi_g5041__6783(csa_tree_add_83_21_pad_groupi_n_688 ,in9[11] ,csa_tree_add_83_21_pad_groupi_n_285);
  or csa_tree_add_83_21_pad_groupi_g5044__3680(csa_tree_add_83_21_pad_groupi_n_685 ,csa_tree_add_83_21_pad_groupi_n_17 ,csa_tree_add_83_21_pad_groupi_n_118);
  or csa_tree_add_83_21_pad_groupi_g5046__1617(csa_tree_add_83_21_pad_groupi_n_683 ,csa_tree_add_83_21_pad_groupi_n_149 ,csa_tree_add_83_21_pad_groupi_n_583);
  and csa_tree_add_83_21_pad_groupi_g5047__2802(csa_tree_add_83_21_pad_groupi_n_682 ,in8[12] ,csa_tree_add_83_21_pad_groupi_n_579);
  and csa_tree_add_83_21_pad_groupi_g5048__1705(csa_tree_add_83_21_pad_groupi_n_681 ,in9[11] ,csa_tree_add_83_21_pad_groupi_n_135);
  and csa_tree_add_83_21_pad_groupi_g5049__5122(csa_tree_add_83_21_pad_groupi_n_680 ,in9[6] ,csa_tree_add_83_21_pad_groupi_n_445);
  nor csa_tree_add_83_21_pad_groupi_g5050__8246(csa_tree_add_83_21_pad_groupi_n_679 ,csa_tree_add_83_21_pad_groupi_n_252 ,csa_tree_add_83_21_pad_groupi_n_223);
  and csa_tree_add_83_21_pad_groupi_g5052__7098(csa_tree_add_83_21_pad_groupi_n_677 ,in9[3] ,csa_tree_add_83_21_pad_groupi_n_139);
  and csa_tree_add_83_21_pad_groupi_g5053__6131(csa_tree_add_83_21_pad_groupi_n_676 ,in9[6] ,csa_tree_add_83_21_pad_groupi_n_136);
  and csa_tree_add_83_21_pad_groupi_g5054__1881(csa_tree_add_83_21_pad_groupi_n_675 ,in9[4] ,csa_tree_add_83_21_pad_groupi_n_144);
  and csa_tree_add_83_21_pad_groupi_g5055__5115(csa_tree_add_83_21_pad_groupi_n_674 ,in9[4] ,csa_tree_add_83_21_pad_groupi_n_138);
  nor csa_tree_add_83_21_pad_groupi_g5056__7482(csa_tree_add_83_21_pad_groupi_n_673 ,csa_tree_add_83_21_pad_groupi_n_369 ,csa_tree_add_83_21_pad_groupi_n_581);
  and csa_tree_add_83_21_pad_groupi_g5057__4733(csa_tree_add_83_21_pad_groupi_n_672 ,in9[12] ,csa_tree_add_83_21_pad_groupi_n_428);
  and csa_tree_add_83_21_pad_groupi_g5058__6161(csa_tree_add_83_21_pad_groupi_n_671 ,in9[4] ,csa_tree_add_83_21_pad_groupi_n_124);
  and csa_tree_add_83_21_pad_groupi_g5059__9315(csa_tree_add_83_21_pad_groupi_n_670 ,in9[9] ,csa_tree_add_83_21_pad_groupi_n_439);
  and csa_tree_add_83_21_pad_groupi_g5060__9945(csa_tree_add_83_21_pad_groupi_n_669 ,in9[14] ,csa_tree_add_83_21_pad_groupi_n_288);
  and csa_tree_add_83_21_pad_groupi_g5062__2883(csa_tree_add_83_21_pad_groupi_n_667 ,in9[14] ,csa_tree_add_83_21_pad_groupi_n_425);
  and csa_tree_add_83_21_pad_groupi_g5063__2346(csa_tree_add_83_21_pad_groupi_n_666 ,in8[12] ,csa_tree_add_83_21_pad_groupi_n_280);
  and csa_tree_add_83_21_pad_groupi_g5064__1666(csa_tree_add_83_21_pad_groupi_n_665 ,in9[7] ,csa_tree_add_83_21_pad_groupi_n_171);
  and csa_tree_add_83_21_pad_groupi_g5066__7410(csa_tree_add_83_21_pad_groupi_n_663 ,csa_tree_add_83_21_pad_groupi_n_406 ,csa_tree_add_83_21_pad_groupi_n_583);
  and csa_tree_add_83_21_pad_groupi_g5067__6417(csa_tree_add_83_21_pad_groupi_n_662 ,in9[7] ,csa_tree_add_83_21_pad_groupi_n_429);
  and csa_tree_add_83_21_pad_groupi_g5068__5477(csa_tree_add_83_21_pad_groupi_n_661 ,in9[9] ,csa_tree_add_83_21_pad_groupi_n_145);
  and csa_tree_add_83_21_pad_groupi_g5069__2398(csa_tree_add_83_21_pad_groupi_n_660 ,in9[14] ,csa_tree_add_83_21_pad_groupi_n_127);
  nor csa_tree_add_83_21_pad_groupi_g5070__5107(csa_tree_add_83_21_pad_groupi_n_659 ,csa_tree_add_83_21_pad_groupi_n_112 ,csa_tree_add_83_21_pad_groupi_n_202);
  and csa_tree_add_83_21_pad_groupi_g5071__6260(csa_tree_add_83_21_pad_groupi_n_658 ,in9[3] ,csa_tree_add_83_21_pad_groupi_n_133);
  nor csa_tree_add_83_21_pad_groupi_g5072__4319(csa_tree_add_83_21_pad_groupi_n_657 ,csa_tree_add_83_21_pad_groupi_n_118 ,csa_tree_add_83_21_pad_groupi_n_215);
  or csa_tree_add_83_21_pad_groupi_g5073__8428(csa_tree_add_83_21_pad_groupi_n_656 ,csa_tree_add_83_21_pad_groupi_n_373 ,csa_tree_add_83_21_pad_groupi_n_357);
  or csa_tree_add_83_21_pad_groupi_g5074__5526(csa_tree_add_83_21_pad_groupi_n_655 ,csa_tree_add_83_21_pad_groupi_n_27 ,csa_tree_add_83_21_pad_groupi_n_427);
  and csa_tree_add_83_21_pad_groupi_g5075__6783(csa_tree_add_83_21_pad_groupi_n_654 ,in9[11] ,csa_tree_add_83_21_pad_groupi_n_130);
  and csa_tree_add_83_21_pad_groupi_g5076__3680(csa_tree_add_83_21_pad_groupi_n_653 ,in9[1] ,csa_tree_add_83_21_pad_groupi_n_147);
  nor csa_tree_add_83_21_pad_groupi_g5077__1617(csa_tree_add_83_21_pad_groupi_n_652 ,csa_tree_add_83_21_pad_groupi_n_93 ,csa_tree_add_83_21_pad_groupi_n_74);
  and csa_tree_add_83_21_pad_groupi_g5078__2802(csa_tree_add_83_21_pad_groupi_n_651 ,in9[13] ,csa_tree_add_83_21_pad_groupi_n_148);
  and csa_tree_add_83_21_pad_groupi_g5079__1705(csa_tree_add_83_21_pad_groupi_n_650 ,in9[6] ,csa_tree_add_83_21_pad_groupi_n_148);
  and csa_tree_add_83_21_pad_groupi_g5080__5122(csa_tree_add_83_21_pad_groupi_n_649 ,in9[12] ,csa_tree_add_83_21_pad_groupi_n_142);
  and csa_tree_add_83_21_pad_groupi_g5081__8246(csa_tree_add_83_21_pad_groupi_n_648 ,in9[3] ,csa_tree_add_83_21_pad_groupi_n_129);
  and csa_tree_add_83_21_pad_groupi_g5082__7098(csa_tree_add_83_21_pad_groupi_n_647 ,in9[4] ,csa_tree_add_83_21_pad_groupi_n_284);
  or csa_tree_add_83_21_pad_groupi_g5084__6131(csa_tree_add_83_21_pad_groupi_n_706 ,csa_tree_add_83_21_pad_groupi_n_24 ,csa_tree_add_83_21_pad_groupi_n_502);
  or csa_tree_add_83_21_pad_groupi_g5085__1881(csa_tree_add_83_21_pad_groupi_n_704 ,csa_tree_add_83_21_pad_groupi_n_24 ,csa_tree_add_83_21_pad_groupi_n_257);
  nor csa_tree_add_83_21_pad_groupi_g5086__5115(csa_tree_add_83_21_pad_groupi_n_644 ,csa_tree_add_83_21_pad_groupi_n_113 ,csa_tree_add_83_21_pad_groupi_n_178);
  nor csa_tree_add_83_21_pad_groupi_g5087__7482(csa_tree_add_83_21_pad_groupi_n_643 ,csa_tree_add_83_21_pad_groupi_n_160 ,csa_tree_add_83_21_pad_groupi_n_578);
  or csa_tree_add_83_21_pad_groupi_g5088__4733(csa_tree_add_83_21_pad_groupi_n_642 ,csa_tree_add_83_21_pad_groupi_n_47 ,csa_tree_add_83_21_pad_groupi_n_497);
  and csa_tree_add_83_21_pad_groupi_g5090__6161(csa_tree_add_83_21_pad_groupi_n_640 ,in9[6] ,csa_tree_add_83_21_pad_groupi_n_130);
  and csa_tree_add_83_21_pad_groupi_g5091__9315(csa_tree_add_83_21_pad_groupi_n_639 ,in9[13] ,csa_tree_add_83_21_pad_groupi_n_171);
  nor csa_tree_add_83_21_pad_groupi_g5092__9945(csa_tree_add_83_21_pad_groupi_n_638 ,csa_tree_add_83_21_pad_groupi_n_87 ,csa_tree_add_83_21_pad_groupi_n_434);
  and csa_tree_add_83_21_pad_groupi_g5093__2883(csa_tree_add_83_21_pad_groupi_n_637 ,in9[10] ,csa_tree_add_83_21_pad_groupi_n_166);
  nor csa_tree_add_83_21_pad_groupi_g5095__2346(csa_tree_add_83_21_pad_groupi_n_635 ,csa_tree_add_83_21_pad_groupi_n_96 ,csa_tree_add_83_21_pad_groupi_n_255);
  and csa_tree_add_83_21_pad_groupi_g5096__1666(csa_tree_add_83_21_pad_groupi_n_634 ,in9[2] ,csa_tree_add_83_21_pad_groupi_n_168);
  and csa_tree_add_83_21_pad_groupi_g5097__7410(csa_tree_add_83_21_pad_groupi_n_633 ,in9[13] ,csa_tree_add_83_21_pad_groupi_n_124);
  nor csa_tree_add_83_21_pad_groupi_g5099__6417(csa_tree_add_83_21_pad_groupi_n_631 ,csa_tree_add_83_21_pad_groupi_n_231 ,csa_tree_add_83_21_pad_groupi_n_257);
  and csa_tree_add_83_21_pad_groupi_g5101__5477(csa_tree_add_83_21_pad_groupi_n_629 ,in9[13] ,csa_tree_add_83_21_pad_groupi_n_287);
  and csa_tree_add_83_21_pad_groupi_g5102__2398(csa_tree_add_83_21_pad_groupi_n_628 ,in9[11] ,csa_tree_add_83_21_pad_groupi_n_145);
  and csa_tree_add_83_21_pad_groupi_g5103__5107(csa_tree_add_83_21_pad_groupi_n_627 ,in9[7] ,csa_tree_add_83_21_pad_groupi_n_141);
  nor csa_tree_add_83_21_pad_groupi_g5104__6260(csa_tree_add_83_21_pad_groupi_n_626 ,csa_tree_add_83_21_pad_groupi_n_71 ,csa_tree_add_83_21_pad_groupi_n_507);
  and csa_tree_add_83_21_pad_groupi_g5105__4319(csa_tree_add_83_21_pad_groupi_n_625 ,in9[7] ,csa_tree_add_83_21_pad_groupi_n_285);
  and csa_tree_add_83_21_pad_groupi_g5106__8428(csa_tree_add_83_21_pad_groupi_n_624 ,in9[5] ,csa_tree_add_83_21_pad_groupi_n_165);
  and csa_tree_add_83_21_pad_groupi_g5107__5526(csa_tree_add_83_21_pad_groupi_n_623 ,in9[10] ,csa_tree_add_83_21_pad_groupi_n_132);
  nor csa_tree_add_83_21_pad_groupi_g5108__6783(csa_tree_add_83_21_pad_groupi_n_622 ,csa_tree_add_83_21_pad_groupi_n_159 ,csa_tree_add_83_21_pad_groupi_n_282);
  nor csa_tree_add_83_21_pad_groupi_g5109__3680(csa_tree_add_83_21_pad_groupi_n_621 ,csa_tree_add_83_21_pad_groupi_n_98 ,csa_tree_add_83_21_pad_groupi_n_430);
  nor csa_tree_add_83_21_pad_groupi_g5110__1617(csa_tree_add_83_21_pad_groupi_n_620 ,csa_tree_add_83_21_pad_groupi_n_194 ,csa_tree_add_83_21_pad_groupi_n_502);
  nor csa_tree_add_83_21_pad_groupi_g5111__2802(csa_tree_add_83_21_pad_groupi_n_619 ,csa_tree_add_83_21_pad_groupi_n_116 ,csa_tree_add_83_21_pad_groupi_n_187);
  and csa_tree_add_83_21_pad_groupi_g5112__1705(csa_tree_add_83_21_pad_groupi_n_618 ,in9[8] ,csa_tree_add_83_21_pad_groupi_n_165);
  and csa_tree_add_83_21_pad_groupi_g5113__5122(csa_tree_add_83_21_pad_groupi_n_617 ,in9[8] ,csa_tree_add_83_21_pad_groupi_n_136);
  nor csa_tree_add_83_21_pad_groupi_g5114__8246(csa_tree_add_83_21_pad_groupi_n_616 ,csa_tree_add_83_21_pad_groupi_n_119 ,csa_tree_add_83_21_pad_groupi_n_181);
  nor csa_tree_add_83_21_pad_groupi_g5117__7098(csa_tree_add_83_21_pad_groupi_n_613 ,csa_tree_add_83_21_pad_groupi_n_204 ,csa_tree_add_83_21_pad_groupi_n_432);
  or csa_tree_add_83_21_pad_groupi_g5118__6131(csa_tree_add_83_21_pad_groupi_n_612 ,csa_tree_add_83_21_pad_groupi_n_64 ,csa_tree_add_83_21_pad_groupi_n_438);
  and csa_tree_add_83_21_pad_groupi_g5119__1881(csa_tree_add_83_21_pad_groupi_n_611 ,in9[8] ,csa_tree_add_83_21_pad_groupi_n_284);
  nor csa_tree_add_83_21_pad_groupi_g5120__5115(csa_tree_add_83_21_pad_groupi_n_610 ,csa_tree_add_83_21_pad_groupi_n_116 ,csa_tree_add_83_21_pad_groupi_n_184);
  nor csa_tree_add_83_21_pad_groupi_g5121__7482(csa_tree_add_83_21_pad_groupi_n_609 ,csa_tree_add_83_21_pad_groupi_n_91 ,csa_tree_add_83_21_pad_groupi_n_501);
  and csa_tree_add_83_21_pad_groupi_g5122__4733(csa_tree_add_83_21_pad_groupi_n_608 ,in9[12] ,csa_tree_add_83_21_pad_groupi_n_166);
  and csa_tree_add_83_21_pad_groupi_g5123__6161(csa_tree_add_83_21_pad_groupi_n_607 ,in9[11] ,csa_tree_add_83_21_pad_groupi_n_431);
  or csa_tree_add_83_21_pad_groupi_g5124__9315(csa_tree_add_83_21_pad_groupi_n_606 ,csa_tree_add_83_21_pad_groupi_n_17 ,csa_tree_add_83_21_pad_groupi_n_255);
  and csa_tree_add_83_21_pad_groupi_g5125__9945(csa_tree_add_83_21_pad_groupi_n_605 ,in9[9] ,csa_tree_add_83_21_pad_groupi_n_127);
  nor csa_tree_add_83_21_pad_groupi_g5126__2883(csa_tree_add_83_21_pad_groupi_n_604 ,csa_tree_add_83_21_pad_groupi_n_211 ,csa_tree_add_83_21_pad_groupi_n_508);
  and csa_tree_add_83_21_pad_groupi_g5127__2346(csa_tree_add_83_21_pad_groupi_n_603 ,in9[12] ,csa_tree_add_83_21_pad_groupi_n_169);
  and csa_tree_add_83_21_pad_groupi_g5128__1666(csa_tree_add_83_21_pad_groupi_n_602 ,in9[1] ,csa_tree_add_83_21_pad_groupi_n_123);
  nor csa_tree_add_83_21_pad_groupi_g5130__7410(csa_tree_add_83_21_pad_groupi_n_600 ,in8[12] ,csa_tree_add_83_21_pad_groupi_n_582);
  and csa_tree_add_83_21_pad_groupi_g5131__6417(csa_tree_add_83_21_pad_groupi_n_599 ,in9[9] ,csa_tree_add_83_21_pad_groupi_n_139);
  nor csa_tree_add_83_21_pad_groupi_g5132__5477(csa_tree_add_83_21_pad_groupi_n_598 ,csa_tree_add_83_21_pad_groupi_n_101 ,csa_tree_add_83_21_pad_groupi_n_508);
  or csa_tree_add_83_21_pad_groupi_g5135__2398(csa_tree_add_83_21_pad_groupi_n_595 ,csa_tree_add_83_21_pad_groupi_n_55 ,csa_tree_add_83_21_pad_groupi_n_115);
  or csa_tree_add_83_21_pad_groupi_g5136__5107(csa_tree_add_83_21_pad_groupi_n_594 ,csa_tree_add_83_21_pad_groupi_n_50 ,csa_tree_add_83_21_pad_groupi_n_426);
  nor csa_tree_add_83_21_pad_groupi_g5137__6260(csa_tree_add_83_21_pad_groupi_n_593 ,in8[11] ,csa_tree_add_83_21_pad_groupi_n_580);
  and csa_tree_add_83_21_pad_groupi_g5139__4319(csa_tree_add_83_21_pad_groupi_n_591 ,in9[10] ,csa_tree_add_83_21_pad_groupi_n_288);
  and csa_tree_add_83_21_pad_groupi_g5140__8428(csa_tree_add_83_21_pad_groupi_n_590 ,in9[13] ,csa_tree_add_83_21_pad_groupi_n_435);
  and csa_tree_add_83_21_pad_groupi_g5141__5526(csa_tree_add_83_21_pad_groupi_n_589 ,in9[10] ,csa_tree_add_83_21_pad_groupi_n_172);
  nor csa_tree_add_83_21_pad_groupi_g5142__6783(csa_tree_add_83_21_pad_groupi_n_588 ,csa_tree_add_83_21_pad_groupi_n_158 ,csa_tree_add_83_21_pad_groupi_n_280);
  or csa_tree_add_83_21_pad_groupi_g5143__3680(csa_tree_add_83_21_pad_groupi_n_587 ,csa_tree_add_83_21_pad_groupi_n_151 ,csa_tree_add_83_21_pad_groupi_n_580);
  or csa_tree_add_83_21_pad_groupi_g5144__1617(csa_tree_add_83_21_pad_groupi_n_586 ,csa_tree_add_83_21_pad_groupi_n_15 ,csa_tree_add_83_21_pad_groupi_n_581);
  or csa_tree_add_83_21_pad_groupi_g5145__2802(csa_tree_add_83_21_pad_groupi_n_646 ,csa_tree_add_83_21_pad_groupi_n_57 ,csa_tree_add_83_21_pad_groupi_n_493);
  or csa_tree_add_83_21_pad_groupi_g5146__1705(csa_tree_add_83_21_pad_groupi_n_645 ,csa_tree_add_83_21_pad_groupi_n_42 ,csa_tree_add_83_21_pad_groupi_n_278);
  nor csa_tree_add_83_21_pad_groupi_g5150__5122(csa_tree_add_83_21_pad_groupi_n_577 ,csa_tree_add_83_21_pad_groupi_n_183 ,csa_tree_add_83_21_pad_groupi_n_332);
  nor csa_tree_add_83_21_pad_groupi_g5151__8246(csa_tree_add_83_21_pad_groupi_n_576 ,csa_tree_add_83_21_pad_groupi_n_42 ,csa_tree_add_83_21_pad_groupi_n_302);
  nor csa_tree_add_83_21_pad_groupi_g5152__7098(csa_tree_add_83_21_pad_groupi_n_575 ,csa_tree_add_83_21_pad_groupi_n_233 ,csa_tree_add_83_21_pad_groupi_n_306);
  nor csa_tree_add_83_21_pad_groupi_g5153__6131(csa_tree_add_83_21_pad_groupi_n_574 ,csa_tree_add_83_21_pad_groupi_n_193 ,csa_tree_add_83_21_pad_groupi_n_341);
  nor csa_tree_add_83_21_pad_groupi_g5154__1881(csa_tree_add_83_21_pad_groupi_n_573 ,csa_tree_add_83_21_pad_groupi_n_84 ,csa_tree_add_83_21_pad_groupi_n_312);
  nor csa_tree_add_83_21_pad_groupi_g5163__5115(csa_tree_add_83_21_pad_groupi_n_564 ,csa_tree_add_83_21_pad_groupi_n_78 ,csa_tree_add_83_21_pad_groupi_n_330);
  nor csa_tree_add_83_21_pad_groupi_g5170__7482(csa_tree_add_83_21_pad_groupi_n_557 ,csa_tree_add_83_21_pad_groupi_n_71 ,csa_tree_add_83_21_pad_groupi_n_335);
  nor csa_tree_add_83_21_pad_groupi_g5171__4733(csa_tree_add_83_21_pad_groupi_n_556 ,csa_tree_add_83_21_pad_groupi_n_101 ,csa_tree_add_83_21_pad_groupi_n_315);
  nor csa_tree_add_83_21_pad_groupi_g5172__6161(csa_tree_add_83_21_pad_groupi_n_555 ,csa_tree_add_83_21_pad_groupi_n_186 ,csa_tree_add_83_21_pad_groupi_n_336);
  nor csa_tree_add_83_21_pad_groupi_g5173__9315(csa_tree_add_83_21_pad_groupi_n_554 ,csa_tree_add_83_21_pad_groupi_n_177 ,csa_tree_add_83_21_pad_groupi_n_309);
  nor csa_tree_add_83_21_pad_groupi_g5174__9945(csa_tree_add_83_21_pad_groupi_n_553 ,csa_tree_add_83_21_pad_groupi_n_244 ,csa_tree_add_83_21_pad_groupi_n_320);
  nor csa_tree_add_83_21_pad_groupi_g5175__2883(csa_tree_add_83_21_pad_groupi_n_552 ,csa_tree_add_83_21_pad_groupi_n_247 ,csa_tree_add_83_21_pad_groupi_n_323);
  nor csa_tree_add_83_21_pad_groupi_g5176__2346(csa_tree_add_83_21_pad_groupi_n_551 ,csa_tree_add_83_21_pad_groupi_n_67 ,csa_tree_add_83_21_pad_groupi_n_317);
  nor csa_tree_add_83_21_pad_groupi_g5177__1666(csa_tree_add_83_21_pad_groupi_n_550 ,csa_tree_add_83_21_pad_groupi_n_175 ,csa_tree_add_83_21_pad_groupi_n_339);
  nor csa_tree_add_83_21_pad_groupi_g5178__7410(csa_tree_add_83_21_pad_groupi_n_549 ,csa_tree_add_83_21_pad_groupi_n_85 ,csa_tree_add_83_21_pad_groupi_n_321);
  nor csa_tree_add_83_21_pad_groupi_g5179__6417(csa_tree_add_83_21_pad_groupi_n_548 ,csa_tree_add_83_21_pad_groupi_n_88 ,csa_tree_add_83_21_pad_groupi_n_305);
  nor csa_tree_add_83_21_pad_groupi_g5180__5477(csa_tree_add_83_21_pad_groupi_n_547 ,csa_tree_add_83_21_pad_groupi_n_197 ,csa_tree_add_83_21_pad_groupi_n_323);
  nor csa_tree_add_83_21_pad_groupi_g5181__2398(csa_tree_add_83_21_pad_groupi_n_546 ,csa_tree_add_83_21_pad_groupi_n_100 ,csa_tree_add_83_21_pad_groupi_n_326);
  nor csa_tree_add_83_21_pad_groupi_g5182__5107(csa_tree_add_83_21_pad_groupi_n_545 ,csa_tree_add_83_21_pad_groupi_n_53 ,csa_tree_add_83_21_pad_groupi_n_327);
  nor csa_tree_add_83_21_pad_groupi_g5183__6260(csa_tree_add_83_21_pad_groupi_n_544 ,csa_tree_add_83_21_pad_groupi_n_187 ,csa_tree_add_83_21_pad_groupi_n_326);
  nor csa_tree_add_83_21_pad_groupi_g5184__4319(csa_tree_add_83_21_pad_groupi_n_543 ,csa_tree_add_83_21_pad_groupi_n_196 ,csa_tree_add_83_21_pad_groupi_n_317);
  nor csa_tree_add_83_21_pad_groupi_g5185__8428(csa_tree_add_83_21_pad_groupi_n_542 ,csa_tree_add_83_21_pad_groupi_n_217 ,csa_tree_add_83_21_pad_groupi_n_318);
  nor csa_tree_add_83_21_pad_groupi_g5186__5526(csa_tree_add_83_21_pad_groupi_n_541 ,csa_tree_add_83_21_pad_groupi_n_209 ,csa_tree_add_83_21_pad_groupi_n_344);
  nor csa_tree_add_83_21_pad_groupi_g5187__6783(csa_tree_add_83_21_pad_groupi_n_540 ,csa_tree_add_83_21_pad_groupi_n_229 ,csa_tree_add_83_21_pad_groupi_n_324);
  nor csa_tree_add_83_21_pad_groupi_g5188__3680(csa_tree_add_83_21_pad_groupi_n_539 ,csa_tree_add_83_21_pad_groupi_n_41 ,csa_tree_add_83_21_pad_groupi_n_335);
  nor csa_tree_add_83_21_pad_groupi_g5189__1617(csa_tree_add_83_21_pad_groupi_n_538 ,csa_tree_add_83_21_pad_groupi_n_36 ,csa_tree_add_83_21_pad_groupi_n_336);
  nor csa_tree_add_83_21_pad_groupi_g5190__2802(csa_tree_add_83_21_pad_groupi_n_537 ,csa_tree_add_83_21_pad_groupi_n_79 ,csa_tree_add_83_21_pad_groupi_n_324);
  nor csa_tree_add_83_21_pad_groupi_g5191__1705(csa_tree_add_83_21_pad_groupi_n_536 ,csa_tree_add_83_21_pad_groupi_n_204 ,csa_tree_add_83_21_pad_groupi_n_345);
  nor csa_tree_add_83_21_pad_groupi_g5192__5122(csa_tree_add_83_21_pad_groupi_n_535 ,csa_tree_add_83_21_pad_groupi_n_28 ,csa_tree_add_83_21_pad_groupi_n_329);
  nor csa_tree_add_83_21_pad_groupi_g5193__8246(csa_tree_add_83_21_pad_groupi_n_534 ,csa_tree_add_83_21_pad_groupi_n_194 ,csa_tree_add_83_21_pad_groupi_n_327);
  nor csa_tree_add_83_21_pad_groupi_g5194__7098(csa_tree_add_83_21_pad_groupi_n_533 ,csa_tree_add_83_21_pad_groupi_n_191 ,csa_tree_add_83_21_pad_groupi_n_338);
  nor csa_tree_add_83_21_pad_groupi_g5195__6131(csa_tree_add_83_21_pad_groupi_n_532 ,csa_tree_add_83_21_pad_groupi_n_184 ,csa_tree_add_83_21_pad_groupi_n_318);
  or csa_tree_add_83_21_pad_groupi_g5196__1881(csa_tree_add_83_21_pad_groupi_n_531 ,csa_tree_add_83_21_pad_groupi_n_174 ,csa_tree_add_83_21_pad_groupi_n_305);
  nor csa_tree_add_83_21_pad_groupi_g5197__5115(csa_tree_add_83_21_pad_groupi_n_530 ,csa_tree_add_83_21_pad_groupi_n_39 ,csa_tree_add_83_21_pad_groupi_n_330);
  nor csa_tree_add_83_21_pad_groupi_g5198__7482(csa_tree_add_83_21_pad_groupi_n_529 ,csa_tree_add_83_21_pad_groupi_n_243 ,csa_tree_add_83_21_pad_groupi_n_344);
  nor csa_tree_add_83_21_pad_groupi_g5199__4733(csa_tree_add_83_21_pad_groupi_n_528 ,csa_tree_add_83_21_pad_groupi_n_91 ,csa_tree_add_83_21_pad_groupi_n_345);
  nor csa_tree_add_83_21_pad_groupi_g5200__6161(csa_tree_add_83_21_pad_groupi_n_527 ,csa_tree_add_83_21_pad_groupi_n_231 ,csa_tree_add_83_21_pad_groupi_n_321);
  nor csa_tree_add_83_21_pad_groupi_g5201__9315(csa_tree_add_83_21_pad_groupi_n_526 ,csa_tree_add_83_21_pad_groupi_n_217 ,csa_tree_add_83_21_pad_groupi_n_265);
  nor csa_tree_add_83_21_pad_groupi_g5202__9945(csa_tree_add_83_21_pad_groupi_n_525 ,csa_tree_add_83_21_pad_groupi_n_64 ,csa_tree_add_83_21_pad_groupi_n_311);
  nor csa_tree_add_83_21_pad_groupi_g5203__2883(csa_tree_add_83_21_pad_groupi_n_524 ,csa_tree_add_83_21_pad_groupi_n_55 ,csa_tree_add_83_21_pad_groupi_n_269);
  nor csa_tree_add_83_21_pad_groupi_g5204__2346(csa_tree_add_83_21_pad_groupi_n_523 ,csa_tree_add_83_21_pad_groupi_n_76 ,csa_tree_add_83_21_pad_groupi_n_312);
  nor csa_tree_add_83_21_pad_groupi_g5205__1666(csa_tree_add_83_21_pad_groupi_n_522 ,csa_tree_add_83_21_pad_groupi_n_201 ,csa_tree_add_83_21_pad_groupi_n_339);
  nor csa_tree_add_83_21_pad_groupi_g5206__7410(csa_tree_add_83_21_pad_groupi_n_521 ,csa_tree_add_83_21_pad_groupi_n_22 ,csa_tree_add_83_21_pad_groupi_n_275);
  nor csa_tree_add_83_21_pad_groupi_g5207__6417(csa_tree_add_83_21_pad_groupi_n_520 ,csa_tree_add_83_21_pad_groupi_n_222 ,csa_tree_add_83_21_pad_groupi_n_262);
  nor csa_tree_add_83_21_pad_groupi_g5208__5477(csa_tree_add_83_21_pad_groupi_n_519 ,csa_tree_add_83_21_pad_groupi_n_50 ,csa_tree_add_83_21_pad_groupi_n_272);
  or csa_tree_add_83_21_pad_groupi_g5209__2398(csa_tree_add_83_21_pad_groupi_n_518 ,csa_tree_add_83_21_pad_groupi_n_21 ,csa_tree_add_83_21_pad_groupi_n_266);
  nor csa_tree_add_83_21_pad_groupi_g5210__5107(csa_tree_add_83_21_pad_groupi_n_517 ,csa_tree_add_83_21_pad_groupi_n_178 ,csa_tree_add_83_21_pad_groupi_n_274);
  nor csa_tree_add_83_21_pad_groupi_g5211__6260(csa_tree_add_83_21_pad_groupi_n_516 ,csa_tree_add_83_21_pad_groupi_n_225 ,csa_tree_add_83_21_pad_groupi_n_263);
  nor csa_tree_add_83_21_pad_groupi_g5212__4319(csa_tree_add_83_21_pad_groupi_n_515 ,csa_tree_add_83_21_pad_groupi_n_47 ,csa_tree_add_83_21_pad_groupi_n_268);
  nor csa_tree_add_83_21_pad_groupi_g5213__8428(csa_tree_add_83_21_pad_groupi_n_514 ,csa_tree_add_83_21_pad_groupi_n_197 ,csa_tree_add_83_21_pad_groupi_n_333);
  nor csa_tree_add_83_21_pad_groupi_g5214__5526(csa_tree_add_83_21_pad_groupi_n_513 ,csa_tree_add_83_21_pad_groupi_n_227 ,csa_tree_add_83_21_pad_groupi_n_320);
  nor csa_tree_add_83_21_pad_groupi_g5215__6783(csa_tree_add_83_21_pad_groupi_n_512 ,csa_tree_add_83_21_pad_groupi_n_59 ,csa_tree_add_83_21_pad_groupi_n_342);
  or csa_tree_add_83_21_pad_groupi_g5217__3680(csa_tree_add_83_21_pad_groupi_n_583 ,csa_tree_add_83_21_pad_groupi_n_121 ,csa_tree_add_83_21_pad_groupi_n_424);
  or csa_tree_add_83_21_pad_groupi_g5218__1617(csa_tree_add_83_21_pad_groupi_n_582 ,csa_tree_add_83_21_pad_groupi_n_162 ,csa_tree_add_83_21_pad_groupi_n_402);
  or csa_tree_add_83_21_pad_groupi_g5219__2802(csa_tree_add_83_21_pad_groupi_n_581 ,csa_tree_add_83_21_pad_groupi_n_121 ,csa_tree_add_83_21_pad_groupi_n_109);
  or csa_tree_add_83_21_pad_groupi_g5220__1705(csa_tree_add_83_21_pad_groupi_n_580 ,csa_tree_add_83_21_pad_groupi_n_162 ,csa_tree_add_83_21_pad_groupi_n_404);
  or csa_tree_add_83_21_pad_groupi_g5221__5122(csa_tree_add_83_21_pad_groupi_n_579 ,csa_tree_add_83_21_pad_groupi_n_163 ,csa_tree_add_83_21_pad_groupi_n_403);
  not csa_tree_add_83_21_pad_groupi_g5223(csa_tree_add_83_21_pad_groupi_n_510 ,csa_tree_add_83_21_pad_groupi_n_505);
  not csa_tree_add_83_21_pad_groupi_g5224(csa_tree_add_83_21_pad_groupi_n_509 ,csa_tree_add_83_21_pad_groupi_n_505);
  not csa_tree_add_83_21_pad_groupi_g5225(csa_tree_add_83_21_pad_groupi_n_508 ,csa_tree_add_83_21_pad_groupi_n_506);
  not csa_tree_add_83_21_pad_groupi_g5226(csa_tree_add_83_21_pad_groupi_n_507 ,csa_tree_add_83_21_pad_groupi_n_506);
  not csa_tree_add_83_21_pad_groupi_g5227(csa_tree_add_83_21_pad_groupi_n_506 ,csa_tree_add_83_21_pad_groupi_n_505);
  not csa_tree_add_83_21_pad_groupi_g5228(csa_tree_add_83_21_pad_groupi_n_504 ,csa_tree_add_83_21_pad_groupi_n_499);
  not csa_tree_add_83_21_pad_groupi_g5229(csa_tree_add_83_21_pad_groupi_n_503 ,csa_tree_add_83_21_pad_groupi_n_499);
  not csa_tree_add_83_21_pad_groupi_g5230(csa_tree_add_83_21_pad_groupi_n_502 ,csa_tree_add_83_21_pad_groupi_n_500);
  not csa_tree_add_83_21_pad_groupi_g5231(csa_tree_add_83_21_pad_groupi_n_501 ,csa_tree_add_83_21_pad_groupi_n_500);
  not csa_tree_add_83_21_pad_groupi_g5232(csa_tree_add_83_21_pad_groupi_n_500 ,csa_tree_add_83_21_pad_groupi_n_499);
  not csa_tree_add_83_21_pad_groupi_g5233(csa_tree_add_83_21_pad_groupi_n_498 ,csa_tree_add_83_21_pad_groupi_n_278);
  not csa_tree_add_83_21_pad_groupi_g5234(csa_tree_add_83_21_pad_groupi_n_496 ,csa_tree_add_83_21_pad_groupi_n_497);
  not csa_tree_add_83_21_pad_groupi_g5235(csa_tree_add_83_21_pad_groupi_n_495 ,csa_tree_add_83_21_pad_groupi_n_493);
  not csa_tree_add_83_21_pad_groupi_g5236(csa_tree_add_83_21_pad_groupi_n_494 ,csa_tree_add_83_21_pad_groupi_n_493);
  or csa_tree_add_83_21_pad_groupi_g5237__8246(csa_tree_add_83_21_pad_groupi_n_492 ,csa_tree_add_83_21_pad_groupi_n_27 ,csa_tree_add_83_21_pad_groupi_n_311);
  nor csa_tree_add_83_21_pad_groupi_g5238__7098(csa_tree_add_83_21_pad_groupi_n_491 ,csa_tree_add_83_21_pad_groupi_n_180 ,csa_tree_add_83_21_pad_groupi_n_329);
  nor csa_tree_add_83_21_pad_groupi_g5239__6131(csa_tree_add_83_21_pad_groupi_n_490 ,csa_tree_add_83_21_pad_groupi_n_220 ,csa_tree_add_83_21_pad_groupi_n_271);
  nor csa_tree_add_83_21_pad_groupi_g5240__1881(csa_tree_add_83_21_pad_groupi_n_489 ,csa_tree_add_83_21_pad_groupi_n_82 ,csa_tree_add_83_21_pad_groupi_n_275);
  nor csa_tree_add_83_21_pad_groupi_g5241__5115(csa_tree_add_83_21_pad_groupi_n_488 ,csa_tree_add_83_21_pad_groupi_n_181 ,csa_tree_add_83_21_pad_groupi_n_309);
  nor csa_tree_add_83_21_pad_groupi_g5242__7482(csa_tree_add_83_21_pad_groupi_n_487 ,csa_tree_add_83_21_pad_groupi_n_88 ,csa_tree_add_83_21_pad_groupi_n_341);
  nor csa_tree_add_83_21_pad_groupi_g5243__4733(csa_tree_add_83_21_pad_groupi_n_486 ,csa_tree_add_83_21_pad_groupi_n_227 ,csa_tree_add_83_21_pad_groupi_n_306);
  or csa_tree_add_83_21_pad_groupi_g5244__6161(csa_tree_add_83_21_pad_groupi_n_485 ,csa_tree_add_83_21_pad_groupi_n_30 ,csa_tree_add_83_21_pad_groupi_n_302);
  nor csa_tree_add_83_21_pad_groupi_g5245(csa_tree_add_83_21_pad_groupi_n_484 ,csa_tree_add_83_21_pad_groupi_n_174 ,csa_tree_add_83_21_pad_groupi_n_315);
  or csa_tree_add_83_21_pad_groupi_g5246(csa_tree_add_83_21_pad_groupi_n_483 ,csa_tree_add_83_21_pad_groupi_n_30 ,csa_tree_add_83_21_pad_groupi_n_263);
  nor csa_tree_add_83_21_pad_groupi_g5247(csa_tree_add_83_21_pad_groupi_n_482 ,csa_tree_add_83_21_pad_groupi_n_96 ,csa_tree_add_83_21_pad_groupi_n_338);
  nor csa_tree_add_83_21_pad_groupi_g5248(csa_tree_add_83_21_pad_groupi_n_481 ,csa_tree_add_83_21_pad_groupi_n_233 ,csa_tree_add_83_21_pad_groupi_n_269);
  nor csa_tree_add_83_21_pad_groupi_g5249(csa_tree_add_83_21_pad_groupi_n_480 ,csa_tree_add_83_21_pad_groupi_n_25 ,csa_tree_add_83_21_pad_groupi_n_272);
  nor csa_tree_add_83_21_pad_groupi_g5250(csa_tree_add_83_21_pad_groupi_n_479 ,csa_tree_add_83_21_pad_groupi_n_214 ,csa_tree_add_83_21_pad_groupi_n_266);
  nor csa_tree_add_83_21_pad_groupi_g5251(csa_tree_add_83_21_pad_groupi_n_478 ,csa_tree_add_83_21_pad_groupi_n_235 ,csa_tree_add_83_21_pad_groupi_n_332);
  nor csa_tree_add_83_21_pad_groupi_g5252(csa_tree_add_83_21_pad_groupi_n_477 ,csa_tree_add_83_21_pad_groupi_n_73 ,csa_tree_add_83_21_pad_groupi_n_342);
  nor csa_tree_add_83_21_pad_groupi_g5253(csa_tree_add_83_21_pad_groupi_n_476 ,csa_tree_add_83_21_pad_groupi_n_206 ,csa_tree_add_83_21_pad_groupi_n_314);
  nor csa_tree_add_83_21_pad_groupi_g5254(csa_tree_add_83_21_pad_groupi_n_475 ,csa_tree_add_83_21_pad_groupi_n_69 ,csa_tree_add_83_21_pad_groupi_n_308);
  nor csa_tree_add_83_21_pad_groupi_g5255(csa_tree_add_83_21_pad_groupi_n_474 ,csa_tree_add_83_21_pad_groupi_n_209 ,csa_tree_add_83_21_pad_groupi_n_303);
  nor csa_tree_add_83_21_pad_groupi_g5256(csa_tree_add_83_21_pad_groupi_n_473 ,csa_tree_add_83_21_pad_groupi_n_76 ,csa_tree_add_83_21_pad_groupi_n_314);
  or csa_tree_add_83_21_pad_groupi_g5257(csa_tree_add_83_21_pad_groupi_n_472 ,csa_tree_add_83_21_pad_groupi_n_45 ,csa_tree_add_83_21_pad_groupi_n_308);
  nor csa_tree_add_83_21_pad_groupi_g5258(csa_tree_add_83_21_pad_groupi_n_471 ,csa_tree_add_83_21_pad_groupi_n_211 ,csa_tree_add_83_21_pad_groupi_n_303);
  nor csa_tree_add_83_21_pad_groupi_g5259(csa_tree_add_83_21_pad_groupi_n_470 ,csa_tree_add_83_21_pad_groupi_n_67 ,csa_tree_add_83_21_pad_groupi_n_333);
  nor csa_tree_add_83_21_pad_groupi_g5260(csa_tree_add_83_21_pad_groupi_n_469 ,csa_tree_add_83_21_pad_groupi_n_180 ,csa_tree_add_83_21_pad_groupi_n_300);
  nor csa_tree_add_83_21_pad_groupi_g5261(csa_tree_add_83_21_pad_groupi_n_468 ,csa_tree_add_83_21_pad_groupi_n_177 ,csa_tree_add_83_21_pad_groupi_n_399);
  nor csa_tree_add_83_21_pad_groupi_g5262(csa_tree_add_83_21_pad_groupi_n_467 ,csa_tree_add_83_21_pad_groupi_n_52 ,csa_tree_add_83_21_pad_groupi_n_291);
  nor csa_tree_add_83_21_pad_groupi_g5263(csa_tree_add_83_21_pad_groupi_n_466 ,csa_tree_add_83_21_pad_groupi_n_45 ,csa_tree_add_83_21_pad_groupi_n_290);
  nor csa_tree_add_83_21_pad_groupi_g5264(csa_tree_add_83_21_pad_groupi_n_465 ,csa_tree_add_83_21_pad_groupi_n_175 ,csa_tree_add_83_21_pad_groupi_n_297);
  or csa_tree_add_83_21_pad_groupi_g5265(csa_tree_add_83_21_pad_groupi_n_464 ,csa_tree_add_83_21_pad_groupi_n_36 ,csa_tree_add_83_21_pad_groupi_n_296);
  nor csa_tree_add_83_21_pad_groupi_g5266(csa_tree_add_83_21_pad_groupi_n_463 ,csa_tree_add_83_21_pad_groupi_n_90 ,csa_tree_add_83_21_pad_groupi_n_260);
  nor csa_tree_add_83_21_pad_groupi_g5267(csa_tree_add_83_21_pad_groupi_n_462 ,csa_tree_add_83_21_pad_groupi_n_212 ,csa_tree_add_83_21_pad_groupi_n_299);
  nor csa_tree_add_83_21_pad_groupi_g5268(csa_tree_add_83_21_pad_groupi_n_461 ,csa_tree_add_83_21_pad_groupi_n_95 ,csa_tree_add_83_21_pad_groupi_n_299);
  or csa_tree_add_83_21_pad_groupi_g5269(csa_tree_add_83_21_pad_groupi_n_460 ,csa_tree_add_83_21_pad_groupi_n_39 ,csa_tree_add_83_21_pad_groupi_n_290);
  nor csa_tree_add_83_21_pad_groupi_g5271(csa_tree_add_83_21_pad_groupi_n_458 ,csa_tree_add_83_21_pad_groupi_n_186 ,csa_tree_add_83_21_pad_groupi_n_300);
  or csa_tree_add_83_21_pad_groupi_g5272(csa_tree_add_83_21_pad_groupi_n_457 ,csa_tree_add_83_21_pad_groupi_n_21 ,csa_tree_add_83_21_pad_groupi_n_291);
  nor csa_tree_add_83_21_pad_groupi_g5273(csa_tree_add_83_21_pad_groupi_n_456 ,csa_tree_add_83_21_pad_groupi_n_98 ,csa_tree_add_83_21_pad_groupi_n_296);
  nor csa_tree_add_83_21_pad_groupi_g5274(csa_tree_add_83_21_pad_groupi_n_455 ,csa_tree_add_83_21_pad_groupi_n_207 ,csa_tree_add_83_21_pad_groupi_n_297);
  nor csa_tree_add_83_21_pad_groupi_g5284(csa_tree_add_83_21_pad_groupi_n_445 ,csa_tree_add_83_21_pad_groupi_n_106 ,csa_tree_add_83_21_pad_groupi_n_294);
  nor csa_tree_add_83_21_pad_groupi_g5290(csa_tree_add_83_21_pad_groupi_n_439 ,csa_tree_add_83_21_pad_groupi_n_109 ,csa_tree_add_83_21_pad_groupi_n_241);
  or csa_tree_add_83_21_pad_groupi_g5291(csa_tree_add_83_21_pad_groupi_n_438 ,csa_tree_add_83_21_pad_groupi_n_32 ,csa_tree_add_83_21_pad_groupi_n_103);
  nor csa_tree_add_83_21_pad_groupi_g5294(csa_tree_add_83_21_pad_groupi_n_435 ,csa_tree_add_83_21_pad_groupi_n_107 ,csa_tree_add_83_21_pad_groupi_n_240);
  or csa_tree_add_83_21_pad_groupi_g5295(csa_tree_add_83_21_pad_groupi_n_434 ,csa_tree_add_83_21_pad_groupi_n_293 ,csa_tree_add_83_21_pad_groupi_n_110);
  nor csa_tree_add_83_21_pad_groupi_g5296(csa_tree_add_83_21_pad_groupi_n_433 ,csa_tree_add_83_21_pad_groupi_n_103 ,csa_tree_add_83_21_pad_groupi_n_294);
  or csa_tree_add_83_21_pad_groupi_g5297(csa_tree_add_83_21_pad_groupi_n_432 ,csa_tree_add_83_21_pad_groupi_n_13 ,csa_tree_add_83_21_pad_groupi_n_61);
  nor csa_tree_add_83_21_pad_groupi_g5298(csa_tree_add_83_21_pad_groupi_n_431 ,csa_tree_add_83_21_pad_groupi_n_110 ,csa_tree_add_83_21_pad_groupi_n_238);
  or csa_tree_add_83_21_pad_groupi_g5299(csa_tree_add_83_21_pad_groupi_n_430 ,csa_tree_add_83_21_pad_groupi_n_13 ,csa_tree_add_83_21_pad_groupi_n_104);
  nor csa_tree_add_83_21_pad_groupi_g5300(csa_tree_add_83_21_pad_groupi_n_429 ,csa_tree_add_83_21_pad_groupi_n_61 ,csa_tree_add_83_21_pad_groupi_n_32);
  nor csa_tree_add_83_21_pad_groupi_g5301(csa_tree_add_83_21_pad_groupi_n_428 ,csa_tree_add_83_21_pad_groupi_n_249 ,csa_tree_add_83_21_pad_groupi_n_34);
  or csa_tree_add_83_21_pad_groupi_g5302(csa_tree_add_83_21_pad_groupi_n_427 ,csa_tree_add_83_21_pad_groupi_n_15 ,csa_tree_add_83_21_pad_groupi_n_106);
  or csa_tree_add_83_21_pad_groupi_g5303(csa_tree_add_83_21_pad_groupi_n_426 ,csa_tree_add_83_21_pad_groupi_n_34 ,csa_tree_add_83_21_pad_groupi_n_107);
  nor csa_tree_add_83_21_pad_groupi_g5304(csa_tree_add_83_21_pad_groupi_n_425 ,csa_tree_add_83_21_pad_groupi_n_104 ,csa_tree_add_83_21_pad_groupi_n_237);
  or csa_tree_add_83_21_pad_groupi_g5305(csa_tree_add_83_21_pad_groupi_n_511 ,csa_tree_add_83_21_pad_groupi_n_154 ,csa_tree_add_83_21_pad_groupi_n_424);
  or csa_tree_add_83_21_pad_groupi_g5306(csa_tree_add_83_21_pad_groupi_n_505 ,csa_tree_add_83_21_pad_groupi_n_150 ,csa_tree_add_83_21_pad_groupi_n_403);
  or csa_tree_add_83_21_pad_groupi_g5307(csa_tree_add_83_21_pad_groupi_n_499 ,csa_tree_add_83_21_pad_groupi_n_155 ,csa_tree_add_83_21_pad_groupi_n_402);
  or csa_tree_add_83_21_pad_groupi_g5309(csa_tree_add_83_21_pad_groupi_n_493 ,csa_tree_add_83_21_pad_groupi_n_152 ,csa_tree_add_83_21_pad_groupi_n_404);
  not csa_tree_add_83_21_pad_groupi_g5311(csa_tree_add_83_21_pad_groupi_n_423 ,csa_tree_add_83_21_pad_groupi_n_158);
  not csa_tree_add_83_21_pad_groupi_g5312(csa_tree_add_83_21_pad_groupi_n_422 ,csa_tree_add_83_21_pad_groupi_n_155);
  not csa_tree_add_83_21_pad_groupi_g5315(csa_tree_add_83_21_pad_groupi_n_419 ,csa_tree_add_83_21_pad_groupi_n_154);
  not csa_tree_add_83_21_pad_groupi_g5317(csa_tree_add_83_21_pad_groupi_n_418 ,csa_tree_add_83_21_pad_groupi_n_149);
  not csa_tree_add_83_21_pad_groupi_g5319(csa_tree_add_83_21_pad_groupi_n_416 ,csa_tree_add_83_21_pad_groupi_n_152);
  not csa_tree_add_83_21_pad_groupi_g5321(csa_tree_add_83_21_pad_groupi_n_415 ,csa_tree_add_83_21_pad_groupi_n_151);
  not csa_tree_add_83_21_pad_groupi_g5323(csa_tree_add_83_21_pad_groupi_n_414 ,csa_tree_add_83_21_pad_groupi_n_160);
  not csa_tree_add_83_21_pad_groupi_g5324(csa_tree_add_83_21_pad_groupi_n_413 ,csa_tree_add_83_21_pad_groupi_n_153);
  not csa_tree_add_83_21_pad_groupi_g5327(csa_tree_add_83_21_pad_groupi_n_411 ,csa_tree_add_83_21_pad_groupi_n_159);
  not csa_tree_add_83_21_pad_groupi_g5328(csa_tree_add_83_21_pad_groupi_n_410 ,csa_tree_add_83_21_pad_groupi_n_150);
  or csa_tree_add_83_21_pad_groupi_g5331(csa_tree_add_83_21_pad_groupi_n_406 ,in8[10] ,in8[9]);
  and csa_tree_add_83_21_pad_groupi_g5332(csa_tree_add_83_21_pad_groupi_n_424 ,csa_tree_add_83_21_pad_groupi_n_375 ,csa_tree_add_83_21_pad_groupi_n_388);
  and csa_tree_add_83_21_pad_groupi_g5333(csa_tree_add_83_21_pad_groupi_n_421 ,n_673 ,n_680);
  and csa_tree_add_83_21_pad_groupi_g5334(csa_tree_add_83_21_pad_groupi_n_420 ,in10[0] ,n_682);
  and csa_tree_add_83_21_pad_groupi_g5335(csa_tree_add_83_21_pad_groupi_n_417 ,n_674 ,n_681);
  and csa_tree_add_83_21_pad_groupi_g5337(csa_tree_add_83_21_pad_groupi_n_409 ,n_672 ,n_679);
  not csa_tree_add_83_21_pad_groupi_g5339(csa_tree_add_83_21_pad_groupi_n_399 ,csa_tree_add_83_21_pad_groupi_n_293);
  not csa_tree_add_83_21_pad_groupi_g5340(csa_tree_add_83_21_pad_groupi_n_398 ,csa_tree_add_83_21_pad_groupi_n_395);
  not csa_tree_add_83_21_pad_groupi_g5341(csa_tree_add_83_21_pad_groupi_n_397 ,csa_tree_add_83_21_pad_groupi_n_258);
  not csa_tree_add_83_21_pad_groupi_g5345(csa_tree_add_83_21_pad_groupi_n_396 ,csa_tree_add_83_21_pad_groupi_n_395);
  and csa_tree_add_83_21_pad_groupi_g5346(csa_tree_add_83_21_pad_groupi_n_394 ,in8[10] ,in8[9]);
  and csa_tree_add_83_21_pad_groupi_g5348(csa_tree_add_83_21_pad_groupi_n_404 ,csa_tree_add_83_21_pad_groupi_n_391 ,csa_tree_add_83_21_pad_groupi_n_393);
  and csa_tree_add_83_21_pad_groupi_g5349(csa_tree_add_83_21_pad_groupi_n_403 ,csa_tree_add_83_21_pad_groupi_n_378 ,csa_tree_add_83_21_pad_groupi_n_377);
  and csa_tree_add_83_21_pad_groupi_g5350(csa_tree_add_83_21_pad_groupi_n_402 ,csa_tree_add_83_21_pad_groupi_n_392 ,csa_tree_add_83_21_pad_groupi_n_376);
  and csa_tree_add_83_21_pad_groupi_g5351(csa_tree_add_83_21_pad_groupi_n_401 ,csa_tree_add_83_21_pad_groupi_n_390 ,csa_tree_add_83_21_pad_groupi_n_389);
  or csa_tree_add_83_21_pad_groupi_g5353(csa_tree_add_83_21_pad_groupi_n_395 ,csa_tree_add_83_21_pad_groupi_n_390 ,csa_tree_add_83_21_pad_groupi_n_389);
  not csa_tree_add_83_21_pad_groupi_g5354(csa_tree_add_83_21_pad_groupi_n_393 ,n_681);
  not csa_tree_add_83_21_pad_groupi_g5355(csa_tree_add_83_21_pad_groupi_n_392 ,n_673);
  not csa_tree_add_83_21_pad_groupi_g5356(csa_tree_add_83_21_pad_groupi_n_391 ,n_674);
  not csa_tree_add_83_21_pad_groupi_g5357(csa_tree_add_83_21_pad_groupi_n_390 ,n_676);
  not csa_tree_add_83_21_pad_groupi_g5358(csa_tree_add_83_21_pad_groupi_n_389 ,n_683);
  not csa_tree_add_83_21_pad_groupi_g5359(csa_tree_add_83_21_pad_groupi_n_388 ,n_682);
  not csa_tree_add_83_21_pad_groupi_g5360(csa_tree_add_83_21_pad_groupi_n_387 ,in8[7]);
  not csa_tree_add_83_21_pad_groupi_g5361(csa_tree_add_83_21_pad_groupi_n_386 ,in9[15]);
  not csa_tree_add_83_21_pad_groupi_g5362(csa_tree_add_83_21_pad_groupi_n_385 ,in9[2]);
  not csa_tree_add_83_21_pad_groupi_g5363(csa_tree_add_83_21_pad_groupi_n_384 ,in9[5]);
  not csa_tree_add_83_21_pad_groupi_g5364(csa_tree_add_83_21_pad_groupi_n_383 ,in9[13]);
  not csa_tree_add_83_21_pad_groupi_g5365(csa_tree_add_83_21_pad_groupi_n_382 ,in9[3]);
  not csa_tree_add_83_21_pad_groupi_g5366(csa_tree_add_83_21_pad_groupi_n_381 ,in9[9]);
  not csa_tree_add_83_21_pad_groupi_g5367(csa_tree_add_83_21_pad_groupi_n_380 ,in9[1]);
  not csa_tree_add_83_21_pad_groupi_g5368(csa_tree_add_83_21_pad_groupi_n_379 ,in9[8]);
  not csa_tree_add_83_21_pad_groupi_g5369(csa_tree_add_83_21_pad_groupi_n_378 ,n_672);
  not csa_tree_add_83_21_pad_groupi_g5370(csa_tree_add_83_21_pad_groupi_n_377 ,n_679);
  not csa_tree_add_83_21_pad_groupi_g5371(csa_tree_add_83_21_pad_groupi_n_376 ,n_680);
  not csa_tree_add_83_21_pad_groupi_g5372(csa_tree_add_83_21_pad_groupi_n_375 ,in10[0]);
  not csa_tree_add_83_21_pad_groupi_g5373(csa_tree_add_83_21_pad_groupi_n_374 ,in8[0]);
  not csa_tree_add_83_21_pad_groupi_g5374(csa_tree_add_83_21_pad_groupi_n_373 ,in8[11]);
  not csa_tree_add_83_21_pad_groupi_g5375(csa_tree_add_83_21_pad_groupi_n_372 ,in8[8]);
  not csa_tree_add_83_21_pad_groupi_g5376(csa_tree_add_83_21_pad_groupi_n_371 ,in8[1]);
  not csa_tree_add_83_21_pad_groupi_g5377(csa_tree_add_83_21_pad_groupi_n_370 ,in8[6]);
  not csa_tree_add_83_21_pad_groupi_g5378(csa_tree_add_83_21_pad_groupi_n_369 ,in8[9]);
  not csa_tree_add_83_21_pad_groupi_g5379(csa_tree_add_83_21_pad_groupi_n_368 ,in9[0]);
  not csa_tree_add_83_21_pad_groupi_g5380(csa_tree_add_83_21_pad_groupi_n_367 ,in9[4]);
  not csa_tree_add_83_21_pad_groupi_g5381(csa_tree_add_83_21_pad_groupi_n_366 ,in9[12]);
  not csa_tree_add_83_21_pad_groupi_g5382(csa_tree_add_83_21_pad_groupi_n_365 ,in9[11]);
  not csa_tree_add_83_21_pad_groupi_g5383(csa_tree_add_83_21_pad_groupi_n_364 ,in9[7]);
  not csa_tree_add_83_21_pad_groupi_g5384(csa_tree_add_83_21_pad_groupi_n_363 ,in9[10]);
  not csa_tree_add_83_21_pad_groupi_g5385(csa_tree_add_83_21_pad_groupi_n_362 ,in9[6]);
  not csa_tree_add_83_21_pad_groupi_g5386(csa_tree_add_83_21_pad_groupi_n_361 ,in9[14]);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5534(csa_tree_add_83_21_pad_groupi_n_345 ,csa_tree_add_83_21_pad_groupi_n_343);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5535(csa_tree_add_83_21_pad_groupi_n_344 ,csa_tree_add_83_21_pad_groupi_n_343);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5536(csa_tree_add_83_21_pad_groupi_n_343 ,csa_tree_add_83_21_pad_groupi_n_356);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5538(csa_tree_add_83_21_pad_groupi_n_342 ,csa_tree_add_83_21_pad_groupi_n_340);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5539(csa_tree_add_83_21_pad_groupi_n_341 ,csa_tree_add_83_21_pad_groupi_n_340);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5540(csa_tree_add_83_21_pad_groupi_n_340 ,csa_tree_add_83_21_pad_groupi_n_422);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5542(csa_tree_add_83_21_pad_groupi_n_339 ,csa_tree_add_83_21_pad_groupi_n_337);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5543(csa_tree_add_83_21_pad_groupi_n_338 ,csa_tree_add_83_21_pad_groupi_n_337);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5544(csa_tree_add_83_21_pad_groupi_n_337 ,csa_tree_add_83_21_pad_groupi_n_413);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5546(csa_tree_add_83_21_pad_groupi_n_336 ,csa_tree_add_83_21_pad_groupi_n_334);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5547(csa_tree_add_83_21_pad_groupi_n_335 ,csa_tree_add_83_21_pad_groupi_n_334);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5548(csa_tree_add_83_21_pad_groupi_n_334 ,csa_tree_add_83_21_pad_groupi_n_348);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5550(csa_tree_add_83_21_pad_groupi_n_333 ,csa_tree_add_83_21_pad_groupi_n_331);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5551(csa_tree_add_83_21_pad_groupi_n_332 ,csa_tree_add_83_21_pad_groupi_n_331);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5552(csa_tree_add_83_21_pad_groupi_n_331 ,csa_tree_add_83_21_pad_groupi_n_411);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5554(csa_tree_add_83_21_pad_groupi_n_330 ,csa_tree_add_83_21_pad_groupi_n_328);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5555(csa_tree_add_83_21_pad_groupi_n_329 ,csa_tree_add_83_21_pad_groupi_n_328);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5556(csa_tree_add_83_21_pad_groupi_n_328 ,csa_tree_add_83_21_pad_groupi_n_410);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5558(csa_tree_add_83_21_pad_groupi_n_327 ,csa_tree_add_83_21_pad_groupi_n_325);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5559(csa_tree_add_83_21_pad_groupi_n_326 ,csa_tree_add_83_21_pad_groupi_n_325);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5560(csa_tree_add_83_21_pad_groupi_n_325 ,csa_tree_add_83_21_pad_groupi_n_350);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5562(csa_tree_add_83_21_pad_groupi_n_324 ,csa_tree_add_83_21_pad_groupi_n_322);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5563(csa_tree_add_83_21_pad_groupi_n_323 ,csa_tree_add_83_21_pad_groupi_n_322);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5564(csa_tree_add_83_21_pad_groupi_n_322 ,csa_tree_add_83_21_pad_groupi_n_419);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5566(csa_tree_add_83_21_pad_groupi_n_321 ,csa_tree_add_83_21_pad_groupi_n_319);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5567(csa_tree_add_83_21_pad_groupi_n_320 ,csa_tree_add_83_21_pad_groupi_n_319);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5568(csa_tree_add_83_21_pad_groupi_n_319 ,csa_tree_add_83_21_pad_groupi_n_416);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5570(csa_tree_add_83_21_pad_groupi_n_318 ,csa_tree_add_83_21_pad_groupi_n_316);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5571(csa_tree_add_83_21_pad_groupi_n_317 ,csa_tree_add_83_21_pad_groupi_n_316);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5572(csa_tree_add_83_21_pad_groupi_n_316 ,csa_tree_add_83_21_pad_groupi_n_351);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5574(csa_tree_add_83_21_pad_groupi_n_315 ,csa_tree_add_83_21_pad_groupi_n_313);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5575(csa_tree_add_83_21_pad_groupi_n_314 ,csa_tree_add_83_21_pad_groupi_n_313);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5576(csa_tree_add_83_21_pad_groupi_n_313 ,csa_tree_add_83_21_pad_groupi_n_415);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5578(csa_tree_add_83_21_pad_groupi_n_312 ,csa_tree_add_83_21_pad_groupi_n_310);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5579(csa_tree_add_83_21_pad_groupi_n_311 ,csa_tree_add_83_21_pad_groupi_n_310);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5580(csa_tree_add_83_21_pad_groupi_n_310 ,csa_tree_add_83_21_pad_groupi_n_423);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5582(csa_tree_add_83_21_pad_groupi_n_309 ,csa_tree_add_83_21_pad_groupi_n_307);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5583(csa_tree_add_83_21_pad_groupi_n_308 ,csa_tree_add_83_21_pad_groupi_n_307);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5584(csa_tree_add_83_21_pad_groupi_n_307 ,csa_tree_add_83_21_pad_groupi_n_414);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5586(csa_tree_add_83_21_pad_groupi_n_306 ,csa_tree_add_83_21_pad_groupi_n_304);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5587(csa_tree_add_83_21_pad_groupi_n_305 ,csa_tree_add_83_21_pad_groupi_n_304);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5588(csa_tree_add_83_21_pad_groupi_n_304 ,csa_tree_add_83_21_pad_groupi_n_353);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5590(csa_tree_add_83_21_pad_groupi_n_303 ,csa_tree_add_83_21_pad_groupi_n_301);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5591(csa_tree_add_83_21_pad_groupi_n_302 ,csa_tree_add_83_21_pad_groupi_n_301);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5592(csa_tree_add_83_21_pad_groupi_n_301 ,csa_tree_add_83_21_pad_groupi_n_418);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5594(csa_tree_add_83_21_pad_groupi_n_300 ,csa_tree_add_83_21_pad_groupi_n_298);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5595(csa_tree_add_83_21_pad_groupi_n_299 ,csa_tree_add_83_21_pad_groupi_n_298);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5596(csa_tree_add_83_21_pad_groupi_n_298 ,csa_tree_add_83_21_pad_groupi_n_397);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5598(csa_tree_add_83_21_pad_groupi_n_297 ,csa_tree_add_83_21_pad_groupi_n_295);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5599(csa_tree_add_83_21_pad_groupi_n_296 ,csa_tree_add_83_21_pad_groupi_n_295);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5600(csa_tree_add_83_21_pad_groupi_n_295 ,csa_tree_add_83_21_pad_groupi_n_346);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5602(csa_tree_add_83_21_pad_groupi_n_294 ,csa_tree_add_83_21_pad_groupi_n_292);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5603(csa_tree_add_83_21_pad_groupi_n_293 ,csa_tree_add_83_21_pad_groupi_n_292);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5604(csa_tree_add_83_21_pad_groupi_n_292 ,csa_tree_add_83_21_pad_groupi_n_398);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5606(csa_tree_add_83_21_pad_groupi_n_291 ,csa_tree_add_83_21_pad_groupi_n_289);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5607(csa_tree_add_83_21_pad_groupi_n_290 ,csa_tree_add_83_21_pad_groupi_n_289);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5608(csa_tree_add_83_21_pad_groupi_n_289 ,csa_tree_add_83_21_pad_groupi_n_397);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5610(csa_tree_add_83_21_pad_groupi_n_288 ,csa_tree_add_83_21_pad_groupi_n_286);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5611(csa_tree_add_83_21_pad_groupi_n_287 ,csa_tree_add_83_21_pad_groupi_n_286);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5612(csa_tree_add_83_21_pad_groupi_n_286 ,csa_tree_add_83_21_pad_groupi_n_509);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5614(csa_tree_add_83_21_pad_groupi_n_285 ,csa_tree_add_83_21_pad_groupi_n_283);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5615(csa_tree_add_83_21_pad_groupi_n_284 ,csa_tree_add_83_21_pad_groupi_n_283);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5616(csa_tree_add_83_21_pad_groupi_n_283 ,csa_tree_add_83_21_pad_groupi_n_503);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5620(csa_tree_add_83_21_pad_groupi_n_358 ,csa_tree_add_83_21_pad_groupi_n_581);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5623(csa_tree_add_83_21_pad_groupi_n_282 ,csa_tree_add_83_21_pad_groupi_n_281);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5624(csa_tree_add_83_21_pad_groupi_n_281 ,csa_tree_add_83_21_pad_groupi_n_579);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5627(csa_tree_add_83_21_pad_groupi_n_280 ,csa_tree_add_83_21_pad_groupi_n_279);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5628(csa_tree_add_83_21_pad_groupi_n_279 ,csa_tree_add_83_21_pad_groupi_n_582);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5632(csa_tree_add_83_21_pad_groupi_n_357 ,csa_tree_add_83_21_pad_groupi_n_580);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5635(csa_tree_add_83_21_pad_groupi_n_278 ,csa_tree_add_83_21_pad_groupi_n_277);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5636(csa_tree_add_83_21_pad_groupi_n_277 ,csa_tree_add_83_21_pad_groupi_n_497);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5639(csa_tree_add_83_21_pad_groupi_n_276 ,csa_tree_add_83_21_pad_groupi_n_359);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5640(csa_tree_add_83_21_pad_groupi_n_359 ,csa_tree_add_83_21_pad_groupi_n_934);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5642(csa_tree_add_83_21_pad_groupi_n_275 ,csa_tree_add_83_21_pad_groupi_n_273);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5643(csa_tree_add_83_21_pad_groupi_n_274 ,csa_tree_add_83_21_pad_groupi_n_273);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5644(csa_tree_add_83_21_pad_groupi_n_273 ,csa_tree_add_83_21_pad_groupi_n_355);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5646(csa_tree_add_83_21_pad_groupi_n_272 ,csa_tree_add_83_21_pad_groupi_n_270);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5647(csa_tree_add_83_21_pad_groupi_n_271 ,csa_tree_add_83_21_pad_groupi_n_270);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5648(csa_tree_add_83_21_pad_groupi_n_270 ,csa_tree_add_83_21_pad_groupi_n_349);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5650(csa_tree_add_83_21_pad_groupi_n_269 ,csa_tree_add_83_21_pad_groupi_n_267);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5651(csa_tree_add_83_21_pad_groupi_n_268 ,csa_tree_add_83_21_pad_groupi_n_267);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5652(csa_tree_add_83_21_pad_groupi_n_267 ,csa_tree_add_83_21_pad_groupi_n_347);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5654(csa_tree_add_83_21_pad_groupi_n_266 ,csa_tree_add_83_21_pad_groupi_n_264);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5655(csa_tree_add_83_21_pad_groupi_n_265 ,csa_tree_add_83_21_pad_groupi_n_264);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5656(csa_tree_add_83_21_pad_groupi_n_264 ,csa_tree_add_83_21_pad_groupi_n_354);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5658(csa_tree_add_83_21_pad_groupi_n_263 ,csa_tree_add_83_21_pad_groupi_n_261);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5659(csa_tree_add_83_21_pad_groupi_n_262 ,csa_tree_add_83_21_pad_groupi_n_261);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5660(csa_tree_add_83_21_pad_groupi_n_261 ,csa_tree_add_83_21_pad_groupi_n_352);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5662(csa_tree_add_83_21_pad_groupi_n_260 ,csa_tree_add_83_21_pad_groupi_n_259);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5664(csa_tree_add_83_21_pad_groupi_n_259 ,csa_tree_add_83_21_pad_groupi_n_399);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5686(csa_tree_add_83_21_pad_groupi_n_258 ,csa_tree_add_83_21_pad_groupi_n_346);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5688(csa_tree_add_83_21_pad_groupi_n_346 ,csa_tree_add_83_21_pad_groupi_n_398);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5690(csa_tree_add_83_21_pad_groupi_n_257 ,csa_tree_add_83_21_pad_groupi_n_256);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5692(csa_tree_add_83_21_pad_groupi_n_256 ,csa_tree_add_83_21_pad_groupi_n_507);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5694(csa_tree_add_83_21_pad_groupi_n_255 ,csa_tree_add_83_21_pad_groupi_n_254);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5696(csa_tree_add_83_21_pad_groupi_n_254 ,csa_tree_add_83_21_pad_groupi_n_501);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5709(csa_tree_add_83_21_pad_groupi_n_253 ,csa_tree_add_83_21_pad_groupi_n_251);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5710(csa_tree_add_83_21_pad_groupi_n_252 ,csa_tree_add_83_21_pad_groupi_n_251);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5711(csa_tree_add_83_21_pad_groupi_n_251 ,csa_tree_add_83_21_pad_groupi_n_511);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5713(csa_tree_add_83_21_pad_groupi_n_250 ,csa_tree_add_83_21_pad_groupi_n_248);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5714(csa_tree_add_83_21_pad_groupi_n_249 ,csa_tree_add_83_21_pad_groupi_n_248);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5715(csa_tree_add_83_21_pad_groupi_n_248 ,csa_tree_add_83_21_pad_groupi_n_401);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5721(csa_tree_add_83_21_pad_groupi_n_247 ,csa_tree_add_83_21_pad_groupi_n_245);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5722(csa_tree_add_83_21_pad_groupi_n_246 ,csa_tree_add_83_21_pad_groupi_n_245);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5723(csa_tree_add_83_21_pad_groupi_n_245 ,csa_tree_add_83_21_pad_groupi_n_385);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5733(csa_tree_add_83_21_pad_groupi_n_244 ,csa_tree_add_83_21_pad_groupi_n_242);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5734(csa_tree_add_83_21_pad_groupi_n_243 ,csa_tree_add_83_21_pad_groupi_n_242);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5735(csa_tree_add_83_21_pad_groupi_n_242 ,csa_tree_add_83_21_pad_groupi_n_368);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5737(csa_tree_add_83_21_pad_groupi_n_241 ,csa_tree_add_83_21_pad_groupi_n_239);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5738(csa_tree_add_83_21_pad_groupi_n_240 ,csa_tree_add_83_21_pad_groupi_n_239);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5739(csa_tree_add_83_21_pad_groupi_n_239 ,csa_tree_add_83_21_pad_groupi_n_396);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5741(csa_tree_add_83_21_pad_groupi_n_238 ,csa_tree_add_83_21_pad_groupi_n_236);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5742(csa_tree_add_83_21_pad_groupi_n_237 ,csa_tree_add_83_21_pad_groupi_n_236);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5743(csa_tree_add_83_21_pad_groupi_n_236 ,csa_tree_add_83_21_pad_groupi_n_396);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5746(csa_tree_add_83_21_pad_groupi_n_235 ,csa_tree_add_83_21_pad_groupi_n_234);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5747(csa_tree_add_83_21_pad_groupi_n_234 ,csa_tree_add_83_21_pad_groupi_n_381);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5750(csa_tree_add_83_21_pad_groupi_n_233 ,csa_tree_add_83_21_pad_groupi_n_232);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5751(csa_tree_add_83_21_pad_groupi_n_232 ,csa_tree_add_83_21_pad_groupi_n_366);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5754(csa_tree_add_83_21_pad_groupi_n_231 ,csa_tree_add_83_21_pad_groupi_n_230);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5755(csa_tree_add_83_21_pad_groupi_n_230 ,csa_tree_add_83_21_pad_groupi_n_382);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5758(csa_tree_add_83_21_pad_groupi_n_229 ,csa_tree_add_83_21_pad_groupi_n_228);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5759(csa_tree_add_83_21_pad_groupi_n_228 ,csa_tree_add_83_21_pad_groupi_n_383);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5762(csa_tree_add_83_21_pad_groupi_n_227 ,csa_tree_add_83_21_pad_groupi_n_226);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5763(csa_tree_add_83_21_pad_groupi_n_226 ,csa_tree_add_83_21_pad_groupi_n_365);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5766(csa_tree_add_83_21_pad_groupi_n_225 ,csa_tree_add_83_21_pad_groupi_n_224);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5767(csa_tree_add_83_21_pad_groupi_n_224 ,csa_tree_add_83_21_pad_groupi_n_363);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5769(csa_tree_add_83_21_pad_groupi_n_223 ,csa_tree_add_83_21_pad_groupi_n_221);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5770(csa_tree_add_83_21_pad_groupi_n_222 ,csa_tree_add_83_21_pad_groupi_n_221);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5771(csa_tree_add_83_21_pad_groupi_n_221 ,csa_tree_add_83_21_pad_groupi_n_366);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5774(csa_tree_add_83_21_pad_groupi_n_220 ,csa_tree_add_83_21_pad_groupi_n_219);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5775(csa_tree_add_83_21_pad_groupi_n_219 ,csa_tree_add_83_21_pad_groupi_n_362);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5777(csa_tree_add_83_21_pad_groupi_n_218 ,csa_tree_add_83_21_pad_groupi_n_216);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5778(csa_tree_add_83_21_pad_groupi_n_217 ,csa_tree_add_83_21_pad_groupi_n_216);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5779(csa_tree_add_83_21_pad_groupi_n_216 ,csa_tree_add_83_21_pad_groupi_n_380);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5781(csa_tree_add_83_21_pad_groupi_n_215 ,csa_tree_add_83_21_pad_groupi_n_213);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5782(csa_tree_add_83_21_pad_groupi_n_214 ,csa_tree_add_83_21_pad_groupi_n_213);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5783(csa_tree_add_83_21_pad_groupi_n_213 ,csa_tree_add_83_21_pad_groupi_n_381);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5785(csa_tree_add_83_21_pad_groupi_n_212 ,csa_tree_add_83_21_pad_groupi_n_210);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5786(csa_tree_add_83_21_pad_groupi_n_211 ,csa_tree_add_83_21_pad_groupi_n_210);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5787(csa_tree_add_83_21_pad_groupi_n_210 ,csa_tree_add_83_21_pad_groupi_n_362);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5790(csa_tree_add_83_21_pad_groupi_n_209 ,csa_tree_add_83_21_pad_groupi_n_208);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5791(csa_tree_add_83_21_pad_groupi_n_208 ,csa_tree_add_83_21_pad_groupi_n_379);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5793(csa_tree_add_83_21_pad_groupi_n_207 ,csa_tree_add_83_21_pad_groupi_n_205);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5794(csa_tree_add_83_21_pad_groupi_n_206 ,csa_tree_add_83_21_pad_groupi_n_205);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5795(csa_tree_add_83_21_pad_groupi_n_205 ,csa_tree_add_83_21_pad_groupi_n_379);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5798(csa_tree_add_83_21_pad_groupi_n_204 ,csa_tree_add_83_21_pad_groupi_n_203);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5799(csa_tree_add_83_21_pad_groupi_n_203 ,csa_tree_add_83_21_pad_groupi_n_384);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5801(csa_tree_add_83_21_pad_groupi_n_202 ,csa_tree_add_83_21_pad_groupi_n_200);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5802(csa_tree_add_83_21_pad_groupi_n_201 ,csa_tree_add_83_21_pad_groupi_n_200);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5803(csa_tree_add_83_21_pad_groupi_n_200 ,csa_tree_add_83_21_pad_groupi_n_382);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5807(csa_tree_add_83_21_pad_groupi_n_198 ,csa_tree_add_83_21_pad_groupi_n_361);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5809(csa_tree_add_83_21_pad_groupi_n_197 ,csa_tree_add_83_21_pad_groupi_n_195);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5810(csa_tree_add_83_21_pad_groupi_n_196 ,csa_tree_add_83_21_pad_groupi_n_195);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5811(csa_tree_add_83_21_pad_groupi_n_195 ,csa_tree_add_83_21_pad_groupi_n_384);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5813(csa_tree_add_83_21_pad_groupi_n_194 ,csa_tree_add_83_21_pad_groupi_n_192);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5814(csa_tree_add_83_21_pad_groupi_n_193 ,csa_tree_add_83_21_pad_groupi_n_192);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5815(csa_tree_add_83_21_pad_groupi_n_192 ,csa_tree_add_83_21_pad_groupi_n_361);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5817(csa_tree_add_83_21_pad_groupi_n_191 ,csa_tree_add_83_21_pad_groupi_n_190);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5819(csa_tree_add_83_21_pad_groupi_n_190 ,csa_tree_add_83_21_pad_groupi_n_364);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5822(csa_tree_add_83_21_pad_groupi_n_189 ,csa_tree_add_83_21_pad_groupi_n_188);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5823(csa_tree_add_83_21_pad_groupi_n_188 ,csa_tree_add_83_21_pad_groupi_n_367);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5825(csa_tree_add_83_21_pad_groupi_n_187 ,csa_tree_add_83_21_pad_groupi_n_185);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5826(csa_tree_add_83_21_pad_groupi_n_186 ,csa_tree_add_83_21_pad_groupi_n_185);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5827(csa_tree_add_83_21_pad_groupi_n_185 ,csa_tree_add_83_21_pad_groupi_n_383);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5829(csa_tree_add_83_21_pad_groupi_n_184 ,csa_tree_add_83_21_pad_groupi_n_182);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5830(csa_tree_add_83_21_pad_groupi_n_183 ,csa_tree_add_83_21_pad_groupi_n_182);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5831(csa_tree_add_83_21_pad_groupi_n_182 ,csa_tree_add_83_21_pad_groupi_n_364);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5833(csa_tree_add_83_21_pad_groupi_n_181 ,csa_tree_add_83_21_pad_groupi_n_179);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5834(csa_tree_add_83_21_pad_groupi_n_180 ,csa_tree_add_83_21_pad_groupi_n_179);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5835(csa_tree_add_83_21_pad_groupi_n_179 ,csa_tree_add_83_21_pad_groupi_n_365);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5837(csa_tree_add_83_21_pad_groupi_n_178 ,csa_tree_add_83_21_pad_groupi_n_176);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5838(csa_tree_add_83_21_pad_groupi_n_177 ,csa_tree_add_83_21_pad_groupi_n_176);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5839(csa_tree_add_83_21_pad_groupi_n_176 ,csa_tree_add_83_21_pad_groupi_n_363);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5841(csa_tree_add_83_21_pad_groupi_n_175 ,csa_tree_add_83_21_pad_groupi_n_173);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5842(csa_tree_add_83_21_pad_groupi_n_174 ,csa_tree_add_83_21_pad_groupi_n_173);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5843(csa_tree_add_83_21_pad_groupi_n_173 ,csa_tree_add_83_21_pad_groupi_n_367);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5845(csa_tree_add_83_21_pad_groupi_n_172 ,csa_tree_add_83_21_pad_groupi_n_170);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5846(csa_tree_add_83_21_pad_groupi_n_171 ,csa_tree_add_83_21_pad_groupi_n_170);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5847(csa_tree_add_83_21_pad_groupi_n_170 ,csa_tree_add_83_21_pad_groupi_n_495);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5849(csa_tree_add_83_21_pad_groupi_n_169 ,csa_tree_add_83_21_pad_groupi_n_167);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5850(csa_tree_add_83_21_pad_groupi_n_168 ,csa_tree_add_83_21_pad_groupi_n_167);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5851(csa_tree_add_83_21_pad_groupi_n_167 ,csa_tree_add_83_21_pad_groupi_n_495);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5853(csa_tree_add_83_21_pad_groupi_n_166 ,csa_tree_add_83_21_pad_groupi_n_164);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5854(csa_tree_add_83_21_pad_groupi_n_165 ,csa_tree_add_83_21_pad_groupi_n_164);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5855(csa_tree_add_83_21_pad_groupi_n_164 ,csa_tree_add_83_21_pad_groupi_n_498);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5857(csa_tree_add_83_21_pad_groupi_n_163 ,csa_tree_add_83_21_pad_groupi_n_161);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5858(csa_tree_add_83_21_pad_groupi_n_162 ,csa_tree_add_83_21_pad_groupi_n_161);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5859(csa_tree_add_83_21_pad_groupi_n_161 ,csa_tree_add_83_21_pad_groupi_n_386);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5861(csa_tree_add_83_21_pad_groupi_n_160 ,csa_tree_add_83_21_pad_groupi_n_350);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5863(csa_tree_add_83_21_pad_groupi_n_350 ,csa_tree_add_83_21_pad_groupi_n_412);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5865(csa_tree_add_83_21_pad_groupi_n_159 ,csa_tree_add_83_21_pad_groupi_n_348);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5867(csa_tree_add_83_21_pad_groupi_n_348 ,csa_tree_add_83_21_pad_groupi_n_409);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5869(csa_tree_add_83_21_pad_groupi_n_158 ,csa_tree_add_83_21_pad_groupi_n_356);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5871(csa_tree_add_83_21_pad_groupi_n_356 ,csa_tree_add_83_21_pad_groupi_n_421);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5877(csa_tree_add_83_21_pad_groupi_n_155 ,csa_tree_add_83_21_pad_groupi_n_355);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5879(csa_tree_add_83_21_pad_groupi_n_355 ,csa_tree_add_83_21_pad_groupi_n_421);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5881(csa_tree_add_83_21_pad_groupi_n_154 ,csa_tree_add_83_21_pad_groupi_n_353);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5883(csa_tree_add_83_21_pad_groupi_n_353 ,csa_tree_add_83_21_pad_groupi_n_420);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5885(csa_tree_add_83_21_pad_groupi_n_153 ,csa_tree_add_83_21_pad_groupi_n_349);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5887(csa_tree_add_83_21_pad_groupi_n_349 ,csa_tree_add_83_21_pad_groupi_n_412);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5889(csa_tree_add_83_21_pad_groupi_n_152 ,csa_tree_add_83_21_pad_groupi_n_351);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5891(csa_tree_add_83_21_pad_groupi_n_351 ,csa_tree_add_83_21_pad_groupi_n_417);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5893(csa_tree_add_83_21_pad_groupi_n_151 ,csa_tree_add_83_21_pad_groupi_n_352);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5895(csa_tree_add_83_21_pad_groupi_n_352 ,csa_tree_add_83_21_pad_groupi_n_417);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5897(csa_tree_add_83_21_pad_groupi_n_150 ,csa_tree_add_83_21_pad_groupi_n_347);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5899(csa_tree_add_83_21_pad_groupi_n_347 ,csa_tree_add_83_21_pad_groupi_n_409);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5901(csa_tree_add_83_21_pad_groupi_n_149 ,csa_tree_add_83_21_pad_groupi_n_354);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5903(csa_tree_add_83_21_pad_groupi_n_354 ,csa_tree_add_83_21_pad_groupi_n_420);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5905(csa_tree_add_83_21_pad_groupi_n_148 ,csa_tree_add_83_21_pad_groupi_n_146);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5906(csa_tree_add_83_21_pad_groupi_n_147 ,csa_tree_add_83_21_pad_groupi_n_146);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5907(csa_tree_add_83_21_pad_groupi_n_146 ,csa_tree_add_83_21_pad_groupi_n_504);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5909(csa_tree_add_83_21_pad_groupi_n_145 ,csa_tree_add_83_21_pad_groupi_n_143);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5910(csa_tree_add_83_21_pad_groupi_n_144 ,csa_tree_add_83_21_pad_groupi_n_143);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5911(csa_tree_add_83_21_pad_groupi_n_143 ,csa_tree_add_83_21_pad_groupi_n_510);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5913(csa_tree_add_83_21_pad_groupi_n_142 ,csa_tree_add_83_21_pad_groupi_n_140);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5914(csa_tree_add_83_21_pad_groupi_n_141 ,csa_tree_add_83_21_pad_groupi_n_140);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5915(csa_tree_add_83_21_pad_groupi_n_140 ,csa_tree_add_83_21_pad_groupi_n_510);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5917(csa_tree_add_83_21_pad_groupi_n_139 ,csa_tree_add_83_21_pad_groupi_n_137);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5918(csa_tree_add_83_21_pad_groupi_n_138 ,csa_tree_add_83_21_pad_groupi_n_137);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5919(csa_tree_add_83_21_pad_groupi_n_137 ,csa_tree_add_83_21_pad_groupi_n_494);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5921(csa_tree_add_83_21_pad_groupi_n_136 ,csa_tree_add_83_21_pad_groupi_n_134);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5922(csa_tree_add_83_21_pad_groupi_n_135 ,csa_tree_add_83_21_pad_groupi_n_134);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5923(csa_tree_add_83_21_pad_groupi_n_134 ,csa_tree_add_83_21_pad_groupi_n_494);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5925(csa_tree_add_83_21_pad_groupi_n_133 ,csa_tree_add_83_21_pad_groupi_n_131);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5926(csa_tree_add_83_21_pad_groupi_n_132 ,csa_tree_add_83_21_pad_groupi_n_131);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5927(csa_tree_add_83_21_pad_groupi_n_131 ,csa_tree_add_83_21_pad_groupi_n_504);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5929(csa_tree_add_83_21_pad_groupi_n_130 ,csa_tree_add_83_21_pad_groupi_n_128);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5930(csa_tree_add_83_21_pad_groupi_n_129 ,csa_tree_add_83_21_pad_groupi_n_128);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5931(csa_tree_add_83_21_pad_groupi_n_128 ,csa_tree_add_83_21_pad_groupi_n_498);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5933(csa_tree_add_83_21_pad_groupi_n_127 ,csa_tree_add_83_21_pad_groupi_n_125);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5934(csa_tree_add_83_21_pad_groupi_n_126 ,csa_tree_add_83_21_pad_groupi_n_125);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5935(csa_tree_add_83_21_pad_groupi_n_125 ,csa_tree_add_83_21_pad_groupi_n_496);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5937(csa_tree_add_83_21_pad_groupi_n_124 ,csa_tree_add_83_21_pad_groupi_n_122);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5938(csa_tree_add_83_21_pad_groupi_n_123 ,csa_tree_add_83_21_pad_groupi_n_122);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5939(csa_tree_add_83_21_pad_groupi_n_122 ,csa_tree_add_83_21_pad_groupi_n_496);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5941(csa_tree_add_83_21_pad_groupi_n_121 ,csa_tree_add_83_21_pad_groupi_n_120);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5943(csa_tree_add_83_21_pad_groupi_n_120 ,csa_tree_add_83_21_pad_groupi_n_386);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5945(csa_tree_add_83_21_pad_groupi_n_119 ,csa_tree_add_83_21_pad_groupi_n_117);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5946(csa_tree_add_83_21_pad_groupi_n_118 ,csa_tree_add_83_21_pad_groupi_n_117);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5947(csa_tree_add_83_21_pad_groupi_n_117 ,csa_tree_add_83_21_pad_groupi_n_511);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5949(csa_tree_add_83_21_pad_groupi_n_116 ,csa_tree_add_83_21_pad_groupi_n_114);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5950(csa_tree_add_83_21_pad_groupi_n_115 ,csa_tree_add_83_21_pad_groupi_n_114);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5951(csa_tree_add_83_21_pad_groupi_n_114 ,csa_tree_add_83_21_pad_groupi_n_511);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5953(csa_tree_add_83_21_pad_groupi_n_113 ,csa_tree_add_83_21_pad_groupi_n_111);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5954(csa_tree_add_83_21_pad_groupi_n_112 ,csa_tree_add_83_21_pad_groupi_n_111);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5955(csa_tree_add_83_21_pad_groupi_n_111 ,csa_tree_add_83_21_pad_groupi_n_253);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5957(csa_tree_add_83_21_pad_groupi_n_110 ,csa_tree_add_83_21_pad_groupi_n_108);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5958(csa_tree_add_83_21_pad_groupi_n_109 ,csa_tree_add_83_21_pad_groupi_n_108);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5959(csa_tree_add_83_21_pad_groupi_n_108 ,csa_tree_add_83_21_pad_groupi_n_401);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5961(csa_tree_add_83_21_pad_groupi_n_107 ,csa_tree_add_83_21_pad_groupi_n_105);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5962(csa_tree_add_83_21_pad_groupi_n_106 ,csa_tree_add_83_21_pad_groupi_n_105);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5963(csa_tree_add_83_21_pad_groupi_n_105 ,csa_tree_add_83_21_pad_groupi_n_401);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5965(csa_tree_add_83_21_pad_groupi_n_104 ,csa_tree_add_83_21_pad_groupi_n_102);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5966(csa_tree_add_83_21_pad_groupi_n_103 ,csa_tree_add_83_21_pad_groupi_n_102);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5967(csa_tree_add_83_21_pad_groupi_n_102 ,csa_tree_add_83_21_pad_groupi_n_250);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5969(csa_tree_add_83_21_pad_groupi_n_101 ,csa_tree_add_83_21_pad_groupi_n_99);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5970(csa_tree_add_83_21_pad_groupi_n_100 ,csa_tree_add_83_21_pad_groupi_n_99);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5971(csa_tree_add_83_21_pad_groupi_n_99 ,csa_tree_add_83_21_pad_groupi_n_385);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5973(csa_tree_add_83_21_pad_groupi_n_98 ,csa_tree_add_83_21_pad_groupi_n_97);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5975(csa_tree_add_83_21_pad_groupi_n_97 ,csa_tree_add_83_21_pad_groupi_n_247);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5977(csa_tree_add_83_21_pad_groupi_n_96 ,csa_tree_add_83_21_pad_groupi_n_94);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5978(csa_tree_add_83_21_pad_groupi_n_95 ,csa_tree_add_83_21_pad_groupi_n_94);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5979(csa_tree_add_83_21_pad_groupi_n_94 ,csa_tree_add_83_21_pad_groupi_n_381);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5981(csa_tree_add_83_21_pad_groupi_n_93 ,csa_tree_add_83_21_pad_groupi_n_92);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5983(csa_tree_add_83_21_pad_groupi_n_92 ,csa_tree_add_83_21_pad_groupi_n_252);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5985(csa_tree_add_83_21_pad_groupi_n_91 ,csa_tree_add_83_21_pad_groupi_n_89);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5986(csa_tree_add_83_21_pad_groupi_n_90 ,csa_tree_add_83_21_pad_groupi_n_89);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5987(csa_tree_add_83_21_pad_groupi_n_89 ,csa_tree_add_83_21_pad_groupi_n_366);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5989(csa_tree_add_83_21_pad_groupi_n_88 ,csa_tree_add_83_21_pad_groupi_n_86);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5990(csa_tree_add_83_21_pad_groupi_n_87 ,csa_tree_add_83_21_pad_groupi_n_86);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5991(csa_tree_add_83_21_pad_groupi_n_86 ,csa_tree_add_83_21_pad_groupi_n_382);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5993(csa_tree_add_83_21_pad_groupi_n_85 ,csa_tree_add_83_21_pad_groupi_n_83);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5994(csa_tree_add_83_21_pad_groupi_n_84 ,csa_tree_add_83_21_pad_groupi_n_83);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5995(csa_tree_add_83_21_pad_groupi_n_83 ,csa_tree_add_83_21_pad_groupi_n_383);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5997(csa_tree_add_83_21_pad_groupi_n_82 ,csa_tree_add_83_21_pad_groupi_n_80);
  not csa_tree_add_83_21_pad_groupi_drc_bufs5999(csa_tree_add_83_21_pad_groupi_n_80 ,csa_tree_add_83_21_pad_groupi_n_365);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6001(csa_tree_add_83_21_pad_groupi_n_79 ,csa_tree_add_83_21_pad_groupi_n_77);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6002(csa_tree_add_83_21_pad_groupi_n_78 ,csa_tree_add_83_21_pad_groupi_n_77);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6003(csa_tree_add_83_21_pad_groupi_n_77 ,csa_tree_add_83_21_pad_groupi_n_363);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6005(csa_tree_add_83_21_pad_groupi_n_76 ,csa_tree_add_83_21_pad_groupi_n_75);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6007(csa_tree_add_83_21_pad_groupi_n_75 ,csa_tree_add_83_21_pad_groupi_n_215);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6009(csa_tree_add_83_21_pad_groupi_n_74 ,csa_tree_add_83_21_pad_groupi_n_72);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6010(csa_tree_add_83_21_pad_groupi_n_73 ,csa_tree_add_83_21_pad_groupi_n_72);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6011(csa_tree_add_83_21_pad_groupi_n_72 ,csa_tree_add_83_21_pad_groupi_n_385);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6013(csa_tree_add_83_21_pad_groupi_n_71 ,csa_tree_add_83_21_pad_groupi_n_70);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6015(csa_tree_add_83_21_pad_groupi_n_70 ,csa_tree_add_83_21_pad_groupi_n_218);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6017(csa_tree_add_83_21_pad_groupi_n_69 ,csa_tree_add_83_21_pad_groupi_n_68);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6019(csa_tree_add_83_21_pad_groupi_n_68 ,csa_tree_add_83_21_pad_groupi_n_223);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6021(csa_tree_add_83_21_pad_groupi_n_67 ,csa_tree_add_83_21_pad_groupi_n_65);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6022(csa_tree_add_83_21_pad_groupi_n_66 ,csa_tree_add_83_21_pad_groupi_n_65);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6023(csa_tree_add_83_21_pad_groupi_n_65 ,csa_tree_add_83_21_pad_groupi_n_362);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6025(csa_tree_add_83_21_pad_groupi_n_64 ,csa_tree_add_83_21_pad_groupi_n_62);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6027(csa_tree_add_83_21_pad_groupi_n_62 ,csa_tree_add_83_21_pad_groupi_n_380);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6029(csa_tree_add_83_21_pad_groupi_n_61 ,csa_tree_add_83_21_pad_groupi_n_60);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6031(csa_tree_add_83_21_pad_groupi_n_60 ,csa_tree_add_83_21_pad_groupi_n_249);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6033(csa_tree_add_83_21_pad_groupi_n_59 ,csa_tree_add_83_21_pad_groupi_n_58);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6035(csa_tree_add_83_21_pad_groupi_n_58 ,csa_tree_add_83_21_pad_groupi_n_212);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6037(csa_tree_add_83_21_pad_groupi_n_57 ,csa_tree_add_83_21_pad_groupi_n_56);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6039(csa_tree_add_83_21_pad_groupi_n_56 ,csa_tree_add_83_21_pad_groupi_n_244);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6041(csa_tree_add_83_21_pad_groupi_n_55 ,csa_tree_add_83_21_pad_groupi_n_54);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6043(csa_tree_add_83_21_pad_groupi_n_54 ,csa_tree_add_83_21_pad_groupi_n_207);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6045(csa_tree_add_83_21_pad_groupi_n_53 ,csa_tree_add_83_21_pad_groupi_n_51);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6046(csa_tree_add_83_21_pad_groupi_n_52 ,csa_tree_add_83_21_pad_groupi_n_51);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6047(csa_tree_add_83_21_pad_groupi_n_51 ,csa_tree_add_83_21_pad_groupi_n_384);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6049(csa_tree_add_83_21_pad_groupi_n_50 ,csa_tree_add_83_21_pad_groupi_n_48);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6051(csa_tree_add_83_21_pad_groupi_n_48 ,csa_tree_add_83_21_pad_groupi_n_379);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6053(csa_tree_add_83_21_pad_groupi_n_47 ,csa_tree_add_83_21_pad_groupi_n_46);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6055(csa_tree_add_83_21_pad_groupi_n_46 ,csa_tree_add_83_21_pad_groupi_n_246);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6057(csa_tree_add_83_21_pad_groupi_n_45 ,csa_tree_add_83_21_pad_groupi_n_43);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6059(csa_tree_add_83_21_pad_groupi_n_43 ,csa_tree_add_83_21_pad_groupi_n_380);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6061(csa_tree_add_83_21_pad_groupi_n_42 ,csa_tree_add_83_21_pad_groupi_n_40);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6062(csa_tree_add_83_21_pad_groupi_n_41 ,csa_tree_add_83_21_pad_groupi_n_40);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6063(csa_tree_add_83_21_pad_groupi_n_40 ,csa_tree_add_83_21_pad_groupi_n_368);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6065(csa_tree_add_83_21_pad_groupi_n_39 ,csa_tree_add_83_21_pad_groupi_n_37);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6066(csa_tree_add_83_21_pad_groupi_n_38 ,csa_tree_add_83_21_pad_groupi_n_37);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6067(csa_tree_add_83_21_pad_groupi_n_37 ,csa_tree_add_83_21_pad_groupi_n_361);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6069(csa_tree_add_83_21_pad_groupi_n_36 ,csa_tree_add_83_21_pad_groupi_n_35);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6071(csa_tree_add_83_21_pad_groupi_n_35 ,csa_tree_add_83_21_pad_groupi_n_202);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6073(csa_tree_add_83_21_pad_groupi_n_34 ,csa_tree_add_83_21_pad_groupi_n_33);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6075(csa_tree_add_83_21_pad_groupi_n_33 ,csa_tree_add_83_21_pad_groupi_n_238);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6077(csa_tree_add_83_21_pad_groupi_n_32 ,csa_tree_add_83_21_pad_groupi_n_31);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6079(csa_tree_add_83_21_pad_groupi_n_31 ,csa_tree_add_83_21_pad_groupi_n_241);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6082(csa_tree_add_83_21_pad_groupi_n_30 ,csa_tree_add_83_21_pad_groupi_n_29);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6083(csa_tree_add_83_21_pad_groupi_n_29 ,csa_tree_add_83_21_pad_groupi_n_193);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6085(csa_tree_add_83_21_pad_groupi_n_28 ,csa_tree_add_83_21_pad_groupi_n_26);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6086(csa_tree_add_83_21_pad_groupi_n_27 ,csa_tree_add_83_21_pad_groupi_n_26);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6087(csa_tree_add_83_21_pad_groupi_n_26 ,csa_tree_add_83_21_pad_groupi_n_367);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6089(csa_tree_add_83_21_pad_groupi_n_25 ,csa_tree_add_83_21_pad_groupi_n_23);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6090(csa_tree_add_83_21_pad_groupi_n_24 ,csa_tree_add_83_21_pad_groupi_n_23);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6091(csa_tree_add_83_21_pad_groupi_n_23 ,csa_tree_add_83_21_pad_groupi_n_368);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6093(csa_tree_add_83_21_pad_groupi_n_22 ,csa_tree_add_83_21_pad_groupi_n_20);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6094(csa_tree_add_83_21_pad_groupi_n_21 ,csa_tree_add_83_21_pad_groupi_n_20);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6095(csa_tree_add_83_21_pad_groupi_n_20 ,csa_tree_add_83_21_pad_groupi_n_364);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6098(csa_tree_add_83_21_pad_groupi_n_19 ,csa_tree_add_83_21_pad_groupi_n_18);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6099(csa_tree_add_83_21_pad_groupi_n_18 ,csa_tree_add_83_21_pad_groupi_n_243);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6102(csa_tree_add_83_21_pad_groupi_n_17 ,csa_tree_add_83_21_pad_groupi_n_16);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6103(csa_tree_add_83_21_pad_groupi_n_16 ,csa_tree_add_83_21_pad_groupi_n_196);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6106(csa_tree_add_83_21_pad_groupi_n_15 ,csa_tree_add_83_21_pad_groupi_n_14);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6107(csa_tree_add_83_21_pad_groupi_n_14 ,csa_tree_add_83_21_pad_groupi_n_237);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6110(csa_tree_add_83_21_pad_groupi_n_13 ,csa_tree_add_83_21_pad_groupi_n_12);
  not csa_tree_add_83_21_pad_groupi_drc_bufs6111(csa_tree_add_83_21_pad_groupi_n_12 ,csa_tree_add_83_21_pad_groupi_n_240);
  xor csa_tree_add_83_21_pad_groupi_g2(n_199 ,csa_tree_add_83_21_pad_groupi_n_1537 ,csa_tree_add_83_21_pad_groupi_n_1520);
  xor csa_tree_add_83_21_pad_groupi_g6113(n_197 ,csa_tree_add_83_21_pad_groupi_n_1532 ,csa_tree_add_83_21_pad_groupi_n_1518);
  xor csa_tree_add_83_21_pad_groupi_g6114(n_194 ,csa_tree_add_83_21_pad_groupi_n_1524 ,csa_tree_add_83_21_pad_groupi_n_1482);
  xor csa_tree_add_83_21_pad_groupi_g6115(n_193 ,csa_tree_add_83_21_pad_groupi_n_1522 ,csa_tree_add_83_21_pad_groupi_n_1502);
  xor csa_tree_add_83_21_pad_groupi_g6116(n_192 ,csa_tree_add_83_21_pad_groupi_n_1515 ,csa_tree_add_83_21_pad_groupi_n_1461);
  xor csa_tree_add_83_21_pad_groupi_g6117(csa_tree_add_83_21_pad_groupi_n_6 ,csa_tree_add_83_21_pad_groupi_n_1368 ,csa_tree_add_83_21_pad_groupi_n_1406);
  xor csa_tree_add_83_21_pad_groupi_g6118(csa_tree_add_83_21_pad_groupi_n_5 ,csa_tree_add_83_21_pad_groupi_n_1332 ,csa_tree_add_83_21_pad_groupi_n_1350);
  xor csa_tree_add_83_21_pad_groupi_g6119(csa_tree_add_83_21_pad_groupi_n_4 ,csa_tree_add_83_21_pad_groupi_n_836 ,csa_tree_add_83_21_pad_groupi_n_0);
  xor csa_tree_add_83_21_pad_groupi_g6120(csa_tree_add_83_21_pad_groupi_n_3 ,csa_tree_add_83_21_pad_groupi_n_835 ,csa_tree_add_83_21_pad_groupi_n_948);
  xor csa_tree_add_83_21_pad_groupi_g6122(csa_tree_add_83_21_pad_groupi_n_1 ,csa_tree_add_83_21_pad_groupi_n_358 ,in8[9]);
  xor csa_tree_add_83_21_pad_groupi_g6123(csa_tree_add_83_21_pad_groupi_n_0 ,csa_tree_add_83_21_pad_groupi_n_357 ,in8[11]);
  xnor csa_tree_add_89_22_pad_groupi_g4151(n_174 ,csa_tree_add_89_22_pad_groupi_n_1336 ,csa_tree_add_89_22_pad_groupi_n_1558);
  or csa_tree_add_89_22_pad_groupi_g4152(csa_tree_add_89_22_pad_groupi_n_1558 ,csa_tree_add_89_22_pad_groupi_n_1393 ,csa_tree_add_89_22_pad_groupi_n_1556);
  xnor csa_tree_add_89_22_pad_groupi_g4153(n_173 ,csa_tree_add_89_22_pad_groupi_n_1555 ,csa_tree_add_89_22_pad_groupi_n_1404);
  and csa_tree_add_89_22_pad_groupi_g4154(csa_tree_add_89_22_pad_groupi_n_1556 ,csa_tree_add_89_22_pad_groupi_n_1389 ,csa_tree_add_89_22_pad_groupi_n_1555);
  or csa_tree_add_89_22_pad_groupi_g4155(csa_tree_add_89_22_pad_groupi_n_1555 ,csa_tree_add_89_22_pad_groupi_n_1407 ,csa_tree_add_89_22_pad_groupi_n_1553);
  xnor csa_tree_add_89_22_pad_groupi_g4156(n_172 ,csa_tree_add_89_22_pad_groupi_n_1552 ,csa_tree_add_89_22_pad_groupi_n_1434);
  and csa_tree_add_89_22_pad_groupi_g4157(csa_tree_add_89_22_pad_groupi_n_1553 ,csa_tree_add_89_22_pad_groupi_n_1410 ,csa_tree_add_89_22_pad_groupi_n_1552);
  or csa_tree_add_89_22_pad_groupi_g4158(csa_tree_add_89_22_pad_groupi_n_1552 ,csa_tree_add_89_22_pad_groupi_n_1453 ,csa_tree_add_89_22_pad_groupi_n_1550);
  xnor csa_tree_add_89_22_pad_groupi_g4159(n_171 ,csa_tree_add_89_22_pad_groupi_n_1549 ,csa_tree_add_89_22_pad_groupi_n_1462);
  and csa_tree_add_89_22_pad_groupi_g4160(csa_tree_add_89_22_pad_groupi_n_1550 ,csa_tree_add_89_22_pad_groupi_n_1459 ,csa_tree_add_89_22_pad_groupi_n_1549);
  or csa_tree_add_89_22_pad_groupi_g4161(csa_tree_add_89_22_pad_groupi_n_1549 ,csa_tree_add_89_22_pad_groupi_n_1463 ,csa_tree_add_89_22_pad_groupi_n_1547);
  xnor csa_tree_add_89_22_pad_groupi_g4162(n_170 ,csa_tree_add_89_22_pad_groupi_n_1546 ,csa_tree_add_89_22_pad_groupi_n_1483);
  nor csa_tree_add_89_22_pad_groupi_g4163(csa_tree_add_89_22_pad_groupi_n_1547 ,csa_tree_add_89_22_pad_groupi_n_1546 ,csa_tree_add_89_22_pad_groupi_n_1464);
  and csa_tree_add_89_22_pad_groupi_g4164(csa_tree_add_89_22_pad_groupi_n_1546 ,csa_tree_add_89_22_pad_groupi_n_1500 ,csa_tree_add_89_22_pad_groupi_n_1544);
  xnor csa_tree_add_89_22_pad_groupi_g4165(n_169 ,csa_tree_add_89_22_pad_groupi_n_1542 ,csa_tree_add_89_22_pad_groupi_n_1501);
  or csa_tree_add_89_22_pad_groupi_g4166(csa_tree_add_89_22_pad_groupi_n_1544 ,csa_tree_add_89_22_pad_groupi_n_1494 ,csa_tree_add_89_22_pad_groupi_n_1543);
  not csa_tree_add_89_22_pad_groupi_g4167(csa_tree_add_89_22_pad_groupi_n_1543 ,csa_tree_add_89_22_pad_groupi_n_1542);
  or csa_tree_add_89_22_pad_groupi_g4168(csa_tree_add_89_22_pad_groupi_n_1542 ,csa_tree_add_89_22_pad_groupi_n_1499 ,csa_tree_add_89_22_pad_groupi_n_1540);
  xnor csa_tree_add_89_22_pad_groupi_g4169(n_168 ,csa_tree_add_89_22_pad_groupi_n_1539 ,csa_tree_add_89_22_pad_groupi_n_1503);
  nor csa_tree_add_89_22_pad_groupi_g4170(csa_tree_add_89_22_pad_groupi_n_1540 ,csa_tree_add_89_22_pad_groupi_n_1496 ,csa_tree_add_89_22_pad_groupi_n_1539);
  and csa_tree_add_89_22_pad_groupi_g4171(csa_tree_add_89_22_pad_groupi_n_1539 ,csa_tree_add_89_22_pad_groupi_n_1538 ,csa_tree_add_89_22_pad_groupi_n_1510);
  or csa_tree_add_89_22_pad_groupi_g4173(csa_tree_add_89_22_pad_groupi_n_1538 ,csa_tree_add_89_22_pad_groupi_n_1513 ,csa_tree_add_89_22_pad_groupi_n_1537);
  and csa_tree_add_89_22_pad_groupi_g4175(csa_tree_add_89_22_pad_groupi_n_1537 ,csa_tree_add_89_22_pad_groupi_n_1512 ,csa_tree_add_89_22_pad_groupi_n_1535);
  xnor csa_tree_add_89_22_pad_groupi_g4176(n_166 ,csa_tree_add_89_22_pad_groupi_n_1534 ,csa_tree_add_89_22_pad_groupi_n_1519);
  or csa_tree_add_89_22_pad_groupi_g4177(csa_tree_add_89_22_pad_groupi_n_1535 ,csa_tree_add_89_22_pad_groupi_n_1514 ,csa_tree_add_89_22_pad_groupi_n_1534);
  and csa_tree_add_89_22_pad_groupi_g4178(csa_tree_add_89_22_pad_groupi_n_1534 ,csa_tree_add_89_22_pad_groupi_n_1533 ,csa_tree_add_89_22_pad_groupi_n_1511);
  or csa_tree_add_89_22_pad_groupi_g4180(csa_tree_add_89_22_pad_groupi_n_1533 ,csa_tree_add_89_22_pad_groupi_n_1505 ,csa_tree_add_89_22_pad_groupi_n_1532);
  and csa_tree_add_89_22_pad_groupi_g4182(csa_tree_add_89_22_pad_groupi_n_1532 ,csa_tree_add_89_22_pad_groupi_n_1506 ,csa_tree_add_89_22_pad_groupi_n_1530);
  xnor csa_tree_add_89_22_pad_groupi_g4183(n_164 ,csa_tree_add_89_22_pad_groupi_n_1529 ,csa_tree_add_89_22_pad_groupi_n_1517);
  or csa_tree_add_89_22_pad_groupi_g4184(csa_tree_add_89_22_pad_groupi_n_1530 ,csa_tree_add_89_22_pad_groupi_n_1507 ,csa_tree_add_89_22_pad_groupi_n_1529);
  and csa_tree_add_89_22_pad_groupi_g4185(csa_tree_add_89_22_pad_groupi_n_1529 ,csa_tree_add_89_22_pad_groupi_n_1508 ,csa_tree_add_89_22_pad_groupi_n_1527);
  xnor csa_tree_add_89_22_pad_groupi_g4186(n_163 ,csa_tree_add_89_22_pad_groupi_n_1526 ,csa_tree_add_89_22_pad_groupi_n_1516);
  or csa_tree_add_89_22_pad_groupi_g4187(csa_tree_add_89_22_pad_groupi_n_1527 ,csa_tree_add_89_22_pad_groupi_n_1526 ,csa_tree_add_89_22_pad_groupi_n_1509);
  and csa_tree_add_89_22_pad_groupi_g4188(csa_tree_add_89_22_pad_groupi_n_1526 ,csa_tree_add_89_22_pad_groupi_n_1471 ,csa_tree_add_89_22_pad_groupi_n_1525);
  or csa_tree_add_89_22_pad_groupi_g4190(csa_tree_add_89_22_pad_groupi_n_1525 ,csa_tree_add_89_22_pad_groupi_n_1470 ,csa_tree_add_89_22_pad_groupi_n_1524);
  and csa_tree_add_89_22_pad_groupi_g4192(csa_tree_add_89_22_pad_groupi_n_1524 ,csa_tree_add_89_22_pad_groupi_n_1498 ,csa_tree_add_89_22_pad_groupi_n_1523);
  or csa_tree_add_89_22_pad_groupi_g4194(csa_tree_add_89_22_pad_groupi_n_1523 ,csa_tree_add_89_22_pad_groupi_n_1497 ,csa_tree_add_89_22_pad_groupi_n_1522);
  and csa_tree_add_89_22_pad_groupi_g4196(csa_tree_add_89_22_pad_groupi_n_1522 ,csa_tree_add_89_22_pad_groupi_n_1452 ,csa_tree_add_89_22_pad_groupi_n_1521);
  or csa_tree_add_89_22_pad_groupi_g4198(csa_tree_add_89_22_pad_groupi_n_1521 ,csa_tree_add_89_22_pad_groupi_n_1451 ,csa_tree_add_89_22_pad_groupi_n_1515);
  xnor csa_tree_add_89_22_pad_groupi_g4199(csa_tree_add_89_22_pad_groupi_n_1520 ,csa_tree_add_89_22_pad_groupi_n_1475 ,csa_tree_add_89_22_pad_groupi_n_1491);
  xnor csa_tree_add_89_22_pad_groupi_g4200(csa_tree_add_89_22_pad_groupi_n_1519 ,csa_tree_add_89_22_pad_groupi_n_1473 ,csa_tree_add_89_22_pad_groupi_n_1489);
  xnor csa_tree_add_89_22_pad_groupi_g4201(csa_tree_add_89_22_pad_groupi_n_1518 ,csa_tree_add_89_22_pad_groupi_n_1480 ,csa_tree_add_89_22_pad_groupi_n_1487);
  xnor csa_tree_add_89_22_pad_groupi_g4202(csa_tree_add_89_22_pad_groupi_n_1517 ,csa_tree_add_89_22_pad_groupi_n_1477 ,csa_tree_add_89_22_pad_groupi_n_1493);
  xnor csa_tree_add_89_22_pad_groupi_g4203(csa_tree_add_89_22_pad_groupi_n_1516 ,csa_tree_add_89_22_pad_groupi_n_1448 ,csa_tree_add_89_22_pad_groupi_n_1485);
  nor csa_tree_add_89_22_pad_groupi_g4205(csa_tree_add_89_22_pad_groupi_n_1514 ,csa_tree_add_89_22_pad_groupi_n_1472 ,csa_tree_add_89_22_pad_groupi_n_1489);
  nor csa_tree_add_89_22_pad_groupi_g4206(csa_tree_add_89_22_pad_groupi_n_1513 ,csa_tree_add_89_22_pad_groupi_n_1475 ,csa_tree_add_89_22_pad_groupi_n_1491);
  or csa_tree_add_89_22_pad_groupi_g4207(csa_tree_add_89_22_pad_groupi_n_1512 ,csa_tree_add_89_22_pad_groupi_n_1473 ,csa_tree_add_89_22_pad_groupi_n_1488);
  or csa_tree_add_89_22_pad_groupi_g4208(csa_tree_add_89_22_pad_groupi_n_1511 ,csa_tree_add_89_22_pad_groupi_n_1479 ,csa_tree_add_89_22_pad_groupi_n_1486);
  or csa_tree_add_89_22_pad_groupi_g4209(csa_tree_add_89_22_pad_groupi_n_1510 ,csa_tree_add_89_22_pad_groupi_n_1474 ,csa_tree_add_89_22_pad_groupi_n_1490);
  nor csa_tree_add_89_22_pad_groupi_g4210(csa_tree_add_89_22_pad_groupi_n_1509 ,csa_tree_add_89_22_pad_groupi_n_1447 ,csa_tree_add_89_22_pad_groupi_n_1485);
  and csa_tree_add_89_22_pad_groupi_g4211(csa_tree_add_89_22_pad_groupi_n_1515 ,csa_tree_add_89_22_pad_groupi_n_1450 ,csa_tree_add_89_22_pad_groupi_n_1495);
  or csa_tree_add_89_22_pad_groupi_g4212(csa_tree_add_89_22_pad_groupi_n_1508 ,csa_tree_add_89_22_pad_groupi_n_1448 ,csa_tree_add_89_22_pad_groupi_n_1484);
  nor csa_tree_add_89_22_pad_groupi_g4213(csa_tree_add_89_22_pad_groupi_n_1507 ,csa_tree_add_89_22_pad_groupi_n_1476 ,csa_tree_add_89_22_pad_groupi_n_1493);
  or csa_tree_add_89_22_pad_groupi_g4214(csa_tree_add_89_22_pad_groupi_n_1506 ,csa_tree_add_89_22_pad_groupi_n_1477 ,csa_tree_add_89_22_pad_groupi_n_1492);
  nor csa_tree_add_89_22_pad_groupi_g4215(csa_tree_add_89_22_pad_groupi_n_1505 ,csa_tree_add_89_22_pad_groupi_n_1480 ,csa_tree_add_89_22_pad_groupi_n_1487);
  xnor csa_tree_add_89_22_pad_groupi_g4216(n_159 ,csa_tree_add_89_22_pad_groupi_n_1481 ,csa_tree_add_89_22_pad_groupi_n_1460);
  xnor csa_tree_add_89_22_pad_groupi_g4217(csa_tree_add_89_22_pad_groupi_n_1503 ,csa_tree_add_89_22_pad_groupi_n_1478 ,csa_tree_add_89_22_pad_groupi_n_1467);
  xnor csa_tree_add_89_22_pad_groupi_g4218(csa_tree_add_89_22_pad_groupi_n_1502 ,csa_tree_add_89_22_pad_groupi_n_1412 ,csa_tree_add_89_22_pad_groupi_n_1466);
  xnor csa_tree_add_89_22_pad_groupi_g4219(csa_tree_add_89_22_pad_groupi_n_1501 ,csa_tree_add_89_22_pad_groupi_n_1442 ,csa_tree_add_89_22_pad_groupi_n_1469);
  or csa_tree_add_89_22_pad_groupi_g4220(csa_tree_add_89_22_pad_groupi_n_1500 ,csa_tree_add_89_22_pad_groupi_n_1441 ,csa_tree_add_89_22_pad_groupi_n_6);
  nor csa_tree_add_89_22_pad_groupi_g4221(csa_tree_add_89_22_pad_groupi_n_1499 ,csa_tree_add_89_22_pad_groupi_n_1478 ,csa_tree_add_89_22_pad_groupi_n_1468);
  or csa_tree_add_89_22_pad_groupi_g4222(csa_tree_add_89_22_pad_groupi_n_1498 ,csa_tree_add_89_22_pad_groupi_n_1411 ,csa_tree_add_89_22_pad_groupi_n_1465);
  nor csa_tree_add_89_22_pad_groupi_g4223(csa_tree_add_89_22_pad_groupi_n_1497 ,csa_tree_add_89_22_pad_groupi_n_1412 ,csa_tree_add_89_22_pad_groupi_n_1466);
  and csa_tree_add_89_22_pad_groupi_g4224(csa_tree_add_89_22_pad_groupi_n_1496 ,csa_tree_add_89_22_pad_groupi_n_1478 ,csa_tree_add_89_22_pad_groupi_n_1468);
  or csa_tree_add_89_22_pad_groupi_g4225(csa_tree_add_89_22_pad_groupi_n_1495 ,csa_tree_add_89_22_pad_groupi_n_1449 ,csa_tree_add_89_22_pad_groupi_n_1481);
  nor csa_tree_add_89_22_pad_groupi_g4226(csa_tree_add_89_22_pad_groupi_n_1494 ,csa_tree_add_89_22_pad_groupi_n_1442 ,csa_tree_add_89_22_pad_groupi_n_1469);
  not csa_tree_add_89_22_pad_groupi_g4227(csa_tree_add_89_22_pad_groupi_n_1493 ,csa_tree_add_89_22_pad_groupi_n_1492);
  not csa_tree_add_89_22_pad_groupi_g4228(csa_tree_add_89_22_pad_groupi_n_1491 ,csa_tree_add_89_22_pad_groupi_n_1490);
  not csa_tree_add_89_22_pad_groupi_g4229(csa_tree_add_89_22_pad_groupi_n_1489 ,csa_tree_add_89_22_pad_groupi_n_1488);
  not csa_tree_add_89_22_pad_groupi_g4230(csa_tree_add_89_22_pad_groupi_n_1487 ,csa_tree_add_89_22_pad_groupi_n_1486);
  not csa_tree_add_89_22_pad_groupi_g4231(csa_tree_add_89_22_pad_groupi_n_1485 ,csa_tree_add_89_22_pad_groupi_n_1484);
  xnor csa_tree_add_89_22_pad_groupi_g4232(csa_tree_add_89_22_pad_groupi_n_1483 ,csa_tree_add_89_22_pad_groupi_n_1440 ,csa_tree_add_89_22_pad_groupi_n_1445);
  xnor csa_tree_add_89_22_pad_groupi_g4233(csa_tree_add_89_22_pad_groupi_n_1482 ,csa_tree_add_89_22_pad_groupi_n_1419 ,csa_tree_add_89_22_pad_groupi_n_1444);
  xnor csa_tree_add_89_22_pad_groupi_g4234(csa_tree_add_89_22_pad_groupi_n_1492 ,csa_tree_add_89_22_pad_groupi_n_1387 ,csa_tree_add_89_22_pad_groupi_n_1438);
  xnor csa_tree_add_89_22_pad_groupi_g4235(csa_tree_add_89_22_pad_groupi_n_1490 ,csa_tree_add_89_22_pad_groupi_n_1400 ,csa_tree_add_89_22_pad_groupi_n_1433);
  xnor csa_tree_add_89_22_pad_groupi_g4236(csa_tree_add_89_22_pad_groupi_n_1488 ,csa_tree_add_89_22_pad_groupi_n_1401 ,csa_tree_add_89_22_pad_groupi_n_1436);
  xnor csa_tree_add_89_22_pad_groupi_g4237(csa_tree_add_89_22_pad_groupi_n_1486 ,csa_tree_add_89_22_pad_groupi_n_1402 ,csa_tree_add_89_22_pad_groupi_n_1437);
  xnor csa_tree_add_89_22_pad_groupi_g4238(csa_tree_add_89_22_pad_groupi_n_1484 ,csa_tree_add_89_22_pad_groupi_n_1403 ,csa_tree_add_89_22_pad_groupi_n_1435);
  not csa_tree_add_89_22_pad_groupi_g4239(csa_tree_add_89_22_pad_groupi_n_1479 ,csa_tree_add_89_22_pad_groupi_n_1480);
  not csa_tree_add_89_22_pad_groupi_g4240(csa_tree_add_89_22_pad_groupi_n_1477 ,csa_tree_add_89_22_pad_groupi_n_1476);
  not csa_tree_add_89_22_pad_groupi_g4241(csa_tree_add_89_22_pad_groupi_n_1474 ,csa_tree_add_89_22_pad_groupi_n_1475);
  not csa_tree_add_89_22_pad_groupi_g4242(csa_tree_add_89_22_pad_groupi_n_1473 ,csa_tree_add_89_22_pad_groupi_n_1472);
  or csa_tree_add_89_22_pad_groupi_g4243(csa_tree_add_89_22_pad_groupi_n_1471 ,csa_tree_add_89_22_pad_groupi_n_1418 ,csa_tree_add_89_22_pad_groupi_n_1443);
  nor csa_tree_add_89_22_pad_groupi_g4244(csa_tree_add_89_22_pad_groupi_n_1470 ,csa_tree_add_89_22_pad_groupi_n_1419 ,csa_tree_add_89_22_pad_groupi_n_1444);
  and csa_tree_add_89_22_pad_groupi_g4245(csa_tree_add_89_22_pad_groupi_n_1481 ,csa_tree_add_89_22_pad_groupi_n_1371 ,csa_tree_add_89_22_pad_groupi_n_1439);
  or csa_tree_add_89_22_pad_groupi_g4246(csa_tree_add_89_22_pad_groupi_n_1480 ,csa_tree_add_89_22_pad_groupi_n_1424 ,csa_tree_add_89_22_pad_groupi_n_1456);
  and csa_tree_add_89_22_pad_groupi_g4247(csa_tree_add_89_22_pad_groupi_n_1478 ,csa_tree_add_89_22_pad_groupi_n_1431 ,csa_tree_add_89_22_pad_groupi_n_1454);
  or csa_tree_add_89_22_pad_groupi_g4248(csa_tree_add_89_22_pad_groupi_n_1476 ,csa_tree_add_89_22_pad_groupi_n_1422 ,csa_tree_add_89_22_pad_groupi_n_1455);
  or csa_tree_add_89_22_pad_groupi_g4249(csa_tree_add_89_22_pad_groupi_n_1475 ,csa_tree_add_89_22_pad_groupi_n_1429 ,csa_tree_add_89_22_pad_groupi_n_1458);
  or csa_tree_add_89_22_pad_groupi_g4250(csa_tree_add_89_22_pad_groupi_n_1472 ,csa_tree_add_89_22_pad_groupi_n_1426 ,csa_tree_add_89_22_pad_groupi_n_1457);
  not csa_tree_add_89_22_pad_groupi_g4251(csa_tree_add_89_22_pad_groupi_n_1469 ,csa_tree_add_89_22_pad_groupi_n_6);
  not csa_tree_add_89_22_pad_groupi_g4252(csa_tree_add_89_22_pad_groupi_n_1468 ,csa_tree_add_89_22_pad_groupi_n_1467);
  not csa_tree_add_89_22_pad_groupi_g4253(csa_tree_add_89_22_pad_groupi_n_1466 ,csa_tree_add_89_22_pad_groupi_n_1465);
  and csa_tree_add_89_22_pad_groupi_g4254(csa_tree_add_89_22_pad_groupi_n_1464 ,csa_tree_add_89_22_pad_groupi_n_1440 ,csa_tree_add_89_22_pad_groupi_n_1446);
  nor csa_tree_add_89_22_pad_groupi_g4255(csa_tree_add_89_22_pad_groupi_n_1463 ,csa_tree_add_89_22_pad_groupi_n_1440 ,csa_tree_add_89_22_pad_groupi_n_1446);
  xnor csa_tree_add_89_22_pad_groupi_g4256(csa_tree_add_89_22_pad_groupi_n_1462 ,csa_tree_add_89_22_pad_groupi_n_1432 ,csa_tree_add_89_22_pad_groupi_n_1413);
  xnor csa_tree_add_89_22_pad_groupi_g4257(csa_tree_add_89_22_pad_groupi_n_1461 ,csa_tree_add_89_22_pad_groupi_n_1397 ,csa_tree_add_89_22_pad_groupi_n_1417);
  xnor csa_tree_add_89_22_pad_groupi_g4258(csa_tree_add_89_22_pad_groupi_n_1460 ,csa_tree_add_89_22_pad_groupi_n_1367 ,csa_tree_add_89_22_pad_groupi_n_1415);
  xnor csa_tree_add_89_22_pad_groupi_g4260(csa_tree_add_89_22_pad_groupi_n_1467 ,csa_tree_add_89_22_pad_groupi_n_1384 ,csa_tree_add_89_22_pad_groupi_n_1405);
  xnor csa_tree_add_89_22_pad_groupi_g4261(csa_tree_add_89_22_pad_groupi_n_1465 ,csa_tree_add_89_22_pad_groupi_n_1295 ,csa_tree_add_89_22_pad_groupi_n_5);
  or csa_tree_add_89_22_pad_groupi_g4262(csa_tree_add_89_22_pad_groupi_n_1459 ,csa_tree_add_89_22_pad_groupi_n_1432 ,csa_tree_add_89_22_pad_groupi_n_1413);
  and csa_tree_add_89_22_pad_groupi_g4263(csa_tree_add_89_22_pad_groupi_n_1458 ,csa_tree_add_89_22_pad_groupi_n_1401 ,csa_tree_add_89_22_pad_groupi_n_1427);
  and csa_tree_add_89_22_pad_groupi_g4264(csa_tree_add_89_22_pad_groupi_n_1457 ,csa_tree_add_89_22_pad_groupi_n_1402 ,csa_tree_add_89_22_pad_groupi_n_1425);
  and csa_tree_add_89_22_pad_groupi_g4265(csa_tree_add_89_22_pad_groupi_n_1456 ,csa_tree_add_89_22_pad_groupi_n_1387 ,csa_tree_add_89_22_pad_groupi_n_1423);
  and csa_tree_add_89_22_pad_groupi_g4266(csa_tree_add_89_22_pad_groupi_n_1455 ,csa_tree_add_89_22_pad_groupi_n_1403 ,csa_tree_add_89_22_pad_groupi_n_1421);
  or csa_tree_add_89_22_pad_groupi_g4267(csa_tree_add_89_22_pad_groupi_n_1454 ,csa_tree_add_89_22_pad_groupi_n_1430 ,csa_tree_add_89_22_pad_groupi_n_1386);
  and csa_tree_add_89_22_pad_groupi_g4268(csa_tree_add_89_22_pad_groupi_n_1453 ,csa_tree_add_89_22_pad_groupi_n_1432 ,csa_tree_add_89_22_pad_groupi_n_1413);
  or csa_tree_add_89_22_pad_groupi_g4269(csa_tree_add_89_22_pad_groupi_n_1452 ,csa_tree_add_89_22_pad_groupi_n_1396 ,csa_tree_add_89_22_pad_groupi_n_1416);
  nor csa_tree_add_89_22_pad_groupi_g4270(csa_tree_add_89_22_pad_groupi_n_1451 ,csa_tree_add_89_22_pad_groupi_n_1397 ,csa_tree_add_89_22_pad_groupi_n_1417);
  or csa_tree_add_89_22_pad_groupi_g4271(csa_tree_add_89_22_pad_groupi_n_1450 ,csa_tree_add_89_22_pad_groupi_n_1367 ,csa_tree_add_89_22_pad_groupi_n_1414);
  nor csa_tree_add_89_22_pad_groupi_g4272(csa_tree_add_89_22_pad_groupi_n_1449 ,csa_tree_add_89_22_pad_groupi_n_1366 ,csa_tree_add_89_22_pad_groupi_n_1415);
  not csa_tree_add_89_22_pad_groupi_g4273(csa_tree_add_89_22_pad_groupi_n_1448 ,csa_tree_add_89_22_pad_groupi_n_1447);
  not csa_tree_add_89_22_pad_groupi_g4274(csa_tree_add_89_22_pad_groupi_n_1446 ,csa_tree_add_89_22_pad_groupi_n_1445);
  not csa_tree_add_89_22_pad_groupi_g4275(csa_tree_add_89_22_pad_groupi_n_1444 ,csa_tree_add_89_22_pad_groupi_n_1443);
  not csa_tree_add_89_22_pad_groupi_g4276(csa_tree_add_89_22_pad_groupi_n_1441 ,csa_tree_add_89_22_pad_groupi_n_1442);
  or csa_tree_add_89_22_pad_groupi_g4277(csa_tree_add_89_22_pad_groupi_n_1439 ,csa_tree_add_89_22_pad_groupi_n_1372 ,csa_tree_add_89_22_pad_groupi_n_1428);
  xnor csa_tree_add_89_22_pad_groupi_g4278(csa_tree_add_89_22_pad_groupi_n_1438 ,csa_tree_add_89_22_pad_groupi_n_1291 ,csa_tree_add_89_22_pad_groupi_n_1379);
  xnor csa_tree_add_89_22_pad_groupi_g4279(csa_tree_add_89_22_pad_groupi_n_1437 ,csa_tree_add_89_22_pad_groupi_n_1293 ,csa_tree_add_89_22_pad_groupi_n_1381);
  xnor csa_tree_add_89_22_pad_groupi_g4280(csa_tree_add_89_22_pad_groupi_n_1436 ,csa_tree_add_89_22_pad_groupi_n_1301 ,csa_tree_add_89_22_pad_groupi_n_1376);
  xnor csa_tree_add_89_22_pad_groupi_g4281(csa_tree_add_89_22_pad_groupi_n_1435 ,csa_tree_add_89_22_pad_groupi_n_1303 ,csa_tree_add_89_22_pad_groupi_n_1383);
  xnor csa_tree_add_89_22_pad_groupi_g4282(csa_tree_add_89_22_pad_groupi_n_1434 ,csa_tree_add_89_22_pad_groupi_n_1377 ,csa_tree_add_89_22_pad_groupi_n_1398);
  xnor csa_tree_add_89_22_pad_groupi_g4283(csa_tree_add_89_22_pad_groupi_n_1433 ,csa_tree_add_89_22_pad_groupi_n_1298 ,csa_tree_add_89_22_pad_groupi_n_1386);
  or csa_tree_add_89_22_pad_groupi_g4284(csa_tree_add_89_22_pad_groupi_n_1447 ,csa_tree_add_89_22_pad_groupi_n_1340 ,csa_tree_add_89_22_pad_groupi_n_1420);
  xnor csa_tree_add_89_22_pad_groupi_g4285(csa_tree_add_89_22_pad_groupi_n_1445 ,csa_tree_add_89_22_pad_groupi_n_1334 ,csa_tree_add_89_22_pad_groupi_n_1370);
  xnor csa_tree_add_89_22_pad_groupi_g4286(csa_tree_add_89_22_pad_groupi_n_1443 ,csa_tree_add_89_22_pad_groupi_n_1385 ,csa_tree_add_89_22_pad_groupi_n_1369);
  or csa_tree_add_89_22_pad_groupi_g4287(csa_tree_add_89_22_pad_groupi_n_1442 ,csa_tree_add_89_22_pad_groupi_n_1374 ,csa_tree_add_89_22_pad_groupi_n_1409);
  and csa_tree_add_89_22_pad_groupi_g4288(csa_tree_add_89_22_pad_groupi_n_1440 ,csa_tree_add_89_22_pad_groupi_n_1395 ,csa_tree_add_89_22_pad_groupi_n_1408);
  or csa_tree_add_89_22_pad_groupi_g4289(csa_tree_add_89_22_pad_groupi_n_1431 ,csa_tree_add_89_22_pad_groupi_n_1297 ,csa_tree_add_89_22_pad_groupi_n_1399);
  nor csa_tree_add_89_22_pad_groupi_g4290(csa_tree_add_89_22_pad_groupi_n_1430 ,csa_tree_add_89_22_pad_groupi_n_1298 ,csa_tree_add_89_22_pad_groupi_n_1400);
  nor csa_tree_add_89_22_pad_groupi_g4291(csa_tree_add_89_22_pad_groupi_n_1429 ,csa_tree_add_89_22_pad_groupi_n_1300 ,csa_tree_add_89_22_pad_groupi_n_1376);
  nor csa_tree_add_89_22_pad_groupi_g4292(csa_tree_add_89_22_pad_groupi_n_1428 ,csa_tree_add_89_22_pad_groupi_n_1363 ,csa_tree_add_89_22_pad_groupi_n_1394);
  or csa_tree_add_89_22_pad_groupi_g4293(csa_tree_add_89_22_pad_groupi_n_1427 ,csa_tree_add_89_22_pad_groupi_n_1301 ,csa_tree_add_89_22_pad_groupi_n_1375);
  nor csa_tree_add_89_22_pad_groupi_g4294(csa_tree_add_89_22_pad_groupi_n_1426 ,csa_tree_add_89_22_pad_groupi_n_1292 ,csa_tree_add_89_22_pad_groupi_n_1381);
  or csa_tree_add_89_22_pad_groupi_g4295(csa_tree_add_89_22_pad_groupi_n_1425 ,csa_tree_add_89_22_pad_groupi_n_1293 ,csa_tree_add_89_22_pad_groupi_n_1380);
  nor csa_tree_add_89_22_pad_groupi_g4296(csa_tree_add_89_22_pad_groupi_n_1424 ,csa_tree_add_89_22_pad_groupi_n_1290 ,csa_tree_add_89_22_pad_groupi_n_1379);
  or csa_tree_add_89_22_pad_groupi_g4297(csa_tree_add_89_22_pad_groupi_n_1423 ,csa_tree_add_89_22_pad_groupi_n_1291 ,csa_tree_add_89_22_pad_groupi_n_1378);
  nor csa_tree_add_89_22_pad_groupi_g4298(csa_tree_add_89_22_pad_groupi_n_1422 ,csa_tree_add_89_22_pad_groupi_n_1302 ,csa_tree_add_89_22_pad_groupi_n_1383);
  or csa_tree_add_89_22_pad_groupi_g4299(csa_tree_add_89_22_pad_groupi_n_1421 ,csa_tree_add_89_22_pad_groupi_n_1303 ,csa_tree_add_89_22_pad_groupi_n_1382);
  nor csa_tree_add_89_22_pad_groupi_g4300(csa_tree_add_89_22_pad_groupi_n_1420 ,csa_tree_add_89_22_pad_groupi_n_1355 ,csa_tree_add_89_22_pad_groupi_n_1385);
  or csa_tree_add_89_22_pad_groupi_g4301(csa_tree_add_89_22_pad_groupi_n_1432 ,csa_tree_add_89_22_pad_groupi_n_1365 ,csa_tree_add_89_22_pad_groupi_n_1391);
  not csa_tree_add_89_22_pad_groupi_g4302(csa_tree_add_89_22_pad_groupi_n_1419 ,csa_tree_add_89_22_pad_groupi_n_1418);
  not csa_tree_add_89_22_pad_groupi_g4303(csa_tree_add_89_22_pad_groupi_n_1417 ,csa_tree_add_89_22_pad_groupi_n_1416);
  not csa_tree_add_89_22_pad_groupi_g4304(csa_tree_add_89_22_pad_groupi_n_1415 ,csa_tree_add_89_22_pad_groupi_n_1414);
  not csa_tree_add_89_22_pad_groupi_g4305(csa_tree_add_89_22_pad_groupi_n_1412 ,csa_tree_add_89_22_pad_groupi_n_1411);
  or csa_tree_add_89_22_pad_groupi_g4306(csa_tree_add_89_22_pad_groupi_n_1410 ,csa_tree_add_89_22_pad_groupi_n_1377 ,csa_tree_add_89_22_pad_groupi_n_1398);
  nor csa_tree_add_89_22_pad_groupi_g4307(csa_tree_add_89_22_pad_groupi_n_1409 ,csa_tree_add_89_22_pad_groupi_n_1384 ,csa_tree_add_89_22_pad_groupi_n_1392);
  or csa_tree_add_89_22_pad_groupi_g4308(csa_tree_add_89_22_pad_groupi_n_1408 ,csa_tree_add_89_22_pad_groupi_n_1368 ,csa_tree_add_89_22_pad_groupi_n_1373);
  and csa_tree_add_89_22_pad_groupi_g4309(csa_tree_add_89_22_pad_groupi_n_1407 ,csa_tree_add_89_22_pad_groupi_n_1377 ,csa_tree_add_89_22_pad_groupi_n_1398);
  xnor csa_tree_add_89_22_pad_groupi_g4310(csa_tree_add_89_22_pad_groupi_n_1406 ,csa_tree_add_89_22_pad_groupi_n_1280 ,csa_tree_add_89_22_pad_groupi_n_1346);
  xnor csa_tree_add_89_22_pad_groupi_g4312(csa_tree_add_89_22_pad_groupi_n_1405 ,csa_tree_add_89_22_pad_groupi_n_1304 ,csa_tree_add_89_22_pad_groupi_n_1348);
  xnor csa_tree_add_89_22_pad_groupi_g4313(csa_tree_add_89_22_pad_groupi_n_1404 ,csa_tree_add_89_22_pad_groupi_n_1309 ,csa_tree_add_89_22_pad_groupi_n_1345);
  and csa_tree_add_89_22_pad_groupi_g4314(csa_tree_add_89_22_pad_groupi_n_1418 ,csa_tree_add_89_22_pad_groupi_n_1354 ,csa_tree_add_89_22_pad_groupi_n_1390);
  xnor csa_tree_add_89_22_pad_groupi_g4315(csa_tree_add_89_22_pad_groupi_n_1416 ,csa_tree_add_89_22_pad_groupi_n_1311 ,csa_tree_add_89_22_pad_groupi_n_1337);
  xnor csa_tree_add_89_22_pad_groupi_g4316(csa_tree_add_89_22_pad_groupi_n_1414 ,csa_tree_add_89_22_pad_groupi_n_1320 ,csa_tree_add_89_22_pad_groupi_n_1335);
  xnor csa_tree_add_89_22_pad_groupi_g4317(csa_tree_add_89_22_pad_groupi_n_1413 ,csa_tree_add_89_22_pad_groupi_n_1333 ,csa_tree_add_89_22_pad_groupi_n_1338);
  and csa_tree_add_89_22_pad_groupi_g4318(csa_tree_add_89_22_pad_groupi_n_1411 ,csa_tree_add_89_22_pad_groupi_n_1356 ,csa_tree_add_89_22_pad_groupi_n_1388);
  not csa_tree_add_89_22_pad_groupi_g4319(csa_tree_add_89_22_pad_groupi_n_1400 ,csa_tree_add_89_22_pad_groupi_n_1399);
  not csa_tree_add_89_22_pad_groupi_g4320(csa_tree_add_89_22_pad_groupi_n_1396 ,csa_tree_add_89_22_pad_groupi_n_1397);
  or csa_tree_add_89_22_pad_groupi_g4321(csa_tree_add_89_22_pad_groupi_n_1395 ,csa_tree_add_89_22_pad_groupi_n_1280 ,csa_tree_add_89_22_pad_groupi_n_1347);
  nor csa_tree_add_89_22_pad_groupi_g4322(csa_tree_add_89_22_pad_groupi_n_1394 ,csa_tree_add_89_22_pad_groupi_n_1362 ,csa_tree_add_89_22_pad_groupi_n_1361);
  and csa_tree_add_89_22_pad_groupi_g4323(csa_tree_add_89_22_pad_groupi_n_1393 ,csa_tree_add_89_22_pad_groupi_n_1309 ,csa_tree_add_89_22_pad_groupi_n_1345);
  and csa_tree_add_89_22_pad_groupi_g4324(csa_tree_add_89_22_pad_groupi_n_1392 ,csa_tree_add_89_22_pad_groupi_n_1304 ,csa_tree_add_89_22_pad_groupi_n_1349);
  and csa_tree_add_89_22_pad_groupi_g4325(csa_tree_add_89_22_pad_groupi_n_1391 ,csa_tree_add_89_22_pad_groupi_n_1334 ,csa_tree_add_89_22_pad_groupi_n_1360);
  or csa_tree_add_89_22_pad_groupi_g4326(csa_tree_add_89_22_pad_groupi_n_1390 ,csa_tree_add_89_22_pad_groupi_n_1353 ,csa_tree_add_89_22_pad_groupi_n_1350);
  or csa_tree_add_89_22_pad_groupi_g4327(csa_tree_add_89_22_pad_groupi_n_1389 ,csa_tree_add_89_22_pad_groupi_n_1309 ,csa_tree_add_89_22_pad_groupi_n_1345);
  or csa_tree_add_89_22_pad_groupi_g4328(csa_tree_add_89_22_pad_groupi_n_1388 ,csa_tree_add_89_22_pad_groupi_n_1305 ,csa_tree_add_89_22_pad_groupi_n_1342);
  or csa_tree_add_89_22_pad_groupi_g4329(csa_tree_add_89_22_pad_groupi_n_1403 ,csa_tree_add_89_22_pad_groupi_n_1246 ,csa_tree_add_89_22_pad_groupi_n_1359);
  or csa_tree_add_89_22_pad_groupi_g4330(csa_tree_add_89_22_pad_groupi_n_1402 ,csa_tree_add_89_22_pad_groupi_n_1230 ,csa_tree_add_89_22_pad_groupi_n_1343);
  or csa_tree_add_89_22_pad_groupi_g4331(csa_tree_add_89_22_pad_groupi_n_1401 ,csa_tree_add_89_22_pad_groupi_n_1232 ,csa_tree_add_89_22_pad_groupi_n_1339);
  and csa_tree_add_89_22_pad_groupi_g4332(csa_tree_add_89_22_pad_groupi_n_1399 ,csa_tree_add_89_22_pad_groupi_n_1254 ,csa_tree_add_89_22_pad_groupi_n_1364);
  or csa_tree_add_89_22_pad_groupi_g4333(csa_tree_add_89_22_pad_groupi_n_1398 ,csa_tree_add_89_22_pad_groupi_n_1329 ,csa_tree_add_89_22_pad_groupi_n_1357);
  or csa_tree_add_89_22_pad_groupi_g4334(csa_tree_add_89_22_pad_groupi_n_1397 ,csa_tree_add_89_22_pad_groupi_n_1323 ,csa_tree_add_89_22_pad_groupi_n_1358);
  not csa_tree_add_89_22_pad_groupi_g4335(csa_tree_add_89_22_pad_groupi_n_1383 ,csa_tree_add_89_22_pad_groupi_n_1382);
  not csa_tree_add_89_22_pad_groupi_g4336(csa_tree_add_89_22_pad_groupi_n_1381 ,csa_tree_add_89_22_pad_groupi_n_1380);
  not csa_tree_add_89_22_pad_groupi_g4337(csa_tree_add_89_22_pad_groupi_n_1379 ,csa_tree_add_89_22_pad_groupi_n_1378);
  not csa_tree_add_89_22_pad_groupi_g4338(csa_tree_add_89_22_pad_groupi_n_1376 ,csa_tree_add_89_22_pad_groupi_n_1375);
  nor csa_tree_add_89_22_pad_groupi_g4339(csa_tree_add_89_22_pad_groupi_n_1374 ,csa_tree_add_89_22_pad_groupi_n_1304 ,csa_tree_add_89_22_pad_groupi_n_1349);
  and csa_tree_add_89_22_pad_groupi_g4340(csa_tree_add_89_22_pad_groupi_n_1373 ,csa_tree_add_89_22_pad_groupi_n_1280 ,csa_tree_add_89_22_pad_groupi_n_1347);
  nor csa_tree_add_89_22_pad_groupi_g4341(csa_tree_add_89_22_pad_groupi_n_1372 ,csa_tree_add_89_22_pad_groupi_n_1306 ,csa_tree_add_89_22_pad_groupi_n_1352);
  or csa_tree_add_89_22_pad_groupi_g4342(csa_tree_add_89_22_pad_groupi_n_1371 ,csa_tree_add_89_22_pad_groupi_n_1307 ,csa_tree_add_89_22_pad_groupi_n_1351);
  xnor csa_tree_add_89_22_pad_groupi_g4343(csa_tree_add_89_22_pad_groupi_n_1370 ,csa_tree_add_89_22_pad_groupi_n_1261 ,csa_tree_add_89_22_pad_groupi_n_1310);
  xnor csa_tree_add_89_22_pad_groupi_g4344(csa_tree_add_89_22_pad_groupi_n_1369 ,csa_tree_add_89_22_pad_groupi_n_1299 ,csa_tree_add_89_22_pad_groupi_n_1330);
  or csa_tree_add_89_22_pad_groupi_g4345(csa_tree_add_89_22_pad_groupi_n_1387 ,csa_tree_add_89_22_pad_groupi_n_1227 ,csa_tree_add_89_22_pad_groupi_n_1341);
  xnor csa_tree_add_89_22_pad_groupi_g4346(csa_tree_add_89_22_pad_groupi_n_1386 ,csa_tree_add_89_22_pad_groupi_n_1317 ,csa_tree_add_89_22_pad_groupi_n_1273);
  xnor csa_tree_add_89_22_pad_groupi_g4347(csa_tree_add_89_22_pad_groupi_n_1385 ,csa_tree_add_89_22_pad_groupi_n_1316 ,csa_tree_add_89_22_pad_groupi_n_1268);
  and csa_tree_add_89_22_pad_groupi_g4348(csa_tree_add_89_22_pad_groupi_n_1384 ,csa_tree_add_89_22_pad_groupi_n_1225 ,csa_tree_add_89_22_pad_groupi_n_1344);
  xnor csa_tree_add_89_22_pad_groupi_g4349(csa_tree_add_89_22_pad_groupi_n_1382 ,csa_tree_add_89_22_pad_groupi_n_1313 ,csa_tree_add_89_22_pad_groupi_n_1266);
  xnor csa_tree_add_89_22_pad_groupi_g4350(csa_tree_add_89_22_pad_groupi_n_1380 ,csa_tree_add_89_22_pad_groupi_n_1315 ,csa_tree_add_89_22_pad_groupi_n_1270);
  xnor csa_tree_add_89_22_pad_groupi_g4351(csa_tree_add_89_22_pad_groupi_n_1378 ,csa_tree_add_89_22_pad_groupi_n_1314 ,csa_tree_add_89_22_pad_groupi_n_1267);
  xnor csa_tree_add_89_22_pad_groupi_g4352(csa_tree_add_89_22_pad_groupi_n_1377 ,csa_tree_add_89_22_pad_groupi_n_1262 ,csa_tree_add_89_22_pad_groupi_n_1308);
  xnor csa_tree_add_89_22_pad_groupi_g4353(csa_tree_add_89_22_pad_groupi_n_1375 ,csa_tree_add_89_22_pad_groupi_n_1318 ,csa_tree_add_89_22_pad_groupi_n_1271);
  not csa_tree_add_89_22_pad_groupi_g4355(csa_tree_add_89_22_pad_groupi_n_1367 ,csa_tree_add_89_22_pad_groupi_n_1366);
  and csa_tree_add_89_22_pad_groupi_g4356(csa_tree_add_89_22_pad_groupi_n_1365 ,csa_tree_add_89_22_pad_groupi_n_1261 ,csa_tree_add_89_22_pad_groupi_n_1310);
  or csa_tree_add_89_22_pad_groupi_g4357(csa_tree_add_89_22_pad_groupi_n_1364 ,csa_tree_add_89_22_pad_groupi_n_1224 ,csa_tree_add_89_22_pad_groupi_n_1319);
  and csa_tree_add_89_22_pad_groupi_g4358(csa_tree_add_89_22_pad_groupi_n_1363 ,csa_tree_add_89_22_pad_groupi_n_1265 ,csa_tree_add_89_22_pad_groupi_n_1321);
  nor csa_tree_add_89_22_pad_groupi_g4359(csa_tree_add_89_22_pad_groupi_n_1362 ,csa_tree_add_89_22_pad_groupi_n_1265 ,csa_tree_add_89_22_pad_groupi_n_1321);
  nor csa_tree_add_89_22_pad_groupi_g4360(csa_tree_add_89_22_pad_groupi_n_1361 ,csa_tree_add_89_22_pad_groupi_n_1285 ,csa_tree_add_89_22_pad_groupi_n_1326);
  or csa_tree_add_89_22_pad_groupi_g4361(csa_tree_add_89_22_pad_groupi_n_1360 ,csa_tree_add_89_22_pad_groupi_n_1261 ,csa_tree_add_89_22_pad_groupi_n_1310);
  nor csa_tree_add_89_22_pad_groupi_g4362(csa_tree_add_89_22_pad_groupi_n_1359 ,csa_tree_add_89_22_pad_groupi_n_1245 ,csa_tree_add_89_22_pad_groupi_n_1316);
  nor csa_tree_add_89_22_pad_groupi_g4363(csa_tree_add_89_22_pad_groupi_n_1358 ,csa_tree_add_89_22_pad_groupi_n_1328 ,csa_tree_add_89_22_pad_groupi_n_1320);
  nor csa_tree_add_89_22_pad_groupi_g4364(csa_tree_add_89_22_pad_groupi_n_1357 ,csa_tree_add_89_22_pad_groupi_n_1333 ,csa_tree_add_89_22_pad_groupi_n_1322);
  or csa_tree_add_89_22_pad_groupi_g4365(csa_tree_add_89_22_pad_groupi_n_1356 ,csa_tree_add_89_22_pad_groupi_n_1278 ,csa_tree_add_89_22_pad_groupi_n_1312);
  nor csa_tree_add_89_22_pad_groupi_g4366(csa_tree_add_89_22_pad_groupi_n_1355 ,csa_tree_add_89_22_pad_groupi_n_1299 ,csa_tree_add_89_22_pad_groupi_n_1330);
  or csa_tree_add_89_22_pad_groupi_g4367(csa_tree_add_89_22_pad_groupi_n_1354 ,csa_tree_add_89_22_pad_groupi_n_1294 ,csa_tree_add_89_22_pad_groupi_n_1332);
  nor csa_tree_add_89_22_pad_groupi_g4368(csa_tree_add_89_22_pad_groupi_n_1353 ,csa_tree_add_89_22_pad_groupi_n_1295 ,csa_tree_add_89_22_pad_groupi_n_1331);
  and csa_tree_add_89_22_pad_groupi_g4369(csa_tree_add_89_22_pad_groupi_n_1368 ,csa_tree_add_89_22_pad_groupi_n_1243 ,csa_tree_add_89_22_pad_groupi_n_1324);
  or csa_tree_add_89_22_pad_groupi_g4370(csa_tree_add_89_22_pad_groupi_n_1366 ,csa_tree_add_89_22_pad_groupi_n_1185 ,csa_tree_add_89_22_pad_groupi_n_1327);
  not csa_tree_add_89_22_pad_groupi_g4371(csa_tree_add_89_22_pad_groupi_n_1352 ,csa_tree_add_89_22_pad_groupi_n_1351);
  not csa_tree_add_89_22_pad_groupi_g4373(csa_tree_add_89_22_pad_groupi_n_1349 ,csa_tree_add_89_22_pad_groupi_n_1348);
  not csa_tree_add_89_22_pad_groupi_g4374(csa_tree_add_89_22_pad_groupi_n_1347 ,csa_tree_add_89_22_pad_groupi_n_1346);
  or csa_tree_add_89_22_pad_groupi_g4375(csa_tree_add_89_22_pad_groupi_n_1344 ,csa_tree_add_89_22_pad_groupi_n_1223 ,csa_tree_add_89_22_pad_groupi_n_1317);
  and csa_tree_add_89_22_pad_groupi_g4376(csa_tree_add_89_22_pad_groupi_n_1343 ,csa_tree_add_89_22_pad_groupi_n_1228 ,csa_tree_add_89_22_pad_groupi_n_1314);
  and csa_tree_add_89_22_pad_groupi_g4377(csa_tree_add_89_22_pad_groupi_n_1342 ,csa_tree_add_89_22_pad_groupi_n_1278 ,csa_tree_add_89_22_pad_groupi_n_1312);
  and csa_tree_add_89_22_pad_groupi_g4378(csa_tree_add_89_22_pad_groupi_n_1341 ,csa_tree_add_89_22_pad_groupi_n_1226 ,csa_tree_add_89_22_pad_groupi_n_1313);
  and csa_tree_add_89_22_pad_groupi_g4379(csa_tree_add_89_22_pad_groupi_n_1340 ,csa_tree_add_89_22_pad_groupi_n_1299 ,csa_tree_add_89_22_pad_groupi_n_1330);
  and csa_tree_add_89_22_pad_groupi_g4380(csa_tree_add_89_22_pad_groupi_n_1339 ,csa_tree_add_89_22_pad_groupi_n_1231 ,csa_tree_add_89_22_pad_groupi_n_1315);
  xnor csa_tree_add_89_22_pad_groupi_g4381(csa_tree_add_89_22_pad_groupi_n_1338 ,csa_tree_add_89_22_pad_groupi_n_1201 ,csa_tree_add_89_22_pad_groupi_n_1279);
  xnor csa_tree_add_89_22_pad_groupi_g4382(csa_tree_add_89_22_pad_groupi_n_1351 ,csa_tree_add_89_22_pad_groupi_n_1281 ,csa_tree_add_89_22_pad_groupi_n_1211);
  xor csa_tree_add_89_22_pad_groupi_g4383(csa_tree_add_89_22_pad_groupi_n_1337 ,csa_tree_add_89_22_pad_groupi_n_1278 ,csa_tree_add_89_22_pad_groupi_n_1305);
  xnor csa_tree_add_89_22_pad_groupi_g4384(csa_tree_add_89_22_pad_groupi_n_1336 ,csa_tree_add_89_22_pad_groupi_n_1075 ,csa_tree_add_89_22_pad_groupi_n_1274);
  xnor csa_tree_add_89_22_pad_groupi_g4385(csa_tree_add_89_22_pad_groupi_n_1335 ,csa_tree_add_89_22_pad_groupi_n_1235 ,csa_tree_add_89_22_pad_groupi_n_1296);
  xnor csa_tree_add_89_22_pad_groupi_g4386(csa_tree_add_89_22_pad_groupi_n_1350 ,csa_tree_add_89_22_pad_groupi_n_1264 ,csa_tree_add_89_22_pad_groupi_n_1272);
  xnor csa_tree_add_89_22_pad_groupi_g4387(csa_tree_add_89_22_pad_groupi_n_1348 ,csa_tree_add_89_22_pad_groupi_n_1282 ,csa_tree_add_89_22_pad_groupi_n_1269);
  xnor csa_tree_add_89_22_pad_groupi_g4388(csa_tree_add_89_22_pad_groupi_n_1346 ,csa_tree_add_89_22_pad_groupi_n_1263 ,csa_tree_add_89_22_pad_groupi_n_1275);
  or csa_tree_add_89_22_pad_groupi_g4389(csa_tree_add_89_22_pad_groupi_n_1345 ,csa_tree_add_89_22_pad_groupi_n_1277 ,csa_tree_add_89_22_pad_groupi_n_1325);
  not csa_tree_add_89_22_pad_groupi_g4390(csa_tree_add_89_22_pad_groupi_n_1332 ,csa_tree_add_89_22_pad_groupi_n_1331);
  nor csa_tree_add_89_22_pad_groupi_g4391(csa_tree_add_89_22_pad_groupi_n_1329 ,csa_tree_add_89_22_pad_groupi_n_1202 ,csa_tree_add_89_22_pad_groupi_n_1279);
  nor csa_tree_add_89_22_pad_groupi_g4392(csa_tree_add_89_22_pad_groupi_n_1328 ,csa_tree_add_89_22_pad_groupi_n_1235 ,csa_tree_add_89_22_pad_groupi_n_1296);
  nor csa_tree_add_89_22_pad_groupi_g4393(csa_tree_add_89_22_pad_groupi_n_1327 ,csa_tree_add_89_22_pad_groupi_n_1184 ,csa_tree_add_89_22_pad_groupi_n_1281);
  nor csa_tree_add_89_22_pad_groupi_g4394(csa_tree_add_89_22_pad_groupi_n_1326 ,csa_tree_add_89_22_pad_groupi_n_1287 ,csa_tree_add_89_22_pad_groupi_n_1288);
  nor csa_tree_add_89_22_pad_groupi_g4395(csa_tree_add_89_22_pad_groupi_n_1325 ,csa_tree_add_89_22_pad_groupi_n_1276 ,csa_tree_add_89_22_pad_groupi_n_1262);
  or csa_tree_add_89_22_pad_groupi_g4396(csa_tree_add_89_22_pad_groupi_n_1324 ,csa_tree_add_89_22_pad_groupi_n_1252 ,csa_tree_add_89_22_pad_groupi_n_1283);
  and csa_tree_add_89_22_pad_groupi_g4397(csa_tree_add_89_22_pad_groupi_n_1323 ,csa_tree_add_89_22_pad_groupi_n_1235 ,csa_tree_add_89_22_pad_groupi_n_1296);
  and csa_tree_add_89_22_pad_groupi_g4398(csa_tree_add_89_22_pad_groupi_n_1322 ,csa_tree_add_89_22_pad_groupi_n_1202 ,csa_tree_add_89_22_pad_groupi_n_1279);
  or csa_tree_add_89_22_pad_groupi_g4399(csa_tree_add_89_22_pad_groupi_n_1334 ,csa_tree_add_89_22_pad_groupi_n_1240 ,csa_tree_add_89_22_pad_groupi_n_1284);
  and csa_tree_add_89_22_pad_groupi_g4400(csa_tree_add_89_22_pad_groupi_n_1333 ,csa_tree_add_89_22_pad_groupi_n_1156 ,csa_tree_add_89_22_pad_groupi_n_1286);
  xnor csa_tree_add_89_22_pad_groupi_g4401(csa_tree_add_89_22_pad_groupi_n_1331 ,csa_tree_add_89_22_pad_groupi_n_1039 ,csa_tree_add_89_22_pad_groupi_n_1216);
  or csa_tree_add_89_22_pad_groupi_g4402(csa_tree_add_89_22_pad_groupi_n_1330 ,csa_tree_add_89_22_pad_groupi_n_1242 ,csa_tree_add_89_22_pad_groupi_n_1289);
  not csa_tree_add_89_22_pad_groupi_g4403(csa_tree_add_89_22_pad_groupi_n_1319 ,csa_tree_add_89_22_pad_groupi_n_1318);
  not csa_tree_add_89_22_pad_groupi_g4404(csa_tree_add_89_22_pad_groupi_n_1312 ,csa_tree_add_89_22_pad_groupi_n_1311);
  xnor csa_tree_add_89_22_pad_groupi_g4405(csa_tree_add_89_22_pad_groupi_n_1321 ,csa_tree_add_89_22_pad_groupi_n_1176 ,csa_tree_add_89_22_pad_groupi_n_1210);
  xnor csa_tree_add_89_22_pad_groupi_g4406(csa_tree_add_89_22_pad_groupi_n_1308 ,csa_tree_add_89_22_pad_groupi_n_1132 ,csa_tree_add_89_22_pad_groupi_n_1233);
  xnor csa_tree_add_89_22_pad_groupi_g4407(csa_tree_add_89_22_pad_groupi_n_1320 ,csa_tree_add_89_22_pad_groupi_n_1084 ,csa_tree_add_89_22_pad_groupi_n_1220);
  xnor csa_tree_add_89_22_pad_groupi_g4408(csa_tree_add_89_22_pad_groupi_n_1318 ,csa_tree_add_89_22_pad_groupi_n_1138 ,csa_tree_add_89_22_pad_groupi_n_1221);
  xnor csa_tree_add_89_22_pad_groupi_g4409(csa_tree_add_89_22_pad_groupi_n_1317 ,csa_tree_add_89_22_pad_groupi_n_1092 ,csa_tree_add_89_22_pad_groupi_n_1213);
  xnor csa_tree_add_89_22_pad_groupi_g4410(csa_tree_add_89_22_pad_groupi_n_1316 ,csa_tree_add_89_22_pad_groupi_n_1088 ,csa_tree_add_89_22_pad_groupi_n_1214);
  xnor csa_tree_add_89_22_pad_groupi_g4411(csa_tree_add_89_22_pad_groupi_n_1315 ,csa_tree_add_89_22_pad_groupi_n_1141 ,csa_tree_add_89_22_pad_groupi_n_1218);
  xnor csa_tree_add_89_22_pad_groupi_g4412(csa_tree_add_89_22_pad_groupi_n_1314 ,csa_tree_add_89_22_pad_groupi_n_1102 ,csa_tree_add_89_22_pad_groupi_n_1217);
  xnor csa_tree_add_89_22_pad_groupi_g4413(csa_tree_add_89_22_pad_groupi_n_1313 ,csa_tree_add_89_22_pad_groupi_n_1107 ,csa_tree_add_89_22_pad_groupi_n_1222);
  xnor csa_tree_add_89_22_pad_groupi_g4414(csa_tree_add_89_22_pad_groupi_n_1311 ,csa_tree_add_89_22_pad_groupi_n_1209 ,csa_tree_add_89_22_pad_groupi_n_1215);
  xnor csa_tree_add_89_22_pad_groupi_g4415(csa_tree_add_89_22_pad_groupi_n_1310 ,csa_tree_add_89_22_pad_groupi_n_1236 ,csa_tree_add_89_22_pad_groupi_n_1212);
  xnor csa_tree_add_89_22_pad_groupi_g4416(csa_tree_add_89_22_pad_groupi_n_1309 ,csa_tree_add_89_22_pad_groupi_n_1175 ,csa_tree_add_89_22_pad_groupi_n_1219);
  not csa_tree_add_89_22_pad_groupi_g4417(csa_tree_add_89_22_pad_groupi_n_1307 ,csa_tree_add_89_22_pad_groupi_n_1306);
  not csa_tree_add_89_22_pad_groupi_g4418(csa_tree_add_89_22_pad_groupi_n_1302 ,csa_tree_add_89_22_pad_groupi_n_1303);
  not csa_tree_add_89_22_pad_groupi_g4419(csa_tree_add_89_22_pad_groupi_n_1300 ,csa_tree_add_89_22_pad_groupi_n_1301);
  not csa_tree_add_89_22_pad_groupi_g4420(csa_tree_add_89_22_pad_groupi_n_1297 ,csa_tree_add_89_22_pad_groupi_n_1298);
  not csa_tree_add_89_22_pad_groupi_g4421(csa_tree_add_89_22_pad_groupi_n_1295 ,csa_tree_add_89_22_pad_groupi_n_1294);
  not csa_tree_add_89_22_pad_groupi_g4422(csa_tree_add_89_22_pad_groupi_n_1292 ,csa_tree_add_89_22_pad_groupi_n_1293);
  not csa_tree_add_89_22_pad_groupi_g4423(csa_tree_add_89_22_pad_groupi_n_1290 ,csa_tree_add_89_22_pad_groupi_n_1291);
  nor csa_tree_add_89_22_pad_groupi_g4424(csa_tree_add_89_22_pad_groupi_n_1289 ,csa_tree_add_89_22_pad_groupi_n_1247 ,csa_tree_add_89_22_pad_groupi_n_1264);
  nor csa_tree_add_89_22_pad_groupi_g4425(csa_tree_add_89_22_pad_groupi_n_1288 ,csa_tree_add_89_22_pad_groupi_n_1048 ,csa_tree_add_89_22_pad_groupi_n_1238);
  nor csa_tree_add_89_22_pad_groupi_g4426(csa_tree_add_89_22_pad_groupi_n_1287 ,csa_tree_add_89_22_pad_groupi_n_1178 ,csa_tree_add_89_22_pad_groupi_n_1251);
  or csa_tree_add_89_22_pad_groupi_g4427(csa_tree_add_89_22_pad_groupi_n_1286 ,csa_tree_add_89_22_pad_groupi_n_1150 ,csa_tree_add_89_22_pad_groupi_n_1237);
  nor csa_tree_add_89_22_pad_groupi_g4428(csa_tree_add_89_22_pad_groupi_n_1285 ,csa_tree_add_89_22_pad_groupi_n_1047 ,csa_tree_add_89_22_pad_groupi_n_1239);
  and csa_tree_add_89_22_pad_groupi_g4429(csa_tree_add_89_22_pad_groupi_n_1284 ,csa_tree_add_89_22_pad_groupi_n_1241 ,csa_tree_add_89_22_pad_groupi_n_1263);
  or csa_tree_add_89_22_pad_groupi_g4430(csa_tree_add_89_22_pad_groupi_n_1306 ,csa_tree_add_89_22_pad_groupi_n_1183 ,csa_tree_add_89_22_pad_groupi_n_1253);
  and csa_tree_add_89_22_pad_groupi_g4431(csa_tree_add_89_22_pad_groupi_n_1305 ,csa_tree_add_89_22_pad_groupi_n_1192 ,csa_tree_add_89_22_pad_groupi_n_1257);
  and csa_tree_add_89_22_pad_groupi_g4432(csa_tree_add_89_22_pad_groupi_n_1304 ,csa_tree_add_89_22_pad_groupi_n_1155 ,csa_tree_add_89_22_pad_groupi_n_1260);
  or csa_tree_add_89_22_pad_groupi_g4433(csa_tree_add_89_22_pad_groupi_n_1303 ,csa_tree_add_89_22_pad_groupi_n_1154 ,csa_tree_add_89_22_pad_groupi_n_1248);
  or csa_tree_add_89_22_pad_groupi_g4434(csa_tree_add_89_22_pad_groupi_n_1301 ,csa_tree_add_89_22_pad_groupi_n_1187 ,csa_tree_add_89_22_pad_groupi_n_1255);
  or csa_tree_add_89_22_pad_groupi_g4435(csa_tree_add_89_22_pad_groupi_n_1299 ,csa_tree_add_89_22_pad_groupi_n_1147 ,csa_tree_add_89_22_pad_groupi_n_1244);
  or csa_tree_add_89_22_pad_groupi_g4436(csa_tree_add_89_22_pad_groupi_n_1298 ,csa_tree_add_89_22_pad_groupi_n_1198 ,csa_tree_add_89_22_pad_groupi_n_1258);
  or csa_tree_add_89_22_pad_groupi_g4437(csa_tree_add_89_22_pad_groupi_n_1296 ,csa_tree_add_89_22_pad_groupi_n_1188 ,csa_tree_add_89_22_pad_groupi_n_1256);
  and csa_tree_add_89_22_pad_groupi_g4438(csa_tree_add_89_22_pad_groupi_n_1294 ,csa_tree_add_89_22_pad_groupi_n_1197 ,csa_tree_add_89_22_pad_groupi_n_1259);
  or csa_tree_add_89_22_pad_groupi_g4439(csa_tree_add_89_22_pad_groupi_n_1293 ,csa_tree_add_89_22_pad_groupi_n_1179 ,csa_tree_add_89_22_pad_groupi_n_1250);
  or csa_tree_add_89_22_pad_groupi_g4440(csa_tree_add_89_22_pad_groupi_n_1291 ,csa_tree_add_89_22_pad_groupi_n_1200 ,csa_tree_add_89_22_pad_groupi_n_1249);
  not csa_tree_add_89_22_pad_groupi_g4441(csa_tree_add_89_22_pad_groupi_n_1283 ,csa_tree_add_89_22_pad_groupi_n_1282);
  nor csa_tree_add_89_22_pad_groupi_g4442(csa_tree_add_89_22_pad_groupi_n_1277 ,csa_tree_add_89_22_pad_groupi_n_1132 ,csa_tree_add_89_22_pad_groupi_n_1234);
  and csa_tree_add_89_22_pad_groupi_g4443(csa_tree_add_89_22_pad_groupi_n_1276 ,csa_tree_add_89_22_pad_groupi_n_1132 ,csa_tree_add_89_22_pad_groupi_n_1234);
  xnor csa_tree_add_89_22_pad_groupi_g4444(csa_tree_add_89_22_pad_groupi_n_1275 ,csa_tree_add_89_22_pad_groupi_n_1207 ,csa_tree_add_89_22_pad_groupi_n_1098);
  nor csa_tree_add_89_22_pad_groupi_g4445(csa_tree_add_89_22_pad_groupi_n_1274 ,csa_tree_add_89_22_pad_groupi_n_1157 ,csa_tree_add_89_22_pad_groupi_n_1229);
  xnor csa_tree_add_89_22_pad_groupi_g4446(csa_tree_add_89_22_pad_groupi_n_1273 ,csa_tree_add_89_22_pad_groupi_n_1163 ,csa_tree_add_89_22_pad_groupi_n_1166);
  xnor csa_tree_add_89_22_pad_groupi_g4447(csa_tree_add_89_22_pad_groupi_n_1272 ,csa_tree_add_89_22_pad_groupi_n_1099 ,csa_tree_add_89_22_pad_groupi_n_1169);
  xnor csa_tree_add_89_22_pad_groupi_g4448(csa_tree_add_89_22_pad_groupi_n_1271 ,csa_tree_add_89_22_pad_groupi_n_1204 ,csa_tree_add_89_22_pad_groupi_n_1160);
  xnor csa_tree_add_89_22_pad_groupi_g4449(csa_tree_add_89_22_pad_groupi_n_1270 ,csa_tree_add_89_22_pad_groupi_n_1208 ,csa_tree_add_89_22_pad_groupi_n_1174);
  xnor csa_tree_add_89_22_pad_groupi_g4450(csa_tree_add_89_22_pad_groupi_n_1269 ,csa_tree_add_89_22_pad_groupi_n_1206 ,csa_tree_add_89_22_pad_groupi_n_1171);
  xnor csa_tree_add_89_22_pad_groupi_g4451(csa_tree_add_89_22_pad_groupi_n_1268 ,csa_tree_add_89_22_pad_groupi_n_1164 ,csa_tree_add_89_22_pad_groupi_n_1167);
  xnor csa_tree_add_89_22_pad_groupi_g4452(csa_tree_add_89_22_pad_groupi_n_1267 ,csa_tree_add_89_22_pad_groupi_n_1173 ,csa_tree_add_89_22_pad_groupi_n_1172);
  xnor csa_tree_add_89_22_pad_groupi_g4453(csa_tree_add_89_22_pad_groupi_n_1266 ,csa_tree_add_89_22_pad_groupi_n_1161 ,csa_tree_add_89_22_pad_groupi_n_1168);
  xnor csa_tree_add_89_22_pad_groupi_g4454(csa_tree_add_89_22_pad_groupi_n_1282 ,csa_tree_add_89_22_pad_groupi_n_1106 ,csa_tree_add_89_22_pad_groupi_n_1143);
  xnor csa_tree_add_89_22_pad_groupi_g4455(csa_tree_add_89_22_pad_groupi_n_1281 ,csa_tree_add_89_22_pad_groupi_n_1080 ,csa_tree_add_89_22_pad_groupi_n_1145);
  xnor csa_tree_add_89_22_pad_groupi_g4456(csa_tree_add_89_22_pad_groupi_n_1280 ,csa_tree_add_89_22_pad_groupi_n_1103 ,csa_tree_add_89_22_pad_groupi_n_1146);
  xnor csa_tree_add_89_22_pad_groupi_g4457(csa_tree_add_89_22_pad_groupi_n_1279 ,csa_tree_add_89_22_pad_groupi_n_1101 ,csa_tree_add_89_22_pad_groupi_n_1142);
  xnor csa_tree_add_89_22_pad_groupi_g4458(csa_tree_add_89_22_pad_groupi_n_1278 ,csa_tree_add_89_22_pad_groupi_n_1105 ,csa_tree_add_89_22_pad_groupi_n_1144);
  or csa_tree_add_89_22_pad_groupi_g4459(csa_tree_add_89_22_pad_groupi_n_1260 ,csa_tree_add_89_22_pad_groupi_n_1104 ,csa_tree_add_89_22_pad_groupi_n_1151);
  or csa_tree_add_89_22_pad_groupi_g4460(csa_tree_add_89_22_pad_groupi_n_1259 ,csa_tree_add_89_22_pad_groupi_n_1209 ,csa_tree_add_89_22_pad_groupi_n_1193);
  nor csa_tree_add_89_22_pad_groupi_g4461(csa_tree_add_89_22_pad_groupi_n_1258 ,csa_tree_add_89_22_pad_groupi_n_1074 ,csa_tree_add_89_22_pad_groupi_n_1195);
  or csa_tree_add_89_22_pad_groupi_g4462(csa_tree_add_89_22_pad_groupi_n_1257 ,csa_tree_add_89_22_pad_groupi_n_1072 ,csa_tree_add_89_22_pad_groupi_n_1190);
  nor csa_tree_add_89_22_pad_groupi_g4463(csa_tree_add_89_22_pad_groupi_n_1256 ,csa_tree_add_89_22_pad_groupi_n_1067 ,csa_tree_add_89_22_pad_groupi_n_1186);
  and csa_tree_add_89_22_pad_groupi_g4464(csa_tree_add_89_22_pad_groupi_n_1255 ,csa_tree_add_89_22_pad_groupi_n_1141 ,csa_tree_add_89_22_pad_groupi_n_1189);
  or csa_tree_add_89_22_pad_groupi_g4465(csa_tree_add_89_22_pad_groupi_n_1254 ,csa_tree_add_89_22_pad_groupi_n_1203 ,csa_tree_add_89_22_pad_groupi_n_1159);
  and csa_tree_add_89_22_pad_groupi_g4466(csa_tree_add_89_22_pad_groupi_n_1253 ,csa_tree_add_89_22_pad_groupi_n_1181 ,csa_tree_add_89_22_pad_groupi_n_1176);
  nor csa_tree_add_89_22_pad_groupi_g4467(csa_tree_add_89_22_pad_groupi_n_1252 ,csa_tree_add_89_22_pad_groupi_n_1206 ,csa_tree_add_89_22_pad_groupi_n_1171);
  nor csa_tree_add_89_22_pad_groupi_g4468(csa_tree_add_89_22_pad_groupi_n_1251 ,csa_tree_add_89_22_pad_groupi_n_1177 ,csa_tree_add_89_22_pad_groupi_n_1191);
  and csa_tree_add_89_22_pad_groupi_g4469(csa_tree_add_89_22_pad_groupi_n_1250 ,csa_tree_add_89_22_pad_groupi_n_1102 ,csa_tree_add_89_22_pad_groupi_n_1194);
  and csa_tree_add_89_22_pad_groupi_g4470(csa_tree_add_89_22_pad_groupi_n_1249 ,csa_tree_add_89_22_pad_groupi_n_1107 ,csa_tree_add_89_22_pad_groupi_n_1158);
  nor csa_tree_add_89_22_pad_groupi_g4471(csa_tree_add_89_22_pad_groupi_n_1248 ,csa_tree_add_89_22_pad_groupi_n_1042 ,csa_tree_add_89_22_pad_groupi_n_1153);
  nor csa_tree_add_89_22_pad_groupi_g4472(csa_tree_add_89_22_pad_groupi_n_1247 ,csa_tree_add_89_22_pad_groupi_n_1099 ,csa_tree_add_89_22_pad_groupi_n_1169);
  and csa_tree_add_89_22_pad_groupi_g4473(csa_tree_add_89_22_pad_groupi_n_1246 ,csa_tree_add_89_22_pad_groupi_n_1164 ,csa_tree_add_89_22_pad_groupi_n_1167);
  nor csa_tree_add_89_22_pad_groupi_g4474(csa_tree_add_89_22_pad_groupi_n_1245 ,csa_tree_add_89_22_pad_groupi_n_1164 ,csa_tree_add_89_22_pad_groupi_n_1167);
  nor csa_tree_add_89_22_pad_groupi_g4475(csa_tree_add_89_22_pad_groupi_n_1244 ,csa_tree_add_89_22_pad_groupi_n_1039 ,csa_tree_add_89_22_pad_groupi_n_1148);
  or csa_tree_add_89_22_pad_groupi_g4476(csa_tree_add_89_22_pad_groupi_n_1243 ,csa_tree_add_89_22_pad_groupi_n_1205 ,csa_tree_add_89_22_pad_groupi_n_1170);
  and csa_tree_add_89_22_pad_groupi_g4477(csa_tree_add_89_22_pad_groupi_n_1242 ,csa_tree_add_89_22_pad_groupi_n_1099 ,csa_tree_add_89_22_pad_groupi_n_1169);
  or csa_tree_add_89_22_pad_groupi_g4478(csa_tree_add_89_22_pad_groupi_n_1241 ,csa_tree_add_89_22_pad_groupi_n_1207 ,csa_tree_add_89_22_pad_groupi_n_1098);
  and csa_tree_add_89_22_pad_groupi_g4479(csa_tree_add_89_22_pad_groupi_n_1240 ,csa_tree_add_89_22_pad_groupi_n_1207 ,csa_tree_add_89_22_pad_groupi_n_1098);
  or csa_tree_add_89_22_pad_groupi_g4480(csa_tree_add_89_22_pad_groupi_n_1265 ,csa_tree_add_89_22_pad_groupi_n_1051 ,csa_tree_add_89_22_pad_groupi_n_1180);
  and csa_tree_add_89_22_pad_groupi_g4481(csa_tree_add_89_22_pad_groupi_n_1264 ,csa_tree_add_89_22_pad_groupi_n_1115 ,csa_tree_add_89_22_pad_groupi_n_1199);
  or csa_tree_add_89_22_pad_groupi_g4482(csa_tree_add_89_22_pad_groupi_n_1263 ,csa_tree_add_89_22_pad_groupi_n_1123 ,csa_tree_add_89_22_pad_groupi_n_1182);
  and csa_tree_add_89_22_pad_groupi_g4483(csa_tree_add_89_22_pad_groupi_n_1262 ,csa_tree_add_89_22_pad_groupi_n_1114 ,csa_tree_add_89_22_pad_groupi_n_1149);
  or csa_tree_add_89_22_pad_groupi_g4484(csa_tree_add_89_22_pad_groupi_n_1261 ,csa_tree_add_89_22_pad_groupi_n_1124 ,csa_tree_add_89_22_pad_groupi_n_1196);
  not csa_tree_add_89_22_pad_groupi_g4485(csa_tree_add_89_22_pad_groupi_n_1239 ,csa_tree_add_89_22_pad_groupi_n_1238);
  not csa_tree_add_89_22_pad_groupi_g4486(csa_tree_add_89_22_pad_groupi_n_1237 ,csa_tree_add_89_22_pad_groupi_n_1236);
  not csa_tree_add_89_22_pad_groupi_g4487(csa_tree_add_89_22_pad_groupi_n_1234 ,csa_tree_add_89_22_pad_groupi_n_1233);
  and csa_tree_add_89_22_pad_groupi_g4488(csa_tree_add_89_22_pad_groupi_n_1232 ,csa_tree_add_89_22_pad_groupi_n_1208 ,csa_tree_add_89_22_pad_groupi_n_1174);
  or csa_tree_add_89_22_pad_groupi_g4489(csa_tree_add_89_22_pad_groupi_n_1231 ,csa_tree_add_89_22_pad_groupi_n_1208 ,csa_tree_add_89_22_pad_groupi_n_1174);
  and csa_tree_add_89_22_pad_groupi_g4490(csa_tree_add_89_22_pad_groupi_n_1230 ,csa_tree_add_89_22_pad_groupi_n_1173 ,csa_tree_add_89_22_pad_groupi_n_1172);
  nor csa_tree_add_89_22_pad_groupi_g4491(csa_tree_add_89_22_pad_groupi_n_1229 ,csa_tree_add_89_22_pad_groupi_n_1152 ,csa_tree_add_89_22_pad_groupi_n_1175);
  or csa_tree_add_89_22_pad_groupi_g4492(csa_tree_add_89_22_pad_groupi_n_1228 ,csa_tree_add_89_22_pad_groupi_n_1173 ,csa_tree_add_89_22_pad_groupi_n_1172);
  and csa_tree_add_89_22_pad_groupi_g4493(csa_tree_add_89_22_pad_groupi_n_1227 ,csa_tree_add_89_22_pad_groupi_n_1161 ,csa_tree_add_89_22_pad_groupi_n_1168);
  or csa_tree_add_89_22_pad_groupi_g4494(csa_tree_add_89_22_pad_groupi_n_1226 ,csa_tree_add_89_22_pad_groupi_n_1161 ,csa_tree_add_89_22_pad_groupi_n_1168);
  or csa_tree_add_89_22_pad_groupi_g4495(csa_tree_add_89_22_pad_groupi_n_1225 ,csa_tree_add_89_22_pad_groupi_n_1162 ,csa_tree_add_89_22_pad_groupi_n_1165);
  nor csa_tree_add_89_22_pad_groupi_g4496(csa_tree_add_89_22_pad_groupi_n_1224 ,csa_tree_add_89_22_pad_groupi_n_1204 ,csa_tree_add_89_22_pad_groupi_n_1160);
  nor csa_tree_add_89_22_pad_groupi_g4497(csa_tree_add_89_22_pad_groupi_n_1223 ,csa_tree_add_89_22_pad_groupi_n_1163 ,csa_tree_add_89_22_pad_groupi_n_1166);
  xnor csa_tree_add_89_22_pad_groupi_g4498(csa_tree_add_89_22_pad_groupi_n_1222 ,csa_tree_add_89_22_pad_groupi_n_1035 ,csa_tree_add_89_22_pad_groupi_n_1094);
  xnor csa_tree_add_89_22_pad_groupi_g4499(csa_tree_add_89_22_pad_groupi_n_1221 ,csa_tree_add_89_22_pad_groupi_n_1100 ,csa_tree_add_89_22_pad_groupi_n_1074);
  xnor csa_tree_add_89_22_pad_groupi_g4500(csa_tree_add_89_22_pad_groupi_n_1220 ,csa_tree_add_89_22_pad_groupi_n_1072 ,csa_tree_add_89_22_pad_groupi_n_1090);
  xnor csa_tree_add_89_22_pad_groupi_g4501(csa_tree_add_89_22_pad_groupi_n_1219 ,csa_tree_add_89_22_pad_groupi_n_1016 ,csa_tree_add_89_22_pad_groupi_n_1097);
  xnor csa_tree_add_89_22_pad_groupi_g4502(csa_tree_add_89_22_pad_groupi_n_1218 ,csa_tree_add_89_22_pad_groupi_n_1056 ,csa_tree_add_89_22_pad_groupi_n_3);
  xnor csa_tree_add_89_22_pad_groupi_g4503(csa_tree_add_89_22_pad_groupi_n_1238 ,csa_tree_add_89_22_pad_groupi_n_1140 ,csa_tree_add_89_22_pad_groupi_n_1076);
  xnor csa_tree_add_89_22_pad_groupi_g4504(csa_tree_add_89_22_pad_groupi_n_1217 ,csa_tree_add_89_22_pad_groupi_n_1055 ,csa_tree_add_89_22_pad_groupi_n_1095);
  xnor csa_tree_add_89_22_pad_groupi_g4505(csa_tree_add_89_22_pad_groupi_n_1216 ,csa_tree_add_89_22_pad_groupi_n_1036 ,csa_tree_add_89_22_pad_groupi_n_1087);
  xnor csa_tree_add_89_22_pad_groupi_g4506(csa_tree_add_89_22_pad_groupi_n_1215 ,csa_tree_add_89_22_pad_groupi_n_1137 ,csa_tree_add_89_22_pad_groupi_n_1086);
  xnor csa_tree_add_89_22_pad_groupi_g4507(csa_tree_add_89_22_pad_groupi_n_1214 ,csa_tree_add_89_22_pad_groupi_n_1042 ,csa_tree_add_89_22_pad_groupi_n_1093);
  xnor csa_tree_add_89_22_pad_groupi_g4508(csa_tree_add_89_22_pad_groupi_n_1213 ,csa_tree_add_89_22_pad_groupi_n_1034 ,csa_tree_add_89_22_pad_groupi_n_1104);
  xnor csa_tree_add_89_22_pad_groupi_g4509(csa_tree_add_89_22_pad_groupi_n_1212 ,csa_tree_add_89_22_pad_groupi_n_1131 ,csa_tree_add_89_22_pad_groupi_n_1082);
  xnor csa_tree_add_89_22_pad_groupi_g4510(csa_tree_add_89_22_pad_groupi_n_1211 ,csa_tree_add_89_22_pad_groupi_n_1134 ,csa_tree_add_89_22_pad_groupi_n_1135);
  xnor csa_tree_add_89_22_pad_groupi_g4511(csa_tree_add_89_22_pad_groupi_n_1210 ,csa_tree_add_89_22_pad_groupi_n_1062 ,csa_tree_add_89_22_pad_groupi_n_1133);
  xnor csa_tree_add_89_22_pad_groupi_g4512(csa_tree_add_89_22_pad_groupi_n_1236 ,csa_tree_add_89_22_pad_groupi_n_1043 ,csa_tree_add_89_22_pad_groupi_n_1078);
  xnor csa_tree_add_89_22_pad_groupi_g4513(csa_tree_add_89_22_pad_groupi_n_1235 ,csa_tree_add_89_22_pad_groupi_n_1070 ,csa_tree_add_89_22_pad_groupi_n_1079);
  xnor csa_tree_add_89_22_pad_groupi_g4514(csa_tree_add_89_22_pad_groupi_n_1233 ,csa_tree_add_89_22_pad_groupi_n_976 ,csa_tree_add_89_22_pad_groupi_n_1077);
  not csa_tree_add_89_22_pad_groupi_g4515(csa_tree_add_89_22_pad_groupi_n_1206 ,csa_tree_add_89_22_pad_groupi_n_1205);
  not csa_tree_add_89_22_pad_groupi_g4516(csa_tree_add_89_22_pad_groupi_n_1204 ,csa_tree_add_89_22_pad_groupi_n_1203);
  not csa_tree_add_89_22_pad_groupi_g4517(csa_tree_add_89_22_pad_groupi_n_1202 ,csa_tree_add_89_22_pad_groupi_n_1201);
  and csa_tree_add_89_22_pad_groupi_g4518(csa_tree_add_89_22_pad_groupi_n_1200 ,csa_tree_add_89_22_pad_groupi_n_1035 ,csa_tree_add_89_22_pad_groupi_n_1094);
  or csa_tree_add_89_22_pad_groupi_g4519(csa_tree_add_89_22_pad_groupi_n_1199 ,csa_tree_add_89_22_pad_groupi_n_1105 ,csa_tree_add_89_22_pad_groupi_n_1128);
  nor csa_tree_add_89_22_pad_groupi_g4520(csa_tree_add_89_22_pad_groupi_n_1198 ,csa_tree_add_89_22_pad_groupi_n_1100 ,csa_tree_add_89_22_pad_groupi_n_1139);
  or csa_tree_add_89_22_pad_groupi_g4521(csa_tree_add_89_22_pad_groupi_n_1197 ,csa_tree_add_89_22_pad_groupi_n_1136 ,csa_tree_add_89_22_pad_groupi_n_1086);
  and csa_tree_add_89_22_pad_groupi_g4522(csa_tree_add_89_22_pad_groupi_n_1196 ,csa_tree_add_89_22_pad_groupi_n_1118 ,csa_tree_add_89_22_pad_groupi_n_1103);
  and csa_tree_add_89_22_pad_groupi_g4523(csa_tree_add_89_22_pad_groupi_n_1195 ,csa_tree_add_89_22_pad_groupi_n_1100 ,csa_tree_add_89_22_pad_groupi_n_1139);
  or csa_tree_add_89_22_pad_groupi_g4524(csa_tree_add_89_22_pad_groupi_n_1194 ,csa_tree_add_89_22_pad_groupi_n_1055 ,csa_tree_add_89_22_pad_groupi_n_1095);
  nor csa_tree_add_89_22_pad_groupi_g4525(csa_tree_add_89_22_pad_groupi_n_1193 ,csa_tree_add_89_22_pad_groupi_n_1137 ,csa_tree_add_89_22_pad_groupi_n_1085);
  or csa_tree_add_89_22_pad_groupi_g4526(csa_tree_add_89_22_pad_groupi_n_1192 ,csa_tree_add_89_22_pad_groupi_n_1083 ,csa_tree_add_89_22_pad_groupi_n_1089);
  nor csa_tree_add_89_22_pad_groupi_g4527(csa_tree_add_89_22_pad_groupi_n_1191 ,csa_tree_add_89_22_pad_groupi_n_1022 ,csa_tree_add_89_22_pad_groupi_n_1109);
  nor csa_tree_add_89_22_pad_groupi_g4528(csa_tree_add_89_22_pad_groupi_n_1190 ,csa_tree_add_89_22_pad_groupi_n_1084 ,csa_tree_add_89_22_pad_groupi_n_1090);
  or csa_tree_add_89_22_pad_groupi_g4529(csa_tree_add_89_22_pad_groupi_n_1189 ,csa_tree_add_89_22_pad_groupi_n_1056 ,csa_tree_add_89_22_pad_groupi_n_3);
  nor csa_tree_add_89_22_pad_groupi_g4530(csa_tree_add_89_22_pad_groupi_n_1188 ,csa_tree_add_89_22_pad_groupi_n_1019 ,csa_tree_add_89_22_pad_groupi_n_1080);
  and csa_tree_add_89_22_pad_groupi_g4531(csa_tree_add_89_22_pad_groupi_n_1187 ,csa_tree_add_89_22_pad_groupi_n_1056 ,csa_tree_add_89_22_pad_groupi_n_3);
  and csa_tree_add_89_22_pad_groupi_g4532(csa_tree_add_89_22_pad_groupi_n_1186 ,csa_tree_add_89_22_pad_groupi_n_1019 ,csa_tree_add_89_22_pad_groupi_n_1080);
  and csa_tree_add_89_22_pad_groupi_g4533(csa_tree_add_89_22_pad_groupi_n_1185 ,csa_tree_add_89_22_pad_groupi_n_1134 ,csa_tree_add_89_22_pad_groupi_n_1135);
  nor csa_tree_add_89_22_pad_groupi_g4534(csa_tree_add_89_22_pad_groupi_n_1184 ,csa_tree_add_89_22_pad_groupi_n_1134 ,csa_tree_add_89_22_pad_groupi_n_1135);
  and csa_tree_add_89_22_pad_groupi_g4535(csa_tree_add_89_22_pad_groupi_n_1183 ,csa_tree_add_89_22_pad_groupi_n_1062 ,csa_tree_add_89_22_pad_groupi_n_1133);
  and csa_tree_add_89_22_pad_groupi_g4536(csa_tree_add_89_22_pad_groupi_n_1182 ,csa_tree_add_89_22_pad_groupi_n_1120 ,csa_tree_add_89_22_pad_groupi_n_1106);
  or csa_tree_add_89_22_pad_groupi_g4537(csa_tree_add_89_22_pad_groupi_n_1181 ,csa_tree_add_89_22_pad_groupi_n_1062 ,csa_tree_add_89_22_pad_groupi_n_1133);
  and csa_tree_add_89_22_pad_groupi_g4538(csa_tree_add_89_22_pad_groupi_n_1180 ,csa_tree_add_89_22_pad_groupi_n_1050 ,csa_tree_add_89_22_pad_groupi_n_1140);
  and csa_tree_add_89_22_pad_groupi_g4539(csa_tree_add_89_22_pad_groupi_n_1179 ,csa_tree_add_89_22_pad_groupi_n_1055 ,csa_tree_add_89_22_pad_groupi_n_1095);
  nor csa_tree_add_89_22_pad_groupi_g4540(csa_tree_add_89_22_pad_groupi_n_1178 ,csa_tree_add_89_22_pad_groupi_n_1023 ,csa_tree_add_89_22_pad_groupi_n_1108);
  nor csa_tree_add_89_22_pad_groupi_g4541(csa_tree_add_89_22_pad_groupi_n_1177 ,csa_tree_add_89_22_pad_groupi_n_1031 ,csa_tree_add_89_22_pad_groupi_n_1119);
  and csa_tree_add_89_22_pad_groupi_g4542(csa_tree_add_89_22_pad_groupi_n_1209 ,csa_tree_add_89_22_pad_groupi_n_1054 ,csa_tree_add_89_22_pad_groupi_n_1127);
  or csa_tree_add_89_22_pad_groupi_g4543(csa_tree_add_89_22_pad_groupi_n_1208 ,csa_tree_add_89_22_pad_groupi_n_901 ,csa_tree_add_89_22_pad_groupi_n_1122);
  or csa_tree_add_89_22_pad_groupi_g4544(csa_tree_add_89_22_pad_groupi_n_1207 ,csa_tree_add_89_22_pad_groupi_n_914 ,csa_tree_add_89_22_pad_groupi_n_1125);
  and csa_tree_add_89_22_pad_groupi_g4545(csa_tree_add_89_22_pad_groupi_n_1205 ,csa_tree_add_89_22_pad_groupi_n_884 ,csa_tree_add_89_22_pad_groupi_n_1116);
  and csa_tree_add_89_22_pad_groupi_g4546(csa_tree_add_89_22_pad_groupi_n_1203 ,csa_tree_add_89_22_pad_groupi_n_921 ,csa_tree_add_89_22_pad_groupi_n_1126);
  or csa_tree_add_89_22_pad_groupi_g4547(csa_tree_add_89_22_pad_groupi_n_1201 ,csa_tree_add_89_22_pad_groupi_n_1049 ,csa_tree_add_89_22_pad_groupi_n_1117);
  not csa_tree_add_89_22_pad_groupi_g4548(csa_tree_add_89_22_pad_groupi_n_1170 ,csa_tree_add_89_22_pad_groupi_n_1171);
  not csa_tree_add_89_22_pad_groupi_g4549(csa_tree_add_89_22_pad_groupi_n_1166 ,csa_tree_add_89_22_pad_groupi_n_1165);
  not csa_tree_add_89_22_pad_groupi_g4550(csa_tree_add_89_22_pad_groupi_n_1163 ,csa_tree_add_89_22_pad_groupi_n_1162);
  not csa_tree_add_89_22_pad_groupi_g4551(csa_tree_add_89_22_pad_groupi_n_1160 ,csa_tree_add_89_22_pad_groupi_n_1159);
  or csa_tree_add_89_22_pad_groupi_g4552(csa_tree_add_89_22_pad_groupi_n_1158 ,csa_tree_add_89_22_pad_groupi_n_1035 ,csa_tree_add_89_22_pad_groupi_n_1094);
  and csa_tree_add_89_22_pad_groupi_g4553(csa_tree_add_89_22_pad_groupi_n_1157 ,csa_tree_add_89_22_pad_groupi_n_1015 ,csa_tree_add_89_22_pad_groupi_n_1097);
  or csa_tree_add_89_22_pad_groupi_g4554(csa_tree_add_89_22_pad_groupi_n_1156 ,csa_tree_add_89_22_pad_groupi_n_1130 ,csa_tree_add_89_22_pad_groupi_n_1081);
  or csa_tree_add_89_22_pad_groupi_g4555(csa_tree_add_89_22_pad_groupi_n_1155 ,csa_tree_add_89_22_pad_groupi_n_1033 ,csa_tree_add_89_22_pad_groupi_n_1091);
  and csa_tree_add_89_22_pad_groupi_g4556(csa_tree_add_89_22_pad_groupi_n_1154 ,csa_tree_add_89_22_pad_groupi_n_1093 ,csa_tree_add_89_22_pad_groupi_n_1088);
  nor csa_tree_add_89_22_pad_groupi_g4557(csa_tree_add_89_22_pad_groupi_n_1153 ,csa_tree_add_89_22_pad_groupi_n_1093 ,csa_tree_add_89_22_pad_groupi_n_1088);
  and csa_tree_add_89_22_pad_groupi_g4558(csa_tree_add_89_22_pad_groupi_n_1152 ,csa_tree_add_89_22_pad_groupi_n_1016 ,csa_tree_add_89_22_pad_groupi_n_1096);
  nor csa_tree_add_89_22_pad_groupi_g4559(csa_tree_add_89_22_pad_groupi_n_1151 ,csa_tree_add_89_22_pad_groupi_n_1034 ,csa_tree_add_89_22_pad_groupi_n_1092);
  nor csa_tree_add_89_22_pad_groupi_g4560(csa_tree_add_89_22_pad_groupi_n_1150 ,csa_tree_add_89_22_pad_groupi_n_1131 ,csa_tree_add_89_22_pad_groupi_n_1082);
  or csa_tree_add_89_22_pad_groupi_g4561(csa_tree_add_89_22_pad_groupi_n_1149 ,csa_tree_add_89_22_pad_groupi_n_1110 ,csa_tree_add_89_22_pad_groupi_n_1101);
  and csa_tree_add_89_22_pad_groupi_g4562(csa_tree_add_89_22_pad_groupi_n_1148 ,csa_tree_add_89_22_pad_groupi_n_1037 ,csa_tree_add_89_22_pad_groupi_n_1087);
  nor csa_tree_add_89_22_pad_groupi_g4563(csa_tree_add_89_22_pad_groupi_n_1147 ,csa_tree_add_89_22_pad_groupi_n_1037 ,csa_tree_add_89_22_pad_groupi_n_1087);
  xnor csa_tree_add_89_22_pad_groupi_g4564(csa_tree_add_89_22_pad_groupi_n_1146 ,csa_tree_add_89_22_pad_groupi_n_1010 ,csa_tree_add_89_22_pad_groupi_n_1064);
  xnor csa_tree_add_89_22_pad_groupi_g4565(csa_tree_add_89_22_pad_groupi_n_1145 ,csa_tree_add_89_22_pad_groupi_n_1067 ,csa_tree_add_89_22_pad_groupi_n_1019);
  xnor csa_tree_add_89_22_pad_groupi_g4566(csa_tree_add_89_22_pad_groupi_n_1144 ,csa_tree_add_89_22_pad_groupi_n_1058 ,csa_tree_add_89_22_pad_groupi_n_1061);
  xnor csa_tree_add_89_22_pad_groupi_g4567(csa_tree_add_89_22_pad_groupi_n_1143 ,csa_tree_add_89_22_pad_groupi_n_1011 ,csa_tree_add_89_22_pad_groupi_n_1059);
  xnor csa_tree_add_89_22_pad_groupi_g4568(csa_tree_add_89_22_pad_groupi_n_1142 ,csa_tree_add_89_22_pad_groupi_n_1018 ,csa_tree_add_89_22_pad_groupi_n_1066);
  xnor csa_tree_add_89_22_pad_groupi_g4569(csa_tree_add_89_22_pad_groupi_n_1176 ,csa_tree_add_89_22_pad_groupi_n_1020 ,csa_tree_add_89_22_pad_groupi_n_1025);
  and csa_tree_add_89_22_pad_groupi_g4570(csa_tree_add_89_22_pad_groupi_n_1175 ,csa_tree_add_89_22_pad_groupi_n_1030 ,csa_tree_add_89_22_pad_groupi_n_1111);
  xnor csa_tree_add_89_22_pad_groupi_g4571(csa_tree_add_89_22_pad_groupi_n_1174 ,csa_tree_add_89_22_pad_groupi_n_1068 ,csa_tree_add_89_22_pad_groupi_n_950);
  or csa_tree_add_89_22_pad_groupi_g4572(csa_tree_add_89_22_pad_groupi_n_1173 ,csa_tree_add_89_22_pad_groupi_n_908 ,csa_tree_add_89_22_pad_groupi_n_1121);
  xnor csa_tree_add_89_22_pad_groupi_g4573(csa_tree_add_89_22_pad_groupi_n_1172 ,csa_tree_add_89_22_pad_groupi_n_1045 ,csa_tree_add_89_22_pad_groupi_n_944);
  xnor csa_tree_add_89_22_pad_groupi_g4574(csa_tree_add_89_22_pad_groupi_n_1171 ,csa_tree_add_89_22_pad_groupi_n_1073 ,csa_tree_add_89_22_pad_groupi_n_941);
  xnor csa_tree_add_89_22_pad_groupi_g4575(csa_tree_add_89_22_pad_groupi_n_1169 ,csa_tree_add_89_22_pad_groupi_n_1041 ,csa_tree_add_89_22_pad_groupi_n_974);
  xnor csa_tree_add_89_22_pad_groupi_g4576(csa_tree_add_89_22_pad_groupi_n_1168 ,csa_tree_add_89_22_pad_groupi_n_1044 ,csa_tree_add_89_22_pad_groupi_n_939);
  xnor csa_tree_add_89_22_pad_groupi_g4577(csa_tree_add_89_22_pad_groupi_n_1167 ,csa_tree_add_89_22_pad_groupi_n_1040 ,csa_tree_add_89_22_pad_groupi_n_969);
  xnor csa_tree_add_89_22_pad_groupi_g4578(csa_tree_add_89_22_pad_groupi_n_1165 ,csa_tree_add_89_22_pad_groupi_n_1038 ,csa_tree_add_89_22_pad_groupi_n_970);
  or csa_tree_add_89_22_pad_groupi_g4579(csa_tree_add_89_22_pad_groupi_n_1164 ,csa_tree_add_89_22_pad_groupi_n_858 ,csa_tree_add_89_22_pad_groupi_n_1113);
  and csa_tree_add_89_22_pad_groupi_g4580(csa_tree_add_89_22_pad_groupi_n_1162 ,csa_tree_add_89_22_pad_groupi_n_857 ,csa_tree_add_89_22_pad_groupi_n_1112);
  or csa_tree_add_89_22_pad_groupi_g4581(csa_tree_add_89_22_pad_groupi_n_1161 ,csa_tree_add_89_22_pad_groupi_n_873 ,csa_tree_add_89_22_pad_groupi_n_1129);
  xnor csa_tree_add_89_22_pad_groupi_g4582(csa_tree_add_89_22_pad_groupi_n_1159 ,csa_tree_add_89_22_pad_groupi_n_1046 ,csa_tree_add_89_22_pad_groupi_n_955);
  not csa_tree_add_89_22_pad_groupi_g4583(csa_tree_add_89_22_pad_groupi_n_1139 ,csa_tree_add_89_22_pad_groupi_n_1138);
  not csa_tree_add_89_22_pad_groupi_g4584(csa_tree_add_89_22_pad_groupi_n_1136 ,csa_tree_add_89_22_pad_groupi_n_1137);
  not csa_tree_add_89_22_pad_groupi_g4585(csa_tree_add_89_22_pad_groupi_n_1130 ,csa_tree_add_89_22_pad_groupi_n_1131);
  and csa_tree_add_89_22_pad_groupi_g4586(csa_tree_add_89_22_pad_groupi_n_1129 ,csa_tree_add_89_22_pad_groupi_n_871 ,csa_tree_add_89_22_pad_groupi_n_1040);
  nor csa_tree_add_89_22_pad_groupi_g4587(csa_tree_add_89_22_pad_groupi_n_1128 ,csa_tree_add_89_22_pad_groupi_n_1058 ,csa_tree_add_89_22_pad_groupi_n_1061);
  or csa_tree_add_89_22_pad_groupi_g4588(csa_tree_add_89_22_pad_groupi_n_1127 ,csa_tree_add_89_22_pad_groupi_n_1053 ,csa_tree_add_89_22_pad_groupi_n_1071);
  or csa_tree_add_89_22_pad_groupi_g4589(csa_tree_add_89_22_pad_groupi_n_1126 ,csa_tree_add_89_22_pad_groupi_n_918 ,csa_tree_add_89_22_pad_groupi_n_1069);
  and csa_tree_add_89_22_pad_groupi_g4590(csa_tree_add_89_22_pad_groupi_n_1125 ,csa_tree_add_89_22_pad_groupi_n_932 ,csa_tree_add_89_22_pad_groupi_n_1073);
  nor csa_tree_add_89_22_pad_groupi_g4591(csa_tree_add_89_22_pad_groupi_n_1124 ,csa_tree_add_89_22_pad_groupi_n_1010 ,csa_tree_add_89_22_pad_groupi_n_1063);
  and csa_tree_add_89_22_pad_groupi_g4592(csa_tree_add_89_22_pad_groupi_n_1123 ,csa_tree_add_89_22_pad_groupi_n_1011 ,csa_tree_add_89_22_pad_groupi_n_1059);
  and csa_tree_add_89_22_pad_groupi_g4593(csa_tree_add_89_22_pad_groupi_n_1122 ,csa_tree_add_89_22_pad_groupi_n_880 ,csa_tree_add_89_22_pad_groupi_n_1045);
  and csa_tree_add_89_22_pad_groupi_g4594(csa_tree_add_89_22_pad_groupi_n_1121 ,csa_tree_add_89_22_pad_groupi_n_867 ,csa_tree_add_89_22_pad_groupi_n_1044);
  or csa_tree_add_89_22_pad_groupi_g4595(csa_tree_add_89_22_pad_groupi_n_1120 ,csa_tree_add_89_22_pad_groupi_n_1011 ,csa_tree_add_89_22_pad_groupi_n_1059);
  nor csa_tree_add_89_22_pad_groupi_g4596(csa_tree_add_89_22_pad_groupi_n_1119 ,csa_tree_add_89_22_pad_groupi_n_1026 ,csa_tree_add_89_22_pad_groupi_n_980);
  or csa_tree_add_89_22_pad_groupi_g4597(csa_tree_add_89_22_pad_groupi_n_1118 ,csa_tree_add_89_22_pad_groupi_n_1009 ,csa_tree_add_89_22_pad_groupi_n_1064);
  and csa_tree_add_89_22_pad_groupi_g4598(csa_tree_add_89_22_pad_groupi_n_1117 ,csa_tree_add_89_22_pad_groupi_n_1029 ,csa_tree_add_89_22_pad_groupi_n_1043);
  or csa_tree_add_89_22_pad_groupi_g4599(csa_tree_add_89_22_pad_groupi_n_1116 ,csa_tree_add_89_22_pad_groupi_n_882 ,csa_tree_add_89_22_pad_groupi_n_1038);
  or csa_tree_add_89_22_pad_groupi_g4600(csa_tree_add_89_22_pad_groupi_n_1115 ,csa_tree_add_89_22_pad_groupi_n_1057 ,csa_tree_add_89_22_pad_groupi_n_1060);
  or csa_tree_add_89_22_pad_groupi_g4601(csa_tree_add_89_22_pad_groupi_n_1114 ,csa_tree_add_89_22_pad_groupi_n_1017 ,csa_tree_add_89_22_pad_groupi_n_1065);
  and csa_tree_add_89_22_pad_groupi_g4602(csa_tree_add_89_22_pad_groupi_n_1113 ,csa_tree_add_89_22_pad_groupi_n_860 ,csa_tree_add_89_22_pad_groupi_n_1041);
  or csa_tree_add_89_22_pad_groupi_g4603(csa_tree_add_89_22_pad_groupi_n_1112 ,csa_tree_add_89_22_pad_groupi_n_854 ,csa_tree_add_89_22_pad_groupi_n_1046);
  or csa_tree_add_89_22_pad_groupi_g4604(csa_tree_add_89_22_pad_groupi_n_1111 ,csa_tree_add_89_22_pad_groupi_n_1028 ,csa_tree_add_89_22_pad_groupi_n_976);
  nor csa_tree_add_89_22_pad_groupi_g4605(csa_tree_add_89_22_pad_groupi_n_1110 ,csa_tree_add_89_22_pad_groupi_n_1018 ,csa_tree_add_89_22_pad_groupi_n_1066);
  xnor csa_tree_add_89_22_pad_groupi_g4606(csa_tree_add_89_22_pad_groupi_n_1141 ,csa_tree_add_89_22_pad_groupi_n_842 ,csa_tree_add_89_22_pad_groupi_n_951);
  xnor csa_tree_add_89_22_pad_groupi_g4607(csa_tree_add_89_22_pad_groupi_n_1140 ,csa_tree_add_89_22_pad_groupi_n_803 ,csa_tree_add_89_22_pad_groupi_n_964);
  xnor csa_tree_add_89_22_pad_groupi_g4608(csa_tree_add_89_22_pad_groupi_n_1138 ,csa_tree_add_89_22_pad_groupi_n_773 ,csa_tree_add_89_22_pad_groupi_n_962);
  xnor csa_tree_add_89_22_pad_groupi_g4609(csa_tree_add_89_22_pad_groupi_n_1137 ,csa_tree_add_89_22_pad_groupi_n_783 ,csa_tree_add_89_22_pad_groupi_n_960);
  xnor csa_tree_add_89_22_pad_groupi_g4610(csa_tree_add_89_22_pad_groupi_n_1135 ,csa_tree_add_89_22_pad_groupi_n_840 ,csa_tree_add_89_22_pad_groupi_n_965);
  or csa_tree_add_89_22_pad_groupi_g4611(csa_tree_add_89_22_pad_groupi_n_1134 ,csa_tree_add_89_22_pad_groupi_n_1000 ,csa_tree_add_89_22_pad_groupi_n_1052);
  xnor csa_tree_add_89_22_pad_groupi_g4612(csa_tree_add_89_22_pad_groupi_n_1133 ,csa_tree_add_89_22_pad_groupi_n_778 ,csa_tree_add_89_22_pad_groupi_n_949);
  and csa_tree_add_89_22_pad_groupi_g4613(csa_tree_add_89_22_pad_groupi_n_1132 ,csa_tree_add_89_22_pad_groupi_n_888 ,csa_tree_add_89_22_pad_groupi_n_1032);
  or csa_tree_add_89_22_pad_groupi_g4614(csa_tree_add_89_22_pad_groupi_n_1131 ,csa_tree_add_89_22_pad_groupi_n_868 ,csa_tree_add_89_22_pad_groupi_n_1027);
  not csa_tree_add_89_22_pad_groupi_g4615(csa_tree_add_89_22_pad_groupi_n_1109 ,csa_tree_add_89_22_pad_groupi_n_1108);
  not csa_tree_add_89_22_pad_groupi_g4616(csa_tree_add_89_22_pad_groupi_n_1097 ,csa_tree_add_89_22_pad_groupi_n_1096);
  not csa_tree_add_89_22_pad_groupi_g4617(csa_tree_add_89_22_pad_groupi_n_1091 ,csa_tree_add_89_22_pad_groupi_n_1092);
  not csa_tree_add_89_22_pad_groupi_g4618(csa_tree_add_89_22_pad_groupi_n_1090 ,csa_tree_add_89_22_pad_groupi_n_1089);
  not csa_tree_add_89_22_pad_groupi_g4619(csa_tree_add_89_22_pad_groupi_n_1085 ,csa_tree_add_89_22_pad_groupi_n_1086);
  not csa_tree_add_89_22_pad_groupi_g4620(csa_tree_add_89_22_pad_groupi_n_1083 ,csa_tree_add_89_22_pad_groupi_n_1084);
  not csa_tree_add_89_22_pad_groupi_g4621(csa_tree_add_89_22_pad_groupi_n_1081 ,csa_tree_add_89_22_pad_groupi_n_1082);
  xnor csa_tree_add_89_22_pad_groupi_g4622(csa_tree_add_89_22_pad_groupi_n_1079 ,csa_tree_add_89_22_pad_groupi_n_975 ,csa_tree_add_89_22_pad_groupi_n_934);
  xnor csa_tree_add_89_22_pad_groupi_g4623(csa_tree_add_89_22_pad_groupi_n_1108 ,csa_tree_add_89_22_pad_groupi_n_892 ,csa_tree_add_89_22_pad_groupi_n_961);
  xnor csa_tree_add_89_22_pad_groupi_g4624(csa_tree_add_89_22_pad_groupi_n_1078 ,csa_tree_add_89_22_pad_groupi_n_797 ,csa_tree_add_89_22_pad_groupi_n_4);
  xnor csa_tree_add_89_22_pad_groupi_g4625(csa_tree_add_89_22_pad_groupi_n_1077 ,csa_tree_add_89_22_pad_groupi_n_746 ,csa_tree_add_89_22_pad_groupi_n_1014);
  xnor csa_tree_add_89_22_pad_groupi_g4626(csa_tree_add_89_22_pad_groupi_n_1076 ,csa_tree_add_89_22_pad_groupi_n_1012 ,csa_tree_add_89_22_pad_groupi_n_933);
  xnor csa_tree_add_89_22_pad_groupi_g4627(csa_tree_add_89_22_pad_groupi_n_1075 ,csa_tree_add_89_22_pad_groupi_n_2 ,csa_tree_add_89_22_pad_groupi_n_978);
  xnor csa_tree_add_89_22_pad_groupi_g4628(csa_tree_add_89_22_pad_groupi_n_1107 ,csa_tree_add_89_22_pad_groupi_n_768 ,csa_tree_add_89_22_pad_groupi_n_942);
  xnor csa_tree_add_89_22_pad_groupi_g4629(csa_tree_add_89_22_pad_groupi_n_1106 ,csa_tree_add_89_22_pad_groupi_n_764 ,csa_tree_add_89_22_pad_groupi_n_968);
  xnor csa_tree_add_89_22_pad_groupi_g4630(csa_tree_add_89_22_pad_groupi_n_1105 ,csa_tree_add_89_22_pad_groupi_n_740 ,csa_tree_add_89_22_pad_groupi_n_963);
  xnor csa_tree_add_89_22_pad_groupi_g4631(csa_tree_add_89_22_pad_groupi_n_1104 ,csa_tree_add_89_22_pad_groupi_n_782 ,csa_tree_add_89_22_pad_groupi_n_967);
  xnor csa_tree_add_89_22_pad_groupi_g4632(csa_tree_add_89_22_pad_groupi_n_1103 ,csa_tree_add_89_22_pad_groupi_n_1021 ,csa_tree_add_89_22_pad_groupi_n_957);
  xnor csa_tree_add_89_22_pad_groupi_g4633(csa_tree_add_89_22_pad_groupi_n_1102 ,csa_tree_add_89_22_pad_groupi_n_769 ,csa_tree_add_89_22_pad_groupi_n_945);
  xnor csa_tree_add_89_22_pad_groupi_g4634(csa_tree_add_89_22_pad_groupi_n_1101 ,csa_tree_add_89_22_pad_groupi_n_977 ,csa_tree_add_89_22_pad_groupi_n_966);
  xnor csa_tree_add_89_22_pad_groupi_g4635(csa_tree_add_89_22_pad_groupi_n_1100 ,csa_tree_add_89_22_pad_groupi_n_838 ,csa_tree_add_89_22_pad_groupi_n_946);
  xnor csa_tree_add_89_22_pad_groupi_g4637(csa_tree_add_89_22_pad_groupi_n_1099 ,csa_tree_add_89_22_pad_groupi_n_750 ,csa_tree_add_89_22_pad_groupi_n_952);
  xnor csa_tree_add_89_22_pad_groupi_g4638(csa_tree_add_89_22_pad_groupi_n_1098 ,csa_tree_add_89_22_pad_groupi_n_743 ,csa_tree_add_89_22_pad_groupi_n_972);
  xnor csa_tree_add_89_22_pad_groupi_g4639(csa_tree_add_89_22_pad_groupi_n_1096 ,csa_tree_add_89_22_pad_groupi_n_971 ,csa_tree_add_89_22_pad_groupi_n_578);
  xnor csa_tree_add_89_22_pad_groupi_g4640(csa_tree_add_89_22_pad_groupi_n_1095 ,csa_tree_add_89_22_pad_groupi_n_770 ,csa_tree_add_89_22_pad_groupi_n_947);
  xnor csa_tree_add_89_22_pad_groupi_g4641(csa_tree_add_89_22_pad_groupi_n_1094 ,csa_tree_add_89_22_pad_groupi_n_830 ,csa_tree_add_89_22_pad_groupi_n_943);
  xnor csa_tree_add_89_22_pad_groupi_g4642(csa_tree_add_89_22_pad_groupi_n_1093 ,csa_tree_add_89_22_pad_groupi_n_780 ,csa_tree_add_89_22_pad_groupi_n_938);
  xnor csa_tree_add_89_22_pad_groupi_g4643(csa_tree_add_89_22_pad_groupi_n_1092 ,csa_tree_add_89_22_pad_groupi_n_775 ,csa_tree_add_89_22_pad_groupi_n_937);
  xnor csa_tree_add_89_22_pad_groupi_g4644(csa_tree_add_89_22_pad_groupi_n_1089 ,csa_tree_add_89_22_pad_groupi_n_827 ,csa_tree_add_89_22_pad_groupi_n_973);
  xnor csa_tree_add_89_22_pad_groupi_g4645(csa_tree_add_89_22_pad_groupi_n_1088 ,csa_tree_add_89_22_pad_groupi_n_777 ,csa_tree_add_89_22_pad_groupi_n_940);
  xnor csa_tree_add_89_22_pad_groupi_g4646(csa_tree_add_89_22_pad_groupi_n_1087 ,csa_tree_add_89_22_pad_groupi_n_774 ,csa_tree_add_89_22_pad_groupi_n_954);
  xnor csa_tree_add_89_22_pad_groupi_g4647(csa_tree_add_89_22_pad_groupi_n_1086 ,csa_tree_add_89_22_pad_groupi_n_893 ,csa_tree_add_89_22_pad_groupi_n_959);
  xnor csa_tree_add_89_22_pad_groupi_g4648(csa_tree_add_89_22_pad_groupi_n_1084 ,csa_tree_add_89_22_pad_groupi_n_785 ,csa_tree_add_89_22_pad_groupi_n_956);
  xnor csa_tree_add_89_22_pad_groupi_g4649(csa_tree_add_89_22_pad_groupi_n_1082 ,csa_tree_add_89_22_pad_groupi_n_839 ,csa_tree_add_89_22_pad_groupi_n_958);
  xnor csa_tree_add_89_22_pad_groupi_g4650(csa_tree_add_89_22_pad_groupi_n_1080 ,csa_tree_add_89_22_pad_groupi_n_936 ,csa_tree_add_89_22_pad_groupi_n_953);
  not csa_tree_add_89_22_pad_groupi_g4651(csa_tree_add_89_22_pad_groupi_n_1071 ,csa_tree_add_89_22_pad_groupi_n_1070);
  not csa_tree_add_89_22_pad_groupi_g4652(csa_tree_add_89_22_pad_groupi_n_1069 ,csa_tree_add_89_22_pad_groupi_n_1068);
  not csa_tree_add_89_22_pad_groupi_g4653(csa_tree_add_89_22_pad_groupi_n_1065 ,csa_tree_add_89_22_pad_groupi_n_1066);
  not csa_tree_add_89_22_pad_groupi_g4654(csa_tree_add_89_22_pad_groupi_n_1063 ,csa_tree_add_89_22_pad_groupi_n_1064);
  not csa_tree_add_89_22_pad_groupi_g4655(csa_tree_add_89_22_pad_groupi_n_1060 ,csa_tree_add_89_22_pad_groupi_n_1061);
  not csa_tree_add_89_22_pad_groupi_g4656(csa_tree_add_89_22_pad_groupi_n_1057 ,csa_tree_add_89_22_pad_groupi_n_1058);
  or csa_tree_add_89_22_pad_groupi_g4657(csa_tree_add_89_22_pad_groupi_n_1054 ,csa_tree_add_89_22_pad_groupi_n_276 ,csa_tree_add_89_22_pad_groupi_n_975);
  and csa_tree_add_89_22_pad_groupi_g4658(csa_tree_add_89_22_pad_groupi_n_1053 ,csa_tree_add_89_22_pad_groupi_n_934 ,csa_tree_add_89_22_pad_groupi_n_975);
  and csa_tree_add_89_22_pad_groupi_g4659(csa_tree_add_89_22_pad_groupi_n_1052 ,csa_tree_add_89_22_pad_groupi_n_998 ,csa_tree_add_89_22_pad_groupi_n_1020);
  and csa_tree_add_89_22_pad_groupi_g4660(csa_tree_add_89_22_pad_groupi_n_1051 ,csa_tree_add_89_22_pad_groupi_n_933 ,csa_tree_add_89_22_pad_groupi_n_1012);
  or csa_tree_add_89_22_pad_groupi_g4661(csa_tree_add_89_22_pad_groupi_n_1050 ,csa_tree_add_89_22_pad_groupi_n_933 ,csa_tree_add_89_22_pad_groupi_n_1012);
  and csa_tree_add_89_22_pad_groupi_g4662(csa_tree_add_89_22_pad_groupi_n_1049 ,csa_tree_add_89_22_pad_groupi_n_797 ,csa_tree_add_89_22_pad_groupi_n_4);
  and csa_tree_add_89_22_pad_groupi_g4663(csa_tree_add_89_22_pad_groupi_n_1074 ,csa_tree_add_89_22_pad_groupi_n_913 ,csa_tree_add_89_22_pad_groupi_n_1007);
  or csa_tree_add_89_22_pad_groupi_g4664(csa_tree_add_89_22_pad_groupi_n_1073 ,csa_tree_add_89_22_pad_groupi_n_910 ,csa_tree_add_89_22_pad_groupi_n_999);
  and csa_tree_add_89_22_pad_groupi_g4665(csa_tree_add_89_22_pad_groupi_n_1072 ,csa_tree_add_89_22_pad_groupi_n_915 ,csa_tree_add_89_22_pad_groupi_n_996);
  or csa_tree_add_89_22_pad_groupi_g4666(csa_tree_add_89_22_pad_groupi_n_1070 ,csa_tree_add_89_22_pad_groupi_n_890 ,csa_tree_add_89_22_pad_groupi_n_1005);
  or csa_tree_add_89_22_pad_groupi_g4667(csa_tree_add_89_22_pad_groupi_n_1068 ,csa_tree_add_89_22_pad_groupi_n_905 ,csa_tree_add_89_22_pad_groupi_n_1003);
  and csa_tree_add_89_22_pad_groupi_g4668(csa_tree_add_89_22_pad_groupi_n_1067 ,csa_tree_add_89_22_pad_groupi_n_912 ,csa_tree_add_89_22_pad_groupi_n_1002);
  or csa_tree_add_89_22_pad_groupi_g4669(csa_tree_add_89_22_pad_groupi_n_1066 ,csa_tree_add_89_22_pad_groupi_n_903 ,csa_tree_add_89_22_pad_groupi_n_1004);
  or csa_tree_add_89_22_pad_groupi_g4670(csa_tree_add_89_22_pad_groupi_n_1064 ,csa_tree_add_89_22_pad_groupi_n_925 ,csa_tree_add_89_22_pad_groupi_n_1006);
  or csa_tree_add_89_22_pad_groupi_g4671(csa_tree_add_89_22_pad_groupi_n_1062 ,csa_tree_add_89_22_pad_groupi_n_874 ,csa_tree_add_89_22_pad_groupi_n_987);
  or csa_tree_add_89_22_pad_groupi_g4672(csa_tree_add_89_22_pad_groupi_n_1061 ,csa_tree_add_89_22_pad_groupi_n_929 ,csa_tree_add_89_22_pad_groupi_n_979);
  or csa_tree_add_89_22_pad_groupi_g4673(csa_tree_add_89_22_pad_groupi_n_1059 ,csa_tree_add_89_22_pad_groupi_n_889 ,csa_tree_add_89_22_pad_groupi_n_995);
  or csa_tree_add_89_22_pad_groupi_g4674(csa_tree_add_89_22_pad_groupi_n_1058 ,csa_tree_add_89_22_pad_groupi_n_911 ,csa_tree_add_89_22_pad_groupi_n_1008);
  or csa_tree_add_89_22_pad_groupi_g4675(csa_tree_add_89_22_pad_groupi_n_1056 ,csa_tree_add_89_22_pad_groupi_n_869 ,csa_tree_add_89_22_pad_groupi_n_1001);
  or csa_tree_add_89_22_pad_groupi_g4676(csa_tree_add_89_22_pad_groupi_n_1055 ,csa_tree_add_89_22_pad_groupi_n_886 ,csa_tree_add_89_22_pad_groupi_n_993);
  not csa_tree_add_89_22_pad_groupi_g4677(csa_tree_add_89_22_pad_groupi_n_1048 ,csa_tree_add_89_22_pad_groupi_n_1047);
  not csa_tree_add_89_22_pad_groupi_g4678(csa_tree_add_89_22_pad_groupi_n_1037 ,csa_tree_add_89_22_pad_groupi_n_1036);
  not csa_tree_add_89_22_pad_groupi_g4679(csa_tree_add_89_22_pad_groupi_n_1033 ,csa_tree_add_89_22_pad_groupi_n_1034);
  or csa_tree_add_89_22_pad_groupi_g4680(csa_tree_add_89_22_pad_groupi_n_1032 ,csa_tree_add_89_22_pad_groupi_n_876 ,csa_tree_add_89_22_pad_groupi_n_977);
  nor csa_tree_add_89_22_pad_groupi_g4681(csa_tree_add_89_22_pad_groupi_n_1031 ,csa_tree_add_89_22_pad_groupi_n_646 ,csa_tree_add_89_22_pad_groupi_n_1024);
  or csa_tree_add_89_22_pad_groupi_g4682(csa_tree_add_89_22_pad_groupi_n_1030 ,csa_tree_add_89_22_pad_groupi_n_745 ,csa_tree_add_89_22_pad_groupi_n_1014);
  or csa_tree_add_89_22_pad_groupi_g4683(csa_tree_add_89_22_pad_groupi_n_1029 ,csa_tree_add_89_22_pad_groupi_n_797 ,csa_tree_add_89_22_pad_groupi_n_4);
  nor csa_tree_add_89_22_pad_groupi_g4684(csa_tree_add_89_22_pad_groupi_n_1028 ,csa_tree_add_89_22_pad_groupi_n_746 ,csa_tree_add_89_22_pad_groupi_n_1013);
  and csa_tree_add_89_22_pad_groupi_g4685(csa_tree_add_89_22_pad_groupi_n_1027 ,csa_tree_add_89_22_pad_groupi_n_865 ,csa_tree_add_89_22_pad_groupi_n_1021);
  and csa_tree_add_89_22_pad_groupi_g4686(csa_tree_add_89_22_pad_groupi_n_1026 ,csa_tree_add_89_22_pad_groupi_n_646 ,csa_tree_add_89_22_pad_groupi_n_1024);
  and csa_tree_add_89_22_pad_groupi_g4687(csa_tree_add_89_22_pad_groupi_n_1047 ,csa_tree_add_89_22_pad_groupi_n_895 ,csa_tree_add_89_22_pad_groupi_n_994);
  xnor csa_tree_add_89_22_pad_groupi_g4688(csa_tree_add_89_22_pad_groupi_n_1025 ,csa_tree_add_89_22_pad_groupi_n_935 ,csa_tree_add_89_22_pad_groupi_n_820);
  and csa_tree_add_89_22_pad_groupi_g4689(csa_tree_add_89_22_pad_groupi_n_1046 ,csa_tree_add_89_22_pad_groupi_n_853 ,csa_tree_add_89_22_pad_groupi_n_982);
  or csa_tree_add_89_22_pad_groupi_g4690(csa_tree_add_89_22_pad_groupi_n_1045 ,csa_tree_add_89_22_pad_groupi_n_906 ,csa_tree_add_89_22_pad_groupi_n_997);
  or csa_tree_add_89_22_pad_groupi_g4691(csa_tree_add_89_22_pad_groupi_n_1044 ,csa_tree_add_89_22_pad_groupi_n_887 ,csa_tree_add_89_22_pad_groupi_n_992);
  or csa_tree_add_89_22_pad_groupi_g4692(csa_tree_add_89_22_pad_groupi_n_1043 ,csa_tree_add_89_22_pad_groupi_n_926 ,csa_tree_add_89_22_pad_groupi_n_991);
  and csa_tree_add_89_22_pad_groupi_g4693(csa_tree_add_89_22_pad_groupi_n_1042 ,csa_tree_add_89_22_pad_groupi_n_864 ,csa_tree_add_89_22_pad_groupi_n_985);
  or csa_tree_add_89_22_pad_groupi_g4694(csa_tree_add_89_22_pad_groupi_n_1041 ,csa_tree_add_89_22_pad_groupi_n_879 ,csa_tree_add_89_22_pad_groupi_n_984);
  or csa_tree_add_89_22_pad_groupi_g4695(csa_tree_add_89_22_pad_groupi_n_1040 ,csa_tree_add_89_22_pad_groupi_n_870 ,csa_tree_add_89_22_pad_groupi_n_988);
  and csa_tree_add_89_22_pad_groupi_g4696(csa_tree_add_89_22_pad_groupi_n_1039 ,csa_tree_add_89_22_pad_groupi_n_852 ,csa_tree_add_89_22_pad_groupi_n_981);
  and csa_tree_add_89_22_pad_groupi_g4697(csa_tree_add_89_22_pad_groupi_n_1038 ,csa_tree_add_89_22_pad_groupi_n_878 ,csa_tree_add_89_22_pad_groupi_n_989);
  or csa_tree_add_89_22_pad_groupi_g4698(csa_tree_add_89_22_pad_groupi_n_1036 ,csa_tree_add_89_22_pad_groupi_n_897 ,csa_tree_add_89_22_pad_groupi_n_983);
  or csa_tree_add_89_22_pad_groupi_g4699(csa_tree_add_89_22_pad_groupi_n_1035 ,csa_tree_add_89_22_pad_groupi_n_907 ,csa_tree_add_89_22_pad_groupi_n_990);
  or csa_tree_add_89_22_pad_groupi_g4700(csa_tree_add_89_22_pad_groupi_n_1034 ,csa_tree_add_89_22_pad_groupi_n_866 ,csa_tree_add_89_22_pad_groupi_n_986);
  not csa_tree_add_89_22_pad_groupi_g4701(csa_tree_add_89_22_pad_groupi_n_1023 ,csa_tree_add_89_22_pad_groupi_n_1022);
  not csa_tree_add_89_22_pad_groupi_g4702(csa_tree_add_89_22_pad_groupi_n_1018 ,csa_tree_add_89_22_pad_groupi_n_1017);
  not csa_tree_add_89_22_pad_groupi_g4703(csa_tree_add_89_22_pad_groupi_n_1016 ,csa_tree_add_89_22_pad_groupi_n_1015);
  not csa_tree_add_89_22_pad_groupi_g4704(csa_tree_add_89_22_pad_groupi_n_1014 ,csa_tree_add_89_22_pad_groupi_n_1013);
  not csa_tree_add_89_22_pad_groupi_g4705(csa_tree_add_89_22_pad_groupi_n_1010 ,csa_tree_add_89_22_pad_groupi_n_1009);
  nor csa_tree_add_89_22_pad_groupi_g4706(csa_tree_add_89_22_pad_groupi_n_1008 ,csa_tree_add_89_22_pad_groupi_n_841 ,csa_tree_add_89_22_pad_groupi_n_930);
  or csa_tree_add_89_22_pad_groupi_g4707(csa_tree_add_89_22_pad_groupi_n_1007 ,csa_tree_add_89_22_pad_groupi_n_843 ,csa_tree_add_89_22_pad_groupi_n_917);
  nor csa_tree_add_89_22_pad_groupi_g4708(csa_tree_add_89_22_pad_groupi_n_1006 ,csa_tree_add_89_22_pad_groupi_n_824 ,csa_tree_add_89_22_pad_groupi_n_872);
  and csa_tree_add_89_22_pad_groupi_g4709(csa_tree_add_89_22_pad_groupi_n_1005 ,csa_tree_add_89_22_pad_groupi_n_840 ,csa_tree_add_89_22_pad_groupi_n_922);
  and csa_tree_add_89_22_pad_groupi_g4710(csa_tree_add_89_22_pad_groupi_n_1004 ,csa_tree_add_89_22_pad_groupi_n_839 ,csa_tree_add_89_22_pad_groupi_n_909);
  and csa_tree_add_89_22_pad_groupi_g4711(csa_tree_add_89_22_pad_groupi_n_1003 ,csa_tree_add_89_22_pad_groupi_n_770 ,csa_tree_add_89_22_pad_groupi_n_916);
  or csa_tree_add_89_22_pad_groupi_g4712(csa_tree_add_89_22_pad_groupi_n_1002 ,csa_tree_add_89_22_pad_groupi_n_779 ,csa_tree_add_89_22_pad_groupi_n_902);
  and csa_tree_add_89_22_pad_groupi_g4713(csa_tree_add_89_22_pad_groupi_n_1001 ,csa_tree_add_89_22_pad_groupi_n_769 ,csa_tree_add_89_22_pad_groupi_n_904);
  and csa_tree_add_89_22_pad_groupi_g4714(csa_tree_add_89_22_pad_groupi_n_1000 ,csa_tree_add_89_22_pad_groupi_n_820 ,csa_tree_add_89_22_pad_groupi_n_935);
  nor csa_tree_add_89_22_pad_groupi_g4715(csa_tree_add_89_22_pad_groupi_n_999 ,csa_tree_add_89_22_pad_groupi_n_834 ,csa_tree_add_89_22_pad_groupi_n_896);
  or csa_tree_add_89_22_pad_groupi_g4716(csa_tree_add_89_22_pad_groupi_n_998 ,csa_tree_add_89_22_pad_groupi_n_820 ,csa_tree_add_89_22_pad_groupi_n_935);
  and csa_tree_add_89_22_pad_groupi_g4717(csa_tree_add_89_22_pad_groupi_n_997 ,csa_tree_add_89_22_pad_groupi_n_830 ,csa_tree_add_89_22_pad_groupi_n_856);
  or csa_tree_add_89_22_pad_groupi_g4718(csa_tree_add_89_22_pad_groupi_n_996 ,csa_tree_add_89_22_pad_groupi_n_936 ,csa_tree_add_89_22_pad_groupi_n_919);
  and csa_tree_add_89_22_pad_groupi_g4719(csa_tree_add_89_22_pad_groupi_n_995 ,csa_tree_add_89_22_pad_groupi_n_775 ,csa_tree_add_89_22_pad_groupi_n_891);
  or csa_tree_add_89_22_pad_groupi_g4720(csa_tree_add_89_22_pad_groupi_n_994 ,csa_tree_add_89_22_pad_groupi_n_892 ,csa_tree_add_89_22_pad_groupi_n_894);
  and csa_tree_add_89_22_pad_groupi_g4721(csa_tree_add_89_22_pad_groupi_n_993 ,csa_tree_add_89_22_pad_groupi_n_768 ,csa_tree_add_89_22_pad_groupi_n_924);
  and csa_tree_add_89_22_pad_groupi_g4722(csa_tree_add_89_22_pad_groupi_n_992 ,csa_tree_add_89_22_pad_groupi_n_780 ,csa_tree_add_89_22_pad_groupi_n_885);
  nor csa_tree_add_89_22_pad_groupi_g4723(csa_tree_add_89_22_pad_groupi_n_991 ,csa_tree_add_89_22_pad_groupi_n_837 ,csa_tree_add_89_22_pad_groupi_n_877);
  and csa_tree_add_89_22_pad_groupi_g4724(csa_tree_add_89_22_pad_groupi_n_990 ,csa_tree_add_89_22_pad_groupi_n_777 ,csa_tree_add_89_22_pad_groupi_n_928);
  or csa_tree_add_89_22_pad_groupi_g4725(csa_tree_add_89_22_pad_groupi_n_989 ,csa_tree_add_89_22_pad_groupi_n_838 ,csa_tree_add_89_22_pad_groupi_n_875);
  nor csa_tree_add_89_22_pad_groupi_g4726(csa_tree_add_89_22_pad_groupi_n_988 ,csa_tree_add_89_22_pad_groupi_n_774 ,csa_tree_add_89_22_pad_groupi_n_855);
  nor csa_tree_add_89_22_pad_groupi_g4727(csa_tree_add_89_22_pad_groupi_n_987 ,csa_tree_add_89_22_pad_groupi_n_776 ,csa_tree_add_89_22_pad_groupi_n_883);
  and csa_tree_add_89_22_pad_groupi_g4728(csa_tree_add_89_22_pad_groupi_n_986 ,csa_tree_add_89_22_pad_groupi_n_773 ,csa_tree_add_89_22_pad_groupi_n_863);
  or csa_tree_add_89_22_pad_groupi_g4729(csa_tree_add_89_22_pad_groupi_n_985 ,csa_tree_add_89_22_pad_groupi_n_823 ,csa_tree_add_89_22_pad_groupi_n_862);
  nor csa_tree_add_89_22_pad_groupi_g4730(csa_tree_add_89_22_pad_groupi_n_984 ,csa_tree_add_89_22_pad_groupi_n_772 ,csa_tree_add_89_22_pad_groupi_n_859);
  nor csa_tree_add_89_22_pad_groupi_g4731(csa_tree_add_89_22_pad_groupi_n_983 ,csa_tree_add_89_22_pad_groupi_n_771 ,csa_tree_add_89_22_pad_groupi_n_900);
  or csa_tree_add_89_22_pad_groupi_g4732(csa_tree_add_89_22_pad_groupi_n_982 ,csa_tree_add_89_22_pad_groupi_n_835 ,csa_tree_add_89_22_pad_groupi_n_851);
  or csa_tree_add_89_22_pad_groupi_g4733(csa_tree_add_89_22_pad_groupi_n_981 ,csa_tree_add_89_22_pad_groupi_n_893 ,csa_tree_add_89_22_pad_groupi_n_920);
  xnor csa_tree_add_89_22_pad_groupi_g4734(csa_tree_add_89_22_pad_groupi_n_980 ,csa_tree_add_89_22_pad_groupi_n_846 ,csa_tree_add_89_22_pad_groupi_n_848);
  and csa_tree_add_89_22_pad_groupi_g4735(csa_tree_add_89_22_pad_groupi_n_979 ,csa_tree_add_89_22_pad_groupi_n_827 ,csa_tree_add_89_22_pad_groupi_n_927);
  or csa_tree_add_89_22_pad_groupi_g4736(csa_tree_add_89_22_pad_groupi_n_1024 ,csa_tree_add_89_22_pad_groupi_n_19 ,csa_tree_add_89_22_pad_groupi_n_898);
  xnor csa_tree_add_89_22_pad_groupi_g4737(csa_tree_add_89_22_pad_groupi_n_1022 ,csa_tree_add_89_22_pad_groupi_n_706 ,csa_tree_add_89_22_pad_groupi_n_844);
  xnor csa_tree_add_89_22_pad_groupi_g4739(csa_tree_add_89_22_pad_groupi_n_1021 ,csa_tree_add_89_22_pad_groupi_n_711 ,in13[9]);
  xnor csa_tree_add_89_22_pad_groupi_g4740(csa_tree_add_89_22_pad_groupi_n_1020 ,csa_tree_add_89_22_pad_groupi_n_645 ,csa_tree_add_89_22_pad_groupi_n_832);
  and csa_tree_add_89_22_pad_groupi_g4741(csa_tree_add_89_22_pad_groupi_n_1019 ,csa_tree_add_89_22_pad_groupi_n_899 ,csa_tree_add_89_22_pad_groupi_n_359);
  and csa_tree_add_89_22_pad_groupi_g4742(csa_tree_add_89_22_pad_groupi_n_1017 ,csa_tree_add_89_22_pad_groupi_n_656 ,csa_tree_add_89_22_pad_groupi_n_923);
  or csa_tree_add_89_22_pad_groupi_g4743(csa_tree_add_89_22_pad_groupi_n_1015 ,csa_tree_add_89_22_pad_groupi_n_682 ,csa_tree_add_89_22_pad_groupi_n_881);
  or csa_tree_add_89_22_pad_groupi_g4744(csa_tree_add_89_22_pad_groupi_n_1013 ,csa_tree_add_89_22_pad_groupi_n_666 ,csa_tree_add_89_22_pad_groupi_n_861);
  xnor csa_tree_add_89_22_pad_groupi_g4745(csa_tree_add_89_22_pad_groupi_n_1012 ,csa_tree_add_89_22_pad_groupi_n_704 ,csa_tree_add_89_22_pad_groupi_n_767);
  xnor csa_tree_add_89_22_pad_groupi_g4746(csa_tree_add_89_22_pad_groupi_n_1011 ,csa_tree_add_89_22_pad_groupi_n_831 ,csa_tree_add_89_22_pad_groupi_n_1);
  or csa_tree_add_89_22_pad_groupi_g4747(csa_tree_add_89_22_pad_groupi_n_1009 ,csa_tree_add_89_22_pad_groupi_n_702 ,csa_tree_add_89_22_pad_groupi_n_931);
  xnor csa_tree_add_89_22_pad_groupi_g4748(csa_tree_add_89_22_pad_groupi_n_974 ,csa_tree_add_89_22_pad_groupi_n_726 ,csa_tree_add_89_22_pad_groupi_n_821);
  xnor csa_tree_add_89_22_pad_groupi_g4749(csa_tree_add_89_22_pad_groupi_n_973 ,csa_tree_add_89_22_pad_groupi_n_802 ,csa_tree_add_89_22_pad_groupi_n_795);
  xnor csa_tree_add_89_22_pad_groupi_g4750(csa_tree_add_89_22_pad_groupi_n_972 ,csa_tree_add_89_22_pad_groupi_n_837 ,csa_tree_add_89_22_pad_groupi_n_766);
  xnor csa_tree_add_89_22_pad_groupi_g4751(csa_tree_add_89_22_pad_groupi_n_971 ,csa_tree_add_89_22_pad_groupi_n_829 ,in13[12]);
  xnor csa_tree_add_89_22_pad_groupi_g4752(csa_tree_add_89_22_pad_groupi_n_970 ,csa_tree_add_89_22_pad_groupi_n_739 ,csa_tree_add_89_22_pad_groupi_n_728);
  xnor csa_tree_add_89_22_pad_groupi_g4753(csa_tree_add_89_22_pad_groupi_n_969 ,csa_tree_add_89_22_pad_groupi_n_758 ,csa_tree_add_89_22_pad_groupi_n_757);
  xor csa_tree_add_89_22_pad_groupi_g4754(csa_tree_add_89_22_pad_groupi_n_968 ,csa_tree_add_89_22_pad_groupi_n_824 ,csa_tree_add_89_22_pad_groupi_n_809);
  xor csa_tree_add_89_22_pad_groupi_g4755(csa_tree_add_89_22_pad_groupi_n_967 ,csa_tree_add_89_22_pad_groupi_n_834 ,in13[8]);
  xnor csa_tree_add_89_22_pad_groupi_g4756(csa_tree_add_89_22_pad_groupi_n_966 ,csa_tree_add_89_22_pad_groupi_n_733 ,csa_tree_add_89_22_pad_groupi_n_755);
  xnor csa_tree_add_89_22_pad_groupi_g4757(csa_tree_add_89_22_pad_groupi_n_965 ,csa_tree_add_89_22_pad_groupi_n_800 ,csa_tree_add_89_22_pad_groupi_n_799);
  xor csa_tree_add_89_22_pad_groupi_g4758(csa_tree_add_89_22_pad_groupi_n_964 ,csa_tree_add_89_22_pad_groupi_n_776 ,csa_tree_add_89_22_pad_groupi_n_721);
  xor csa_tree_add_89_22_pad_groupi_g4759(csa_tree_add_89_22_pad_groupi_n_963 ,csa_tree_add_89_22_pad_groupi_n_772 ,in13[1]);
  xnor csa_tree_add_89_22_pad_groupi_g4760(csa_tree_add_89_22_pad_groupi_n_962 ,csa_tree_add_89_22_pad_groupi_n_765 ,csa_tree_add_89_22_pad_groupi_n_751);
  xnor csa_tree_add_89_22_pad_groupi_g4761(csa_tree_add_89_22_pad_groupi_n_961 ,csa_tree_add_89_22_pad_groupi_n_735 ,csa_tree_add_89_22_pad_groupi_n_792);
  xor csa_tree_add_89_22_pad_groupi_g4762(csa_tree_add_89_22_pad_groupi_n_960 ,csa_tree_add_89_22_pad_groupi_n_771 ,csa_tree_add_89_22_pad_groupi_n_729);
  xnor csa_tree_add_89_22_pad_groupi_g4763(csa_tree_add_89_22_pad_groupi_n_959 ,csa_tree_add_89_22_pad_groupi_n_725 ,csa_tree_add_89_22_pad_groupi_n_723);
  xnor csa_tree_add_89_22_pad_groupi_g4764(csa_tree_add_89_22_pad_groupi_n_958 ,csa_tree_add_89_22_pad_groupi_n_814 ,csa_tree_add_89_22_pad_groupi_n_796);
  xnor csa_tree_add_89_22_pad_groupi_g4765(csa_tree_add_89_22_pad_groupi_n_957 ,csa_tree_add_89_22_pad_groupi_n_784 ,csa_tree_add_89_22_pad_groupi_n_747);
  xor csa_tree_add_89_22_pad_groupi_g4766(csa_tree_add_89_22_pad_groupi_n_956 ,csa_tree_add_89_22_pad_groupi_n_841 ,csa_tree_add_89_22_pad_groupi_n_748);
  xnor csa_tree_add_89_22_pad_groupi_g4767(csa_tree_add_89_22_pad_groupi_n_955 ,csa_tree_add_89_22_pad_groupi_n_760 ,csa_tree_add_89_22_pad_groupi_n_737);
  xnor csa_tree_add_89_22_pad_groupi_g4768(csa_tree_add_89_22_pad_groupi_n_954 ,csa_tree_add_89_22_pad_groupi_n_756 ,in13[2]);
  xnor csa_tree_add_89_22_pad_groupi_g4769(csa_tree_add_89_22_pad_groupi_n_953 ,csa_tree_add_89_22_pad_groupi_n_763 ,csa_tree_add_89_22_pad_groupi_n_817);
  xor csa_tree_add_89_22_pad_groupi_g4770(csa_tree_add_89_22_pad_groupi_n_952 ,csa_tree_add_89_22_pad_groupi_n_823 ,csa_tree_add_89_22_pad_groupi_n_742);
  xnor csa_tree_add_89_22_pad_groupi_g4771(csa_tree_add_89_22_pad_groupi_n_951 ,csa_tree_add_89_22_pad_groupi_n_806 ,csa_tree_add_89_22_pad_groupi_n_753);
  xnor csa_tree_add_89_22_pad_groupi_g4772(csa_tree_add_89_22_pad_groupi_n_950 ,csa_tree_add_89_22_pad_groupi_n_790 ,csa_tree_add_89_22_pad_groupi_n_819);
  xnor csa_tree_add_89_22_pad_groupi_g4773(csa_tree_add_89_22_pad_groupi_n_949 ,csa_tree_add_89_22_pad_groupi_n_813 ,csa_tree_add_89_22_pad_groupi_n_716);
  xnor csa_tree_add_89_22_pad_groupi_g4774(csa_tree_add_89_22_pad_groupi_n_948 ,csa_tree_add_89_22_pad_groupi_n_731 ,in13[6]);
  xnor csa_tree_add_89_22_pad_groupi_g4775(csa_tree_add_89_22_pad_groupi_n_947 ,csa_tree_add_89_22_pad_groupi_n_787 ,in13[5]);
  xnor csa_tree_add_89_22_pad_groupi_g4776(csa_tree_add_89_22_pad_groupi_n_946 ,csa_tree_add_89_22_pad_groupi_n_713 ,in13[7]);
  xnor csa_tree_add_89_22_pad_groupi_g4777(csa_tree_add_89_22_pad_groupi_n_945 ,csa_tree_add_89_22_pad_groupi_n_808 ,csa_tree_add_89_22_pad_groupi_n_788);
  xnor csa_tree_add_89_22_pad_groupi_g4778(csa_tree_add_89_22_pad_groupi_n_944 ,csa_tree_add_89_22_pad_groupi_n_761 ,csa_tree_add_89_22_pad_groupi_n_786);
  xnor csa_tree_add_89_22_pad_groupi_g4779(csa_tree_add_89_22_pad_groupi_n_943 ,csa_tree_add_89_22_pad_groupi_n_798 ,in13[4]);
  xnor csa_tree_add_89_22_pad_groupi_g4780(csa_tree_add_89_22_pad_groupi_n_942 ,csa_tree_add_89_22_pad_groupi_n_719 ,csa_tree_add_89_22_pad_groupi_n_720);
  xnor csa_tree_add_89_22_pad_groupi_g4781(csa_tree_add_89_22_pad_groupi_n_941 ,csa_tree_add_89_22_pad_groupi_n_815 ,csa_tree_add_89_22_pad_groupi_n_717);
  xnor csa_tree_add_89_22_pad_groupi_g4782(csa_tree_add_89_22_pad_groupi_n_940 ,csa_tree_add_89_22_pad_groupi_n_807 ,csa_tree_add_89_22_pad_groupi_n_714);
  xnor csa_tree_add_89_22_pad_groupi_g4783(csa_tree_add_89_22_pad_groupi_n_939 ,csa_tree_add_89_22_pad_groupi_n_810 ,csa_tree_add_89_22_pad_groupi_n_811);
  xnor csa_tree_add_89_22_pad_groupi_g4784(csa_tree_add_89_22_pad_groupi_n_938 ,csa_tree_add_89_22_pad_groupi_n_804 ,in13[3]);
  xnor csa_tree_add_89_22_pad_groupi_g4785(csa_tree_add_89_22_pad_groupi_n_937 ,csa_tree_add_89_22_pad_groupi_n_718 ,csa_tree_add_89_22_pad_groupi_n_793);
  xnor csa_tree_add_89_22_pad_groupi_g4786(csa_tree_add_89_22_pad_groupi_n_977 ,csa_tree_add_89_22_pad_groupi_n_822 ,csa_tree_add_89_22_pad_groupi_n_709);
  xnor csa_tree_add_89_22_pad_groupi_g4787(csa_tree_add_89_22_pad_groupi_n_976 ,csa_tree_add_89_22_pad_groupi_n_828 ,csa_tree_add_89_22_pad_groupi_n_710);
  xnor csa_tree_add_89_22_pad_groupi_g4788(csa_tree_add_89_22_pad_groupi_n_975 ,csa_tree_add_89_22_pad_groupi_n_825 ,in13[0]);
  or csa_tree_add_89_22_pad_groupi_g4791(csa_tree_add_89_22_pad_groupi_n_932 ,csa_tree_add_89_22_pad_groupi_n_815 ,csa_tree_add_89_22_pad_groupi_n_717);
  nor csa_tree_add_89_22_pad_groupi_g4792(csa_tree_add_89_22_pad_groupi_n_931 ,csa_tree_add_89_22_pad_groupi_n_673 ,csa_tree_add_89_22_pad_groupi_n_831);
  nor csa_tree_add_89_22_pad_groupi_g4793(csa_tree_add_89_22_pad_groupi_n_930 ,csa_tree_add_89_22_pad_groupi_n_748 ,csa_tree_add_89_22_pad_groupi_n_785);
  nor csa_tree_add_89_22_pad_groupi_g4794(csa_tree_add_89_22_pad_groupi_n_929 ,csa_tree_add_89_22_pad_groupi_n_802 ,csa_tree_add_89_22_pad_groupi_n_794);
  or csa_tree_add_89_22_pad_groupi_g4795(csa_tree_add_89_22_pad_groupi_n_928 ,csa_tree_add_89_22_pad_groupi_n_807 ,csa_tree_add_89_22_pad_groupi_n_714);
  or csa_tree_add_89_22_pad_groupi_g4796(csa_tree_add_89_22_pad_groupi_n_927 ,csa_tree_add_89_22_pad_groupi_n_801 ,csa_tree_add_89_22_pad_groupi_n_795);
  nor csa_tree_add_89_22_pad_groupi_g4797(csa_tree_add_89_22_pad_groupi_n_926 ,csa_tree_add_89_22_pad_groupi_n_766 ,csa_tree_add_89_22_pad_groupi_n_744);
  and csa_tree_add_89_22_pad_groupi_g4798(csa_tree_add_89_22_pad_groupi_n_925 ,csa_tree_add_89_22_pad_groupi_n_764 ,csa_tree_add_89_22_pad_groupi_n_809);
  or csa_tree_add_89_22_pad_groupi_g4799(csa_tree_add_89_22_pad_groupi_n_924 ,csa_tree_add_89_22_pad_groupi_n_719 ,csa_tree_add_89_22_pad_groupi_n_720);
  or csa_tree_add_89_22_pad_groupi_g4800(csa_tree_add_89_22_pad_groupi_n_923 ,csa_tree_add_89_22_pad_groupi_n_593 ,csa_tree_add_89_22_pad_groupi_n_836);
  or csa_tree_add_89_22_pad_groupi_g4801(csa_tree_add_89_22_pad_groupi_n_922 ,csa_tree_add_89_22_pad_groupi_n_800 ,csa_tree_add_89_22_pad_groupi_n_799);
  or csa_tree_add_89_22_pad_groupi_g4802(csa_tree_add_89_22_pad_groupi_n_921 ,csa_tree_add_89_22_pad_groupi_n_789 ,csa_tree_add_89_22_pad_groupi_n_818);
  nor csa_tree_add_89_22_pad_groupi_g4803(csa_tree_add_89_22_pad_groupi_n_920 ,csa_tree_add_89_22_pad_groupi_n_725 ,csa_tree_add_89_22_pad_groupi_n_723);
  nor csa_tree_add_89_22_pad_groupi_g4804(csa_tree_add_89_22_pad_groupi_n_919 ,csa_tree_add_89_22_pad_groupi_n_763 ,csa_tree_add_89_22_pad_groupi_n_817);
  nor csa_tree_add_89_22_pad_groupi_g4805(csa_tree_add_89_22_pad_groupi_n_918 ,csa_tree_add_89_22_pad_groupi_n_790 ,csa_tree_add_89_22_pad_groupi_n_819);
  nor csa_tree_add_89_22_pad_groupi_g4806(csa_tree_add_89_22_pad_groupi_n_917 ,csa_tree_add_89_22_pad_groupi_n_806 ,csa_tree_add_89_22_pad_groupi_n_753);
  or csa_tree_add_89_22_pad_groupi_g4807(csa_tree_add_89_22_pad_groupi_n_916 ,in13[5] ,csa_tree_add_89_22_pad_groupi_n_787);
  or csa_tree_add_89_22_pad_groupi_g4808(csa_tree_add_89_22_pad_groupi_n_915 ,csa_tree_add_89_22_pad_groupi_n_762 ,csa_tree_add_89_22_pad_groupi_n_816);
  and csa_tree_add_89_22_pad_groupi_g4809(csa_tree_add_89_22_pad_groupi_n_914 ,csa_tree_add_89_22_pad_groupi_n_815 ,csa_tree_add_89_22_pad_groupi_n_717);
  or csa_tree_add_89_22_pad_groupi_g4810(csa_tree_add_89_22_pad_groupi_n_913 ,csa_tree_add_89_22_pad_groupi_n_805 ,csa_tree_add_89_22_pad_groupi_n_752);
  or csa_tree_add_89_22_pad_groupi_g4811(csa_tree_add_89_22_pad_groupi_n_912 ,csa_tree_add_89_22_pad_groupi_n_812 ,csa_tree_add_89_22_pad_groupi_n_715);
  and csa_tree_add_89_22_pad_groupi_g4812(csa_tree_add_89_22_pad_groupi_n_911 ,csa_tree_add_89_22_pad_groupi_n_748 ,csa_tree_add_89_22_pad_groupi_n_785);
  nor csa_tree_add_89_22_pad_groupi_g4813(csa_tree_add_89_22_pad_groupi_n_910 ,csa_tree_add_89_22_pad_groupi_n_372 ,csa_tree_add_89_22_pad_groupi_n_782);
  or csa_tree_add_89_22_pad_groupi_g4814(csa_tree_add_89_22_pad_groupi_n_909 ,csa_tree_add_89_22_pad_groupi_n_814 ,csa_tree_add_89_22_pad_groupi_n_796);
  and csa_tree_add_89_22_pad_groupi_g4815(csa_tree_add_89_22_pad_groupi_n_908 ,csa_tree_add_89_22_pad_groupi_n_810 ,csa_tree_add_89_22_pad_groupi_n_811);
  and csa_tree_add_89_22_pad_groupi_g4816(csa_tree_add_89_22_pad_groupi_n_907 ,csa_tree_add_89_22_pad_groupi_n_807 ,csa_tree_add_89_22_pad_groupi_n_714);
  and csa_tree_add_89_22_pad_groupi_g4817(csa_tree_add_89_22_pad_groupi_n_906 ,in13[4] ,csa_tree_add_89_22_pad_groupi_n_798);
  and csa_tree_add_89_22_pad_groupi_g4818(csa_tree_add_89_22_pad_groupi_n_905 ,in13[5] ,csa_tree_add_89_22_pad_groupi_n_787);
  or csa_tree_add_89_22_pad_groupi_g4819(csa_tree_add_89_22_pad_groupi_n_904 ,csa_tree_add_89_22_pad_groupi_n_808 ,csa_tree_add_89_22_pad_groupi_n_788);
  and csa_tree_add_89_22_pad_groupi_g4820(csa_tree_add_89_22_pad_groupi_n_903 ,csa_tree_add_89_22_pad_groupi_n_814 ,csa_tree_add_89_22_pad_groupi_n_796);
  nor csa_tree_add_89_22_pad_groupi_g4821(csa_tree_add_89_22_pad_groupi_n_902 ,csa_tree_add_89_22_pad_groupi_n_813 ,csa_tree_add_89_22_pad_groupi_n_716);
  and csa_tree_add_89_22_pad_groupi_g4822(csa_tree_add_89_22_pad_groupi_n_901 ,csa_tree_add_89_22_pad_groupi_n_761 ,csa_tree_add_89_22_pad_groupi_n_786);
  nor csa_tree_add_89_22_pad_groupi_g4823(csa_tree_add_89_22_pad_groupi_n_900 ,csa_tree_add_89_22_pad_groupi_n_783 ,csa_tree_add_89_22_pad_groupi_n_729);
  or csa_tree_add_89_22_pad_groupi_g4824(csa_tree_add_89_22_pad_groupi_n_899 ,csa_tree_add_89_22_pad_groupi_n_708 ,csa_tree_add_89_22_pad_groupi_n_845);
  or csa_tree_add_89_22_pad_groupi_g4825(csa_tree_add_89_22_pad_groupi_n_898 ,csa_tree_add_89_22_pad_groupi_n_112 ,csa_tree_add_89_22_pad_groupi_n_781);
  and csa_tree_add_89_22_pad_groupi_g4826(csa_tree_add_89_22_pad_groupi_n_897 ,csa_tree_add_89_22_pad_groupi_n_783 ,csa_tree_add_89_22_pad_groupi_n_729);
  and csa_tree_add_89_22_pad_groupi_g4827(csa_tree_add_89_22_pad_groupi_n_896 ,csa_tree_add_89_22_pad_groupi_n_372 ,csa_tree_add_89_22_pad_groupi_n_782);
  or csa_tree_add_89_22_pad_groupi_g4828(csa_tree_add_89_22_pad_groupi_n_895 ,csa_tree_add_89_22_pad_groupi_n_734 ,csa_tree_add_89_22_pad_groupi_n_791);
  nor csa_tree_add_89_22_pad_groupi_g4829(csa_tree_add_89_22_pad_groupi_n_894 ,csa_tree_add_89_22_pad_groupi_n_735 ,csa_tree_add_89_22_pad_groupi_n_792);
  or csa_tree_add_89_22_pad_groupi_g4830(csa_tree_add_89_22_pad_groupi_n_936 ,csa_tree_add_89_22_pad_groupi_n_645 ,csa_tree_add_89_22_pad_groupi_n_833);
  and csa_tree_add_89_22_pad_groupi_g4831(csa_tree_add_89_22_pad_groupi_n_935 ,csa_tree_add_89_22_pad_groupi_n_705 ,csa_tree_add_89_22_pad_groupi_n_767);
  and csa_tree_add_89_22_pad_groupi_g4832(csa_tree_add_89_22_pad_groupi_n_934 ,csa_tree_add_89_22_pad_groupi_n_708 ,csa_tree_add_89_22_pad_groupi_n_845);
  and csa_tree_add_89_22_pad_groupi_g4833(csa_tree_add_89_22_pad_groupi_n_933 ,csa_tree_add_89_22_pad_groupi_n_707 ,csa_tree_add_89_22_pad_groupi_n_844);
  or csa_tree_add_89_22_pad_groupi_g4834(csa_tree_add_89_22_pad_groupi_n_891 ,csa_tree_add_89_22_pad_groupi_n_718 ,csa_tree_add_89_22_pad_groupi_n_793);
  and csa_tree_add_89_22_pad_groupi_g4835(csa_tree_add_89_22_pad_groupi_n_890 ,csa_tree_add_89_22_pad_groupi_n_800 ,csa_tree_add_89_22_pad_groupi_n_799);
  and csa_tree_add_89_22_pad_groupi_g4836(csa_tree_add_89_22_pad_groupi_n_889 ,csa_tree_add_89_22_pad_groupi_n_718 ,csa_tree_add_89_22_pad_groupi_n_793);
  or csa_tree_add_89_22_pad_groupi_g4837(csa_tree_add_89_22_pad_groupi_n_888 ,csa_tree_add_89_22_pad_groupi_n_732 ,csa_tree_add_89_22_pad_groupi_n_754);
  and csa_tree_add_89_22_pad_groupi_g4838(csa_tree_add_89_22_pad_groupi_n_887 ,in13[3] ,csa_tree_add_89_22_pad_groupi_n_804);
  and csa_tree_add_89_22_pad_groupi_g4839(csa_tree_add_89_22_pad_groupi_n_886 ,csa_tree_add_89_22_pad_groupi_n_719 ,csa_tree_add_89_22_pad_groupi_n_720);
  or csa_tree_add_89_22_pad_groupi_g4840(csa_tree_add_89_22_pad_groupi_n_885 ,in13[3] ,csa_tree_add_89_22_pad_groupi_n_804);
  or csa_tree_add_89_22_pad_groupi_g4841(csa_tree_add_89_22_pad_groupi_n_884 ,csa_tree_add_89_22_pad_groupi_n_738 ,csa_tree_add_89_22_pad_groupi_n_727);
  nor csa_tree_add_89_22_pad_groupi_g4842(csa_tree_add_89_22_pad_groupi_n_883 ,csa_tree_add_89_22_pad_groupi_n_803 ,csa_tree_add_89_22_pad_groupi_n_721);
  nor csa_tree_add_89_22_pad_groupi_g4843(csa_tree_add_89_22_pad_groupi_n_882 ,csa_tree_add_89_22_pad_groupi_n_739 ,csa_tree_add_89_22_pad_groupi_n_728);
  nor csa_tree_add_89_22_pad_groupi_g4844(csa_tree_add_89_22_pad_groupi_n_881 ,csa_tree_add_89_22_pad_groupi_n_700 ,csa_tree_add_89_22_pad_groupi_n_828);
  or csa_tree_add_89_22_pad_groupi_g4845(csa_tree_add_89_22_pad_groupi_n_880 ,csa_tree_add_89_22_pad_groupi_n_761 ,csa_tree_add_89_22_pad_groupi_n_786);
  nor csa_tree_add_89_22_pad_groupi_g4846(csa_tree_add_89_22_pad_groupi_n_879 ,csa_tree_add_89_22_pad_groupi_n_371 ,csa_tree_add_89_22_pad_groupi_n_740);
  or csa_tree_add_89_22_pad_groupi_g4847(csa_tree_add_89_22_pad_groupi_n_878 ,csa_tree_add_89_22_pad_groupi_n_387 ,csa_tree_add_89_22_pad_groupi_n_712);
  and csa_tree_add_89_22_pad_groupi_g4848(csa_tree_add_89_22_pad_groupi_n_877 ,csa_tree_add_89_22_pad_groupi_n_766 ,csa_tree_add_89_22_pad_groupi_n_744);
  nor csa_tree_add_89_22_pad_groupi_g4849(csa_tree_add_89_22_pad_groupi_n_876 ,csa_tree_add_89_22_pad_groupi_n_733 ,csa_tree_add_89_22_pad_groupi_n_755);
  nor csa_tree_add_89_22_pad_groupi_g4850(csa_tree_add_89_22_pad_groupi_n_875 ,in13[7] ,csa_tree_add_89_22_pad_groupi_n_713);
  and csa_tree_add_89_22_pad_groupi_g4851(csa_tree_add_89_22_pad_groupi_n_874 ,csa_tree_add_89_22_pad_groupi_n_803 ,csa_tree_add_89_22_pad_groupi_n_721);
  and csa_tree_add_89_22_pad_groupi_g4852(csa_tree_add_89_22_pad_groupi_n_873 ,csa_tree_add_89_22_pad_groupi_n_758 ,csa_tree_add_89_22_pad_groupi_n_757);
  nor csa_tree_add_89_22_pad_groupi_g4853(csa_tree_add_89_22_pad_groupi_n_872 ,csa_tree_add_89_22_pad_groupi_n_764 ,csa_tree_add_89_22_pad_groupi_n_809);
  or csa_tree_add_89_22_pad_groupi_g4854(csa_tree_add_89_22_pad_groupi_n_871 ,csa_tree_add_89_22_pad_groupi_n_758 ,csa_tree_add_89_22_pad_groupi_n_757);
  and csa_tree_add_89_22_pad_groupi_g4855(csa_tree_add_89_22_pad_groupi_n_870 ,in13[2] ,csa_tree_add_89_22_pad_groupi_n_756);
  and csa_tree_add_89_22_pad_groupi_g4856(csa_tree_add_89_22_pad_groupi_n_869 ,csa_tree_add_89_22_pad_groupi_n_808 ,csa_tree_add_89_22_pad_groupi_n_788);
  and csa_tree_add_89_22_pad_groupi_g4857(csa_tree_add_89_22_pad_groupi_n_868 ,csa_tree_add_89_22_pad_groupi_n_784 ,csa_tree_add_89_22_pad_groupi_n_747);
  or csa_tree_add_89_22_pad_groupi_g4858(csa_tree_add_89_22_pad_groupi_n_867 ,csa_tree_add_89_22_pad_groupi_n_810 ,csa_tree_add_89_22_pad_groupi_n_811);
  and csa_tree_add_89_22_pad_groupi_g4859(csa_tree_add_89_22_pad_groupi_n_866 ,csa_tree_add_89_22_pad_groupi_n_765 ,csa_tree_add_89_22_pad_groupi_n_751);
  or csa_tree_add_89_22_pad_groupi_g4860(csa_tree_add_89_22_pad_groupi_n_865 ,csa_tree_add_89_22_pad_groupi_n_784 ,csa_tree_add_89_22_pad_groupi_n_747);
  or csa_tree_add_89_22_pad_groupi_g4861(csa_tree_add_89_22_pad_groupi_n_864 ,csa_tree_add_89_22_pad_groupi_n_749 ,csa_tree_add_89_22_pad_groupi_n_741);
  or csa_tree_add_89_22_pad_groupi_g4862(csa_tree_add_89_22_pad_groupi_n_863 ,csa_tree_add_89_22_pad_groupi_n_765 ,csa_tree_add_89_22_pad_groupi_n_751);
  nor csa_tree_add_89_22_pad_groupi_g4863(csa_tree_add_89_22_pad_groupi_n_862 ,csa_tree_add_89_22_pad_groupi_n_750 ,csa_tree_add_89_22_pad_groupi_n_742);
  nor csa_tree_add_89_22_pad_groupi_g4864(csa_tree_add_89_22_pad_groupi_n_861 ,csa_tree_add_89_22_pad_groupi_n_600 ,csa_tree_add_89_22_pad_groupi_n_822);
  or csa_tree_add_89_22_pad_groupi_g4865(csa_tree_add_89_22_pad_groupi_n_860 ,csa_tree_add_89_22_pad_groupi_n_726 ,csa_tree_add_89_22_pad_groupi_n_821);
  and csa_tree_add_89_22_pad_groupi_g4866(csa_tree_add_89_22_pad_groupi_n_859 ,csa_tree_add_89_22_pad_groupi_n_371 ,csa_tree_add_89_22_pad_groupi_n_740);
  and csa_tree_add_89_22_pad_groupi_g4867(csa_tree_add_89_22_pad_groupi_n_858 ,csa_tree_add_89_22_pad_groupi_n_726 ,csa_tree_add_89_22_pad_groupi_n_821);
  or csa_tree_add_89_22_pad_groupi_g4868(csa_tree_add_89_22_pad_groupi_n_857 ,csa_tree_add_89_22_pad_groupi_n_759 ,csa_tree_add_89_22_pad_groupi_n_736);
  or csa_tree_add_89_22_pad_groupi_g4869(csa_tree_add_89_22_pad_groupi_n_856 ,in13[4] ,csa_tree_add_89_22_pad_groupi_n_798);
  nor csa_tree_add_89_22_pad_groupi_g4870(csa_tree_add_89_22_pad_groupi_n_855 ,in13[2] ,csa_tree_add_89_22_pad_groupi_n_756);
  nor csa_tree_add_89_22_pad_groupi_g4871(csa_tree_add_89_22_pad_groupi_n_854 ,csa_tree_add_89_22_pad_groupi_n_760 ,csa_tree_add_89_22_pad_groupi_n_737);
  or csa_tree_add_89_22_pad_groupi_g4872(csa_tree_add_89_22_pad_groupi_n_853 ,csa_tree_add_89_22_pad_groupi_n_370 ,csa_tree_add_89_22_pad_groupi_n_730);
  or csa_tree_add_89_22_pad_groupi_g4873(csa_tree_add_89_22_pad_groupi_n_852 ,csa_tree_add_89_22_pad_groupi_n_724 ,csa_tree_add_89_22_pad_groupi_n_722);
  nor csa_tree_add_89_22_pad_groupi_g4874(csa_tree_add_89_22_pad_groupi_n_851 ,in13[6] ,csa_tree_add_89_22_pad_groupi_n_731);
  or csa_tree_add_89_22_pad_groupi_g4876(csa_tree_add_89_22_pad_groupi_n_893 ,csa_tree_add_89_22_pad_groupi_n_374 ,csa_tree_add_89_22_pad_groupi_n_826);
  or csa_tree_add_89_22_pad_groupi_g4877(csa_tree_add_89_22_pad_groupi_n_892 ,csa_tree_add_89_22_pad_groupi_n_847 ,csa_tree_add_89_22_pad_groupi_n_849);
  not csa_tree_add_89_22_pad_groupi_g4878(csa_tree_add_89_22_pad_groupi_n_849 ,csa_tree_add_89_22_pad_groupi_n_848);
  not csa_tree_add_89_22_pad_groupi_g4879(csa_tree_add_89_22_pad_groupi_n_847 ,csa_tree_add_89_22_pad_groupi_n_846);
  not csa_tree_add_89_22_pad_groupi_g4880(csa_tree_add_89_22_pad_groupi_n_843 ,csa_tree_add_89_22_pad_groupi_n_842);
  not csa_tree_add_89_22_pad_groupi_g4883(csa_tree_add_89_22_pad_groupi_n_833 ,csa_tree_add_89_22_pad_groupi_n_832);
  not csa_tree_add_89_22_pad_groupi_g4884(csa_tree_add_89_22_pad_groupi_n_826 ,csa_tree_add_89_22_pad_groupi_n_825);
  not csa_tree_add_89_22_pad_groupi_g4885(csa_tree_add_89_22_pad_groupi_n_818 ,csa_tree_add_89_22_pad_groupi_n_819);
  not csa_tree_add_89_22_pad_groupi_g4886(csa_tree_add_89_22_pad_groupi_n_816 ,csa_tree_add_89_22_pad_groupi_n_817);
  not csa_tree_add_89_22_pad_groupi_g4887(csa_tree_add_89_22_pad_groupi_n_812 ,csa_tree_add_89_22_pad_groupi_n_813);
  not csa_tree_add_89_22_pad_groupi_g4888(csa_tree_add_89_22_pad_groupi_n_805 ,csa_tree_add_89_22_pad_groupi_n_806);
  not csa_tree_add_89_22_pad_groupi_g4889(csa_tree_add_89_22_pad_groupi_n_801 ,csa_tree_add_89_22_pad_groupi_n_802);
  not csa_tree_add_89_22_pad_groupi_g4890(csa_tree_add_89_22_pad_groupi_n_794 ,csa_tree_add_89_22_pad_groupi_n_795);
  not csa_tree_add_89_22_pad_groupi_g4891(csa_tree_add_89_22_pad_groupi_n_791 ,csa_tree_add_89_22_pad_groupi_n_792);
  not csa_tree_add_89_22_pad_groupi_g4892(csa_tree_add_89_22_pad_groupi_n_789 ,csa_tree_add_89_22_pad_groupi_n_790);
  and csa_tree_add_89_22_pad_groupi_g4893(csa_tree_add_89_22_pad_groupi_n_781 ,csa_tree_add_89_22_pad_groupi_n_459 ,csa_tree_add_89_22_pad_groupi_n_612);
  or csa_tree_add_89_22_pad_groupi_g4894(csa_tree_add_89_22_pad_groupi_n_848 ,csa_tree_add_89_22_pad_groupi_n_466 ,csa_tree_add_89_22_pad_groupi_n_621);
  or csa_tree_add_89_22_pad_groupi_g4895(csa_tree_add_89_22_pad_groupi_n_846 ,csa_tree_add_89_22_pad_groupi_n_576 ,csa_tree_add_89_22_pad_groupi_n_703);
  and csa_tree_add_89_22_pad_groupi_g4896(csa_tree_add_89_22_pad_groupi_n_845 ,csa_tree_add_89_22_pad_groupi_n_531 ,csa_tree_add_89_22_pad_groupi_n_685);
  or csa_tree_add_89_22_pad_groupi_g4897(csa_tree_add_89_22_pad_groupi_n_844 ,csa_tree_add_89_22_pad_groupi_n_526 ,csa_tree_add_89_22_pad_groupi_n_652);
  or csa_tree_add_89_22_pad_groupi_g4898(csa_tree_add_89_22_pad_groupi_n_842 ,csa_tree_add_89_22_pad_groupi_n_533 ,csa_tree_add_89_22_pad_groupi_n_618);
  and csa_tree_add_89_22_pad_groupi_g4899(csa_tree_add_89_22_pad_groupi_n_841 ,csa_tree_add_89_22_pad_groupi_n_472 ,csa_tree_add_89_22_pad_groupi_n_642);
  or csa_tree_add_89_22_pad_groupi_g4900(csa_tree_add_89_22_pad_groupi_n_840 ,csa_tree_add_89_22_pad_groupi_n_557 ,csa_tree_add_89_22_pad_groupi_n_598);
  or csa_tree_add_89_22_pad_groupi_g4901(csa_tree_add_89_22_pad_groupi_n_839 ,csa_tree_add_89_22_pad_groupi_n_574 ,csa_tree_add_89_22_pad_groupi_n_588);
  and csa_tree_add_89_22_pad_groupi_g4903(csa_tree_add_89_22_pad_groupi_n_837 ,csa_tree_add_89_22_pad_groupi_n_483 ,csa_tree_add_89_22_pad_groupi_n_587);
  and csa_tree_add_89_22_pad_groupi_g4906(csa_tree_add_89_22_pad_groupi_n_834 ,csa_tree_add_89_22_pad_groupi_n_460 ,csa_tree_add_89_22_pad_groupi_n_586);
  or csa_tree_add_89_22_pad_groupi_g4907(csa_tree_add_89_22_pad_groupi_n_832 ,csa_tree_add_89_22_pad_groupi_n_548 ,csa_tree_add_89_22_pad_groupi_n_699);
  or csa_tree_add_89_22_pad_groupi_g4912(csa_tree_add_89_22_pad_groupi_n_827 ,csa_tree_add_89_22_pad_groupi_n_487 ,csa_tree_add_89_22_pad_groupi_n_647);
  or csa_tree_add_89_22_pad_groupi_g4913(csa_tree_add_89_22_pad_groupi_n_825 ,csa_tree_add_89_22_pad_groupi_n_462 ,csa_tree_add_89_22_pad_groupi_n_662);
  and csa_tree_add_89_22_pad_groupi_g4914(csa_tree_add_89_22_pad_groupi_n_824 ,csa_tree_add_89_22_pad_groupi_n_485 ,csa_tree_add_89_22_pad_groupi_n_683);
  and csa_tree_add_89_22_pad_groupi_g4915(csa_tree_add_89_22_pad_groupi_n_823 ,csa_tree_add_89_22_pad_groupi_n_518 ,csa_tree_add_89_22_pad_groupi_n_595);
  or csa_tree_add_89_22_pad_groupi_g4917(csa_tree_add_89_22_pad_groupi_n_821 ,csa_tree_add_89_22_pad_groupi_n_551 ,csa_tree_add_89_22_pad_groupi_n_665);
  or csa_tree_add_89_22_pad_groupi_g4918(csa_tree_add_89_22_pad_groupi_n_820 ,csa_tree_add_89_22_pad_groupi_n_556 ,csa_tree_add_89_22_pad_groupi_n_677);
  or csa_tree_add_89_22_pad_groupi_g4919(csa_tree_add_89_22_pad_groupi_n_819 ,csa_tree_add_89_22_pad_groupi_n_516 ,csa_tree_add_89_22_pad_groupi_n_681);
  or csa_tree_add_89_22_pad_groupi_g4920(csa_tree_add_89_22_pad_groupi_n_817 ,csa_tree_add_89_22_pad_groupi_n_527 ,csa_tree_add_89_22_pad_groupi_n_674);
  or csa_tree_add_89_22_pad_groupi_g4921(csa_tree_add_89_22_pad_groupi_n_815 ,csa_tree_add_89_22_pad_groupi_n_491 ,csa_tree_add_89_22_pad_groupi_n_649);
  or csa_tree_add_89_22_pad_groupi_g4922(csa_tree_add_89_22_pad_groupi_n_814 ,csa_tree_add_89_22_pad_groupi_n_475 ,csa_tree_add_89_22_pad_groupi_n_633);
  or csa_tree_add_89_22_pad_groupi_g4923(csa_tree_add_89_22_pad_groupi_n_813 ,csa_tree_add_89_22_pad_groupi_n_525 ,csa_tree_add_89_22_pad_groupi_n_695);
  or csa_tree_add_89_22_pad_groupi_g4924(csa_tree_add_89_22_pad_groupi_n_811 ,csa_tree_add_89_22_pad_groupi_n_476 ,csa_tree_add_89_22_pad_groupi_n_599);
  or csa_tree_add_89_22_pad_groupi_g4925(csa_tree_add_89_22_pad_groupi_n_810 ,csa_tree_add_89_22_pad_groupi_n_470 ,csa_tree_add_89_22_pad_groupi_n_627);
  or csa_tree_add_89_22_pad_groupi_g4926(csa_tree_add_89_22_pad_groupi_n_809 ,csa_tree_add_89_22_pad_groupi_n_528 ,csa_tree_add_89_22_pad_groupi_n_651);
  or csa_tree_add_89_22_pad_groupi_g4927(csa_tree_add_89_22_pad_groupi_n_808 ,csa_tree_add_89_22_pad_groupi_n_541 ,csa_tree_add_89_22_pad_groupi_n_635);
  or csa_tree_add_89_22_pad_groupi_g4928(csa_tree_add_89_22_pad_groupi_n_807 ,csa_tree_add_89_22_pad_groupi_n_512 ,csa_tree_add_89_22_pad_groupi_n_625);
  or csa_tree_add_89_22_pad_groupi_g4929(csa_tree_add_89_22_pad_groupi_n_806 ,csa_tree_add_89_22_pad_groupi_n_523 ,csa_tree_add_89_22_pad_groupi_n_623);
  or csa_tree_add_89_22_pad_groupi_g4930(csa_tree_add_89_22_pad_groupi_n_804 ,csa_tree_add_89_22_pad_groupi_n_461 ,csa_tree_add_89_22_pad_groupi_n_694);
  or csa_tree_add_89_22_pad_groupi_g4931(csa_tree_add_89_22_pad_groupi_n_803 ,csa_tree_add_89_22_pad_groupi_n_529 ,csa_tree_add_89_22_pad_groupi_n_653);
  or csa_tree_add_89_22_pad_groupi_g4933(csa_tree_add_89_22_pad_groupi_n_800 ,csa_tree_add_89_22_pad_groupi_n_477 ,csa_tree_add_89_22_pad_groupi_n_658);
  or csa_tree_add_89_22_pad_groupi_g4934(csa_tree_add_89_22_pad_groupi_n_799 ,csa_tree_add_89_22_pad_groupi_n_467 ,csa_tree_add_89_22_pad_groupi_n_680);
  or csa_tree_add_89_22_pad_groupi_g4935(csa_tree_add_89_22_pad_groupi_n_798 ,csa_tree_add_89_22_pad_groupi_n_468 ,csa_tree_add_89_22_pad_groupi_n_607);
  or csa_tree_add_89_22_pad_groupi_g4936(csa_tree_add_89_22_pad_groupi_n_797 ,csa_tree_add_89_22_pad_groupi_n_394 ,csa_tree_add_89_22_pad_groupi_n_663);
  or csa_tree_add_89_22_pad_groupi_g4937(csa_tree_add_89_22_pad_groupi_n_796 ,csa_tree_add_89_22_pad_groupi_n_555 ,csa_tree_add_89_22_pad_groupi_n_669);
  or csa_tree_add_89_22_pad_groupi_g4938(csa_tree_add_89_22_pad_groupi_n_795 ,csa_tree_add_89_22_pad_groupi_n_547 ,csa_tree_add_89_22_pad_groupi_n_696);
  or csa_tree_add_89_22_pad_groupi_g4939(csa_tree_add_89_22_pad_groupi_n_793 ,csa_tree_add_89_22_pad_groupi_n_540 ,csa_tree_add_89_22_pad_groupi_n_697);
  or csa_tree_add_89_22_pad_groupi_g4940(csa_tree_add_89_22_pad_groupi_n_792 ,csa_tree_add_89_22_pad_groupi_n_456 ,csa_tree_add_89_22_pad_groupi_n_638);
  or csa_tree_add_89_22_pad_groupi_g4941(csa_tree_add_89_22_pad_groupi_n_790 ,csa_tree_add_89_22_pad_groupi_n_524 ,csa_tree_add_89_22_pad_groupi_n_661);
  or csa_tree_add_89_22_pad_groupi_g4942(csa_tree_add_89_22_pad_groupi_n_788 ,csa_tree_add_89_22_pad_groupi_n_537 ,csa_tree_add_89_22_pad_groupi_n_616);
  or csa_tree_add_89_22_pad_groupi_g4943(csa_tree_add_89_22_pad_groupi_n_787 ,csa_tree_add_89_22_pad_groupi_n_469 ,csa_tree_add_89_22_pad_groupi_n_672);
  or csa_tree_add_89_22_pad_groupi_g4944(csa_tree_add_89_22_pad_groupi_n_786 ,csa_tree_add_89_22_pad_groupi_n_473 ,csa_tree_add_89_22_pad_groupi_n_589);
  or csa_tree_add_89_22_pad_groupi_g4945(csa_tree_add_89_22_pad_groupi_n_785 ,csa_tree_add_89_22_pad_groupi_n_484 ,csa_tree_add_89_22_pad_groupi_n_698);
  or csa_tree_add_89_22_pad_groupi_g4946(csa_tree_add_89_22_pad_groupi_n_784 ,csa_tree_add_89_22_pad_groupi_n_488 ,csa_tree_add_89_22_pad_groupi_n_608);
  or csa_tree_add_89_22_pad_groupi_g4947(csa_tree_add_89_22_pad_groupi_n_783 ,csa_tree_add_89_22_pad_groupi_n_546 ,csa_tree_add_89_22_pad_groupi_n_648);
  not csa_tree_add_89_22_pad_groupi_g4949(csa_tree_add_89_22_pad_groupi_n_779 ,csa_tree_add_89_22_pad_groupi_n_778);
  not csa_tree_add_89_22_pad_groupi_g4950(csa_tree_add_89_22_pad_groupi_n_762 ,csa_tree_add_89_22_pad_groupi_n_763);
  not csa_tree_add_89_22_pad_groupi_g4951(csa_tree_add_89_22_pad_groupi_n_759 ,csa_tree_add_89_22_pad_groupi_n_760);
  not csa_tree_add_89_22_pad_groupi_g4952(csa_tree_add_89_22_pad_groupi_n_754 ,csa_tree_add_89_22_pad_groupi_n_755);
  not csa_tree_add_89_22_pad_groupi_g4953(csa_tree_add_89_22_pad_groupi_n_752 ,csa_tree_add_89_22_pad_groupi_n_753);
  not csa_tree_add_89_22_pad_groupi_g4954(csa_tree_add_89_22_pad_groupi_n_749 ,csa_tree_add_89_22_pad_groupi_n_750);
  not csa_tree_add_89_22_pad_groupi_g4955(csa_tree_add_89_22_pad_groupi_n_745 ,csa_tree_add_89_22_pad_groupi_n_746);
  not csa_tree_add_89_22_pad_groupi_g4956(csa_tree_add_89_22_pad_groupi_n_744 ,csa_tree_add_89_22_pad_groupi_n_743);
  not csa_tree_add_89_22_pad_groupi_g4957(csa_tree_add_89_22_pad_groupi_n_741 ,csa_tree_add_89_22_pad_groupi_n_742);
  not csa_tree_add_89_22_pad_groupi_g4958(csa_tree_add_89_22_pad_groupi_n_738 ,csa_tree_add_89_22_pad_groupi_n_739);
  not csa_tree_add_89_22_pad_groupi_g4959(csa_tree_add_89_22_pad_groupi_n_736 ,csa_tree_add_89_22_pad_groupi_n_737);
  not csa_tree_add_89_22_pad_groupi_g4960(csa_tree_add_89_22_pad_groupi_n_734 ,csa_tree_add_89_22_pad_groupi_n_735);
  not csa_tree_add_89_22_pad_groupi_g4961(csa_tree_add_89_22_pad_groupi_n_732 ,csa_tree_add_89_22_pad_groupi_n_733);
  not csa_tree_add_89_22_pad_groupi_g4962(csa_tree_add_89_22_pad_groupi_n_730 ,csa_tree_add_89_22_pad_groupi_n_731);
  not csa_tree_add_89_22_pad_groupi_g4963(csa_tree_add_89_22_pad_groupi_n_727 ,csa_tree_add_89_22_pad_groupi_n_728);
  not csa_tree_add_89_22_pad_groupi_g4964(csa_tree_add_89_22_pad_groupi_n_724 ,csa_tree_add_89_22_pad_groupi_n_725);
  not csa_tree_add_89_22_pad_groupi_g4965(csa_tree_add_89_22_pad_groupi_n_722 ,csa_tree_add_89_22_pad_groupi_n_723);
  not csa_tree_add_89_22_pad_groupi_g4966(csa_tree_add_89_22_pad_groupi_n_715 ,csa_tree_add_89_22_pad_groupi_n_716);
  not csa_tree_add_89_22_pad_groupi_g4967(csa_tree_add_89_22_pad_groupi_n_712 ,csa_tree_add_89_22_pad_groupi_n_713);
  xnor csa_tree_add_89_22_pad_groupi_g4968(csa_tree_add_89_22_pad_groupi_n_711 ,csa_tree_add_89_22_pad_groupi_n_583 ,in13[10]);
  xnor csa_tree_add_89_22_pad_groupi_g4970(csa_tree_add_89_22_pad_groupi_n_710 ,csa_tree_add_89_22_pad_groupi_n_282 ,in13[12]);
  xnor csa_tree_add_89_22_pad_groupi_g4972(csa_tree_add_89_22_pad_groupi_n_709 ,csa_tree_add_89_22_pad_groupi_n_582 ,in13[12]);
  or csa_tree_add_89_22_pad_groupi_g4975(csa_tree_add_89_22_pad_groupi_n_778 ,csa_tree_add_89_22_pad_groupi_n_539 ,csa_tree_add_89_22_pad_groupi_n_626);
  or csa_tree_add_89_22_pad_groupi_g4976(csa_tree_add_89_22_pad_groupi_n_777 ,csa_tree_add_89_22_pad_groupi_n_550 ,csa_tree_add_89_22_pad_groupi_n_624);
  and csa_tree_add_89_22_pad_groupi_g4977(csa_tree_add_89_22_pad_groupi_n_776 ,csa_tree_add_89_22_pad_groupi_n_464 ,csa_tree_add_89_22_pad_groupi_n_655);
  or csa_tree_add_89_22_pad_groupi_g4978(csa_tree_add_89_22_pad_groupi_n_775 ,csa_tree_add_89_22_pad_groupi_n_482 ,csa_tree_add_89_22_pad_groupi_n_637);
  or csa_tree_add_89_22_pad_groupi_g4980(csa_tree_add_89_22_pad_groupi_n_773 ,csa_tree_add_89_22_pad_groupi_n_519 ,csa_tree_add_89_22_pad_groupi_n_605);
  and csa_tree_add_89_22_pad_groupi_g4981(csa_tree_add_89_22_pad_groupi_n_772 ,csa_tree_add_89_22_pad_groupi_n_457 ,csa_tree_add_89_22_pad_groupi_n_594);
  and csa_tree_add_89_22_pad_groupi_g4982(csa_tree_add_89_22_pad_groupi_n_771 ,csa_tree_add_89_22_pad_groupi_n_492 ,csa_tree_add_89_22_pad_groupi_n_606);
  or csa_tree_add_89_22_pad_groupi_g4984(csa_tree_add_89_22_pad_groupi_n_769 ,csa_tree_add_89_22_pad_groupi_n_490 ,csa_tree_add_89_22_pad_groupi_n_689);
  or csa_tree_add_89_22_pad_groupi_g4985(csa_tree_add_89_22_pad_groupi_n_768 ,csa_tree_add_89_22_pad_groupi_n_545 ,csa_tree_add_89_22_pad_groupi_n_640);
  or csa_tree_add_89_22_pad_groupi_g4986(csa_tree_add_89_22_pad_groupi_n_767 ,csa_tree_add_89_22_pad_groupi_n_552 ,csa_tree_add_89_22_pad_groupi_n_659);
  or csa_tree_add_89_22_pad_groupi_g4988(csa_tree_add_89_22_pad_groupi_n_765 ,csa_tree_add_89_22_pad_groupi_n_517 ,csa_tree_add_89_22_pad_groupi_n_688);
  or csa_tree_add_89_22_pad_groupi_g4989(csa_tree_add_89_22_pad_groupi_n_764 ,csa_tree_add_89_22_pad_groupi_n_554 ,csa_tree_add_89_22_pad_groupi_n_654);
  or csa_tree_add_89_22_pad_groupi_g4990(csa_tree_add_89_22_pad_groupi_n_763 ,csa_tree_add_89_22_pad_groupi_n_480 ,csa_tree_add_89_22_pad_groupi_n_602);
  or csa_tree_add_89_22_pad_groupi_g4991(csa_tree_add_89_22_pad_groupi_n_761 ,csa_tree_add_89_22_pad_groupi_n_577 ,csa_tree_add_89_22_pad_groupi_n_693);
  or csa_tree_add_89_22_pad_groupi_g4992(csa_tree_add_89_22_pad_groupi_n_760 ,csa_tree_add_89_22_pad_groupi_n_478 ,csa_tree_add_89_22_pad_groupi_n_591);
  or csa_tree_add_89_22_pad_groupi_g4993(csa_tree_add_89_22_pad_groupi_n_758 ,csa_tree_add_89_22_pad_groupi_n_514 ,csa_tree_add_89_22_pad_groupi_n_604);
  or csa_tree_add_89_22_pad_groupi_g4994(csa_tree_add_89_22_pad_groupi_n_757 ,csa_tree_add_89_22_pad_groupi_n_532 ,csa_tree_add_89_22_pad_groupi_n_617);
  or csa_tree_add_89_22_pad_groupi_g4995(csa_tree_add_89_22_pad_groupi_n_756 ,csa_tree_add_89_22_pad_groupi_n_455 ,csa_tree_add_89_22_pad_groupi_n_670);
  or csa_tree_add_89_22_pad_groupi_g4996(csa_tree_add_89_22_pad_groupi_n_755 ,csa_tree_add_89_22_pad_groupi_n_544 ,csa_tree_add_89_22_pad_groupi_n_660);
  or csa_tree_add_89_22_pad_groupi_g4997(csa_tree_add_89_22_pad_groupi_n_753 ,csa_tree_add_89_22_pad_groupi_n_486 ,csa_tree_add_89_22_pad_groupi_n_679);
  or csa_tree_add_89_22_pad_groupi_g4998(csa_tree_add_89_22_pad_groupi_n_751 ,csa_tree_add_89_22_pad_groupi_n_575 ,csa_tree_add_89_22_pad_groupi_n_619);
  or csa_tree_add_89_22_pad_groupi_g4999(csa_tree_add_89_22_pad_groupi_n_750 ,csa_tree_add_89_22_pad_groupi_n_522 ,csa_tree_add_89_22_pad_groupi_n_671);
  or csa_tree_add_89_22_pad_groupi_g5000(csa_tree_add_89_22_pad_groupi_n_748 ,csa_tree_add_89_22_pad_groupi_n_515 ,csa_tree_add_89_22_pad_groupi_n_631);
  or csa_tree_add_89_22_pad_groupi_g5001(csa_tree_add_89_22_pad_groupi_n_747 ,csa_tree_add_89_22_pad_groupi_n_573 ,csa_tree_add_89_22_pad_groupi_n_620);
  or csa_tree_add_89_22_pad_groupi_g5002(csa_tree_add_89_22_pad_groupi_n_746 ,csa_tree_add_89_22_pad_groupi_n_534 ,csa_tree_add_89_22_pad_groupi_n_643);
  or csa_tree_add_89_22_pad_groupi_g5003(csa_tree_add_89_22_pad_groupi_n_743 ,csa_tree_add_89_22_pad_groupi_n_481 ,csa_tree_add_89_22_pad_groupi_n_629);
  or csa_tree_add_89_22_pad_groupi_g5004(csa_tree_add_89_22_pad_groupi_n_742 ,csa_tree_add_89_22_pad_groupi_n_536 ,csa_tree_add_89_22_pad_groupi_n_650);
  or csa_tree_add_89_22_pad_groupi_g5006(csa_tree_add_89_22_pad_groupi_n_739 ,csa_tree_add_89_22_pad_groupi_n_564 ,csa_tree_add_89_22_pad_groupi_n_628);
  or csa_tree_add_89_22_pad_groupi_g5007(csa_tree_add_89_22_pad_groupi_n_737 ,csa_tree_add_89_22_pad_groupi_n_513 ,csa_tree_add_89_22_pad_groupi_n_603);
  or csa_tree_add_89_22_pad_groupi_g5008(csa_tree_add_89_22_pad_groupi_n_735 ,csa_tree_add_89_22_pad_groupi_n_553 ,csa_tree_add_89_22_pad_groupi_n_691);
  or csa_tree_add_89_22_pad_groupi_g5009(csa_tree_add_89_22_pad_groupi_n_733 ,csa_tree_add_89_22_pad_groupi_n_530 ,csa_tree_add_89_22_pad_groupi_n_622);
  or csa_tree_add_89_22_pad_groupi_g5010(csa_tree_add_89_22_pad_groupi_n_731 ,csa_tree_add_89_22_pad_groupi_n_463 ,csa_tree_add_89_22_pad_groupi_n_590);
  or csa_tree_add_89_22_pad_groupi_g5011(csa_tree_add_89_22_pad_groupi_n_729 ,csa_tree_add_89_22_pad_groupi_n_471 ,csa_tree_add_89_22_pad_groupi_n_610);
  or csa_tree_add_89_22_pad_groupi_g5012(csa_tree_add_89_22_pad_groupi_n_728 ,csa_tree_add_89_22_pad_groupi_n_520 ,csa_tree_add_89_22_pad_groupi_n_639);
  or csa_tree_add_89_22_pad_groupi_g5013(csa_tree_add_89_22_pad_groupi_n_726 ,csa_tree_add_89_22_pad_groupi_n_535 ,csa_tree_add_89_22_pad_groupi_n_690);
  or csa_tree_add_89_22_pad_groupi_g5014(csa_tree_add_89_22_pad_groupi_n_725 ,csa_tree_add_89_22_pad_groupi_n_538 ,csa_tree_add_89_22_pad_groupi_n_675);
  or csa_tree_add_89_22_pad_groupi_g5015(csa_tree_add_89_22_pad_groupi_n_723 ,csa_tree_add_89_22_pad_groupi_n_543 ,csa_tree_add_89_22_pad_groupi_n_676);
  or csa_tree_add_89_22_pad_groupi_g5016(csa_tree_add_89_22_pad_groupi_n_721 ,csa_tree_add_89_22_pad_groupi_n_542 ,csa_tree_add_89_22_pad_groupi_n_634);
  or csa_tree_add_89_22_pad_groupi_g5017(csa_tree_add_89_22_pad_groupi_n_720 ,csa_tree_add_89_22_pad_groupi_n_479 ,csa_tree_add_89_22_pad_groupi_n_644);
  or csa_tree_add_89_22_pad_groupi_g5018(csa_tree_add_89_22_pad_groupi_n_719 ,csa_tree_add_89_22_pad_groupi_n_521 ,csa_tree_add_89_22_pad_groupi_n_611);
  or csa_tree_add_89_22_pad_groupi_g5019(csa_tree_add_89_22_pad_groupi_n_718 ,csa_tree_add_89_22_pad_groupi_n_489 ,csa_tree_add_89_22_pad_groupi_n_609);
  or csa_tree_add_89_22_pad_groupi_g5020(csa_tree_add_89_22_pad_groupi_n_717 ,csa_tree_add_89_22_pad_groupi_n_549 ,csa_tree_add_89_22_pad_groupi_n_692);
  or csa_tree_add_89_22_pad_groupi_g5021(csa_tree_add_89_22_pad_groupi_n_716 ,csa_tree_add_89_22_pad_groupi_n_465 ,csa_tree_add_89_22_pad_groupi_n_613);
  or csa_tree_add_89_22_pad_groupi_g5022(csa_tree_add_89_22_pad_groupi_n_714 ,csa_tree_add_89_22_pad_groupi_n_474 ,csa_tree_add_89_22_pad_groupi_n_657);
  or csa_tree_add_89_22_pad_groupi_g5023(csa_tree_add_89_22_pad_groupi_n_713 ,csa_tree_add_89_22_pad_groupi_n_458 ,csa_tree_add_89_22_pad_groupi_n_667);
  not csa_tree_add_89_22_pad_groupi_g5024(csa_tree_add_89_22_pad_groupi_n_707 ,csa_tree_add_89_22_pad_groupi_n_706);
  not csa_tree_add_89_22_pad_groupi_g5025(csa_tree_add_89_22_pad_groupi_n_705 ,csa_tree_add_89_22_pad_groupi_n_704);
  nor csa_tree_add_89_22_pad_groupi_g5026(csa_tree_add_89_22_pad_groupi_n_703 ,csa_tree_add_89_22_pad_groupi_n_113 ,csa_tree_add_89_22_pad_groupi_n_218);
  nor csa_tree_add_89_22_pad_groupi_g5027(csa_tree_add_89_22_pad_groupi_n_702 ,in13[9] ,csa_tree_add_89_22_pad_groupi_n_358);
  nor csa_tree_add_89_22_pad_groupi_g5029(csa_tree_add_89_22_pad_groupi_n_700 ,in13[12] ,csa_tree_add_89_22_pad_groupi_n_579);
  nor csa_tree_add_89_22_pad_groupi_g5030(csa_tree_add_89_22_pad_groupi_n_699 ,csa_tree_add_89_22_pad_groupi_n_115 ,csa_tree_add_89_22_pad_groupi_n_189);
  and csa_tree_add_89_22_pad_groupi_g5031(csa_tree_add_89_22_pad_groupi_n_698 ,in9[5] ,csa_tree_add_89_22_pad_groupi_n_172);
  nor csa_tree_add_89_22_pad_groupi_g5032(csa_tree_add_89_22_pad_groupi_n_697 ,csa_tree_add_89_22_pad_groupi_n_119 ,csa_tree_add_89_22_pad_groupi_n_38);
  nor csa_tree_add_89_22_pad_groupi_g5033(csa_tree_add_89_22_pad_groupi_n_696 ,csa_tree_add_89_22_pad_groupi_n_93 ,csa_tree_add_89_22_pad_groupi_n_66);
  and csa_tree_add_89_22_pad_groupi_g5034(csa_tree_add_89_22_pad_groupi_n_695 ,in9[2] ,csa_tree_add_89_22_pad_groupi_n_133);
  and csa_tree_add_89_22_pad_groupi_g5035(csa_tree_add_89_22_pad_groupi_n_694 ,in9[10] ,csa_tree_add_89_22_pad_groupi_n_433);
  and csa_tree_add_89_22_pad_groupi_g5036(csa_tree_add_89_22_pad_groupi_n_693 ,in9[8] ,csa_tree_add_89_22_pad_groupi_n_287);
  and csa_tree_add_89_22_pad_groupi_g5037(csa_tree_add_89_22_pad_groupi_n_692 ,in9[14] ,csa_tree_add_89_22_pad_groupi_n_169);
  and csa_tree_add_89_22_pad_groupi_g5038(csa_tree_add_89_22_pad_groupi_n_691 ,in9[1] ,csa_tree_add_89_22_pad_groupi_n_168);
  and csa_tree_add_89_22_pad_groupi_g5039(csa_tree_add_89_22_pad_groupi_n_690 ,in9[5] ,csa_tree_add_89_22_pad_groupi_n_142);
  and csa_tree_add_89_22_pad_groupi_g5040(csa_tree_add_89_22_pad_groupi_n_689 ,in9[7] ,csa_tree_add_89_22_pad_groupi_n_126);
  and csa_tree_add_89_22_pad_groupi_g5041(csa_tree_add_89_22_pad_groupi_n_688 ,in9[11] ,csa_tree_add_89_22_pad_groupi_n_285);
  or csa_tree_add_89_22_pad_groupi_g5044(csa_tree_add_89_22_pad_groupi_n_685 ,csa_tree_add_89_22_pad_groupi_n_17 ,csa_tree_add_89_22_pad_groupi_n_118);
  or csa_tree_add_89_22_pad_groupi_g5046(csa_tree_add_89_22_pad_groupi_n_683 ,csa_tree_add_89_22_pad_groupi_n_149 ,csa_tree_add_89_22_pad_groupi_n_583);
  and csa_tree_add_89_22_pad_groupi_g5047(csa_tree_add_89_22_pad_groupi_n_682 ,in13[12] ,csa_tree_add_89_22_pad_groupi_n_579);
  and csa_tree_add_89_22_pad_groupi_g5048(csa_tree_add_89_22_pad_groupi_n_681 ,in9[11] ,csa_tree_add_89_22_pad_groupi_n_135);
  and csa_tree_add_89_22_pad_groupi_g5049(csa_tree_add_89_22_pad_groupi_n_680 ,in9[6] ,csa_tree_add_89_22_pad_groupi_n_445);
  nor csa_tree_add_89_22_pad_groupi_g5050(csa_tree_add_89_22_pad_groupi_n_679 ,csa_tree_add_89_22_pad_groupi_n_252 ,csa_tree_add_89_22_pad_groupi_n_223);
  and csa_tree_add_89_22_pad_groupi_g5052(csa_tree_add_89_22_pad_groupi_n_677 ,in9[3] ,csa_tree_add_89_22_pad_groupi_n_139);
  and csa_tree_add_89_22_pad_groupi_g5053(csa_tree_add_89_22_pad_groupi_n_676 ,in9[6] ,csa_tree_add_89_22_pad_groupi_n_136);
  and csa_tree_add_89_22_pad_groupi_g5054(csa_tree_add_89_22_pad_groupi_n_675 ,in9[4] ,csa_tree_add_89_22_pad_groupi_n_144);
  and csa_tree_add_89_22_pad_groupi_g5055(csa_tree_add_89_22_pad_groupi_n_674 ,in9[4] ,csa_tree_add_89_22_pad_groupi_n_138);
  nor csa_tree_add_89_22_pad_groupi_g5056(csa_tree_add_89_22_pad_groupi_n_673 ,csa_tree_add_89_22_pad_groupi_n_369 ,csa_tree_add_89_22_pad_groupi_n_581);
  and csa_tree_add_89_22_pad_groupi_g5057(csa_tree_add_89_22_pad_groupi_n_672 ,in9[12] ,csa_tree_add_89_22_pad_groupi_n_428);
  and csa_tree_add_89_22_pad_groupi_g5058(csa_tree_add_89_22_pad_groupi_n_671 ,in9[4] ,csa_tree_add_89_22_pad_groupi_n_124);
  and csa_tree_add_89_22_pad_groupi_g5059(csa_tree_add_89_22_pad_groupi_n_670 ,in9[9] ,csa_tree_add_89_22_pad_groupi_n_439);
  and csa_tree_add_89_22_pad_groupi_g5060(csa_tree_add_89_22_pad_groupi_n_669 ,in9[14] ,csa_tree_add_89_22_pad_groupi_n_288);
  and csa_tree_add_89_22_pad_groupi_g5062(csa_tree_add_89_22_pad_groupi_n_667 ,in9[14] ,csa_tree_add_89_22_pad_groupi_n_425);
  and csa_tree_add_89_22_pad_groupi_g5063(csa_tree_add_89_22_pad_groupi_n_666 ,in13[12] ,csa_tree_add_89_22_pad_groupi_n_280);
  and csa_tree_add_89_22_pad_groupi_g5064(csa_tree_add_89_22_pad_groupi_n_665 ,in9[7] ,csa_tree_add_89_22_pad_groupi_n_171);
  and csa_tree_add_89_22_pad_groupi_g5066(csa_tree_add_89_22_pad_groupi_n_663 ,csa_tree_add_89_22_pad_groupi_n_406 ,csa_tree_add_89_22_pad_groupi_n_583);
  and csa_tree_add_89_22_pad_groupi_g5067(csa_tree_add_89_22_pad_groupi_n_662 ,in9[7] ,csa_tree_add_89_22_pad_groupi_n_429);
  and csa_tree_add_89_22_pad_groupi_g5068(csa_tree_add_89_22_pad_groupi_n_661 ,in9[9] ,csa_tree_add_89_22_pad_groupi_n_145);
  and csa_tree_add_89_22_pad_groupi_g5069(csa_tree_add_89_22_pad_groupi_n_660 ,in9[14] ,csa_tree_add_89_22_pad_groupi_n_127);
  nor csa_tree_add_89_22_pad_groupi_g5070(csa_tree_add_89_22_pad_groupi_n_659 ,csa_tree_add_89_22_pad_groupi_n_112 ,csa_tree_add_89_22_pad_groupi_n_202);
  and csa_tree_add_89_22_pad_groupi_g5071(csa_tree_add_89_22_pad_groupi_n_658 ,in9[3] ,csa_tree_add_89_22_pad_groupi_n_133);
  nor csa_tree_add_89_22_pad_groupi_g5072(csa_tree_add_89_22_pad_groupi_n_657 ,csa_tree_add_89_22_pad_groupi_n_118 ,csa_tree_add_89_22_pad_groupi_n_215);
  or csa_tree_add_89_22_pad_groupi_g5073(csa_tree_add_89_22_pad_groupi_n_656 ,csa_tree_add_89_22_pad_groupi_n_373 ,csa_tree_add_89_22_pad_groupi_n_357);
  or csa_tree_add_89_22_pad_groupi_g5074(csa_tree_add_89_22_pad_groupi_n_655 ,csa_tree_add_89_22_pad_groupi_n_27 ,csa_tree_add_89_22_pad_groupi_n_427);
  and csa_tree_add_89_22_pad_groupi_g5075(csa_tree_add_89_22_pad_groupi_n_654 ,in9[11] ,csa_tree_add_89_22_pad_groupi_n_130);
  and csa_tree_add_89_22_pad_groupi_g5076(csa_tree_add_89_22_pad_groupi_n_653 ,in9[1] ,csa_tree_add_89_22_pad_groupi_n_147);
  nor csa_tree_add_89_22_pad_groupi_g5077(csa_tree_add_89_22_pad_groupi_n_652 ,csa_tree_add_89_22_pad_groupi_n_93 ,csa_tree_add_89_22_pad_groupi_n_74);
  and csa_tree_add_89_22_pad_groupi_g5078(csa_tree_add_89_22_pad_groupi_n_651 ,in9[13] ,csa_tree_add_89_22_pad_groupi_n_148);
  and csa_tree_add_89_22_pad_groupi_g5079(csa_tree_add_89_22_pad_groupi_n_650 ,in9[6] ,csa_tree_add_89_22_pad_groupi_n_148);
  and csa_tree_add_89_22_pad_groupi_g5080(csa_tree_add_89_22_pad_groupi_n_649 ,in9[12] ,csa_tree_add_89_22_pad_groupi_n_142);
  and csa_tree_add_89_22_pad_groupi_g5081(csa_tree_add_89_22_pad_groupi_n_648 ,in9[3] ,csa_tree_add_89_22_pad_groupi_n_129);
  and csa_tree_add_89_22_pad_groupi_g5082(csa_tree_add_89_22_pad_groupi_n_647 ,in9[4] ,csa_tree_add_89_22_pad_groupi_n_284);
  or csa_tree_add_89_22_pad_groupi_g5084(csa_tree_add_89_22_pad_groupi_n_706 ,csa_tree_add_89_22_pad_groupi_n_24 ,csa_tree_add_89_22_pad_groupi_n_502);
  or csa_tree_add_89_22_pad_groupi_g5085(csa_tree_add_89_22_pad_groupi_n_704 ,csa_tree_add_89_22_pad_groupi_n_24 ,csa_tree_add_89_22_pad_groupi_n_257);
  nor csa_tree_add_89_22_pad_groupi_g5086(csa_tree_add_89_22_pad_groupi_n_644 ,csa_tree_add_89_22_pad_groupi_n_113 ,csa_tree_add_89_22_pad_groupi_n_178);
  nor csa_tree_add_89_22_pad_groupi_g5087(csa_tree_add_89_22_pad_groupi_n_643 ,csa_tree_add_89_22_pad_groupi_n_160 ,csa_tree_add_89_22_pad_groupi_n_578);
  or csa_tree_add_89_22_pad_groupi_g5088(csa_tree_add_89_22_pad_groupi_n_642 ,csa_tree_add_89_22_pad_groupi_n_47 ,csa_tree_add_89_22_pad_groupi_n_497);
  and csa_tree_add_89_22_pad_groupi_g5090(csa_tree_add_89_22_pad_groupi_n_640 ,in9[6] ,csa_tree_add_89_22_pad_groupi_n_130);
  and csa_tree_add_89_22_pad_groupi_g5091(csa_tree_add_89_22_pad_groupi_n_639 ,in9[13] ,csa_tree_add_89_22_pad_groupi_n_171);
  nor csa_tree_add_89_22_pad_groupi_g5092(csa_tree_add_89_22_pad_groupi_n_638 ,csa_tree_add_89_22_pad_groupi_n_87 ,csa_tree_add_89_22_pad_groupi_n_434);
  and csa_tree_add_89_22_pad_groupi_g5093(csa_tree_add_89_22_pad_groupi_n_637 ,in9[10] ,csa_tree_add_89_22_pad_groupi_n_166);
  nor csa_tree_add_89_22_pad_groupi_g5095(csa_tree_add_89_22_pad_groupi_n_635 ,csa_tree_add_89_22_pad_groupi_n_96 ,csa_tree_add_89_22_pad_groupi_n_255);
  and csa_tree_add_89_22_pad_groupi_g5096(csa_tree_add_89_22_pad_groupi_n_634 ,in9[2] ,csa_tree_add_89_22_pad_groupi_n_168);
  and csa_tree_add_89_22_pad_groupi_g5097(csa_tree_add_89_22_pad_groupi_n_633 ,in9[13] ,csa_tree_add_89_22_pad_groupi_n_124);
  nor csa_tree_add_89_22_pad_groupi_g5099(csa_tree_add_89_22_pad_groupi_n_631 ,csa_tree_add_89_22_pad_groupi_n_231 ,csa_tree_add_89_22_pad_groupi_n_257);
  and csa_tree_add_89_22_pad_groupi_g5101(csa_tree_add_89_22_pad_groupi_n_629 ,in9[13] ,csa_tree_add_89_22_pad_groupi_n_287);
  and csa_tree_add_89_22_pad_groupi_g5102(csa_tree_add_89_22_pad_groupi_n_628 ,in9[11] ,csa_tree_add_89_22_pad_groupi_n_145);
  and csa_tree_add_89_22_pad_groupi_g5103(csa_tree_add_89_22_pad_groupi_n_627 ,in9[7] ,csa_tree_add_89_22_pad_groupi_n_141);
  nor csa_tree_add_89_22_pad_groupi_g5104(csa_tree_add_89_22_pad_groupi_n_626 ,csa_tree_add_89_22_pad_groupi_n_71 ,csa_tree_add_89_22_pad_groupi_n_507);
  and csa_tree_add_89_22_pad_groupi_g5105(csa_tree_add_89_22_pad_groupi_n_625 ,in9[7] ,csa_tree_add_89_22_pad_groupi_n_285);
  and csa_tree_add_89_22_pad_groupi_g5106(csa_tree_add_89_22_pad_groupi_n_624 ,in9[5] ,csa_tree_add_89_22_pad_groupi_n_165);
  and csa_tree_add_89_22_pad_groupi_g5107(csa_tree_add_89_22_pad_groupi_n_623 ,in9[10] ,csa_tree_add_89_22_pad_groupi_n_132);
  nor csa_tree_add_89_22_pad_groupi_g5108(csa_tree_add_89_22_pad_groupi_n_622 ,csa_tree_add_89_22_pad_groupi_n_159 ,csa_tree_add_89_22_pad_groupi_n_282);
  nor csa_tree_add_89_22_pad_groupi_g5109(csa_tree_add_89_22_pad_groupi_n_621 ,csa_tree_add_89_22_pad_groupi_n_98 ,csa_tree_add_89_22_pad_groupi_n_430);
  nor csa_tree_add_89_22_pad_groupi_g5110(csa_tree_add_89_22_pad_groupi_n_620 ,csa_tree_add_89_22_pad_groupi_n_194 ,csa_tree_add_89_22_pad_groupi_n_502);
  nor csa_tree_add_89_22_pad_groupi_g5111(csa_tree_add_89_22_pad_groupi_n_619 ,csa_tree_add_89_22_pad_groupi_n_116 ,csa_tree_add_89_22_pad_groupi_n_187);
  and csa_tree_add_89_22_pad_groupi_g5112(csa_tree_add_89_22_pad_groupi_n_618 ,in9[8] ,csa_tree_add_89_22_pad_groupi_n_165);
  and csa_tree_add_89_22_pad_groupi_g5113(csa_tree_add_89_22_pad_groupi_n_617 ,in9[8] ,csa_tree_add_89_22_pad_groupi_n_136);
  nor csa_tree_add_89_22_pad_groupi_g5114(csa_tree_add_89_22_pad_groupi_n_616 ,csa_tree_add_89_22_pad_groupi_n_119 ,csa_tree_add_89_22_pad_groupi_n_181);
  nor csa_tree_add_89_22_pad_groupi_g5117(csa_tree_add_89_22_pad_groupi_n_613 ,csa_tree_add_89_22_pad_groupi_n_204 ,csa_tree_add_89_22_pad_groupi_n_432);
  or csa_tree_add_89_22_pad_groupi_g5118(csa_tree_add_89_22_pad_groupi_n_612 ,csa_tree_add_89_22_pad_groupi_n_64 ,csa_tree_add_89_22_pad_groupi_n_438);
  and csa_tree_add_89_22_pad_groupi_g5119(csa_tree_add_89_22_pad_groupi_n_611 ,in9[8] ,csa_tree_add_89_22_pad_groupi_n_284);
  nor csa_tree_add_89_22_pad_groupi_g5120(csa_tree_add_89_22_pad_groupi_n_610 ,csa_tree_add_89_22_pad_groupi_n_116 ,csa_tree_add_89_22_pad_groupi_n_184);
  nor csa_tree_add_89_22_pad_groupi_g5121(csa_tree_add_89_22_pad_groupi_n_609 ,csa_tree_add_89_22_pad_groupi_n_91 ,csa_tree_add_89_22_pad_groupi_n_501);
  and csa_tree_add_89_22_pad_groupi_g5122(csa_tree_add_89_22_pad_groupi_n_608 ,in9[12] ,csa_tree_add_89_22_pad_groupi_n_166);
  and csa_tree_add_89_22_pad_groupi_g5123(csa_tree_add_89_22_pad_groupi_n_607 ,in9[11] ,csa_tree_add_89_22_pad_groupi_n_431);
  or csa_tree_add_89_22_pad_groupi_g5124(csa_tree_add_89_22_pad_groupi_n_606 ,csa_tree_add_89_22_pad_groupi_n_17 ,csa_tree_add_89_22_pad_groupi_n_255);
  and csa_tree_add_89_22_pad_groupi_g5125(csa_tree_add_89_22_pad_groupi_n_605 ,in9[9] ,csa_tree_add_89_22_pad_groupi_n_127);
  nor csa_tree_add_89_22_pad_groupi_g5126(csa_tree_add_89_22_pad_groupi_n_604 ,csa_tree_add_89_22_pad_groupi_n_211 ,csa_tree_add_89_22_pad_groupi_n_508);
  and csa_tree_add_89_22_pad_groupi_g5127(csa_tree_add_89_22_pad_groupi_n_603 ,in9[12] ,csa_tree_add_89_22_pad_groupi_n_169);
  and csa_tree_add_89_22_pad_groupi_g5128(csa_tree_add_89_22_pad_groupi_n_602 ,in9[1] ,csa_tree_add_89_22_pad_groupi_n_123);
  nor csa_tree_add_89_22_pad_groupi_g5130(csa_tree_add_89_22_pad_groupi_n_600 ,in13[12] ,csa_tree_add_89_22_pad_groupi_n_582);
  and csa_tree_add_89_22_pad_groupi_g5131(csa_tree_add_89_22_pad_groupi_n_599 ,in9[9] ,csa_tree_add_89_22_pad_groupi_n_139);
  nor csa_tree_add_89_22_pad_groupi_g5132(csa_tree_add_89_22_pad_groupi_n_598 ,csa_tree_add_89_22_pad_groupi_n_101 ,csa_tree_add_89_22_pad_groupi_n_508);
  or csa_tree_add_89_22_pad_groupi_g5135(csa_tree_add_89_22_pad_groupi_n_595 ,csa_tree_add_89_22_pad_groupi_n_55 ,csa_tree_add_89_22_pad_groupi_n_115);
  or csa_tree_add_89_22_pad_groupi_g5136(csa_tree_add_89_22_pad_groupi_n_594 ,csa_tree_add_89_22_pad_groupi_n_50 ,csa_tree_add_89_22_pad_groupi_n_426);
  nor csa_tree_add_89_22_pad_groupi_g5137(csa_tree_add_89_22_pad_groupi_n_593 ,in13[11] ,csa_tree_add_89_22_pad_groupi_n_580);
  and csa_tree_add_89_22_pad_groupi_g5139(csa_tree_add_89_22_pad_groupi_n_591 ,in9[10] ,csa_tree_add_89_22_pad_groupi_n_288);
  and csa_tree_add_89_22_pad_groupi_g5140(csa_tree_add_89_22_pad_groupi_n_590 ,in9[13] ,csa_tree_add_89_22_pad_groupi_n_435);
  and csa_tree_add_89_22_pad_groupi_g5141(csa_tree_add_89_22_pad_groupi_n_589 ,in9[10] ,csa_tree_add_89_22_pad_groupi_n_172);
  nor csa_tree_add_89_22_pad_groupi_g5142(csa_tree_add_89_22_pad_groupi_n_588 ,csa_tree_add_89_22_pad_groupi_n_158 ,csa_tree_add_89_22_pad_groupi_n_280);
  or csa_tree_add_89_22_pad_groupi_g5143(csa_tree_add_89_22_pad_groupi_n_587 ,csa_tree_add_89_22_pad_groupi_n_151 ,csa_tree_add_89_22_pad_groupi_n_580);
  or csa_tree_add_89_22_pad_groupi_g5144(csa_tree_add_89_22_pad_groupi_n_586 ,csa_tree_add_89_22_pad_groupi_n_15 ,csa_tree_add_89_22_pad_groupi_n_581);
  or csa_tree_add_89_22_pad_groupi_g5145(csa_tree_add_89_22_pad_groupi_n_646 ,csa_tree_add_89_22_pad_groupi_n_57 ,csa_tree_add_89_22_pad_groupi_n_493);
  or csa_tree_add_89_22_pad_groupi_g5146(csa_tree_add_89_22_pad_groupi_n_645 ,csa_tree_add_89_22_pad_groupi_n_42 ,csa_tree_add_89_22_pad_groupi_n_278);
  nor csa_tree_add_89_22_pad_groupi_g5150(csa_tree_add_89_22_pad_groupi_n_577 ,csa_tree_add_89_22_pad_groupi_n_183 ,csa_tree_add_89_22_pad_groupi_n_332);
  nor csa_tree_add_89_22_pad_groupi_g5151(csa_tree_add_89_22_pad_groupi_n_576 ,csa_tree_add_89_22_pad_groupi_n_42 ,csa_tree_add_89_22_pad_groupi_n_302);
  nor csa_tree_add_89_22_pad_groupi_g5152(csa_tree_add_89_22_pad_groupi_n_575 ,csa_tree_add_89_22_pad_groupi_n_233 ,csa_tree_add_89_22_pad_groupi_n_306);
  nor csa_tree_add_89_22_pad_groupi_g5153(csa_tree_add_89_22_pad_groupi_n_574 ,csa_tree_add_89_22_pad_groupi_n_193 ,csa_tree_add_89_22_pad_groupi_n_341);
  nor csa_tree_add_89_22_pad_groupi_g5154(csa_tree_add_89_22_pad_groupi_n_573 ,csa_tree_add_89_22_pad_groupi_n_84 ,csa_tree_add_89_22_pad_groupi_n_312);
  nor csa_tree_add_89_22_pad_groupi_g5163(csa_tree_add_89_22_pad_groupi_n_564 ,csa_tree_add_89_22_pad_groupi_n_78 ,csa_tree_add_89_22_pad_groupi_n_330);
  nor csa_tree_add_89_22_pad_groupi_g5170(csa_tree_add_89_22_pad_groupi_n_557 ,csa_tree_add_89_22_pad_groupi_n_71 ,csa_tree_add_89_22_pad_groupi_n_335);
  nor csa_tree_add_89_22_pad_groupi_g5171(csa_tree_add_89_22_pad_groupi_n_556 ,csa_tree_add_89_22_pad_groupi_n_101 ,csa_tree_add_89_22_pad_groupi_n_315);
  nor csa_tree_add_89_22_pad_groupi_g5172(csa_tree_add_89_22_pad_groupi_n_555 ,csa_tree_add_89_22_pad_groupi_n_186 ,csa_tree_add_89_22_pad_groupi_n_336);
  nor csa_tree_add_89_22_pad_groupi_g5173(csa_tree_add_89_22_pad_groupi_n_554 ,csa_tree_add_89_22_pad_groupi_n_177 ,csa_tree_add_89_22_pad_groupi_n_309);
  nor csa_tree_add_89_22_pad_groupi_g5174(csa_tree_add_89_22_pad_groupi_n_553 ,csa_tree_add_89_22_pad_groupi_n_244 ,csa_tree_add_89_22_pad_groupi_n_320);
  nor csa_tree_add_89_22_pad_groupi_g5175(csa_tree_add_89_22_pad_groupi_n_552 ,csa_tree_add_89_22_pad_groupi_n_247 ,csa_tree_add_89_22_pad_groupi_n_323);
  nor csa_tree_add_89_22_pad_groupi_g5176(csa_tree_add_89_22_pad_groupi_n_551 ,csa_tree_add_89_22_pad_groupi_n_67 ,csa_tree_add_89_22_pad_groupi_n_317);
  nor csa_tree_add_89_22_pad_groupi_g5177(csa_tree_add_89_22_pad_groupi_n_550 ,csa_tree_add_89_22_pad_groupi_n_175 ,csa_tree_add_89_22_pad_groupi_n_339);
  nor csa_tree_add_89_22_pad_groupi_g5178(csa_tree_add_89_22_pad_groupi_n_549 ,csa_tree_add_89_22_pad_groupi_n_85 ,csa_tree_add_89_22_pad_groupi_n_321);
  nor csa_tree_add_89_22_pad_groupi_g5179(csa_tree_add_89_22_pad_groupi_n_548 ,csa_tree_add_89_22_pad_groupi_n_88 ,csa_tree_add_89_22_pad_groupi_n_305);
  nor csa_tree_add_89_22_pad_groupi_g5180(csa_tree_add_89_22_pad_groupi_n_547 ,csa_tree_add_89_22_pad_groupi_n_197 ,csa_tree_add_89_22_pad_groupi_n_323);
  nor csa_tree_add_89_22_pad_groupi_g5181(csa_tree_add_89_22_pad_groupi_n_546 ,csa_tree_add_89_22_pad_groupi_n_100 ,csa_tree_add_89_22_pad_groupi_n_326);
  nor csa_tree_add_89_22_pad_groupi_g5182(csa_tree_add_89_22_pad_groupi_n_545 ,csa_tree_add_89_22_pad_groupi_n_53 ,csa_tree_add_89_22_pad_groupi_n_327);
  nor csa_tree_add_89_22_pad_groupi_g5183(csa_tree_add_89_22_pad_groupi_n_544 ,csa_tree_add_89_22_pad_groupi_n_187 ,csa_tree_add_89_22_pad_groupi_n_326);
  nor csa_tree_add_89_22_pad_groupi_g5184(csa_tree_add_89_22_pad_groupi_n_543 ,csa_tree_add_89_22_pad_groupi_n_196 ,csa_tree_add_89_22_pad_groupi_n_317);
  nor csa_tree_add_89_22_pad_groupi_g5185(csa_tree_add_89_22_pad_groupi_n_542 ,csa_tree_add_89_22_pad_groupi_n_217 ,csa_tree_add_89_22_pad_groupi_n_318);
  nor csa_tree_add_89_22_pad_groupi_g5186(csa_tree_add_89_22_pad_groupi_n_541 ,csa_tree_add_89_22_pad_groupi_n_209 ,csa_tree_add_89_22_pad_groupi_n_344);
  nor csa_tree_add_89_22_pad_groupi_g5187(csa_tree_add_89_22_pad_groupi_n_540 ,csa_tree_add_89_22_pad_groupi_n_229 ,csa_tree_add_89_22_pad_groupi_n_324);
  nor csa_tree_add_89_22_pad_groupi_g5188(csa_tree_add_89_22_pad_groupi_n_539 ,csa_tree_add_89_22_pad_groupi_n_41 ,csa_tree_add_89_22_pad_groupi_n_335);
  nor csa_tree_add_89_22_pad_groupi_g5189(csa_tree_add_89_22_pad_groupi_n_538 ,csa_tree_add_89_22_pad_groupi_n_36 ,csa_tree_add_89_22_pad_groupi_n_336);
  nor csa_tree_add_89_22_pad_groupi_g5190(csa_tree_add_89_22_pad_groupi_n_537 ,csa_tree_add_89_22_pad_groupi_n_79 ,csa_tree_add_89_22_pad_groupi_n_324);
  nor csa_tree_add_89_22_pad_groupi_g5191(csa_tree_add_89_22_pad_groupi_n_536 ,csa_tree_add_89_22_pad_groupi_n_204 ,csa_tree_add_89_22_pad_groupi_n_345);
  nor csa_tree_add_89_22_pad_groupi_g5192(csa_tree_add_89_22_pad_groupi_n_535 ,csa_tree_add_89_22_pad_groupi_n_28 ,csa_tree_add_89_22_pad_groupi_n_329);
  nor csa_tree_add_89_22_pad_groupi_g5193(csa_tree_add_89_22_pad_groupi_n_534 ,csa_tree_add_89_22_pad_groupi_n_194 ,csa_tree_add_89_22_pad_groupi_n_327);
  nor csa_tree_add_89_22_pad_groupi_g5194(csa_tree_add_89_22_pad_groupi_n_533 ,csa_tree_add_89_22_pad_groupi_n_191 ,csa_tree_add_89_22_pad_groupi_n_338);
  nor csa_tree_add_89_22_pad_groupi_g5195(csa_tree_add_89_22_pad_groupi_n_532 ,csa_tree_add_89_22_pad_groupi_n_184 ,csa_tree_add_89_22_pad_groupi_n_318);
  or csa_tree_add_89_22_pad_groupi_g5196(csa_tree_add_89_22_pad_groupi_n_531 ,csa_tree_add_89_22_pad_groupi_n_174 ,csa_tree_add_89_22_pad_groupi_n_305);
  nor csa_tree_add_89_22_pad_groupi_g5197(csa_tree_add_89_22_pad_groupi_n_530 ,csa_tree_add_89_22_pad_groupi_n_39 ,csa_tree_add_89_22_pad_groupi_n_330);
  nor csa_tree_add_89_22_pad_groupi_g5198(csa_tree_add_89_22_pad_groupi_n_529 ,csa_tree_add_89_22_pad_groupi_n_243 ,csa_tree_add_89_22_pad_groupi_n_344);
  nor csa_tree_add_89_22_pad_groupi_g5199(csa_tree_add_89_22_pad_groupi_n_528 ,csa_tree_add_89_22_pad_groupi_n_91 ,csa_tree_add_89_22_pad_groupi_n_345);
  nor csa_tree_add_89_22_pad_groupi_g5200(csa_tree_add_89_22_pad_groupi_n_527 ,csa_tree_add_89_22_pad_groupi_n_231 ,csa_tree_add_89_22_pad_groupi_n_321);
  nor csa_tree_add_89_22_pad_groupi_g5201(csa_tree_add_89_22_pad_groupi_n_526 ,csa_tree_add_89_22_pad_groupi_n_217 ,csa_tree_add_89_22_pad_groupi_n_265);
  nor csa_tree_add_89_22_pad_groupi_g5202(csa_tree_add_89_22_pad_groupi_n_525 ,csa_tree_add_89_22_pad_groupi_n_64 ,csa_tree_add_89_22_pad_groupi_n_311);
  nor csa_tree_add_89_22_pad_groupi_g5203(csa_tree_add_89_22_pad_groupi_n_524 ,csa_tree_add_89_22_pad_groupi_n_55 ,csa_tree_add_89_22_pad_groupi_n_269);
  nor csa_tree_add_89_22_pad_groupi_g5204(csa_tree_add_89_22_pad_groupi_n_523 ,csa_tree_add_89_22_pad_groupi_n_76 ,csa_tree_add_89_22_pad_groupi_n_312);
  nor csa_tree_add_89_22_pad_groupi_g5205(csa_tree_add_89_22_pad_groupi_n_522 ,csa_tree_add_89_22_pad_groupi_n_201 ,csa_tree_add_89_22_pad_groupi_n_339);
  nor csa_tree_add_89_22_pad_groupi_g5206(csa_tree_add_89_22_pad_groupi_n_521 ,csa_tree_add_89_22_pad_groupi_n_22 ,csa_tree_add_89_22_pad_groupi_n_275);
  nor csa_tree_add_89_22_pad_groupi_g5207(csa_tree_add_89_22_pad_groupi_n_520 ,csa_tree_add_89_22_pad_groupi_n_222 ,csa_tree_add_89_22_pad_groupi_n_262);
  nor csa_tree_add_89_22_pad_groupi_g5208(csa_tree_add_89_22_pad_groupi_n_519 ,csa_tree_add_89_22_pad_groupi_n_50 ,csa_tree_add_89_22_pad_groupi_n_272);
  or csa_tree_add_89_22_pad_groupi_g5209(csa_tree_add_89_22_pad_groupi_n_518 ,csa_tree_add_89_22_pad_groupi_n_21 ,csa_tree_add_89_22_pad_groupi_n_266);
  nor csa_tree_add_89_22_pad_groupi_g5210(csa_tree_add_89_22_pad_groupi_n_517 ,csa_tree_add_89_22_pad_groupi_n_178 ,csa_tree_add_89_22_pad_groupi_n_274);
  nor csa_tree_add_89_22_pad_groupi_g5211(csa_tree_add_89_22_pad_groupi_n_516 ,csa_tree_add_89_22_pad_groupi_n_225 ,csa_tree_add_89_22_pad_groupi_n_263);
  nor csa_tree_add_89_22_pad_groupi_g5212(csa_tree_add_89_22_pad_groupi_n_515 ,csa_tree_add_89_22_pad_groupi_n_47 ,csa_tree_add_89_22_pad_groupi_n_268);
  nor csa_tree_add_89_22_pad_groupi_g5213(csa_tree_add_89_22_pad_groupi_n_514 ,csa_tree_add_89_22_pad_groupi_n_197 ,csa_tree_add_89_22_pad_groupi_n_333);
  nor csa_tree_add_89_22_pad_groupi_g5214(csa_tree_add_89_22_pad_groupi_n_513 ,csa_tree_add_89_22_pad_groupi_n_227 ,csa_tree_add_89_22_pad_groupi_n_320);
  nor csa_tree_add_89_22_pad_groupi_g5215(csa_tree_add_89_22_pad_groupi_n_512 ,csa_tree_add_89_22_pad_groupi_n_59 ,csa_tree_add_89_22_pad_groupi_n_342);
  or csa_tree_add_89_22_pad_groupi_g5217(csa_tree_add_89_22_pad_groupi_n_583 ,csa_tree_add_89_22_pad_groupi_n_121 ,csa_tree_add_89_22_pad_groupi_n_424);
  or csa_tree_add_89_22_pad_groupi_g5218(csa_tree_add_89_22_pad_groupi_n_582 ,csa_tree_add_89_22_pad_groupi_n_162 ,csa_tree_add_89_22_pad_groupi_n_402);
  or csa_tree_add_89_22_pad_groupi_g5219(csa_tree_add_89_22_pad_groupi_n_581 ,csa_tree_add_89_22_pad_groupi_n_121 ,csa_tree_add_89_22_pad_groupi_n_109);
  or csa_tree_add_89_22_pad_groupi_g5220(csa_tree_add_89_22_pad_groupi_n_580 ,csa_tree_add_89_22_pad_groupi_n_162 ,csa_tree_add_89_22_pad_groupi_n_404);
  or csa_tree_add_89_22_pad_groupi_g5221(csa_tree_add_89_22_pad_groupi_n_579 ,csa_tree_add_89_22_pad_groupi_n_163 ,csa_tree_add_89_22_pad_groupi_n_403);
  not csa_tree_add_89_22_pad_groupi_g5223(csa_tree_add_89_22_pad_groupi_n_510 ,csa_tree_add_89_22_pad_groupi_n_505);
  not csa_tree_add_89_22_pad_groupi_g5224(csa_tree_add_89_22_pad_groupi_n_509 ,csa_tree_add_89_22_pad_groupi_n_505);
  not csa_tree_add_89_22_pad_groupi_g5225(csa_tree_add_89_22_pad_groupi_n_508 ,csa_tree_add_89_22_pad_groupi_n_506);
  not csa_tree_add_89_22_pad_groupi_g5226(csa_tree_add_89_22_pad_groupi_n_507 ,csa_tree_add_89_22_pad_groupi_n_506);
  not csa_tree_add_89_22_pad_groupi_g5227(csa_tree_add_89_22_pad_groupi_n_506 ,csa_tree_add_89_22_pad_groupi_n_505);
  not csa_tree_add_89_22_pad_groupi_g5228(csa_tree_add_89_22_pad_groupi_n_504 ,csa_tree_add_89_22_pad_groupi_n_499);
  not csa_tree_add_89_22_pad_groupi_g5229(csa_tree_add_89_22_pad_groupi_n_503 ,csa_tree_add_89_22_pad_groupi_n_499);
  not csa_tree_add_89_22_pad_groupi_g5230(csa_tree_add_89_22_pad_groupi_n_502 ,csa_tree_add_89_22_pad_groupi_n_500);
  not csa_tree_add_89_22_pad_groupi_g5231(csa_tree_add_89_22_pad_groupi_n_501 ,csa_tree_add_89_22_pad_groupi_n_500);
  not csa_tree_add_89_22_pad_groupi_g5232(csa_tree_add_89_22_pad_groupi_n_500 ,csa_tree_add_89_22_pad_groupi_n_499);
  not csa_tree_add_89_22_pad_groupi_g5233(csa_tree_add_89_22_pad_groupi_n_498 ,csa_tree_add_89_22_pad_groupi_n_278);
  not csa_tree_add_89_22_pad_groupi_g5234(csa_tree_add_89_22_pad_groupi_n_496 ,csa_tree_add_89_22_pad_groupi_n_497);
  not csa_tree_add_89_22_pad_groupi_g5235(csa_tree_add_89_22_pad_groupi_n_495 ,csa_tree_add_89_22_pad_groupi_n_493);
  not csa_tree_add_89_22_pad_groupi_g5236(csa_tree_add_89_22_pad_groupi_n_494 ,csa_tree_add_89_22_pad_groupi_n_493);
  or csa_tree_add_89_22_pad_groupi_g5237(csa_tree_add_89_22_pad_groupi_n_492 ,csa_tree_add_89_22_pad_groupi_n_27 ,csa_tree_add_89_22_pad_groupi_n_311);
  nor csa_tree_add_89_22_pad_groupi_g5238(csa_tree_add_89_22_pad_groupi_n_491 ,csa_tree_add_89_22_pad_groupi_n_180 ,csa_tree_add_89_22_pad_groupi_n_329);
  nor csa_tree_add_89_22_pad_groupi_g5239(csa_tree_add_89_22_pad_groupi_n_490 ,csa_tree_add_89_22_pad_groupi_n_220 ,csa_tree_add_89_22_pad_groupi_n_271);
  nor csa_tree_add_89_22_pad_groupi_g5240(csa_tree_add_89_22_pad_groupi_n_489 ,csa_tree_add_89_22_pad_groupi_n_82 ,csa_tree_add_89_22_pad_groupi_n_275);
  nor csa_tree_add_89_22_pad_groupi_g5241(csa_tree_add_89_22_pad_groupi_n_488 ,csa_tree_add_89_22_pad_groupi_n_181 ,csa_tree_add_89_22_pad_groupi_n_309);
  nor csa_tree_add_89_22_pad_groupi_g5242(csa_tree_add_89_22_pad_groupi_n_487 ,csa_tree_add_89_22_pad_groupi_n_88 ,csa_tree_add_89_22_pad_groupi_n_341);
  nor csa_tree_add_89_22_pad_groupi_g5243(csa_tree_add_89_22_pad_groupi_n_486 ,csa_tree_add_89_22_pad_groupi_n_227 ,csa_tree_add_89_22_pad_groupi_n_306);
  or csa_tree_add_89_22_pad_groupi_g5244(csa_tree_add_89_22_pad_groupi_n_485 ,csa_tree_add_89_22_pad_groupi_n_30 ,csa_tree_add_89_22_pad_groupi_n_302);
  nor csa_tree_add_89_22_pad_groupi_g5245(csa_tree_add_89_22_pad_groupi_n_484 ,csa_tree_add_89_22_pad_groupi_n_174 ,csa_tree_add_89_22_pad_groupi_n_315);
  or csa_tree_add_89_22_pad_groupi_g5246(csa_tree_add_89_22_pad_groupi_n_483 ,csa_tree_add_89_22_pad_groupi_n_30 ,csa_tree_add_89_22_pad_groupi_n_263);
  nor csa_tree_add_89_22_pad_groupi_g5247(csa_tree_add_89_22_pad_groupi_n_482 ,csa_tree_add_89_22_pad_groupi_n_96 ,csa_tree_add_89_22_pad_groupi_n_338);
  nor csa_tree_add_89_22_pad_groupi_g5248(csa_tree_add_89_22_pad_groupi_n_481 ,csa_tree_add_89_22_pad_groupi_n_233 ,csa_tree_add_89_22_pad_groupi_n_269);
  nor csa_tree_add_89_22_pad_groupi_g5249(csa_tree_add_89_22_pad_groupi_n_480 ,csa_tree_add_89_22_pad_groupi_n_25 ,csa_tree_add_89_22_pad_groupi_n_272);
  nor csa_tree_add_89_22_pad_groupi_g5250(csa_tree_add_89_22_pad_groupi_n_479 ,csa_tree_add_89_22_pad_groupi_n_214 ,csa_tree_add_89_22_pad_groupi_n_266);
  nor csa_tree_add_89_22_pad_groupi_g5251(csa_tree_add_89_22_pad_groupi_n_478 ,csa_tree_add_89_22_pad_groupi_n_235 ,csa_tree_add_89_22_pad_groupi_n_332);
  nor csa_tree_add_89_22_pad_groupi_g5252(csa_tree_add_89_22_pad_groupi_n_477 ,csa_tree_add_89_22_pad_groupi_n_73 ,csa_tree_add_89_22_pad_groupi_n_342);
  nor csa_tree_add_89_22_pad_groupi_g5253(csa_tree_add_89_22_pad_groupi_n_476 ,csa_tree_add_89_22_pad_groupi_n_206 ,csa_tree_add_89_22_pad_groupi_n_314);
  nor csa_tree_add_89_22_pad_groupi_g5254(csa_tree_add_89_22_pad_groupi_n_475 ,csa_tree_add_89_22_pad_groupi_n_69 ,csa_tree_add_89_22_pad_groupi_n_308);
  nor csa_tree_add_89_22_pad_groupi_g5255(csa_tree_add_89_22_pad_groupi_n_474 ,csa_tree_add_89_22_pad_groupi_n_209 ,csa_tree_add_89_22_pad_groupi_n_303);
  nor csa_tree_add_89_22_pad_groupi_g5256(csa_tree_add_89_22_pad_groupi_n_473 ,csa_tree_add_89_22_pad_groupi_n_76 ,csa_tree_add_89_22_pad_groupi_n_314);
  or csa_tree_add_89_22_pad_groupi_g5257(csa_tree_add_89_22_pad_groupi_n_472 ,csa_tree_add_89_22_pad_groupi_n_45 ,csa_tree_add_89_22_pad_groupi_n_308);
  nor csa_tree_add_89_22_pad_groupi_g5258(csa_tree_add_89_22_pad_groupi_n_471 ,csa_tree_add_89_22_pad_groupi_n_211 ,csa_tree_add_89_22_pad_groupi_n_303);
  nor csa_tree_add_89_22_pad_groupi_g5259(csa_tree_add_89_22_pad_groupi_n_470 ,csa_tree_add_89_22_pad_groupi_n_67 ,csa_tree_add_89_22_pad_groupi_n_333);
  nor csa_tree_add_89_22_pad_groupi_g5260(csa_tree_add_89_22_pad_groupi_n_469 ,csa_tree_add_89_22_pad_groupi_n_180 ,csa_tree_add_89_22_pad_groupi_n_300);
  nor csa_tree_add_89_22_pad_groupi_g5261(csa_tree_add_89_22_pad_groupi_n_468 ,csa_tree_add_89_22_pad_groupi_n_177 ,csa_tree_add_89_22_pad_groupi_n_399);
  nor csa_tree_add_89_22_pad_groupi_g5262(csa_tree_add_89_22_pad_groupi_n_467 ,csa_tree_add_89_22_pad_groupi_n_52 ,csa_tree_add_89_22_pad_groupi_n_291);
  nor csa_tree_add_89_22_pad_groupi_g5263(csa_tree_add_89_22_pad_groupi_n_466 ,csa_tree_add_89_22_pad_groupi_n_45 ,csa_tree_add_89_22_pad_groupi_n_290);
  nor csa_tree_add_89_22_pad_groupi_g5264(csa_tree_add_89_22_pad_groupi_n_465 ,csa_tree_add_89_22_pad_groupi_n_175 ,csa_tree_add_89_22_pad_groupi_n_297);
  or csa_tree_add_89_22_pad_groupi_g5265(csa_tree_add_89_22_pad_groupi_n_464 ,csa_tree_add_89_22_pad_groupi_n_36 ,csa_tree_add_89_22_pad_groupi_n_296);
  nor csa_tree_add_89_22_pad_groupi_g5266(csa_tree_add_89_22_pad_groupi_n_463 ,csa_tree_add_89_22_pad_groupi_n_90 ,csa_tree_add_89_22_pad_groupi_n_260);
  nor csa_tree_add_89_22_pad_groupi_g5267(csa_tree_add_89_22_pad_groupi_n_462 ,csa_tree_add_89_22_pad_groupi_n_212 ,csa_tree_add_89_22_pad_groupi_n_299);
  nor csa_tree_add_89_22_pad_groupi_g5268(csa_tree_add_89_22_pad_groupi_n_461 ,csa_tree_add_89_22_pad_groupi_n_95 ,csa_tree_add_89_22_pad_groupi_n_299);
  or csa_tree_add_89_22_pad_groupi_g5269(csa_tree_add_89_22_pad_groupi_n_460 ,csa_tree_add_89_22_pad_groupi_n_39 ,csa_tree_add_89_22_pad_groupi_n_290);
  nor csa_tree_add_89_22_pad_groupi_g5271(csa_tree_add_89_22_pad_groupi_n_458 ,csa_tree_add_89_22_pad_groupi_n_186 ,csa_tree_add_89_22_pad_groupi_n_300);
  or csa_tree_add_89_22_pad_groupi_g5272(csa_tree_add_89_22_pad_groupi_n_457 ,csa_tree_add_89_22_pad_groupi_n_21 ,csa_tree_add_89_22_pad_groupi_n_291);
  nor csa_tree_add_89_22_pad_groupi_g5273(csa_tree_add_89_22_pad_groupi_n_456 ,csa_tree_add_89_22_pad_groupi_n_98 ,csa_tree_add_89_22_pad_groupi_n_296);
  nor csa_tree_add_89_22_pad_groupi_g5274(csa_tree_add_89_22_pad_groupi_n_455 ,csa_tree_add_89_22_pad_groupi_n_207 ,csa_tree_add_89_22_pad_groupi_n_297);
  nor csa_tree_add_89_22_pad_groupi_g5284(csa_tree_add_89_22_pad_groupi_n_445 ,csa_tree_add_89_22_pad_groupi_n_106 ,csa_tree_add_89_22_pad_groupi_n_294);
  nor csa_tree_add_89_22_pad_groupi_g5290(csa_tree_add_89_22_pad_groupi_n_439 ,csa_tree_add_89_22_pad_groupi_n_109 ,csa_tree_add_89_22_pad_groupi_n_241);
  or csa_tree_add_89_22_pad_groupi_g5291(csa_tree_add_89_22_pad_groupi_n_438 ,csa_tree_add_89_22_pad_groupi_n_32 ,csa_tree_add_89_22_pad_groupi_n_103);
  nor csa_tree_add_89_22_pad_groupi_g5294(csa_tree_add_89_22_pad_groupi_n_435 ,csa_tree_add_89_22_pad_groupi_n_107 ,csa_tree_add_89_22_pad_groupi_n_240);
  or csa_tree_add_89_22_pad_groupi_g5295(csa_tree_add_89_22_pad_groupi_n_434 ,csa_tree_add_89_22_pad_groupi_n_293 ,csa_tree_add_89_22_pad_groupi_n_110);
  nor csa_tree_add_89_22_pad_groupi_g5296(csa_tree_add_89_22_pad_groupi_n_433 ,csa_tree_add_89_22_pad_groupi_n_103 ,csa_tree_add_89_22_pad_groupi_n_294);
  or csa_tree_add_89_22_pad_groupi_g5297(csa_tree_add_89_22_pad_groupi_n_432 ,csa_tree_add_89_22_pad_groupi_n_13 ,csa_tree_add_89_22_pad_groupi_n_61);
  nor csa_tree_add_89_22_pad_groupi_g5298(csa_tree_add_89_22_pad_groupi_n_431 ,csa_tree_add_89_22_pad_groupi_n_110 ,csa_tree_add_89_22_pad_groupi_n_238);
  or csa_tree_add_89_22_pad_groupi_g5299(csa_tree_add_89_22_pad_groupi_n_430 ,csa_tree_add_89_22_pad_groupi_n_13 ,csa_tree_add_89_22_pad_groupi_n_104);
  nor csa_tree_add_89_22_pad_groupi_g5300(csa_tree_add_89_22_pad_groupi_n_429 ,csa_tree_add_89_22_pad_groupi_n_61 ,csa_tree_add_89_22_pad_groupi_n_32);
  nor csa_tree_add_89_22_pad_groupi_g5301(csa_tree_add_89_22_pad_groupi_n_428 ,csa_tree_add_89_22_pad_groupi_n_249 ,csa_tree_add_89_22_pad_groupi_n_34);
  or csa_tree_add_89_22_pad_groupi_g5302(csa_tree_add_89_22_pad_groupi_n_427 ,csa_tree_add_89_22_pad_groupi_n_15 ,csa_tree_add_89_22_pad_groupi_n_106);
  or csa_tree_add_89_22_pad_groupi_g5303(csa_tree_add_89_22_pad_groupi_n_426 ,csa_tree_add_89_22_pad_groupi_n_34 ,csa_tree_add_89_22_pad_groupi_n_107);
  nor csa_tree_add_89_22_pad_groupi_g5304(csa_tree_add_89_22_pad_groupi_n_425 ,csa_tree_add_89_22_pad_groupi_n_104 ,csa_tree_add_89_22_pad_groupi_n_237);
  or csa_tree_add_89_22_pad_groupi_g5305(csa_tree_add_89_22_pad_groupi_n_511 ,csa_tree_add_89_22_pad_groupi_n_154 ,csa_tree_add_89_22_pad_groupi_n_424);
  or csa_tree_add_89_22_pad_groupi_g5306(csa_tree_add_89_22_pad_groupi_n_505 ,csa_tree_add_89_22_pad_groupi_n_150 ,csa_tree_add_89_22_pad_groupi_n_403);
  or csa_tree_add_89_22_pad_groupi_g5307(csa_tree_add_89_22_pad_groupi_n_499 ,csa_tree_add_89_22_pad_groupi_n_155 ,csa_tree_add_89_22_pad_groupi_n_402);
  or csa_tree_add_89_22_pad_groupi_g5309(csa_tree_add_89_22_pad_groupi_n_493 ,csa_tree_add_89_22_pad_groupi_n_152 ,csa_tree_add_89_22_pad_groupi_n_404);
  not csa_tree_add_89_22_pad_groupi_g5311(csa_tree_add_89_22_pad_groupi_n_423 ,csa_tree_add_89_22_pad_groupi_n_158);
  not csa_tree_add_89_22_pad_groupi_g5312(csa_tree_add_89_22_pad_groupi_n_422 ,csa_tree_add_89_22_pad_groupi_n_155);
  not csa_tree_add_89_22_pad_groupi_g5315(csa_tree_add_89_22_pad_groupi_n_419 ,csa_tree_add_89_22_pad_groupi_n_154);
  not csa_tree_add_89_22_pad_groupi_g5317(csa_tree_add_89_22_pad_groupi_n_418 ,csa_tree_add_89_22_pad_groupi_n_149);
  not csa_tree_add_89_22_pad_groupi_g5319(csa_tree_add_89_22_pad_groupi_n_416 ,csa_tree_add_89_22_pad_groupi_n_152);
  not csa_tree_add_89_22_pad_groupi_g5321(csa_tree_add_89_22_pad_groupi_n_415 ,csa_tree_add_89_22_pad_groupi_n_151);
  not csa_tree_add_89_22_pad_groupi_g5323(csa_tree_add_89_22_pad_groupi_n_414 ,csa_tree_add_89_22_pad_groupi_n_160);
  not csa_tree_add_89_22_pad_groupi_g5324(csa_tree_add_89_22_pad_groupi_n_413 ,csa_tree_add_89_22_pad_groupi_n_153);
  not csa_tree_add_89_22_pad_groupi_g5327(csa_tree_add_89_22_pad_groupi_n_411 ,csa_tree_add_89_22_pad_groupi_n_159);
  not csa_tree_add_89_22_pad_groupi_g5328(csa_tree_add_89_22_pad_groupi_n_410 ,csa_tree_add_89_22_pad_groupi_n_150);
  or csa_tree_add_89_22_pad_groupi_g5331(csa_tree_add_89_22_pad_groupi_n_406 ,in13[10] ,in13[9]);
  and csa_tree_add_89_22_pad_groupi_g5332(csa_tree_add_89_22_pad_groupi_n_424 ,csa_tree_add_89_22_pad_groupi_n_375 ,csa_tree_add_89_22_pad_groupi_n_388);
  and csa_tree_add_89_22_pad_groupi_g5333(csa_tree_add_89_22_pad_groupi_n_421 ,n_719 ,n_726);
  and csa_tree_add_89_22_pad_groupi_g5334(csa_tree_add_89_22_pad_groupi_n_420 ,in14[0] ,n_728);
  and csa_tree_add_89_22_pad_groupi_g5335(csa_tree_add_89_22_pad_groupi_n_417 ,n_720 ,n_727);
  and csa_tree_add_89_22_pad_groupi_g5337(csa_tree_add_89_22_pad_groupi_n_409 ,n_718 ,n_725);
  not csa_tree_add_89_22_pad_groupi_g5339(csa_tree_add_89_22_pad_groupi_n_399 ,csa_tree_add_89_22_pad_groupi_n_293);
  not csa_tree_add_89_22_pad_groupi_g5340(csa_tree_add_89_22_pad_groupi_n_398 ,csa_tree_add_89_22_pad_groupi_n_395);
  not csa_tree_add_89_22_pad_groupi_g5341(csa_tree_add_89_22_pad_groupi_n_397 ,csa_tree_add_89_22_pad_groupi_n_258);
  not csa_tree_add_89_22_pad_groupi_g5345(csa_tree_add_89_22_pad_groupi_n_396 ,csa_tree_add_89_22_pad_groupi_n_395);
  and csa_tree_add_89_22_pad_groupi_g5346(csa_tree_add_89_22_pad_groupi_n_394 ,in13[10] ,in13[9]);
  and csa_tree_add_89_22_pad_groupi_g5348(csa_tree_add_89_22_pad_groupi_n_404 ,csa_tree_add_89_22_pad_groupi_n_391 ,csa_tree_add_89_22_pad_groupi_n_393);
  and csa_tree_add_89_22_pad_groupi_g5349(csa_tree_add_89_22_pad_groupi_n_403 ,csa_tree_add_89_22_pad_groupi_n_378 ,csa_tree_add_89_22_pad_groupi_n_377);
  and csa_tree_add_89_22_pad_groupi_g5350(csa_tree_add_89_22_pad_groupi_n_402 ,csa_tree_add_89_22_pad_groupi_n_392 ,csa_tree_add_89_22_pad_groupi_n_376);
  and csa_tree_add_89_22_pad_groupi_g5351(csa_tree_add_89_22_pad_groupi_n_401 ,csa_tree_add_89_22_pad_groupi_n_390 ,csa_tree_add_89_22_pad_groupi_n_389);
  or csa_tree_add_89_22_pad_groupi_g5353(csa_tree_add_89_22_pad_groupi_n_395 ,csa_tree_add_89_22_pad_groupi_n_390 ,csa_tree_add_89_22_pad_groupi_n_389);
  not csa_tree_add_89_22_pad_groupi_g5354(csa_tree_add_89_22_pad_groupi_n_393 ,n_727);
  not csa_tree_add_89_22_pad_groupi_g5355(csa_tree_add_89_22_pad_groupi_n_392 ,n_719);
  not csa_tree_add_89_22_pad_groupi_g5356(csa_tree_add_89_22_pad_groupi_n_391 ,n_720);
  not csa_tree_add_89_22_pad_groupi_g5357(csa_tree_add_89_22_pad_groupi_n_390 ,n_722);
  not csa_tree_add_89_22_pad_groupi_g5358(csa_tree_add_89_22_pad_groupi_n_389 ,n_729);
  not csa_tree_add_89_22_pad_groupi_g5359(csa_tree_add_89_22_pad_groupi_n_388 ,n_728);
  not csa_tree_add_89_22_pad_groupi_g5360(csa_tree_add_89_22_pad_groupi_n_387 ,in13[7]);
  not csa_tree_add_89_22_pad_groupi_g5361(csa_tree_add_89_22_pad_groupi_n_386 ,in9[15]);
  not csa_tree_add_89_22_pad_groupi_g5362(csa_tree_add_89_22_pad_groupi_n_385 ,in9[2]);
  not csa_tree_add_89_22_pad_groupi_g5363(csa_tree_add_89_22_pad_groupi_n_384 ,in9[5]);
  not csa_tree_add_89_22_pad_groupi_g5364(csa_tree_add_89_22_pad_groupi_n_383 ,in9[13]);
  not csa_tree_add_89_22_pad_groupi_g5365(csa_tree_add_89_22_pad_groupi_n_382 ,in9[3]);
  not csa_tree_add_89_22_pad_groupi_g5366(csa_tree_add_89_22_pad_groupi_n_381 ,in9[9]);
  not csa_tree_add_89_22_pad_groupi_g5367(csa_tree_add_89_22_pad_groupi_n_380 ,in9[1]);
  not csa_tree_add_89_22_pad_groupi_g5368(csa_tree_add_89_22_pad_groupi_n_379 ,in9[8]);
  not csa_tree_add_89_22_pad_groupi_g5369(csa_tree_add_89_22_pad_groupi_n_378 ,n_718);
  not csa_tree_add_89_22_pad_groupi_g5370(csa_tree_add_89_22_pad_groupi_n_377 ,n_725);
  not csa_tree_add_89_22_pad_groupi_g5371(csa_tree_add_89_22_pad_groupi_n_376 ,n_726);
  not csa_tree_add_89_22_pad_groupi_g5372(csa_tree_add_89_22_pad_groupi_n_375 ,in14[0]);
  not csa_tree_add_89_22_pad_groupi_g5373(csa_tree_add_89_22_pad_groupi_n_374 ,in13[0]);
  not csa_tree_add_89_22_pad_groupi_g5374(csa_tree_add_89_22_pad_groupi_n_373 ,in13[11]);
  not csa_tree_add_89_22_pad_groupi_g5375(csa_tree_add_89_22_pad_groupi_n_372 ,in13[8]);
  not csa_tree_add_89_22_pad_groupi_g5376(csa_tree_add_89_22_pad_groupi_n_371 ,in13[1]);
  not csa_tree_add_89_22_pad_groupi_g5377(csa_tree_add_89_22_pad_groupi_n_370 ,in13[6]);
  not csa_tree_add_89_22_pad_groupi_g5378(csa_tree_add_89_22_pad_groupi_n_369 ,in13[9]);
  not csa_tree_add_89_22_pad_groupi_g5379(csa_tree_add_89_22_pad_groupi_n_368 ,in9[0]);
  not csa_tree_add_89_22_pad_groupi_g5380(csa_tree_add_89_22_pad_groupi_n_367 ,in9[4]);
  not csa_tree_add_89_22_pad_groupi_g5381(csa_tree_add_89_22_pad_groupi_n_366 ,in9[12]);
  not csa_tree_add_89_22_pad_groupi_g5382(csa_tree_add_89_22_pad_groupi_n_365 ,in9[11]);
  not csa_tree_add_89_22_pad_groupi_g5383(csa_tree_add_89_22_pad_groupi_n_364 ,in9[7]);
  not csa_tree_add_89_22_pad_groupi_g5384(csa_tree_add_89_22_pad_groupi_n_363 ,in9[10]);
  not csa_tree_add_89_22_pad_groupi_g5385(csa_tree_add_89_22_pad_groupi_n_362 ,in9[6]);
  not csa_tree_add_89_22_pad_groupi_g5386(csa_tree_add_89_22_pad_groupi_n_361 ,in9[14]);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5534(csa_tree_add_89_22_pad_groupi_n_345 ,csa_tree_add_89_22_pad_groupi_n_343);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5535(csa_tree_add_89_22_pad_groupi_n_344 ,csa_tree_add_89_22_pad_groupi_n_343);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5536(csa_tree_add_89_22_pad_groupi_n_343 ,csa_tree_add_89_22_pad_groupi_n_356);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5538(csa_tree_add_89_22_pad_groupi_n_342 ,csa_tree_add_89_22_pad_groupi_n_340);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5539(csa_tree_add_89_22_pad_groupi_n_341 ,csa_tree_add_89_22_pad_groupi_n_340);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5540(csa_tree_add_89_22_pad_groupi_n_340 ,csa_tree_add_89_22_pad_groupi_n_422);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5542(csa_tree_add_89_22_pad_groupi_n_339 ,csa_tree_add_89_22_pad_groupi_n_337);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5543(csa_tree_add_89_22_pad_groupi_n_338 ,csa_tree_add_89_22_pad_groupi_n_337);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5544(csa_tree_add_89_22_pad_groupi_n_337 ,csa_tree_add_89_22_pad_groupi_n_413);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5546(csa_tree_add_89_22_pad_groupi_n_336 ,csa_tree_add_89_22_pad_groupi_n_334);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5547(csa_tree_add_89_22_pad_groupi_n_335 ,csa_tree_add_89_22_pad_groupi_n_334);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5548(csa_tree_add_89_22_pad_groupi_n_334 ,csa_tree_add_89_22_pad_groupi_n_348);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5550(csa_tree_add_89_22_pad_groupi_n_333 ,csa_tree_add_89_22_pad_groupi_n_331);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5551(csa_tree_add_89_22_pad_groupi_n_332 ,csa_tree_add_89_22_pad_groupi_n_331);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5552(csa_tree_add_89_22_pad_groupi_n_331 ,csa_tree_add_89_22_pad_groupi_n_411);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5554(csa_tree_add_89_22_pad_groupi_n_330 ,csa_tree_add_89_22_pad_groupi_n_328);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5555(csa_tree_add_89_22_pad_groupi_n_329 ,csa_tree_add_89_22_pad_groupi_n_328);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5556(csa_tree_add_89_22_pad_groupi_n_328 ,csa_tree_add_89_22_pad_groupi_n_410);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5558(csa_tree_add_89_22_pad_groupi_n_327 ,csa_tree_add_89_22_pad_groupi_n_325);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5559(csa_tree_add_89_22_pad_groupi_n_326 ,csa_tree_add_89_22_pad_groupi_n_325);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5560(csa_tree_add_89_22_pad_groupi_n_325 ,csa_tree_add_89_22_pad_groupi_n_350);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5562(csa_tree_add_89_22_pad_groupi_n_324 ,csa_tree_add_89_22_pad_groupi_n_322);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5563(csa_tree_add_89_22_pad_groupi_n_323 ,csa_tree_add_89_22_pad_groupi_n_322);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5564(csa_tree_add_89_22_pad_groupi_n_322 ,csa_tree_add_89_22_pad_groupi_n_419);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5566(csa_tree_add_89_22_pad_groupi_n_321 ,csa_tree_add_89_22_pad_groupi_n_319);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5567(csa_tree_add_89_22_pad_groupi_n_320 ,csa_tree_add_89_22_pad_groupi_n_319);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5568(csa_tree_add_89_22_pad_groupi_n_319 ,csa_tree_add_89_22_pad_groupi_n_416);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5570(csa_tree_add_89_22_pad_groupi_n_318 ,csa_tree_add_89_22_pad_groupi_n_316);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5571(csa_tree_add_89_22_pad_groupi_n_317 ,csa_tree_add_89_22_pad_groupi_n_316);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5572(csa_tree_add_89_22_pad_groupi_n_316 ,csa_tree_add_89_22_pad_groupi_n_351);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5574(csa_tree_add_89_22_pad_groupi_n_315 ,csa_tree_add_89_22_pad_groupi_n_313);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5575(csa_tree_add_89_22_pad_groupi_n_314 ,csa_tree_add_89_22_pad_groupi_n_313);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5576(csa_tree_add_89_22_pad_groupi_n_313 ,csa_tree_add_89_22_pad_groupi_n_415);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5578(csa_tree_add_89_22_pad_groupi_n_312 ,csa_tree_add_89_22_pad_groupi_n_310);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5579(csa_tree_add_89_22_pad_groupi_n_311 ,csa_tree_add_89_22_pad_groupi_n_310);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5580(csa_tree_add_89_22_pad_groupi_n_310 ,csa_tree_add_89_22_pad_groupi_n_423);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5582(csa_tree_add_89_22_pad_groupi_n_309 ,csa_tree_add_89_22_pad_groupi_n_307);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5583(csa_tree_add_89_22_pad_groupi_n_308 ,csa_tree_add_89_22_pad_groupi_n_307);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5584(csa_tree_add_89_22_pad_groupi_n_307 ,csa_tree_add_89_22_pad_groupi_n_414);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5586(csa_tree_add_89_22_pad_groupi_n_306 ,csa_tree_add_89_22_pad_groupi_n_304);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5587(csa_tree_add_89_22_pad_groupi_n_305 ,csa_tree_add_89_22_pad_groupi_n_304);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5588(csa_tree_add_89_22_pad_groupi_n_304 ,csa_tree_add_89_22_pad_groupi_n_353);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5590(csa_tree_add_89_22_pad_groupi_n_303 ,csa_tree_add_89_22_pad_groupi_n_301);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5591(csa_tree_add_89_22_pad_groupi_n_302 ,csa_tree_add_89_22_pad_groupi_n_301);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5592(csa_tree_add_89_22_pad_groupi_n_301 ,csa_tree_add_89_22_pad_groupi_n_418);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5594(csa_tree_add_89_22_pad_groupi_n_300 ,csa_tree_add_89_22_pad_groupi_n_298);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5595(csa_tree_add_89_22_pad_groupi_n_299 ,csa_tree_add_89_22_pad_groupi_n_298);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5596(csa_tree_add_89_22_pad_groupi_n_298 ,csa_tree_add_89_22_pad_groupi_n_397);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5598(csa_tree_add_89_22_pad_groupi_n_297 ,csa_tree_add_89_22_pad_groupi_n_295);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5599(csa_tree_add_89_22_pad_groupi_n_296 ,csa_tree_add_89_22_pad_groupi_n_295);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5600(csa_tree_add_89_22_pad_groupi_n_295 ,csa_tree_add_89_22_pad_groupi_n_346);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5602(csa_tree_add_89_22_pad_groupi_n_294 ,csa_tree_add_89_22_pad_groupi_n_292);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5603(csa_tree_add_89_22_pad_groupi_n_293 ,csa_tree_add_89_22_pad_groupi_n_292);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5604(csa_tree_add_89_22_pad_groupi_n_292 ,csa_tree_add_89_22_pad_groupi_n_398);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5606(csa_tree_add_89_22_pad_groupi_n_291 ,csa_tree_add_89_22_pad_groupi_n_289);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5607(csa_tree_add_89_22_pad_groupi_n_290 ,csa_tree_add_89_22_pad_groupi_n_289);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5608(csa_tree_add_89_22_pad_groupi_n_289 ,csa_tree_add_89_22_pad_groupi_n_397);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5610(csa_tree_add_89_22_pad_groupi_n_288 ,csa_tree_add_89_22_pad_groupi_n_286);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5611(csa_tree_add_89_22_pad_groupi_n_287 ,csa_tree_add_89_22_pad_groupi_n_286);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5612(csa_tree_add_89_22_pad_groupi_n_286 ,csa_tree_add_89_22_pad_groupi_n_509);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5614(csa_tree_add_89_22_pad_groupi_n_285 ,csa_tree_add_89_22_pad_groupi_n_283);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5615(csa_tree_add_89_22_pad_groupi_n_284 ,csa_tree_add_89_22_pad_groupi_n_283);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5616(csa_tree_add_89_22_pad_groupi_n_283 ,csa_tree_add_89_22_pad_groupi_n_503);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5620(csa_tree_add_89_22_pad_groupi_n_358 ,csa_tree_add_89_22_pad_groupi_n_581);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5623(csa_tree_add_89_22_pad_groupi_n_282 ,csa_tree_add_89_22_pad_groupi_n_281);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5624(csa_tree_add_89_22_pad_groupi_n_281 ,csa_tree_add_89_22_pad_groupi_n_579);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5627(csa_tree_add_89_22_pad_groupi_n_280 ,csa_tree_add_89_22_pad_groupi_n_279);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5628(csa_tree_add_89_22_pad_groupi_n_279 ,csa_tree_add_89_22_pad_groupi_n_582);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5632(csa_tree_add_89_22_pad_groupi_n_357 ,csa_tree_add_89_22_pad_groupi_n_580);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5635(csa_tree_add_89_22_pad_groupi_n_278 ,csa_tree_add_89_22_pad_groupi_n_277);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5636(csa_tree_add_89_22_pad_groupi_n_277 ,csa_tree_add_89_22_pad_groupi_n_497);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5639(csa_tree_add_89_22_pad_groupi_n_276 ,csa_tree_add_89_22_pad_groupi_n_359);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5640(csa_tree_add_89_22_pad_groupi_n_359 ,csa_tree_add_89_22_pad_groupi_n_934);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5642(csa_tree_add_89_22_pad_groupi_n_275 ,csa_tree_add_89_22_pad_groupi_n_273);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5643(csa_tree_add_89_22_pad_groupi_n_274 ,csa_tree_add_89_22_pad_groupi_n_273);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5644(csa_tree_add_89_22_pad_groupi_n_273 ,csa_tree_add_89_22_pad_groupi_n_355);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5646(csa_tree_add_89_22_pad_groupi_n_272 ,csa_tree_add_89_22_pad_groupi_n_270);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5647(csa_tree_add_89_22_pad_groupi_n_271 ,csa_tree_add_89_22_pad_groupi_n_270);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5648(csa_tree_add_89_22_pad_groupi_n_270 ,csa_tree_add_89_22_pad_groupi_n_349);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5650(csa_tree_add_89_22_pad_groupi_n_269 ,csa_tree_add_89_22_pad_groupi_n_267);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5651(csa_tree_add_89_22_pad_groupi_n_268 ,csa_tree_add_89_22_pad_groupi_n_267);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5652(csa_tree_add_89_22_pad_groupi_n_267 ,csa_tree_add_89_22_pad_groupi_n_347);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5654(csa_tree_add_89_22_pad_groupi_n_266 ,csa_tree_add_89_22_pad_groupi_n_264);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5655(csa_tree_add_89_22_pad_groupi_n_265 ,csa_tree_add_89_22_pad_groupi_n_264);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5656(csa_tree_add_89_22_pad_groupi_n_264 ,csa_tree_add_89_22_pad_groupi_n_354);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5658(csa_tree_add_89_22_pad_groupi_n_263 ,csa_tree_add_89_22_pad_groupi_n_261);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5659(csa_tree_add_89_22_pad_groupi_n_262 ,csa_tree_add_89_22_pad_groupi_n_261);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5660(csa_tree_add_89_22_pad_groupi_n_261 ,csa_tree_add_89_22_pad_groupi_n_352);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5662(csa_tree_add_89_22_pad_groupi_n_260 ,csa_tree_add_89_22_pad_groupi_n_259);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5664(csa_tree_add_89_22_pad_groupi_n_259 ,csa_tree_add_89_22_pad_groupi_n_399);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5686(csa_tree_add_89_22_pad_groupi_n_258 ,csa_tree_add_89_22_pad_groupi_n_346);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5688(csa_tree_add_89_22_pad_groupi_n_346 ,csa_tree_add_89_22_pad_groupi_n_398);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5690(csa_tree_add_89_22_pad_groupi_n_257 ,csa_tree_add_89_22_pad_groupi_n_256);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5692(csa_tree_add_89_22_pad_groupi_n_256 ,csa_tree_add_89_22_pad_groupi_n_507);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5694(csa_tree_add_89_22_pad_groupi_n_255 ,csa_tree_add_89_22_pad_groupi_n_254);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5696(csa_tree_add_89_22_pad_groupi_n_254 ,csa_tree_add_89_22_pad_groupi_n_501);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5709(csa_tree_add_89_22_pad_groupi_n_253 ,csa_tree_add_89_22_pad_groupi_n_251);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5710(csa_tree_add_89_22_pad_groupi_n_252 ,csa_tree_add_89_22_pad_groupi_n_251);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5711(csa_tree_add_89_22_pad_groupi_n_251 ,csa_tree_add_89_22_pad_groupi_n_511);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5713(csa_tree_add_89_22_pad_groupi_n_250 ,csa_tree_add_89_22_pad_groupi_n_248);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5714(csa_tree_add_89_22_pad_groupi_n_249 ,csa_tree_add_89_22_pad_groupi_n_248);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5715(csa_tree_add_89_22_pad_groupi_n_248 ,csa_tree_add_89_22_pad_groupi_n_401);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5721(csa_tree_add_89_22_pad_groupi_n_247 ,csa_tree_add_89_22_pad_groupi_n_245);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5722(csa_tree_add_89_22_pad_groupi_n_246 ,csa_tree_add_89_22_pad_groupi_n_245);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5723(csa_tree_add_89_22_pad_groupi_n_245 ,csa_tree_add_89_22_pad_groupi_n_385);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5733(csa_tree_add_89_22_pad_groupi_n_244 ,csa_tree_add_89_22_pad_groupi_n_242);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5734(csa_tree_add_89_22_pad_groupi_n_243 ,csa_tree_add_89_22_pad_groupi_n_242);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5735(csa_tree_add_89_22_pad_groupi_n_242 ,csa_tree_add_89_22_pad_groupi_n_368);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5737(csa_tree_add_89_22_pad_groupi_n_241 ,csa_tree_add_89_22_pad_groupi_n_239);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5738(csa_tree_add_89_22_pad_groupi_n_240 ,csa_tree_add_89_22_pad_groupi_n_239);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5739(csa_tree_add_89_22_pad_groupi_n_239 ,csa_tree_add_89_22_pad_groupi_n_396);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5741(csa_tree_add_89_22_pad_groupi_n_238 ,csa_tree_add_89_22_pad_groupi_n_236);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5742(csa_tree_add_89_22_pad_groupi_n_237 ,csa_tree_add_89_22_pad_groupi_n_236);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5743(csa_tree_add_89_22_pad_groupi_n_236 ,csa_tree_add_89_22_pad_groupi_n_396);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5746(csa_tree_add_89_22_pad_groupi_n_235 ,csa_tree_add_89_22_pad_groupi_n_234);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5747(csa_tree_add_89_22_pad_groupi_n_234 ,csa_tree_add_89_22_pad_groupi_n_381);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5750(csa_tree_add_89_22_pad_groupi_n_233 ,csa_tree_add_89_22_pad_groupi_n_232);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5751(csa_tree_add_89_22_pad_groupi_n_232 ,csa_tree_add_89_22_pad_groupi_n_366);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5754(csa_tree_add_89_22_pad_groupi_n_231 ,csa_tree_add_89_22_pad_groupi_n_230);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5755(csa_tree_add_89_22_pad_groupi_n_230 ,csa_tree_add_89_22_pad_groupi_n_382);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5758(csa_tree_add_89_22_pad_groupi_n_229 ,csa_tree_add_89_22_pad_groupi_n_228);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5759(csa_tree_add_89_22_pad_groupi_n_228 ,csa_tree_add_89_22_pad_groupi_n_383);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5762(csa_tree_add_89_22_pad_groupi_n_227 ,csa_tree_add_89_22_pad_groupi_n_226);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5763(csa_tree_add_89_22_pad_groupi_n_226 ,csa_tree_add_89_22_pad_groupi_n_365);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5766(csa_tree_add_89_22_pad_groupi_n_225 ,csa_tree_add_89_22_pad_groupi_n_224);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5767(csa_tree_add_89_22_pad_groupi_n_224 ,csa_tree_add_89_22_pad_groupi_n_363);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5769(csa_tree_add_89_22_pad_groupi_n_223 ,csa_tree_add_89_22_pad_groupi_n_221);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5770(csa_tree_add_89_22_pad_groupi_n_222 ,csa_tree_add_89_22_pad_groupi_n_221);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5771(csa_tree_add_89_22_pad_groupi_n_221 ,csa_tree_add_89_22_pad_groupi_n_366);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5774(csa_tree_add_89_22_pad_groupi_n_220 ,csa_tree_add_89_22_pad_groupi_n_219);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5775(csa_tree_add_89_22_pad_groupi_n_219 ,csa_tree_add_89_22_pad_groupi_n_362);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5777(csa_tree_add_89_22_pad_groupi_n_218 ,csa_tree_add_89_22_pad_groupi_n_216);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5778(csa_tree_add_89_22_pad_groupi_n_217 ,csa_tree_add_89_22_pad_groupi_n_216);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5779(csa_tree_add_89_22_pad_groupi_n_216 ,csa_tree_add_89_22_pad_groupi_n_380);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5781(csa_tree_add_89_22_pad_groupi_n_215 ,csa_tree_add_89_22_pad_groupi_n_213);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5782(csa_tree_add_89_22_pad_groupi_n_214 ,csa_tree_add_89_22_pad_groupi_n_213);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5783(csa_tree_add_89_22_pad_groupi_n_213 ,csa_tree_add_89_22_pad_groupi_n_381);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5785(csa_tree_add_89_22_pad_groupi_n_212 ,csa_tree_add_89_22_pad_groupi_n_210);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5786(csa_tree_add_89_22_pad_groupi_n_211 ,csa_tree_add_89_22_pad_groupi_n_210);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5787(csa_tree_add_89_22_pad_groupi_n_210 ,csa_tree_add_89_22_pad_groupi_n_362);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5790(csa_tree_add_89_22_pad_groupi_n_209 ,csa_tree_add_89_22_pad_groupi_n_208);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5791(csa_tree_add_89_22_pad_groupi_n_208 ,csa_tree_add_89_22_pad_groupi_n_379);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5793(csa_tree_add_89_22_pad_groupi_n_207 ,csa_tree_add_89_22_pad_groupi_n_205);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5794(csa_tree_add_89_22_pad_groupi_n_206 ,csa_tree_add_89_22_pad_groupi_n_205);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5795(csa_tree_add_89_22_pad_groupi_n_205 ,csa_tree_add_89_22_pad_groupi_n_379);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5798(csa_tree_add_89_22_pad_groupi_n_204 ,csa_tree_add_89_22_pad_groupi_n_203);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5799(csa_tree_add_89_22_pad_groupi_n_203 ,csa_tree_add_89_22_pad_groupi_n_384);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5801(csa_tree_add_89_22_pad_groupi_n_202 ,csa_tree_add_89_22_pad_groupi_n_200);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5802(csa_tree_add_89_22_pad_groupi_n_201 ,csa_tree_add_89_22_pad_groupi_n_200);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5803(csa_tree_add_89_22_pad_groupi_n_200 ,csa_tree_add_89_22_pad_groupi_n_382);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5807(csa_tree_add_89_22_pad_groupi_n_198 ,csa_tree_add_89_22_pad_groupi_n_361);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5809(csa_tree_add_89_22_pad_groupi_n_197 ,csa_tree_add_89_22_pad_groupi_n_195);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5810(csa_tree_add_89_22_pad_groupi_n_196 ,csa_tree_add_89_22_pad_groupi_n_195);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5811(csa_tree_add_89_22_pad_groupi_n_195 ,csa_tree_add_89_22_pad_groupi_n_384);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5813(csa_tree_add_89_22_pad_groupi_n_194 ,csa_tree_add_89_22_pad_groupi_n_192);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5814(csa_tree_add_89_22_pad_groupi_n_193 ,csa_tree_add_89_22_pad_groupi_n_192);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5815(csa_tree_add_89_22_pad_groupi_n_192 ,csa_tree_add_89_22_pad_groupi_n_361);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5817(csa_tree_add_89_22_pad_groupi_n_191 ,csa_tree_add_89_22_pad_groupi_n_190);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5819(csa_tree_add_89_22_pad_groupi_n_190 ,csa_tree_add_89_22_pad_groupi_n_364);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5822(csa_tree_add_89_22_pad_groupi_n_189 ,csa_tree_add_89_22_pad_groupi_n_188);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5823(csa_tree_add_89_22_pad_groupi_n_188 ,csa_tree_add_89_22_pad_groupi_n_367);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5825(csa_tree_add_89_22_pad_groupi_n_187 ,csa_tree_add_89_22_pad_groupi_n_185);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5826(csa_tree_add_89_22_pad_groupi_n_186 ,csa_tree_add_89_22_pad_groupi_n_185);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5827(csa_tree_add_89_22_pad_groupi_n_185 ,csa_tree_add_89_22_pad_groupi_n_383);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5829(csa_tree_add_89_22_pad_groupi_n_184 ,csa_tree_add_89_22_pad_groupi_n_182);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5830(csa_tree_add_89_22_pad_groupi_n_183 ,csa_tree_add_89_22_pad_groupi_n_182);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5831(csa_tree_add_89_22_pad_groupi_n_182 ,csa_tree_add_89_22_pad_groupi_n_364);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5833(csa_tree_add_89_22_pad_groupi_n_181 ,csa_tree_add_89_22_pad_groupi_n_179);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5834(csa_tree_add_89_22_pad_groupi_n_180 ,csa_tree_add_89_22_pad_groupi_n_179);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5835(csa_tree_add_89_22_pad_groupi_n_179 ,csa_tree_add_89_22_pad_groupi_n_365);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5837(csa_tree_add_89_22_pad_groupi_n_178 ,csa_tree_add_89_22_pad_groupi_n_176);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5838(csa_tree_add_89_22_pad_groupi_n_177 ,csa_tree_add_89_22_pad_groupi_n_176);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5839(csa_tree_add_89_22_pad_groupi_n_176 ,csa_tree_add_89_22_pad_groupi_n_363);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5841(csa_tree_add_89_22_pad_groupi_n_175 ,csa_tree_add_89_22_pad_groupi_n_173);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5842(csa_tree_add_89_22_pad_groupi_n_174 ,csa_tree_add_89_22_pad_groupi_n_173);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5843(csa_tree_add_89_22_pad_groupi_n_173 ,csa_tree_add_89_22_pad_groupi_n_367);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5845(csa_tree_add_89_22_pad_groupi_n_172 ,csa_tree_add_89_22_pad_groupi_n_170);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5846(csa_tree_add_89_22_pad_groupi_n_171 ,csa_tree_add_89_22_pad_groupi_n_170);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5847(csa_tree_add_89_22_pad_groupi_n_170 ,csa_tree_add_89_22_pad_groupi_n_495);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5849(csa_tree_add_89_22_pad_groupi_n_169 ,csa_tree_add_89_22_pad_groupi_n_167);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5850(csa_tree_add_89_22_pad_groupi_n_168 ,csa_tree_add_89_22_pad_groupi_n_167);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5851(csa_tree_add_89_22_pad_groupi_n_167 ,csa_tree_add_89_22_pad_groupi_n_495);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5853(csa_tree_add_89_22_pad_groupi_n_166 ,csa_tree_add_89_22_pad_groupi_n_164);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5854(csa_tree_add_89_22_pad_groupi_n_165 ,csa_tree_add_89_22_pad_groupi_n_164);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5855(csa_tree_add_89_22_pad_groupi_n_164 ,csa_tree_add_89_22_pad_groupi_n_498);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5857(csa_tree_add_89_22_pad_groupi_n_163 ,csa_tree_add_89_22_pad_groupi_n_161);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5858(csa_tree_add_89_22_pad_groupi_n_162 ,csa_tree_add_89_22_pad_groupi_n_161);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5859(csa_tree_add_89_22_pad_groupi_n_161 ,csa_tree_add_89_22_pad_groupi_n_386);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5861(csa_tree_add_89_22_pad_groupi_n_160 ,csa_tree_add_89_22_pad_groupi_n_350);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5863(csa_tree_add_89_22_pad_groupi_n_350 ,csa_tree_add_89_22_pad_groupi_n_412);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5865(csa_tree_add_89_22_pad_groupi_n_159 ,csa_tree_add_89_22_pad_groupi_n_348);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5867(csa_tree_add_89_22_pad_groupi_n_348 ,csa_tree_add_89_22_pad_groupi_n_409);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5869(csa_tree_add_89_22_pad_groupi_n_158 ,csa_tree_add_89_22_pad_groupi_n_356);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5871(csa_tree_add_89_22_pad_groupi_n_356 ,csa_tree_add_89_22_pad_groupi_n_421);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5875(csa_tree_add_89_22_pad_groupi_n_156 ,csa_tree_add_89_22_pad_groupi_n_578);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5877(csa_tree_add_89_22_pad_groupi_n_155 ,csa_tree_add_89_22_pad_groupi_n_355);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5879(csa_tree_add_89_22_pad_groupi_n_355 ,csa_tree_add_89_22_pad_groupi_n_421);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5881(csa_tree_add_89_22_pad_groupi_n_154 ,csa_tree_add_89_22_pad_groupi_n_353);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5883(csa_tree_add_89_22_pad_groupi_n_353 ,csa_tree_add_89_22_pad_groupi_n_420);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5885(csa_tree_add_89_22_pad_groupi_n_153 ,csa_tree_add_89_22_pad_groupi_n_349);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5887(csa_tree_add_89_22_pad_groupi_n_349 ,csa_tree_add_89_22_pad_groupi_n_412);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5889(csa_tree_add_89_22_pad_groupi_n_152 ,csa_tree_add_89_22_pad_groupi_n_351);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5891(csa_tree_add_89_22_pad_groupi_n_351 ,csa_tree_add_89_22_pad_groupi_n_417);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5893(csa_tree_add_89_22_pad_groupi_n_151 ,csa_tree_add_89_22_pad_groupi_n_352);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5895(csa_tree_add_89_22_pad_groupi_n_352 ,csa_tree_add_89_22_pad_groupi_n_417);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5897(csa_tree_add_89_22_pad_groupi_n_150 ,csa_tree_add_89_22_pad_groupi_n_347);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5899(csa_tree_add_89_22_pad_groupi_n_347 ,csa_tree_add_89_22_pad_groupi_n_409);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5901(csa_tree_add_89_22_pad_groupi_n_149 ,csa_tree_add_89_22_pad_groupi_n_354);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5903(csa_tree_add_89_22_pad_groupi_n_354 ,csa_tree_add_89_22_pad_groupi_n_420);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5905(csa_tree_add_89_22_pad_groupi_n_148 ,csa_tree_add_89_22_pad_groupi_n_146);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5906(csa_tree_add_89_22_pad_groupi_n_147 ,csa_tree_add_89_22_pad_groupi_n_146);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5907(csa_tree_add_89_22_pad_groupi_n_146 ,csa_tree_add_89_22_pad_groupi_n_504);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5909(csa_tree_add_89_22_pad_groupi_n_145 ,csa_tree_add_89_22_pad_groupi_n_143);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5910(csa_tree_add_89_22_pad_groupi_n_144 ,csa_tree_add_89_22_pad_groupi_n_143);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5911(csa_tree_add_89_22_pad_groupi_n_143 ,csa_tree_add_89_22_pad_groupi_n_510);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5913(csa_tree_add_89_22_pad_groupi_n_142 ,csa_tree_add_89_22_pad_groupi_n_140);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5914(csa_tree_add_89_22_pad_groupi_n_141 ,csa_tree_add_89_22_pad_groupi_n_140);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5915(csa_tree_add_89_22_pad_groupi_n_140 ,csa_tree_add_89_22_pad_groupi_n_510);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5917(csa_tree_add_89_22_pad_groupi_n_139 ,csa_tree_add_89_22_pad_groupi_n_137);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5918(csa_tree_add_89_22_pad_groupi_n_138 ,csa_tree_add_89_22_pad_groupi_n_137);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5919(csa_tree_add_89_22_pad_groupi_n_137 ,csa_tree_add_89_22_pad_groupi_n_494);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5921(csa_tree_add_89_22_pad_groupi_n_136 ,csa_tree_add_89_22_pad_groupi_n_134);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5922(csa_tree_add_89_22_pad_groupi_n_135 ,csa_tree_add_89_22_pad_groupi_n_134);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5923(csa_tree_add_89_22_pad_groupi_n_134 ,csa_tree_add_89_22_pad_groupi_n_494);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5925(csa_tree_add_89_22_pad_groupi_n_133 ,csa_tree_add_89_22_pad_groupi_n_131);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5926(csa_tree_add_89_22_pad_groupi_n_132 ,csa_tree_add_89_22_pad_groupi_n_131);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5927(csa_tree_add_89_22_pad_groupi_n_131 ,csa_tree_add_89_22_pad_groupi_n_504);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5929(csa_tree_add_89_22_pad_groupi_n_130 ,csa_tree_add_89_22_pad_groupi_n_128);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5930(csa_tree_add_89_22_pad_groupi_n_129 ,csa_tree_add_89_22_pad_groupi_n_128);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5931(csa_tree_add_89_22_pad_groupi_n_128 ,csa_tree_add_89_22_pad_groupi_n_498);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5933(csa_tree_add_89_22_pad_groupi_n_127 ,csa_tree_add_89_22_pad_groupi_n_125);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5934(csa_tree_add_89_22_pad_groupi_n_126 ,csa_tree_add_89_22_pad_groupi_n_125);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5935(csa_tree_add_89_22_pad_groupi_n_125 ,csa_tree_add_89_22_pad_groupi_n_496);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5937(csa_tree_add_89_22_pad_groupi_n_124 ,csa_tree_add_89_22_pad_groupi_n_122);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5938(csa_tree_add_89_22_pad_groupi_n_123 ,csa_tree_add_89_22_pad_groupi_n_122);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5939(csa_tree_add_89_22_pad_groupi_n_122 ,csa_tree_add_89_22_pad_groupi_n_496);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5941(csa_tree_add_89_22_pad_groupi_n_121 ,csa_tree_add_89_22_pad_groupi_n_120);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5943(csa_tree_add_89_22_pad_groupi_n_120 ,csa_tree_add_89_22_pad_groupi_n_386);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5945(csa_tree_add_89_22_pad_groupi_n_119 ,csa_tree_add_89_22_pad_groupi_n_117);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5946(csa_tree_add_89_22_pad_groupi_n_118 ,csa_tree_add_89_22_pad_groupi_n_117);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5947(csa_tree_add_89_22_pad_groupi_n_117 ,csa_tree_add_89_22_pad_groupi_n_511);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5949(csa_tree_add_89_22_pad_groupi_n_116 ,csa_tree_add_89_22_pad_groupi_n_114);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5950(csa_tree_add_89_22_pad_groupi_n_115 ,csa_tree_add_89_22_pad_groupi_n_114);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5951(csa_tree_add_89_22_pad_groupi_n_114 ,csa_tree_add_89_22_pad_groupi_n_511);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5953(csa_tree_add_89_22_pad_groupi_n_113 ,csa_tree_add_89_22_pad_groupi_n_111);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5954(csa_tree_add_89_22_pad_groupi_n_112 ,csa_tree_add_89_22_pad_groupi_n_111);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5955(csa_tree_add_89_22_pad_groupi_n_111 ,csa_tree_add_89_22_pad_groupi_n_253);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5957(csa_tree_add_89_22_pad_groupi_n_110 ,csa_tree_add_89_22_pad_groupi_n_108);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5958(csa_tree_add_89_22_pad_groupi_n_109 ,csa_tree_add_89_22_pad_groupi_n_108);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5959(csa_tree_add_89_22_pad_groupi_n_108 ,csa_tree_add_89_22_pad_groupi_n_401);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5961(csa_tree_add_89_22_pad_groupi_n_107 ,csa_tree_add_89_22_pad_groupi_n_105);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5962(csa_tree_add_89_22_pad_groupi_n_106 ,csa_tree_add_89_22_pad_groupi_n_105);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5963(csa_tree_add_89_22_pad_groupi_n_105 ,csa_tree_add_89_22_pad_groupi_n_401);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5965(csa_tree_add_89_22_pad_groupi_n_104 ,csa_tree_add_89_22_pad_groupi_n_102);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5966(csa_tree_add_89_22_pad_groupi_n_103 ,csa_tree_add_89_22_pad_groupi_n_102);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5967(csa_tree_add_89_22_pad_groupi_n_102 ,csa_tree_add_89_22_pad_groupi_n_250);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5969(csa_tree_add_89_22_pad_groupi_n_101 ,csa_tree_add_89_22_pad_groupi_n_99);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5970(csa_tree_add_89_22_pad_groupi_n_100 ,csa_tree_add_89_22_pad_groupi_n_99);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5971(csa_tree_add_89_22_pad_groupi_n_99 ,csa_tree_add_89_22_pad_groupi_n_385);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5973(csa_tree_add_89_22_pad_groupi_n_98 ,csa_tree_add_89_22_pad_groupi_n_97);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5975(csa_tree_add_89_22_pad_groupi_n_97 ,csa_tree_add_89_22_pad_groupi_n_247);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5977(csa_tree_add_89_22_pad_groupi_n_96 ,csa_tree_add_89_22_pad_groupi_n_94);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5978(csa_tree_add_89_22_pad_groupi_n_95 ,csa_tree_add_89_22_pad_groupi_n_94);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5979(csa_tree_add_89_22_pad_groupi_n_94 ,csa_tree_add_89_22_pad_groupi_n_381);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5981(csa_tree_add_89_22_pad_groupi_n_93 ,csa_tree_add_89_22_pad_groupi_n_92);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5983(csa_tree_add_89_22_pad_groupi_n_92 ,csa_tree_add_89_22_pad_groupi_n_252);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5985(csa_tree_add_89_22_pad_groupi_n_91 ,csa_tree_add_89_22_pad_groupi_n_89);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5986(csa_tree_add_89_22_pad_groupi_n_90 ,csa_tree_add_89_22_pad_groupi_n_89);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5987(csa_tree_add_89_22_pad_groupi_n_89 ,csa_tree_add_89_22_pad_groupi_n_366);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5989(csa_tree_add_89_22_pad_groupi_n_88 ,csa_tree_add_89_22_pad_groupi_n_86);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5990(csa_tree_add_89_22_pad_groupi_n_87 ,csa_tree_add_89_22_pad_groupi_n_86);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5991(csa_tree_add_89_22_pad_groupi_n_86 ,csa_tree_add_89_22_pad_groupi_n_382);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5993(csa_tree_add_89_22_pad_groupi_n_85 ,csa_tree_add_89_22_pad_groupi_n_83);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5994(csa_tree_add_89_22_pad_groupi_n_84 ,csa_tree_add_89_22_pad_groupi_n_83);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5995(csa_tree_add_89_22_pad_groupi_n_83 ,csa_tree_add_89_22_pad_groupi_n_383);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5997(csa_tree_add_89_22_pad_groupi_n_82 ,csa_tree_add_89_22_pad_groupi_n_80);
  not csa_tree_add_89_22_pad_groupi_drc_bufs5999(csa_tree_add_89_22_pad_groupi_n_80 ,csa_tree_add_89_22_pad_groupi_n_365);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6001(csa_tree_add_89_22_pad_groupi_n_79 ,csa_tree_add_89_22_pad_groupi_n_77);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6002(csa_tree_add_89_22_pad_groupi_n_78 ,csa_tree_add_89_22_pad_groupi_n_77);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6003(csa_tree_add_89_22_pad_groupi_n_77 ,csa_tree_add_89_22_pad_groupi_n_363);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6005(csa_tree_add_89_22_pad_groupi_n_76 ,csa_tree_add_89_22_pad_groupi_n_75);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6007(csa_tree_add_89_22_pad_groupi_n_75 ,csa_tree_add_89_22_pad_groupi_n_215);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6009(csa_tree_add_89_22_pad_groupi_n_74 ,csa_tree_add_89_22_pad_groupi_n_72);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6010(csa_tree_add_89_22_pad_groupi_n_73 ,csa_tree_add_89_22_pad_groupi_n_72);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6011(csa_tree_add_89_22_pad_groupi_n_72 ,csa_tree_add_89_22_pad_groupi_n_385);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6013(csa_tree_add_89_22_pad_groupi_n_71 ,csa_tree_add_89_22_pad_groupi_n_70);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6015(csa_tree_add_89_22_pad_groupi_n_70 ,csa_tree_add_89_22_pad_groupi_n_218);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6017(csa_tree_add_89_22_pad_groupi_n_69 ,csa_tree_add_89_22_pad_groupi_n_68);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6019(csa_tree_add_89_22_pad_groupi_n_68 ,csa_tree_add_89_22_pad_groupi_n_223);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6021(csa_tree_add_89_22_pad_groupi_n_67 ,csa_tree_add_89_22_pad_groupi_n_65);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6022(csa_tree_add_89_22_pad_groupi_n_66 ,csa_tree_add_89_22_pad_groupi_n_65);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6023(csa_tree_add_89_22_pad_groupi_n_65 ,csa_tree_add_89_22_pad_groupi_n_362);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6025(csa_tree_add_89_22_pad_groupi_n_64 ,csa_tree_add_89_22_pad_groupi_n_62);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6027(csa_tree_add_89_22_pad_groupi_n_62 ,csa_tree_add_89_22_pad_groupi_n_380);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6029(csa_tree_add_89_22_pad_groupi_n_61 ,csa_tree_add_89_22_pad_groupi_n_60);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6031(csa_tree_add_89_22_pad_groupi_n_60 ,csa_tree_add_89_22_pad_groupi_n_249);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6033(csa_tree_add_89_22_pad_groupi_n_59 ,csa_tree_add_89_22_pad_groupi_n_58);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6035(csa_tree_add_89_22_pad_groupi_n_58 ,csa_tree_add_89_22_pad_groupi_n_212);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6037(csa_tree_add_89_22_pad_groupi_n_57 ,csa_tree_add_89_22_pad_groupi_n_56);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6039(csa_tree_add_89_22_pad_groupi_n_56 ,csa_tree_add_89_22_pad_groupi_n_244);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6041(csa_tree_add_89_22_pad_groupi_n_55 ,csa_tree_add_89_22_pad_groupi_n_54);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6043(csa_tree_add_89_22_pad_groupi_n_54 ,csa_tree_add_89_22_pad_groupi_n_207);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6045(csa_tree_add_89_22_pad_groupi_n_53 ,csa_tree_add_89_22_pad_groupi_n_51);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6046(csa_tree_add_89_22_pad_groupi_n_52 ,csa_tree_add_89_22_pad_groupi_n_51);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6047(csa_tree_add_89_22_pad_groupi_n_51 ,csa_tree_add_89_22_pad_groupi_n_384);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6049(csa_tree_add_89_22_pad_groupi_n_50 ,csa_tree_add_89_22_pad_groupi_n_48);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6051(csa_tree_add_89_22_pad_groupi_n_48 ,csa_tree_add_89_22_pad_groupi_n_379);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6053(csa_tree_add_89_22_pad_groupi_n_47 ,csa_tree_add_89_22_pad_groupi_n_46);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6055(csa_tree_add_89_22_pad_groupi_n_46 ,csa_tree_add_89_22_pad_groupi_n_246);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6057(csa_tree_add_89_22_pad_groupi_n_45 ,csa_tree_add_89_22_pad_groupi_n_43);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6059(csa_tree_add_89_22_pad_groupi_n_43 ,csa_tree_add_89_22_pad_groupi_n_380);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6061(csa_tree_add_89_22_pad_groupi_n_42 ,csa_tree_add_89_22_pad_groupi_n_40);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6062(csa_tree_add_89_22_pad_groupi_n_41 ,csa_tree_add_89_22_pad_groupi_n_40);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6063(csa_tree_add_89_22_pad_groupi_n_40 ,csa_tree_add_89_22_pad_groupi_n_368);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6065(csa_tree_add_89_22_pad_groupi_n_39 ,csa_tree_add_89_22_pad_groupi_n_37);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6066(csa_tree_add_89_22_pad_groupi_n_38 ,csa_tree_add_89_22_pad_groupi_n_37);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6067(csa_tree_add_89_22_pad_groupi_n_37 ,csa_tree_add_89_22_pad_groupi_n_361);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6069(csa_tree_add_89_22_pad_groupi_n_36 ,csa_tree_add_89_22_pad_groupi_n_35);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6071(csa_tree_add_89_22_pad_groupi_n_35 ,csa_tree_add_89_22_pad_groupi_n_202);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6073(csa_tree_add_89_22_pad_groupi_n_34 ,csa_tree_add_89_22_pad_groupi_n_33);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6075(csa_tree_add_89_22_pad_groupi_n_33 ,csa_tree_add_89_22_pad_groupi_n_238);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6077(csa_tree_add_89_22_pad_groupi_n_32 ,csa_tree_add_89_22_pad_groupi_n_31);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6079(csa_tree_add_89_22_pad_groupi_n_31 ,csa_tree_add_89_22_pad_groupi_n_241);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6082(csa_tree_add_89_22_pad_groupi_n_30 ,csa_tree_add_89_22_pad_groupi_n_29);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6083(csa_tree_add_89_22_pad_groupi_n_29 ,csa_tree_add_89_22_pad_groupi_n_193);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6085(csa_tree_add_89_22_pad_groupi_n_28 ,csa_tree_add_89_22_pad_groupi_n_26);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6086(csa_tree_add_89_22_pad_groupi_n_27 ,csa_tree_add_89_22_pad_groupi_n_26);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6087(csa_tree_add_89_22_pad_groupi_n_26 ,csa_tree_add_89_22_pad_groupi_n_367);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6089(csa_tree_add_89_22_pad_groupi_n_25 ,csa_tree_add_89_22_pad_groupi_n_23);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6090(csa_tree_add_89_22_pad_groupi_n_24 ,csa_tree_add_89_22_pad_groupi_n_23);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6091(csa_tree_add_89_22_pad_groupi_n_23 ,csa_tree_add_89_22_pad_groupi_n_368);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6093(csa_tree_add_89_22_pad_groupi_n_22 ,csa_tree_add_89_22_pad_groupi_n_20);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6094(csa_tree_add_89_22_pad_groupi_n_21 ,csa_tree_add_89_22_pad_groupi_n_20);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6095(csa_tree_add_89_22_pad_groupi_n_20 ,csa_tree_add_89_22_pad_groupi_n_364);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6098(csa_tree_add_89_22_pad_groupi_n_19 ,csa_tree_add_89_22_pad_groupi_n_18);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6099(csa_tree_add_89_22_pad_groupi_n_18 ,csa_tree_add_89_22_pad_groupi_n_243);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6102(csa_tree_add_89_22_pad_groupi_n_17 ,csa_tree_add_89_22_pad_groupi_n_16);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6103(csa_tree_add_89_22_pad_groupi_n_16 ,csa_tree_add_89_22_pad_groupi_n_196);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6106(csa_tree_add_89_22_pad_groupi_n_15 ,csa_tree_add_89_22_pad_groupi_n_14);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6107(csa_tree_add_89_22_pad_groupi_n_14 ,csa_tree_add_89_22_pad_groupi_n_237);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6110(csa_tree_add_89_22_pad_groupi_n_13 ,csa_tree_add_89_22_pad_groupi_n_12);
  not csa_tree_add_89_22_pad_groupi_drc_bufs6111(csa_tree_add_89_22_pad_groupi_n_12 ,csa_tree_add_89_22_pad_groupi_n_240);
  xor csa_tree_add_89_22_pad_groupi_g2(n_167 ,csa_tree_add_89_22_pad_groupi_n_1537 ,csa_tree_add_89_22_pad_groupi_n_1520);
  xor csa_tree_add_89_22_pad_groupi_g6113(n_165 ,csa_tree_add_89_22_pad_groupi_n_1532 ,csa_tree_add_89_22_pad_groupi_n_1518);
  xor csa_tree_add_89_22_pad_groupi_g6114(n_162 ,csa_tree_add_89_22_pad_groupi_n_1524 ,csa_tree_add_89_22_pad_groupi_n_1482);
  xor csa_tree_add_89_22_pad_groupi_g6115(n_161 ,csa_tree_add_89_22_pad_groupi_n_1522 ,csa_tree_add_89_22_pad_groupi_n_1502);
  xor csa_tree_add_89_22_pad_groupi_g6116(n_160 ,csa_tree_add_89_22_pad_groupi_n_1515 ,csa_tree_add_89_22_pad_groupi_n_1461);
  xor csa_tree_add_89_22_pad_groupi_g6117(csa_tree_add_89_22_pad_groupi_n_6 ,csa_tree_add_89_22_pad_groupi_n_1368 ,csa_tree_add_89_22_pad_groupi_n_1406);
  xor csa_tree_add_89_22_pad_groupi_g6118(csa_tree_add_89_22_pad_groupi_n_5 ,csa_tree_add_89_22_pad_groupi_n_1332 ,csa_tree_add_89_22_pad_groupi_n_1350);
  xor csa_tree_add_89_22_pad_groupi_g6119(csa_tree_add_89_22_pad_groupi_n_4 ,csa_tree_add_89_22_pad_groupi_n_836 ,csa_tree_add_89_22_pad_groupi_n_0);
  xor csa_tree_add_89_22_pad_groupi_g6120(csa_tree_add_89_22_pad_groupi_n_3 ,csa_tree_add_89_22_pad_groupi_n_835 ,csa_tree_add_89_22_pad_groupi_n_948);
  xor csa_tree_add_89_22_pad_groupi_g6121(csa_tree_add_89_22_pad_groupi_n_2 ,csa_tree_add_89_22_pad_groupi_n_584 ,csa_tree_add_89_22_pad_groupi_n_156);
  xor csa_tree_add_89_22_pad_groupi_g6122(csa_tree_add_89_22_pad_groupi_n_1 ,csa_tree_add_89_22_pad_groupi_n_358 ,in13[9]);
  xor csa_tree_add_89_22_pad_groupi_g6123(csa_tree_add_89_22_pad_groupi_n_0 ,csa_tree_add_89_22_pad_groupi_n_357 ,in13[11]);
  xnor csa_tree_add_95_22_pad_groupi_g4151(n_286 ,csa_tree_add_95_22_pad_groupi_n_1336 ,csa_tree_add_95_22_pad_groupi_n_1558);
  or csa_tree_add_95_22_pad_groupi_g4152(csa_tree_add_95_22_pad_groupi_n_1558 ,csa_tree_add_95_22_pad_groupi_n_1393 ,csa_tree_add_95_22_pad_groupi_n_1556);
  xnor csa_tree_add_95_22_pad_groupi_g4153(n_285 ,csa_tree_add_95_22_pad_groupi_n_1555 ,csa_tree_add_95_22_pad_groupi_n_1404);
  and csa_tree_add_95_22_pad_groupi_g4154(csa_tree_add_95_22_pad_groupi_n_1556 ,csa_tree_add_95_22_pad_groupi_n_1389 ,csa_tree_add_95_22_pad_groupi_n_1555);
  or csa_tree_add_95_22_pad_groupi_g4155(csa_tree_add_95_22_pad_groupi_n_1555 ,csa_tree_add_95_22_pad_groupi_n_1407 ,csa_tree_add_95_22_pad_groupi_n_1553);
  xnor csa_tree_add_95_22_pad_groupi_g4156(n_284 ,csa_tree_add_95_22_pad_groupi_n_1552 ,csa_tree_add_95_22_pad_groupi_n_1434);
  and csa_tree_add_95_22_pad_groupi_g4157(csa_tree_add_95_22_pad_groupi_n_1553 ,csa_tree_add_95_22_pad_groupi_n_1410 ,csa_tree_add_95_22_pad_groupi_n_1552);
  or csa_tree_add_95_22_pad_groupi_g4158(csa_tree_add_95_22_pad_groupi_n_1552 ,csa_tree_add_95_22_pad_groupi_n_1453 ,csa_tree_add_95_22_pad_groupi_n_1550);
  xnor csa_tree_add_95_22_pad_groupi_g4159(n_283 ,csa_tree_add_95_22_pad_groupi_n_1549 ,csa_tree_add_95_22_pad_groupi_n_1462);
  and csa_tree_add_95_22_pad_groupi_g4160(csa_tree_add_95_22_pad_groupi_n_1550 ,csa_tree_add_95_22_pad_groupi_n_1459 ,csa_tree_add_95_22_pad_groupi_n_1549);
  or csa_tree_add_95_22_pad_groupi_g4161(csa_tree_add_95_22_pad_groupi_n_1549 ,csa_tree_add_95_22_pad_groupi_n_1463 ,csa_tree_add_95_22_pad_groupi_n_1547);
  xnor csa_tree_add_95_22_pad_groupi_g4162(n_282 ,csa_tree_add_95_22_pad_groupi_n_1546 ,csa_tree_add_95_22_pad_groupi_n_1483);
  nor csa_tree_add_95_22_pad_groupi_g4163(csa_tree_add_95_22_pad_groupi_n_1547 ,csa_tree_add_95_22_pad_groupi_n_1546 ,csa_tree_add_95_22_pad_groupi_n_1464);
  and csa_tree_add_95_22_pad_groupi_g4164(csa_tree_add_95_22_pad_groupi_n_1546 ,csa_tree_add_95_22_pad_groupi_n_1500 ,csa_tree_add_95_22_pad_groupi_n_1544);
  xnor csa_tree_add_95_22_pad_groupi_g4165(n_281 ,csa_tree_add_95_22_pad_groupi_n_1542 ,csa_tree_add_95_22_pad_groupi_n_1501);
  or csa_tree_add_95_22_pad_groupi_g4166(csa_tree_add_95_22_pad_groupi_n_1544 ,csa_tree_add_95_22_pad_groupi_n_1494 ,csa_tree_add_95_22_pad_groupi_n_1543);
  not csa_tree_add_95_22_pad_groupi_g4167(csa_tree_add_95_22_pad_groupi_n_1543 ,csa_tree_add_95_22_pad_groupi_n_1542);
  or csa_tree_add_95_22_pad_groupi_g4168(csa_tree_add_95_22_pad_groupi_n_1542 ,csa_tree_add_95_22_pad_groupi_n_1499 ,csa_tree_add_95_22_pad_groupi_n_1540);
  xnor csa_tree_add_95_22_pad_groupi_g4169(n_280 ,csa_tree_add_95_22_pad_groupi_n_1539 ,csa_tree_add_95_22_pad_groupi_n_1503);
  nor csa_tree_add_95_22_pad_groupi_g4170(csa_tree_add_95_22_pad_groupi_n_1540 ,csa_tree_add_95_22_pad_groupi_n_1496 ,csa_tree_add_95_22_pad_groupi_n_1539);
  and csa_tree_add_95_22_pad_groupi_g4171(csa_tree_add_95_22_pad_groupi_n_1539 ,csa_tree_add_95_22_pad_groupi_n_1538 ,csa_tree_add_95_22_pad_groupi_n_1510);
  or csa_tree_add_95_22_pad_groupi_g4173(csa_tree_add_95_22_pad_groupi_n_1538 ,csa_tree_add_95_22_pad_groupi_n_1513 ,csa_tree_add_95_22_pad_groupi_n_1537);
  and csa_tree_add_95_22_pad_groupi_g4175(csa_tree_add_95_22_pad_groupi_n_1537 ,csa_tree_add_95_22_pad_groupi_n_1512 ,csa_tree_add_95_22_pad_groupi_n_1535);
  xnor csa_tree_add_95_22_pad_groupi_g4176(n_278 ,csa_tree_add_95_22_pad_groupi_n_1534 ,csa_tree_add_95_22_pad_groupi_n_1519);
  or csa_tree_add_95_22_pad_groupi_g4177(csa_tree_add_95_22_pad_groupi_n_1535 ,csa_tree_add_95_22_pad_groupi_n_1514 ,csa_tree_add_95_22_pad_groupi_n_1534);
  and csa_tree_add_95_22_pad_groupi_g4178(csa_tree_add_95_22_pad_groupi_n_1534 ,csa_tree_add_95_22_pad_groupi_n_1533 ,csa_tree_add_95_22_pad_groupi_n_1511);
  or csa_tree_add_95_22_pad_groupi_g4180(csa_tree_add_95_22_pad_groupi_n_1533 ,csa_tree_add_95_22_pad_groupi_n_1505 ,csa_tree_add_95_22_pad_groupi_n_1532);
  and csa_tree_add_95_22_pad_groupi_g4182(csa_tree_add_95_22_pad_groupi_n_1532 ,csa_tree_add_95_22_pad_groupi_n_1506 ,csa_tree_add_95_22_pad_groupi_n_1530);
  xnor csa_tree_add_95_22_pad_groupi_g4183(n_276 ,csa_tree_add_95_22_pad_groupi_n_1529 ,csa_tree_add_95_22_pad_groupi_n_1517);
  or csa_tree_add_95_22_pad_groupi_g4184(csa_tree_add_95_22_pad_groupi_n_1530 ,csa_tree_add_95_22_pad_groupi_n_1507 ,csa_tree_add_95_22_pad_groupi_n_1529);
  and csa_tree_add_95_22_pad_groupi_g4185(csa_tree_add_95_22_pad_groupi_n_1529 ,csa_tree_add_95_22_pad_groupi_n_1508 ,csa_tree_add_95_22_pad_groupi_n_1527);
  xnor csa_tree_add_95_22_pad_groupi_g4186(n_275 ,csa_tree_add_95_22_pad_groupi_n_1526 ,csa_tree_add_95_22_pad_groupi_n_1516);
  or csa_tree_add_95_22_pad_groupi_g4187(csa_tree_add_95_22_pad_groupi_n_1527 ,csa_tree_add_95_22_pad_groupi_n_1526 ,csa_tree_add_95_22_pad_groupi_n_1509);
  and csa_tree_add_95_22_pad_groupi_g4188(csa_tree_add_95_22_pad_groupi_n_1526 ,csa_tree_add_95_22_pad_groupi_n_1471 ,csa_tree_add_95_22_pad_groupi_n_1525);
  or csa_tree_add_95_22_pad_groupi_g4190(csa_tree_add_95_22_pad_groupi_n_1525 ,csa_tree_add_95_22_pad_groupi_n_1470 ,csa_tree_add_95_22_pad_groupi_n_1524);
  and csa_tree_add_95_22_pad_groupi_g4192(csa_tree_add_95_22_pad_groupi_n_1524 ,csa_tree_add_95_22_pad_groupi_n_1498 ,csa_tree_add_95_22_pad_groupi_n_1523);
  or csa_tree_add_95_22_pad_groupi_g4194(csa_tree_add_95_22_pad_groupi_n_1523 ,csa_tree_add_95_22_pad_groupi_n_1497 ,csa_tree_add_95_22_pad_groupi_n_1522);
  and csa_tree_add_95_22_pad_groupi_g4196(csa_tree_add_95_22_pad_groupi_n_1522 ,csa_tree_add_95_22_pad_groupi_n_1452 ,csa_tree_add_95_22_pad_groupi_n_1521);
  or csa_tree_add_95_22_pad_groupi_g4198(csa_tree_add_95_22_pad_groupi_n_1521 ,csa_tree_add_95_22_pad_groupi_n_1451 ,csa_tree_add_95_22_pad_groupi_n_1515);
  xnor csa_tree_add_95_22_pad_groupi_g4199(csa_tree_add_95_22_pad_groupi_n_1520 ,csa_tree_add_95_22_pad_groupi_n_1475 ,csa_tree_add_95_22_pad_groupi_n_1491);
  xnor csa_tree_add_95_22_pad_groupi_g4200(csa_tree_add_95_22_pad_groupi_n_1519 ,csa_tree_add_95_22_pad_groupi_n_1473 ,csa_tree_add_95_22_pad_groupi_n_1489);
  xnor csa_tree_add_95_22_pad_groupi_g4201(csa_tree_add_95_22_pad_groupi_n_1518 ,csa_tree_add_95_22_pad_groupi_n_1480 ,csa_tree_add_95_22_pad_groupi_n_1487);
  xnor csa_tree_add_95_22_pad_groupi_g4202(csa_tree_add_95_22_pad_groupi_n_1517 ,csa_tree_add_95_22_pad_groupi_n_1477 ,csa_tree_add_95_22_pad_groupi_n_1493);
  xnor csa_tree_add_95_22_pad_groupi_g4203(csa_tree_add_95_22_pad_groupi_n_1516 ,csa_tree_add_95_22_pad_groupi_n_1448 ,csa_tree_add_95_22_pad_groupi_n_1485);
  nor csa_tree_add_95_22_pad_groupi_g4205(csa_tree_add_95_22_pad_groupi_n_1514 ,csa_tree_add_95_22_pad_groupi_n_1472 ,csa_tree_add_95_22_pad_groupi_n_1489);
  nor csa_tree_add_95_22_pad_groupi_g4206(csa_tree_add_95_22_pad_groupi_n_1513 ,csa_tree_add_95_22_pad_groupi_n_1475 ,csa_tree_add_95_22_pad_groupi_n_1491);
  or csa_tree_add_95_22_pad_groupi_g4207(csa_tree_add_95_22_pad_groupi_n_1512 ,csa_tree_add_95_22_pad_groupi_n_1473 ,csa_tree_add_95_22_pad_groupi_n_1488);
  or csa_tree_add_95_22_pad_groupi_g4208(csa_tree_add_95_22_pad_groupi_n_1511 ,csa_tree_add_95_22_pad_groupi_n_1479 ,csa_tree_add_95_22_pad_groupi_n_1486);
  or csa_tree_add_95_22_pad_groupi_g4209(csa_tree_add_95_22_pad_groupi_n_1510 ,csa_tree_add_95_22_pad_groupi_n_1474 ,csa_tree_add_95_22_pad_groupi_n_1490);
  nor csa_tree_add_95_22_pad_groupi_g4210(csa_tree_add_95_22_pad_groupi_n_1509 ,csa_tree_add_95_22_pad_groupi_n_1447 ,csa_tree_add_95_22_pad_groupi_n_1485);
  and csa_tree_add_95_22_pad_groupi_g4211(csa_tree_add_95_22_pad_groupi_n_1515 ,csa_tree_add_95_22_pad_groupi_n_1450 ,csa_tree_add_95_22_pad_groupi_n_1495);
  or csa_tree_add_95_22_pad_groupi_g4212(csa_tree_add_95_22_pad_groupi_n_1508 ,csa_tree_add_95_22_pad_groupi_n_1448 ,csa_tree_add_95_22_pad_groupi_n_1484);
  nor csa_tree_add_95_22_pad_groupi_g4213(csa_tree_add_95_22_pad_groupi_n_1507 ,csa_tree_add_95_22_pad_groupi_n_1476 ,csa_tree_add_95_22_pad_groupi_n_1493);
  or csa_tree_add_95_22_pad_groupi_g4214(csa_tree_add_95_22_pad_groupi_n_1506 ,csa_tree_add_95_22_pad_groupi_n_1477 ,csa_tree_add_95_22_pad_groupi_n_1492);
  nor csa_tree_add_95_22_pad_groupi_g4215(csa_tree_add_95_22_pad_groupi_n_1505 ,csa_tree_add_95_22_pad_groupi_n_1480 ,csa_tree_add_95_22_pad_groupi_n_1487);
  xnor csa_tree_add_95_22_pad_groupi_g4216(n_271 ,csa_tree_add_95_22_pad_groupi_n_1481 ,csa_tree_add_95_22_pad_groupi_n_1460);
  xnor csa_tree_add_95_22_pad_groupi_g4217(csa_tree_add_95_22_pad_groupi_n_1503 ,csa_tree_add_95_22_pad_groupi_n_1478 ,csa_tree_add_95_22_pad_groupi_n_1467);
  xnor csa_tree_add_95_22_pad_groupi_g4218(csa_tree_add_95_22_pad_groupi_n_1502 ,csa_tree_add_95_22_pad_groupi_n_1412 ,csa_tree_add_95_22_pad_groupi_n_1466);
  xnor csa_tree_add_95_22_pad_groupi_g4219(csa_tree_add_95_22_pad_groupi_n_1501 ,csa_tree_add_95_22_pad_groupi_n_1442 ,csa_tree_add_95_22_pad_groupi_n_1469);
  or csa_tree_add_95_22_pad_groupi_g4220(csa_tree_add_95_22_pad_groupi_n_1500 ,csa_tree_add_95_22_pad_groupi_n_1441 ,csa_tree_add_95_22_pad_groupi_n_6);
  nor csa_tree_add_95_22_pad_groupi_g4221(csa_tree_add_95_22_pad_groupi_n_1499 ,csa_tree_add_95_22_pad_groupi_n_1478 ,csa_tree_add_95_22_pad_groupi_n_1468);
  or csa_tree_add_95_22_pad_groupi_g4222(csa_tree_add_95_22_pad_groupi_n_1498 ,csa_tree_add_95_22_pad_groupi_n_1411 ,csa_tree_add_95_22_pad_groupi_n_1465);
  nor csa_tree_add_95_22_pad_groupi_g4223(csa_tree_add_95_22_pad_groupi_n_1497 ,csa_tree_add_95_22_pad_groupi_n_1412 ,csa_tree_add_95_22_pad_groupi_n_1466);
  and csa_tree_add_95_22_pad_groupi_g4224(csa_tree_add_95_22_pad_groupi_n_1496 ,csa_tree_add_95_22_pad_groupi_n_1478 ,csa_tree_add_95_22_pad_groupi_n_1468);
  or csa_tree_add_95_22_pad_groupi_g4225(csa_tree_add_95_22_pad_groupi_n_1495 ,csa_tree_add_95_22_pad_groupi_n_1449 ,csa_tree_add_95_22_pad_groupi_n_1481);
  nor csa_tree_add_95_22_pad_groupi_g4226(csa_tree_add_95_22_pad_groupi_n_1494 ,csa_tree_add_95_22_pad_groupi_n_1442 ,csa_tree_add_95_22_pad_groupi_n_1469);
  not csa_tree_add_95_22_pad_groupi_g4227(csa_tree_add_95_22_pad_groupi_n_1493 ,csa_tree_add_95_22_pad_groupi_n_1492);
  not csa_tree_add_95_22_pad_groupi_g4228(csa_tree_add_95_22_pad_groupi_n_1491 ,csa_tree_add_95_22_pad_groupi_n_1490);
  not csa_tree_add_95_22_pad_groupi_g4229(csa_tree_add_95_22_pad_groupi_n_1489 ,csa_tree_add_95_22_pad_groupi_n_1488);
  not csa_tree_add_95_22_pad_groupi_g4230(csa_tree_add_95_22_pad_groupi_n_1487 ,csa_tree_add_95_22_pad_groupi_n_1486);
  not csa_tree_add_95_22_pad_groupi_g4231(csa_tree_add_95_22_pad_groupi_n_1485 ,csa_tree_add_95_22_pad_groupi_n_1484);
  xnor csa_tree_add_95_22_pad_groupi_g4232(csa_tree_add_95_22_pad_groupi_n_1483 ,csa_tree_add_95_22_pad_groupi_n_1440 ,csa_tree_add_95_22_pad_groupi_n_1445);
  xnor csa_tree_add_95_22_pad_groupi_g4233(csa_tree_add_95_22_pad_groupi_n_1482 ,csa_tree_add_95_22_pad_groupi_n_1419 ,csa_tree_add_95_22_pad_groupi_n_1444);
  xnor csa_tree_add_95_22_pad_groupi_g4234(csa_tree_add_95_22_pad_groupi_n_1492 ,csa_tree_add_95_22_pad_groupi_n_1387 ,csa_tree_add_95_22_pad_groupi_n_1438);
  xnor csa_tree_add_95_22_pad_groupi_g4235(csa_tree_add_95_22_pad_groupi_n_1490 ,csa_tree_add_95_22_pad_groupi_n_1400 ,csa_tree_add_95_22_pad_groupi_n_1433);
  xnor csa_tree_add_95_22_pad_groupi_g4236(csa_tree_add_95_22_pad_groupi_n_1488 ,csa_tree_add_95_22_pad_groupi_n_1401 ,csa_tree_add_95_22_pad_groupi_n_1436);
  xnor csa_tree_add_95_22_pad_groupi_g4237(csa_tree_add_95_22_pad_groupi_n_1486 ,csa_tree_add_95_22_pad_groupi_n_1402 ,csa_tree_add_95_22_pad_groupi_n_1437);
  xnor csa_tree_add_95_22_pad_groupi_g4238(csa_tree_add_95_22_pad_groupi_n_1484 ,csa_tree_add_95_22_pad_groupi_n_1403 ,csa_tree_add_95_22_pad_groupi_n_1435);
  not csa_tree_add_95_22_pad_groupi_g4239(csa_tree_add_95_22_pad_groupi_n_1479 ,csa_tree_add_95_22_pad_groupi_n_1480);
  not csa_tree_add_95_22_pad_groupi_g4240(csa_tree_add_95_22_pad_groupi_n_1477 ,csa_tree_add_95_22_pad_groupi_n_1476);
  not csa_tree_add_95_22_pad_groupi_g4241(csa_tree_add_95_22_pad_groupi_n_1474 ,csa_tree_add_95_22_pad_groupi_n_1475);
  not csa_tree_add_95_22_pad_groupi_g4242(csa_tree_add_95_22_pad_groupi_n_1473 ,csa_tree_add_95_22_pad_groupi_n_1472);
  or csa_tree_add_95_22_pad_groupi_g4243(csa_tree_add_95_22_pad_groupi_n_1471 ,csa_tree_add_95_22_pad_groupi_n_1418 ,csa_tree_add_95_22_pad_groupi_n_1443);
  nor csa_tree_add_95_22_pad_groupi_g4244(csa_tree_add_95_22_pad_groupi_n_1470 ,csa_tree_add_95_22_pad_groupi_n_1419 ,csa_tree_add_95_22_pad_groupi_n_1444);
  and csa_tree_add_95_22_pad_groupi_g4245(csa_tree_add_95_22_pad_groupi_n_1481 ,csa_tree_add_95_22_pad_groupi_n_1371 ,csa_tree_add_95_22_pad_groupi_n_1439);
  or csa_tree_add_95_22_pad_groupi_g4246(csa_tree_add_95_22_pad_groupi_n_1480 ,csa_tree_add_95_22_pad_groupi_n_1424 ,csa_tree_add_95_22_pad_groupi_n_1456);
  and csa_tree_add_95_22_pad_groupi_g4247(csa_tree_add_95_22_pad_groupi_n_1478 ,csa_tree_add_95_22_pad_groupi_n_1431 ,csa_tree_add_95_22_pad_groupi_n_1454);
  or csa_tree_add_95_22_pad_groupi_g4248(csa_tree_add_95_22_pad_groupi_n_1476 ,csa_tree_add_95_22_pad_groupi_n_1422 ,csa_tree_add_95_22_pad_groupi_n_1455);
  or csa_tree_add_95_22_pad_groupi_g4249(csa_tree_add_95_22_pad_groupi_n_1475 ,csa_tree_add_95_22_pad_groupi_n_1429 ,csa_tree_add_95_22_pad_groupi_n_1458);
  or csa_tree_add_95_22_pad_groupi_g4250(csa_tree_add_95_22_pad_groupi_n_1472 ,csa_tree_add_95_22_pad_groupi_n_1426 ,csa_tree_add_95_22_pad_groupi_n_1457);
  not csa_tree_add_95_22_pad_groupi_g4251(csa_tree_add_95_22_pad_groupi_n_1469 ,csa_tree_add_95_22_pad_groupi_n_6);
  not csa_tree_add_95_22_pad_groupi_g4252(csa_tree_add_95_22_pad_groupi_n_1468 ,csa_tree_add_95_22_pad_groupi_n_1467);
  not csa_tree_add_95_22_pad_groupi_g4253(csa_tree_add_95_22_pad_groupi_n_1466 ,csa_tree_add_95_22_pad_groupi_n_1465);
  and csa_tree_add_95_22_pad_groupi_g4254(csa_tree_add_95_22_pad_groupi_n_1464 ,csa_tree_add_95_22_pad_groupi_n_1440 ,csa_tree_add_95_22_pad_groupi_n_1446);
  nor csa_tree_add_95_22_pad_groupi_g4255(csa_tree_add_95_22_pad_groupi_n_1463 ,csa_tree_add_95_22_pad_groupi_n_1440 ,csa_tree_add_95_22_pad_groupi_n_1446);
  xnor csa_tree_add_95_22_pad_groupi_g4256(csa_tree_add_95_22_pad_groupi_n_1462 ,csa_tree_add_95_22_pad_groupi_n_1432 ,csa_tree_add_95_22_pad_groupi_n_1413);
  xnor csa_tree_add_95_22_pad_groupi_g4257(csa_tree_add_95_22_pad_groupi_n_1461 ,csa_tree_add_95_22_pad_groupi_n_1397 ,csa_tree_add_95_22_pad_groupi_n_1417);
  xnor csa_tree_add_95_22_pad_groupi_g4258(csa_tree_add_95_22_pad_groupi_n_1460 ,csa_tree_add_95_22_pad_groupi_n_1367 ,csa_tree_add_95_22_pad_groupi_n_1415);
  xnor csa_tree_add_95_22_pad_groupi_g4260(csa_tree_add_95_22_pad_groupi_n_1467 ,csa_tree_add_95_22_pad_groupi_n_1384 ,csa_tree_add_95_22_pad_groupi_n_1405);
  xnor csa_tree_add_95_22_pad_groupi_g4261(csa_tree_add_95_22_pad_groupi_n_1465 ,csa_tree_add_95_22_pad_groupi_n_1295 ,csa_tree_add_95_22_pad_groupi_n_5);
  or csa_tree_add_95_22_pad_groupi_g4262(csa_tree_add_95_22_pad_groupi_n_1459 ,csa_tree_add_95_22_pad_groupi_n_1432 ,csa_tree_add_95_22_pad_groupi_n_1413);
  and csa_tree_add_95_22_pad_groupi_g4263(csa_tree_add_95_22_pad_groupi_n_1458 ,csa_tree_add_95_22_pad_groupi_n_1401 ,csa_tree_add_95_22_pad_groupi_n_1427);
  and csa_tree_add_95_22_pad_groupi_g4264(csa_tree_add_95_22_pad_groupi_n_1457 ,csa_tree_add_95_22_pad_groupi_n_1402 ,csa_tree_add_95_22_pad_groupi_n_1425);
  and csa_tree_add_95_22_pad_groupi_g4265(csa_tree_add_95_22_pad_groupi_n_1456 ,csa_tree_add_95_22_pad_groupi_n_1387 ,csa_tree_add_95_22_pad_groupi_n_1423);
  and csa_tree_add_95_22_pad_groupi_g4266(csa_tree_add_95_22_pad_groupi_n_1455 ,csa_tree_add_95_22_pad_groupi_n_1403 ,csa_tree_add_95_22_pad_groupi_n_1421);
  or csa_tree_add_95_22_pad_groupi_g4267(csa_tree_add_95_22_pad_groupi_n_1454 ,csa_tree_add_95_22_pad_groupi_n_1430 ,csa_tree_add_95_22_pad_groupi_n_1386);
  and csa_tree_add_95_22_pad_groupi_g4268(csa_tree_add_95_22_pad_groupi_n_1453 ,csa_tree_add_95_22_pad_groupi_n_1432 ,csa_tree_add_95_22_pad_groupi_n_1413);
  or csa_tree_add_95_22_pad_groupi_g4269(csa_tree_add_95_22_pad_groupi_n_1452 ,csa_tree_add_95_22_pad_groupi_n_1396 ,csa_tree_add_95_22_pad_groupi_n_1416);
  nor csa_tree_add_95_22_pad_groupi_g4270(csa_tree_add_95_22_pad_groupi_n_1451 ,csa_tree_add_95_22_pad_groupi_n_1397 ,csa_tree_add_95_22_pad_groupi_n_1417);
  or csa_tree_add_95_22_pad_groupi_g4271(csa_tree_add_95_22_pad_groupi_n_1450 ,csa_tree_add_95_22_pad_groupi_n_1367 ,csa_tree_add_95_22_pad_groupi_n_1414);
  nor csa_tree_add_95_22_pad_groupi_g4272(csa_tree_add_95_22_pad_groupi_n_1449 ,csa_tree_add_95_22_pad_groupi_n_1366 ,csa_tree_add_95_22_pad_groupi_n_1415);
  not csa_tree_add_95_22_pad_groupi_g4273(csa_tree_add_95_22_pad_groupi_n_1448 ,csa_tree_add_95_22_pad_groupi_n_1447);
  not csa_tree_add_95_22_pad_groupi_g4274(csa_tree_add_95_22_pad_groupi_n_1446 ,csa_tree_add_95_22_pad_groupi_n_1445);
  not csa_tree_add_95_22_pad_groupi_g4275(csa_tree_add_95_22_pad_groupi_n_1444 ,csa_tree_add_95_22_pad_groupi_n_1443);
  not csa_tree_add_95_22_pad_groupi_g4276(csa_tree_add_95_22_pad_groupi_n_1441 ,csa_tree_add_95_22_pad_groupi_n_1442);
  or csa_tree_add_95_22_pad_groupi_g4277(csa_tree_add_95_22_pad_groupi_n_1439 ,csa_tree_add_95_22_pad_groupi_n_1372 ,csa_tree_add_95_22_pad_groupi_n_1428);
  xnor csa_tree_add_95_22_pad_groupi_g4278(csa_tree_add_95_22_pad_groupi_n_1438 ,csa_tree_add_95_22_pad_groupi_n_1291 ,csa_tree_add_95_22_pad_groupi_n_1379);
  xnor csa_tree_add_95_22_pad_groupi_g4279(csa_tree_add_95_22_pad_groupi_n_1437 ,csa_tree_add_95_22_pad_groupi_n_1293 ,csa_tree_add_95_22_pad_groupi_n_1381);
  xnor csa_tree_add_95_22_pad_groupi_g4280(csa_tree_add_95_22_pad_groupi_n_1436 ,csa_tree_add_95_22_pad_groupi_n_1301 ,csa_tree_add_95_22_pad_groupi_n_1376);
  xnor csa_tree_add_95_22_pad_groupi_g4281(csa_tree_add_95_22_pad_groupi_n_1435 ,csa_tree_add_95_22_pad_groupi_n_1303 ,csa_tree_add_95_22_pad_groupi_n_1383);
  xnor csa_tree_add_95_22_pad_groupi_g4282(csa_tree_add_95_22_pad_groupi_n_1434 ,csa_tree_add_95_22_pad_groupi_n_1377 ,csa_tree_add_95_22_pad_groupi_n_1398);
  xnor csa_tree_add_95_22_pad_groupi_g4283(csa_tree_add_95_22_pad_groupi_n_1433 ,csa_tree_add_95_22_pad_groupi_n_1298 ,csa_tree_add_95_22_pad_groupi_n_1386);
  or csa_tree_add_95_22_pad_groupi_g4284(csa_tree_add_95_22_pad_groupi_n_1447 ,csa_tree_add_95_22_pad_groupi_n_1340 ,csa_tree_add_95_22_pad_groupi_n_1420);
  xnor csa_tree_add_95_22_pad_groupi_g4285(csa_tree_add_95_22_pad_groupi_n_1445 ,csa_tree_add_95_22_pad_groupi_n_1334 ,csa_tree_add_95_22_pad_groupi_n_1370);
  xnor csa_tree_add_95_22_pad_groupi_g4286(csa_tree_add_95_22_pad_groupi_n_1443 ,csa_tree_add_95_22_pad_groupi_n_1385 ,csa_tree_add_95_22_pad_groupi_n_1369);
  or csa_tree_add_95_22_pad_groupi_g4287(csa_tree_add_95_22_pad_groupi_n_1442 ,csa_tree_add_95_22_pad_groupi_n_1374 ,csa_tree_add_95_22_pad_groupi_n_1409);
  and csa_tree_add_95_22_pad_groupi_g4288(csa_tree_add_95_22_pad_groupi_n_1440 ,csa_tree_add_95_22_pad_groupi_n_1395 ,csa_tree_add_95_22_pad_groupi_n_1408);
  or csa_tree_add_95_22_pad_groupi_g4289(csa_tree_add_95_22_pad_groupi_n_1431 ,csa_tree_add_95_22_pad_groupi_n_1297 ,csa_tree_add_95_22_pad_groupi_n_1399);
  nor csa_tree_add_95_22_pad_groupi_g4290(csa_tree_add_95_22_pad_groupi_n_1430 ,csa_tree_add_95_22_pad_groupi_n_1298 ,csa_tree_add_95_22_pad_groupi_n_1400);
  nor csa_tree_add_95_22_pad_groupi_g4291(csa_tree_add_95_22_pad_groupi_n_1429 ,csa_tree_add_95_22_pad_groupi_n_1300 ,csa_tree_add_95_22_pad_groupi_n_1376);
  nor csa_tree_add_95_22_pad_groupi_g4292(csa_tree_add_95_22_pad_groupi_n_1428 ,csa_tree_add_95_22_pad_groupi_n_1363 ,csa_tree_add_95_22_pad_groupi_n_1394);
  or csa_tree_add_95_22_pad_groupi_g4293(csa_tree_add_95_22_pad_groupi_n_1427 ,csa_tree_add_95_22_pad_groupi_n_1301 ,csa_tree_add_95_22_pad_groupi_n_1375);
  nor csa_tree_add_95_22_pad_groupi_g4294(csa_tree_add_95_22_pad_groupi_n_1426 ,csa_tree_add_95_22_pad_groupi_n_1292 ,csa_tree_add_95_22_pad_groupi_n_1381);
  or csa_tree_add_95_22_pad_groupi_g4295(csa_tree_add_95_22_pad_groupi_n_1425 ,csa_tree_add_95_22_pad_groupi_n_1293 ,csa_tree_add_95_22_pad_groupi_n_1380);
  nor csa_tree_add_95_22_pad_groupi_g4296(csa_tree_add_95_22_pad_groupi_n_1424 ,csa_tree_add_95_22_pad_groupi_n_1290 ,csa_tree_add_95_22_pad_groupi_n_1379);
  or csa_tree_add_95_22_pad_groupi_g4297(csa_tree_add_95_22_pad_groupi_n_1423 ,csa_tree_add_95_22_pad_groupi_n_1291 ,csa_tree_add_95_22_pad_groupi_n_1378);
  nor csa_tree_add_95_22_pad_groupi_g4298(csa_tree_add_95_22_pad_groupi_n_1422 ,csa_tree_add_95_22_pad_groupi_n_1302 ,csa_tree_add_95_22_pad_groupi_n_1383);
  or csa_tree_add_95_22_pad_groupi_g4299(csa_tree_add_95_22_pad_groupi_n_1421 ,csa_tree_add_95_22_pad_groupi_n_1303 ,csa_tree_add_95_22_pad_groupi_n_1382);
  nor csa_tree_add_95_22_pad_groupi_g4300(csa_tree_add_95_22_pad_groupi_n_1420 ,csa_tree_add_95_22_pad_groupi_n_1355 ,csa_tree_add_95_22_pad_groupi_n_1385);
  or csa_tree_add_95_22_pad_groupi_g4301(csa_tree_add_95_22_pad_groupi_n_1432 ,csa_tree_add_95_22_pad_groupi_n_1365 ,csa_tree_add_95_22_pad_groupi_n_1391);
  not csa_tree_add_95_22_pad_groupi_g4302(csa_tree_add_95_22_pad_groupi_n_1419 ,csa_tree_add_95_22_pad_groupi_n_1418);
  not csa_tree_add_95_22_pad_groupi_g4303(csa_tree_add_95_22_pad_groupi_n_1417 ,csa_tree_add_95_22_pad_groupi_n_1416);
  not csa_tree_add_95_22_pad_groupi_g4304(csa_tree_add_95_22_pad_groupi_n_1415 ,csa_tree_add_95_22_pad_groupi_n_1414);
  not csa_tree_add_95_22_pad_groupi_g4305(csa_tree_add_95_22_pad_groupi_n_1412 ,csa_tree_add_95_22_pad_groupi_n_1411);
  or csa_tree_add_95_22_pad_groupi_g4306(csa_tree_add_95_22_pad_groupi_n_1410 ,csa_tree_add_95_22_pad_groupi_n_1377 ,csa_tree_add_95_22_pad_groupi_n_1398);
  nor csa_tree_add_95_22_pad_groupi_g4307(csa_tree_add_95_22_pad_groupi_n_1409 ,csa_tree_add_95_22_pad_groupi_n_1384 ,csa_tree_add_95_22_pad_groupi_n_1392);
  or csa_tree_add_95_22_pad_groupi_g4308(csa_tree_add_95_22_pad_groupi_n_1408 ,csa_tree_add_95_22_pad_groupi_n_1368 ,csa_tree_add_95_22_pad_groupi_n_1373);
  and csa_tree_add_95_22_pad_groupi_g4309(csa_tree_add_95_22_pad_groupi_n_1407 ,csa_tree_add_95_22_pad_groupi_n_1377 ,csa_tree_add_95_22_pad_groupi_n_1398);
  xnor csa_tree_add_95_22_pad_groupi_g4310(csa_tree_add_95_22_pad_groupi_n_1406 ,csa_tree_add_95_22_pad_groupi_n_1280 ,csa_tree_add_95_22_pad_groupi_n_1346);
  xnor csa_tree_add_95_22_pad_groupi_g4312(csa_tree_add_95_22_pad_groupi_n_1405 ,csa_tree_add_95_22_pad_groupi_n_1304 ,csa_tree_add_95_22_pad_groupi_n_1348);
  xnor csa_tree_add_95_22_pad_groupi_g4313(csa_tree_add_95_22_pad_groupi_n_1404 ,csa_tree_add_95_22_pad_groupi_n_1309 ,csa_tree_add_95_22_pad_groupi_n_1345);
  and csa_tree_add_95_22_pad_groupi_g4314(csa_tree_add_95_22_pad_groupi_n_1418 ,csa_tree_add_95_22_pad_groupi_n_1354 ,csa_tree_add_95_22_pad_groupi_n_1390);
  xnor csa_tree_add_95_22_pad_groupi_g4315(csa_tree_add_95_22_pad_groupi_n_1416 ,csa_tree_add_95_22_pad_groupi_n_1311 ,csa_tree_add_95_22_pad_groupi_n_1337);
  xnor csa_tree_add_95_22_pad_groupi_g4316(csa_tree_add_95_22_pad_groupi_n_1414 ,csa_tree_add_95_22_pad_groupi_n_1320 ,csa_tree_add_95_22_pad_groupi_n_1335);
  xnor csa_tree_add_95_22_pad_groupi_g4317(csa_tree_add_95_22_pad_groupi_n_1413 ,csa_tree_add_95_22_pad_groupi_n_1333 ,csa_tree_add_95_22_pad_groupi_n_1338);
  and csa_tree_add_95_22_pad_groupi_g4318(csa_tree_add_95_22_pad_groupi_n_1411 ,csa_tree_add_95_22_pad_groupi_n_1356 ,csa_tree_add_95_22_pad_groupi_n_1388);
  not csa_tree_add_95_22_pad_groupi_g4319(csa_tree_add_95_22_pad_groupi_n_1400 ,csa_tree_add_95_22_pad_groupi_n_1399);
  not csa_tree_add_95_22_pad_groupi_g4320(csa_tree_add_95_22_pad_groupi_n_1396 ,csa_tree_add_95_22_pad_groupi_n_1397);
  or csa_tree_add_95_22_pad_groupi_g4321(csa_tree_add_95_22_pad_groupi_n_1395 ,csa_tree_add_95_22_pad_groupi_n_1280 ,csa_tree_add_95_22_pad_groupi_n_1347);
  nor csa_tree_add_95_22_pad_groupi_g4322(csa_tree_add_95_22_pad_groupi_n_1394 ,csa_tree_add_95_22_pad_groupi_n_1362 ,csa_tree_add_95_22_pad_groupi_n_1361);
  and csa_tree_add_95_22_pad_groupi_g4323(csa_tree_add_95_22_pad_groupi_n_1393 ,csa_tree_add_95_22_pad_groupi_n_1309 ,csa_tree_add_95_22_pad_groupi_n_1345);
  and csa_tree_add_95_22_pad_groupi_g4324(csa_tree_add_95_22_pad_groupi_n_1392 ,csa_tree_add_95_22_pad_groupi_n_1304 ,csa_tree_add_95_22_pad_groupi_n_1349);
  and csa_tree_add_95_22_pad_groupi_g4325(csa_tree_add_95_22_pad_groupi_n_1391 ,csa_tree_add_95_22_pad_groupi_n_1334 ,csa_tree_add_95_22_pad_groupi_n_1360);
  or csa_tree_add_95_22_pad_groupi_g4326(csa_tree_add_95_22_pad_groupi_n_1390 ,csa_tree_add_95_22_pad_groupi_n_1353 ,csa_tree_add_95_22_pad_groupi_n_1350);
  or csa_tree_add_95_22_pad_groupi_g4327(csa_tree_add_95_22_pad_groupi_n_1389 ,csa_tree_add_95_22_pad_groupi_n_1309 ,csa_tree_add_95_22_pad_groupi_n_1345);
  or csa_tree_add_95_22_pad_groupi_g4328(csa_tree_add_95_22_pad_groupi_n_1388 ,csa_tree_add_95_22_pad_groupi_n_1305 ,csa_tree_add_95_22_pad_groupi_n_1342);
  or csa_tree_add_95_22_pad_groupi_g4329(csa_tree_add_95_22_pad_groupi_n_1403 ,csa_tree_add_95_22_pad_groupi_n_1246 ,csa_tree_add_95_22_pad_groupi_n_1359);
  or csa_tree_add_95_22_pad_groupi_g4330(csa_tree_add_95_22_pad_groupi_n_1402 ,csa_tree_add_95_22_pad_groupi_n_1230 ,csa_tree_add_95_22_pad_groupi_n_1343);
  or csa_tree_add_95_22_pad_groupi_g4331(csa_tree_add_95_22_pad_groupi_n_1401 ,csa_tree_add_95_22_pad_groupi_n_1232 ,csa_tree_add_95_22_pad_groupi_n_1339);
  and csa_tree_add_95_22_pad_groupi_g4332(csa_tree_add_95_22_pad_groupi_n_1399 ,csa_tree_add_95_22_pad_groupi_n_1254 ,csa_tree_add_95_22_pad_groupi_n_1364);
  or csa_tree_add_95_22_pad_groupi_g4333(csa_tree_add_95_22_pad_groupi_n_1398 ,csa_tree_add_95_22_pad_groupi_n_1329 ,csa_tree_add_95_22_pad_groupi_n_1357);
  or csa_tree_add_95_22_pad_groupi_g4334(csa_tree_add_95_22_pad_groupi_n_1397 ,csa_tree_add_95_22_pad_groupi_n_1323 ,csa_tree_add_95_22_pad_groupi_n_1358);
  not csa_tree_add_95_22_pad_groupi_g4335(csa_tree_add_95_22_pad_groupi_n_1383 ,csa_tree_add_95_22_pad_groupi_n_1382);
  not csa_tree_add_95_22_pad_groupi_g4336(csa_tree_add_95_22_pad_groupi_n_1381 ,csa_tree_add_95_22_pad_groupi_n_1380);
  not csa_tree_add_95_22_pad_groupi_g4337(csa_tree_add_95_22_pad_groupi_n_1379 ,csa_tree_add_95_22_pad_groupi_n_1378);
  not csa_tree_add_95_22_pad_groupi_g4338(csa_tree_add_95_22_pad_groupi_n_1376 ,csa_tree_add_95_22_pad_groupi_n_1375);
  nor csa_tree_add_95_22_pad_groupi_g4339(csa_tree_add_95_22_pad_groupi_n_1374 ,csa_tree_add_95_22_pad_groupi_n_1304 ,csa_tree_add_95_22_pad_groupi_n_1349);
  and csa_tree_add_95_22_pad_groupi_g4340(csa_tree_add_95_22_pad_groupi_n_1373 ,csa_tree_add_95_22_pad_groupi_n_1280 ,csa_tree_add_95_22_pad_groupi_n_1347);
  nor csa_tree_add_95_22_pad_groupi_g4341(csa_tree_add_95_22_pad_groupi_n_1372 ,csa_tree_add_95_22_pad_groupi_n_1306 ,csa_tree_add_95_22_pad_groupi_n_1352);
  or csa_tree_add_95_22_pad_groupi_g4342(csa_tree_add_95_22_pad_groupi_n_1371 ,csa_tree_add_95_22_pad_groupi_n_1307 ,csa_tree_add_95_22_pad_groupi_n_1351);
  xnor csa_tree_add_95_22_pad_groupi_g4343(csa_tree_add_95_22_pad_groupi_n_1370 ,csa_tree_add_95_22_pad_groupi_n_1261 ,csa_tree_add_95_22_pad_groupi_n_1310);
  xnor csa_tree_add_95_22_pad_groupi_g4344(csa_tree_add_95_22_pad_groupi_n_1369 ,csa_tree_add_95_22_pad_groupi_n_1299 ,csa_tree_add_95_22_pad_groupi_n_1330);
  or csa_tree_add_95_22_pad_groupi_g4345(csa_tree_add_95_22_pad_groupi_n_1387 ,csa_tree_add_95_22_pad_groupi_n_1227 ,csa_tree_add_95_22_pad_groupi_n_1341);
  xnor csa_tree_add_95_22_pad_groupi_g4346(csa_tree_add_95_22_pad_groupi_n_1386 ,csa_tree_add_95_22_pad_groupi_n_1317 ,csa_tree_add_95_22_pad_groupi_n_1273);
  xnor csa_tree_add_95_22_pad_groupi_g4347(csa_tree_add_95_22_pad_groupi_n_1385 ,csa_tree_add_95_22_pad_groupi_n_1316 ,csa_tree_add_95_22_pad_groupi_n_1268);
  and csa_tree_add_95_22_pad_groupi_g4348(csa_tree_add_95_22_pad_groupi_n_1384 ,csa_tree_add_95_22_pad_groupi_n_1225 ,csa_tree_add_95_22_pad_groupi_n_1344);
  xnor csa_tree_add_95_22_pad_groupi_g4349(csa_tree_add_95_22_pad_groupi_n_1382 ,csa_tree_add_95_22_pad_groupi_n_1313 ,csa_tree_add_95_22_pad_groupi_n_1266);
  xnor csa_tree_add_95_22_pad_groupi_g4350(csa_tree_add_95_22_pad_groupi_n_1380 ,csa_tree_add_95_22_pad_groupi_n_1315 ,csa_tree_add_95_22_pad_groupi_n_1270);
  xnor csa_tree_add_95_22_pad_groupi_g4351(csa_tree_add_95_22_pad_groupi_n_1378 ,csa_tree_add_95_22_pad_groupi_n_1314 ,csa_tree_add_95_22_pad_groupi_n_1267);
  xnor csa_tree_add_95_22_pad_groupi_g4352(csa_tree_add_95_22_pad_groupi_n_1377 ,csa_tree_add_95_22_pad_groupi_n_1262 ,csa_tree_add_95_22_pad_groupi_n_1308);
  xnor csa_tree_add_95_22_pad_groupi_g4353(csa_tree_add_95_22_pad_groupi_n_1375 ,csa_tree_add_95_22_pad_groupi_n_1318 ,csa_tree_add_95_22_pad_groupi_n_1271);
  not csa_tree_add_95_22_pad_groupi_g4355(csa_tree_add_95_22_pad_groupi_n_1367 ,csa_tree_add_95_22_pad_groupi_n_1366);
  and csa_tree_add_95_22_pad_groupi_g4356(csa_tree_add_95_22_pad_groupi_n_1365 ,csa_tree_add_95_22_pad_groupi_n_1261 ,csa_tree_add_95_22_pad_groupi_n_1310);
  or csa_tree_add_95_22_pad_groupi_g4357(csa_tree_add_95_22_pad_groupi_n_1364 ,csa_tree_add_95_22_pad_groupi_n_1224 ,csa_tree_add_95_22_pad_groupi_n_1319);
  and csa_tree_add_95_22_pad_groupi_g4358(csa_tree_add_95_22_pad_groupi_n_1363 ,csa_tree_add_95_22_pad_groupi_n_1265 ,csa_tree_add_95_22_pad_groupi_n_1321);
  nor csa_tree_add_95_22_pad_groupi_g4359(csa_tree_add_95_22_pad_groupi_n_1362 ,csa_tree_add_95_22_pad_groupi_n_1265 ,csa_tree_add_95_22_pad_groupi_n_1321);
  nor csa_tree_add_95_22_pad_groupi_g4360(csa_tree_add_95_22_pad_groupi_n_1361 ,csa_tree_add_95_22_pad_groupi_n_1285 ,csa_tree_add_95_22_pad_groupi_n_1326);
  or csa_tree_add_95_22_pad_groupi_g4361(csa_tree_add_95_22_pad_groupi_n_1360 ,csa_tree_add_95_22_pad_groupi_n_1261 ,csa_tree_add_95_22_pad_groupi_n_1310);
  nor csa_tree_add_95_22_pad_groupi_g4362(csa_tree_add_95_22_pad_groupi_n_1359 ,csa_tree_add_95_22_pad_groupi_n_1245 ,csa_tree_add_95_22_pad_groupi_n_1316);
  nor csa_tree_add_95_22_pad_groupi_g4363(csa_tree_add_95_22_pad_groupi_n_1358 ,csa_tree_add_95_22_pad_groupi_n_1328 ,csa_tree_add_95_22_pad_groupi_n_1320);
  nor csa_tree_add_95_22_pad_groupi_g4364(csa_tree_add_95_22_pad_groupi_n_1357 ,csa_tree_add_95_22_pad_groupi_n_1333 ,csa_tree_add_95_22_pad_groupi_n_1322);
  or csa_tree_add_95_22_pad_groupi_g4365(csa_tree_add_95_22_pad_groupi_n_1356 ,csa_tree_add_95_22_pad_groupi_n_1278 ,csa_tree_add_95_22_pad_groupi_n_1312);
  nor csa_tree_add_95_22_pad_groupi_g4366(csa_tree_add_95_22_pad_groupi_n_1355 ,csa_tree_add_95_22_pad_groupi_n_1299 ,csa_tree_add_95_22_pad_groupi_n_1330);
  or csa_tree_add_95_22_pad_groupi_g4367(csa_tree_add_95_22_pad_groupi_n_1354 ,csa_tree_add_95_22_pad_groupi_n_1294 ,csa_tree_add_95_22_pad_groupi_n_1332);
  nor csa_tree_add_95_22_pad_groupi_g4368(csa_tree_add_95_22_pad_groupi_n_1353 ,csa_tree_add_95_22_pad_groupi_n_1295 ,csa_tree_add_95_22_pad_groupi_n_1331);
  and csa_tree_add_95_22_pad_groupi_g4369(csa_tree_add_95_22_pad_groupi_n_1368 ,csa_tree_add_95_22_pad_groupi_n_1243 ,csa_tree_add_95_22_pad_groupi_n_1324);
  or csa_tree_add_95_22_pad_groupi_g4370(csa_tree_add_95_22_pad_groupi_n_1366 ,csa_tree_add_95_22_pad_groupi_n_1185 ,csa_tree_add_95_22_pad_groupi_n_1327);
  not csa_tree_add_95_22_pad_groupi_g4371(csa_tree_add_95_22_pad_groupi_n_1352 ,csa_tree_add_95_22_pad_groupi_n_1351);
  not csa_tree_add_95_22_pad_groupi_g4373(csa_tree_add_95_22_pad_groupi_n_1349 ,csa_tree_add_95_22_pad_groupi_n_1348);
  not csa_tree_add_95_22_pad_groupi_g4374(csa_tree_add_95_22_pad_groupi_n_1347 ,csa_tree_add_95_22_pad_groupi_n_1346);
  or csa_tree_add_95_22_pad_groupi_g4375(csa_tree_add_95_22_pad_groupi_n_1344 ,csa_tree_add_95_22_pad_groupi_n_1223 ,csa_tree_add_95_22_pad_groupi_n_1317);
  and csa_tree_add_95_22_pad_groupi_g4376(csa_tree_add_95_22_pad_groupi_n_1343 ,csa_tree_add_95_22_pad_groupi_n_1228 ,csa_tree_add_95_22_pad_groupi_n_1314);
  and csa_tree_add_95_22_pad_groupi_g4377(csa_tree_add_95_22_pad_groupi_n_1342 ,csa_tree_add_95_22_pad_groupi_n_1278 ,csa_tree_add_95_22_pad_groupi_n_1312);
  and csa_tree_add_95_22_pad_groupi_g4378(csa_tree_add_95_22_pad_groupi_n_1341 ,csa_tree_add_95_22_pad_groupi_n_1226 ,csa_tree_add_95_22_pad_groupi_n_1313);
  and csa_tree_add_95_22_pad_groupi_g4379(csa_tree_add_95_22_pad_groupi_n_1340 ,csa_tree_add_95_22_pad_groupi_n_1299 ,csa_tree_add_95_22_pad_groupi_n_1330);
  and csa_tree_add_95_22_pad_groupi_g4380(csa_tree_add_95_22_pad_groupi_n_1339 ,csa_tree_add_95_22_pad_groupi_n_1231 ,csa_tree_add_95_22_pad_groupi_n_1315);
  xnor csa_tree_add_95_22_pad_groupi_g4381(csa_tree_add_95_22_pad_groupi_n_1338 ,csa_tree_add_95_22_pad_groupi_n_1201 ,csa_tree_add_95_22_pad_groupi_n_1279);
  xnor csa_tree_add_95_22_pad_groupi_g4382(csa_tree_add_95_22_pad_groupi_n_1351 ,csa_tree_add_95_22_pad_groupi_n_1281 ,csa_tree_add_95_22_pad_groupi_n_1211);
  xor csa_tree_add_95_22_pad_groupi_g4383(csa_tree_add_95_22_pad_groupi_n_1337 ,csa_tree_add_95_22_pad_groupi_n_1278 ,csa_tree_add_95_22_pad_groupi_n_1305);
  xnor csa_tree_add_95_22_pad_groupi_g4384(csa_tree_add_95_22_pad_groupi_n_1336 ,csa_tree_add_95_22_pad_groupi_n_1075 ,csa_tree_add_95_22_pad_groupi_n_1274);
  xnor csa_tree_add_95_22_pad_groupi_g4385(csa_tree_add_95_22_pad_groupi_n_1335 ,csa_tree_add_95_22_pad_groupi_n_1235 ,csa_tree_add_95_22_pad_groupi_n_1296);
  xnor csa_tree_add_95_22_pad_groupi_g4386(csa_tree_add_95_22_pad_groupi_n_1350 ,csa_tree_add_95_22_pad_groupi_n_1264 ,csa_tree_add_95_22_pad_groupi_n_1272);
  xnor csa_tree_add_95_22_pad_groupi_g4387(csa_tree_add_95_22_pad_groupi_n_1348 ,csa_tree_add_95_22_pad_groupi_n_1282 ,csa_tree_add_95_22_pad_groupi_n_1269);
  xnor csa_tree_add_95_22_pad_groupi_g4388(csa_tree_add_95_22_pad_groupi_n_1346 ,csa_tree_add_95_22_pad_groupi_n_1263 ,csa_tree_add_95_22_pad_groupi_n_1275);
  or csa_tree_add_95_22_pad_groupi_g4389(csa_tree_add_95_22_pad_groupi_n_1345 ,csa_tree_add_95_22_pad_groupi_n_1277 ,csa_tree_add_95_22_pad_groupi_n_1325);
  not csa_tree_add_95_22_pad_groupi_g4390(csa_tree_add_95_22_pad_groupi_n_1332 ,csa_tree_add_95_22_pad_groupi_n_1331);
  nor csa_tree_add_95_22_pad_groupi_g4391(csa_tree_add_95_22_pad_groupi_n_1329 ,csa_tree_add_95_22_pad_groupi_n_1202 ,csa_tree_add_95_22_pad_groupi_n_1279);
  nor csa_tree_add_95_22_pad_groupi_g4392(csa_tree_add_95_22_pad_groupi_n_1328 ,csa_tree_add_95_22_pad_groupi_n_1235 ,csa_tree_add_95_22_pad_groupi_n_1296);
  nor csa_tree_add_95_22_pad_groupi_g4393(csa_tree_add_95_22_pad_groupi_n_1327 ,csa_tree_add_95_22_pad_groupi_n_1184 ,csa_tree_add_95_22_pad_groupi_n_1281);
  nor csa_tree_add_95_22_pad_groupi_g4394(csa_tree_add_95_22_pad_groupi_n_1326 ,csa_tree_add_95_22_pad_groupi_n_1287 ,csa_tree_add_95_22_pad_groupi_n_1288);
  nor csa_tree_add_95_22_pad_groupi_g4395(csa_tree_add_95_22_pad_groupi_n_1325 ,csa_tree_add_95_22_pad_groupi_n_1276 ,csa_tree_add_95_22_pad_groupi_n_1262);
  or csa_tree_add_95_22_pad_groupi_g4396(csa_tree_add_95_22_pad_groupi_n_1324 ,csa_tree_add_95_22_pad_groupi_n_1252 ,csa_tree_add_95_22_pad_groupi_n_1283);
  and csa_tree_add_95_22_pad_groupi_g4397(csa_tree_add_95_22_pad_groupi_n_1323 ,csa_tree_add_95_22_pad_groupi_n_1235 ,csa_tree_add_95_22_pad_groupi_n_1296);
  and csa_tree_add_95_22_pad_groupi_g4398(csa_tree_add_95_22_pad_groupi_n_1322 ,csa_tree_add_95_22_pad_groupi_n_1202 ,csa_tree_add_95_22_pad_groupi_n_1279);
  or csa_tree_add_95_22_pad_groupi_g4399(csa_tree_add_95_22_pad_groupi_n_1334 ,csa_tree_add_95_22_pad_groupi_n_1240 ,csa_tree_add_95_22_pad_groupi_n_1284);
  and csa_tree_add_95_22_pad_groupi_g4400(csa_tree_add_95_22_pad_groupi_n_1333 ,csa_tree_add_95_22_pad_groupi_n_1156 ,csa_tree_add_95_22_pad_groupi_n_1286);
  xnor csa_tree_add_95_22_pad_groupi_g4401(csa_tree_add_95_22_pad_groupi_n_1331 ,csa_tree_add_95_22_pad_groupi_n_1039 ,csa_tree_add_95_22_pad_groupi_n_1216);
  or csa_tree_add_95_22_pad_groupi_g4402(csa_tree_add_95_22_pad_groupi_n_1330 ,csa_tree_add_95_22_pad_groupi_n_1242 ,csa_tree_add_95_22_pad_groupi_n_1289);
  not csa_tree_add_95_22_pad_groupi_g4403(csa_tree_add_95_22_pad_groupi_n_1319 ,csa_tree_add_95_22_pad_groupi_n_1318);
  not csa_tree_add_95_22_pad_groupi_g4404(csa_tree_add_95_22_pad_groupi_n_1312 ,csa_tree_add_95_22_pad_groupi_n_1311);
  xnor csa_tree_add_95_22_pad_groupi_g4405(csa_tree_add_95_22_pad_groupi_n_1321 ,csa_tree_add_95_22_pad_groupi_n_1176 ,csa_tree_add_95_22_pad_groupi_n_1210);
  xnor csa_tree_add_95_22_pad_groupi_g4406(csa_tree_add_95_22_pad_groupi_n_1308 ,csa_tree_add_95_22_pad_groupi_n_1132 ,csa_tree_add_95_22_pad_groupi_n_1233);
  xnor csa_tree_add_95_22_pad_groupi_g4407(csa_tree_add_95_22_pad_groupi_n_1320 ,csa_tree_add_95_22_pad_groupi_n_1084 ,csa_tree_add_95_22_pad_groupi_n_1220);
  xnor csa_tree_add_95_22_pad_groupi_g4408(csa_tree_add_95_22_pad_groupi_n_1318 ,csa_tree_add_95_22_pad_groupi_n_1138 ,csa_tree_add_95_22_pad_groupi_n_1221);
  xnor csa_tree_add_95_22_pad_groupi_g4409(csa_tree_add_95_22_pad_groupi_n_1317 ,csa_tree_add_95_22_pad_groupi_n_1092 ,csa_tree_add_95_22_pad_groupi_n_1213);
  xnor csa_tree_add_95_22_pad_groupi_g4410(csa_tree_add_95_22_pad_groupi_n_1316 ,csa_tree_add_95_22_pad_groupi_n_1088 ,csa_tree_add_95_22_pad_groupi_n_1214);
  xnor csa_tree_add_95_22_pad_groupi_g4411(csa_tree_add_95_22_pad_groupi_n_1315 ,csa_tree_add_95_22_pad_groupi_n_1141 ,csa_tree_add_95_22_pad_groupi_n_1218);
  xnor csa_tree_add_95_22_pad_groupi_g4412(csa_tree_add_95_22_pad_groupi_n_1314 ,csa_tree_add_95_22_pad_groupi_n_1102 ,csa_tree_add_95_22_pad_groupi_n_1217);
  xnor csa_tree_add_95_22_pad_groupi_g4413(csa_tree_add_95_22_pad_groupi_n_1313 ,csa_tree_add_95_22_pad_groupi_n_1107 ,csa_tree_add_95_22_pad_groupi_n_1222);
  xnor csa_tree_add_95_22_pad_groupi_g4414(csa_tree_add_95_22_pad_groupi_n_1311 ,csa_tree_add_95_22_pad_groupi_n_1209 ,csa_tree_add_95_22_pad_groupi_n_1215);
  xnor csa_tree_add_95_22_pad_groupi_g4415(csa_tree_add_95_22_pad_groupi_n_1310 ,csa_tree_add_95_22_pad_groupi_n_1236 ,csa_tree_add_95_22_pad_groupi_n_1212);
  xnor csa_tree_add_95_22_pad_groupi_g4416(csa_tree_add_95_22_pad_groupi_n_1309 ,csa_tree_add_95_22_pad_groupi_n_1175 ,csa_tree_add_95_22_pad_groupi_n_1219);
  not csa_tree_add_95_22_pad_groupi_g4417(csa_tree_add_95_22_pad_groupi_n_1307 ,csa_tree_add_95_22_pad_groupi_n_1306);
  not csa_tree_add_95_22_pad_groupi_g4418(csa_tree_add_95_22_pad_groupi_n_1302 ,csa_tree_add_95_22_pad_groupi_n_1303);
  not csa_tree_add_95_22_pad_groupi_g4419(csa_tree_add_95_22_pad_groupi_n_1300 ,csa_tree_add_95_22_pad_groupi_n_1301);
  not csa_tree_add_95_22_pad_groupi_g4420(csa_tree_add_95_22_pad_groupi_n_1297 ,csa_tree_add_95_22_pad_groupi_n_1298);
  not csa_tree_add_95_22_pad_groupi_g4421(csa_tree_add_95_22_pad_groupi_n_1295 ,csa_tree_add_95_22_pad_groupi_n_1294);
  not csa_tree_add_95_22_pad_groupi_g4422(csa_tree_add_95_22_pad_groupi_n_1292 ,csa_tree_add_95_22_pad_groupi_n_1293);
  not csa_tree_add_95_22_pad_groupi_g4423(csa_tree_add_95_22_pad_groupi_n_1290 ,csa_tree_add_95_22_pad_groupi_n_1291);
  nor csa_tree_add_95_22_pad_groupi_g4424(csa_tree_add_95_22_pad_groupi_n_1289 ,csa_tree_add_95_22_pad_groupi_n_1247 ,csa_tree_add_95_22_pad_groupi_n_1264);
  nor csa_tree_add_95_22_pad_groupi_g4425(csa_tree_add_95_22_pad_groupi_n_1288 ,csa_tree_add_95_22_pad_groupi_n_1048 ,csa_tree_add_95_22_pad_groupi_n_1238);
  nor csa_tree_add_95_22_pad_groupi_g4426(csa_tree_add_95_22_pad_groupi_n_1287 ,csa_tree_add_95_22_pad_groupi_n_1178 ,csa_tree_add_95_22_pad_groupi_n_1251);
  or csa_tree_add_95_22_pad_groupi_g4427(csa_tree_add_95_22_pad_groupi_n_1286 ,csa_tree_add_95_22_pad_groupi_n_1150 ,csa_tree_add_95_22_pad_groupi_n_1237);
  nor csa_tree_add_95_22_pad_groupi_g4428(csa_tree_add_95_22_pad_groupi_n_1285 ,csa_tree_add_95_22_pad_groupi_n_1047 ,csa_tree_add_95_22_pad_groupi_n_1239);
  and csa_tree_add_95_22_pad_groupi_g4429(csa_tree_add_95_22_pad_groupi_n_1284 ,csa_tree_add_95_22_pad_groupi_n_1241 ,csa_tree_add_95_22_pad_groupi_n_1263);
  or csa_tree_add_95_22_pad_groupi_g4430(csa_tree_add_95_22_pad_groupi_n_1306 ,csa_tree_add_95_22_pad_groupi_n_1183 ,csa_tree_add_95_22_pad_groupi_n_1253);
  and csa_tree_add_95_22_pad_groupi_g4431(csa_tree_add_95_22_pad_groupi_n_1305 ,csa_tree_add_95_22_pad_groupi_n_1192 ,csa_tree_add_95_22_pad_groupi_n_1257);
  and csa_tree_add_95_22_pad_groupi_g4432(csa_tree_add_95_22_pad_groupi_n_1304 ,csa_tree_add_95_22_pad_groupi_n_1155 ,csa_tree_add_95_22_pad_groupi_n_1260);
  or csa_tree_add_95_22_pad_groupi_g4433(csa_tree_add_95_22_pad_groupi_n_1303 ,csa_tree_add_95_22_pad_groupi_n_1154 ,csa_tree_add_95_22_pad_groupi_n_1248);
  or csa_tree_add_95_22_pad_groupi_g4434(csa_tree_add_95_22_pad_groupi_n_1301 ,csa_tree_add_95_22_pad_groupi_n_1187 ,csa_tree_add_95_22_pad_groupi_n_1255);
  or csa_tree_add_95_22_pad_groupi_g4435(csa_tree_add_95_22_pad_groupi_n_1299 ,csa_tree_add_95_22_pad_groupi_n_1147 ,csa_tree_add_95_22_pad_groupi_n_1244);
  or csa_tree_add_95_22_pad_groupi_g4436(csa_tree_add_95_22_pad_groupi_n_1298 ,csa_tree_add_95_22_pad_groupi_n_1198 ,csa_tree_add_95_22_pad_groupi_n_1258);
  or csa_tree_add_95_22_pad_groupi_g4437(csa_tree_add_95_22_pad_groupi_n_1296 ,csa_tree_add_95_22_pad_groupi_n_1188 ,csa_tree_add_95_22_pad_groupi_n_1256);
  and csa_tree_add_95_22_pad_groupi_g4438(csa_tree_add_95_22_pad_groupi_n_1294 ,csa_tree_add_95_22_pad_groupi_n_1197 ,csa_tree_add_95_22_pad_groupi_n_1259);
  or csa_tree_add_95_22_pad_groupi_g4439(csa_tree_add_95_22_pad_groupi_n_1293 ,csa_tree_add_95_22_pad_groupi_n_1179 ,csa_tree_add_95_22_pad_groupi_n_1250);
  or csa_tree_add_95_22_pad_groupi_g4440(csa_tree_add_95_22_pad_groupi_n_1291 ,csa_tree_add_95_22_pad_groupi_n_1200 ,csa_tree_add_95_22_pad_groupi_n_1249);
  not csa_tree_add_95_22_pad_groupi_g4441(csa_tree_add_95_22_pad_groupi_n_1283 ,csa_tree_add_95_22_pad_groupi_n_1282);
  nor csa_tree_add_95_22_pad_groupi_g4442(csa_tree_add_95_22_pad_groupi_n_1277 ,csa_tree_add_95_22_pad_groupi_n_1132 ,csa_tree_add_95_22_pad_groupi_n_1234);
  and csa_tree_add_95_22_pad_groupi_g4443(csa_tree_add_95_22_pad_groupi_n_1276 ,csa_tree_add_95_22_pad_groupi_n_1132 ,csa_tree_add_95_22_pad_groupi_n_1234);
  xnor csa_tree_add_95_22_pad_groupi_g4444(csa_tree_add_95_22_pad_groupi_n_1275 ,csa_tree_add_95_22_pad_groupi_n_1207 ,csa_tree_add_95_22_pad_groupi_n_1098);
  nor csa_tree_add_95_22_pad_groupi_g4445(csa_tree_add_95_22_pad_groupi_n_1274 ,csa_tree_add_95_22_pad_groupi_n_1157 ,csa_tree_add_95_22_pad_groupi_n_1229);
  xnor csa_tree_add_95_22_pad_groupi_g4446(csa_tree_add_95_22_pad_groupi_n_1273 ,csa_tree_add_95_22_pad_groupi_n_1163 ,csa_tree_add_95_22_pad_groupi_n_1166);
  xnor csa_tree_add_95_22_pad_groupi_g4447(csa_tree_add_95_22_pad_groupi_n_1272 ,csa_tree_add_95_22_pad_groupi_n_1099 ,csa_tree_add_95_22_pad_groupi_n_1169);
  xnor csa_tree_add_95_22_pad_groupi_g4448(csa_tree_add_95_22_pad_groupi_n_1271 ,csa_tree_add_95_22_pad_groupi_n_1204 ,csa_tree_add_95_22_pad_groupi_n_1160);
  xnor csa_tree_add_95_22_pad_groupi_g4449(csa_tree_add_95_22_pad_groupi_n_1270 ,csa_tree_add_95_22_pad_groupi_n_1208 ,csa_tree_add_95_22_pad_groupi_n_1174);
  xnor csa_tree_add_95_22_pad_groupi_g4450(csa_tree_add_95_22_pad_groupi_n_1269 ,csa_tree_add_95_22_pad_groupi_n_1206 ,csa_tree_add_95_22_pad_groupi_n_1171);
  xnor csa_tree_add_95_22_pad_groupi_g4451(csa_tree_add_95_22_pad_groupi_n_1268 ,csa_tree_add_95_22_pad_groupi_n_1164 ,csa_tree_add_95_22_pad_groupi_n_1167);
  xnor csa_tree_add_95_22_pad_groupi_g4452(csa_tree_add_95_22_pad_groupi_n_1267 ,csa_tree_add_95_22_pad_groupi_n_1173 ,csa_tree_add_95_22_pad_groupi_n_1172);
  xnor csa_tree_add_95_22_pad_groupi_g4453(csa_tree_add_95_22_pad_groupi_n_1266 ,csa_tree_add_95_22_pad_groupi_n_1161 ,csa_tree_add_95_22_pad_groupi_n_1168);
  xnor csa_tree_add_95_22_pad_groupi_g4454(csa_tree_add_95_22_pad_groupi_n_1282 ,csa_tree_add_95_22_pad_groupi_n_1106 ,csa_tree_add_95_22_pad_groupi_n_1143);
  xnor csa_tree_add_95_22_pad_groupi_g4455(csa_tree_add_95_22_pad_groupi_n_1281 ,csa_tree_add_95_22_pad_groupi_n_1080 ,csa_tree_add_95_22_pad_groupi_n_1145);
  xnor csa_tree_add_95_22_pad_groupi_g4456(csa_tree_add_95_22_pad_groupi_n_1280 ,csa_tree_add_95_22_pad_groupi_n_1103 ,csa_tree_add_95_22_pad_groupi_n_1146);
  xnor csa_tree_add_95_22_pad_groupi_g4457(csa_tree_add_95_22_pad_groupi_n_1279 ,csa_tree_add_95_22_pad_groupi_n_1101 ,csa_tree_add_95_22_pad_groupi_n_1142);
  xnor csa_tree_add_95_22_pad_groupi_g4458(csa_tree_add_95_22_pad_groupi_n_1278 ,csa_tree_add_95_22_pad_groupi_n_1105 ,csa_tree_add_95_22_pad_groupi_n_1144);
  or csa_tree_add_95_22_pad_groupi_g4459(csa_tree_add_95_22_pad_groupi_n_1260 ,csa_tree_add_95_22_pad_groupi_n_1104 ,csa_tree_add_95_22_pad_groupi_n_1151);
  or csa_tree_add_95_22_pad_groupi_g4460(csa_tree_add_95_22_pad_groupi_n_1259 ,csa_tree_add_95_22_pad_groupi_n_1209 ,csa_tree_add_95_22_pad_groupi_n_1193);
  nor csa_tree_add_95_22_pad_groupi_g4461(csa_tree_add_95_22_pad_groupi_n_1258 ,csa_tree_add_95_22_pad_groupi_n_1074 ,csa_tree_add_95_22_pad_groupi_n_1195);
  or csa_tree_add_95_22_pad_groupi_g4462(csa_tree_add_95_22_pad_groupi_n_1257 ,csa_tree_add_95_22_pad_groupi_n_1072 ,csa_tree_add_95_22_pad_groupi_n_1190);
  nor csa_tree_add_95_22_pad_groupi_g4463(csa_tree_add_95_22_pad_groupi_n_1256 ,csa_tree_add_95_22_pad_groupi_n_1067 ,csa_tree_add_95_22_pad_groupi_n_1186);
  and csa_tree_add_95_22_pad_groupi_g4464(csa_tree_add_95_22_pad_groupi_n_1255 ,csa_tree_add_95_22_pad_groupi_n_1141 ,csa_tree_add_95_22_pad_groupi_n_1189);
  or csa_tree_add_95_22_pad_groupi_g4465(csa_tree_add_95_22_pad_groupi_n_1254 ,csa_tree_add_95_22_pad_groupi_n_1203 ,csa_tree_add_95_22_pad_groupi_n_1159);
  and csa_tree_add_95_22_pad_groupi_g4466(csa_tree_add_95_22_pad_groupi_n_1253 ,csa_tree_add_95_22_pad_groupi_n_1181 ,csa_tree_add_95_22_pad_groupi_n_1176);
  nor csa_tree_add_95_22_pad_groupi_g4467(csa_tree_add_95_22_pad_groupi_n_1252 ,csa_tree_add_95_22_pad_groupi_n_1206 ,csa_tree_add_95_22_pad_groupi_n_1171);
  nor csa_tree_add_95_22_pad_groupi_g4468(csa_tree_add_95_22_pad_groupi_n_1251 ,csa_tree_add_95_22_pad_groupi_n_1177 ,csa_tree_add_95_22_pad_groupi_n_1191);
  and csa_tree_add_95_22_pad_groupi_g4469(csa_tree_add_95_22_pad_groupi_n_1250 ,csa_tree_add_95_22_pad_groupi_n_1102 ,csa_tree_add_95_22_pad_groupi_n_1194);
  and csa_tree_add_95_22_pad_groupi_g4470(csa_tree_add_95_22_pad_groupi_n_1249 ,csa_tree_add_95_22_pad_groupi_n_1107 ,csa_tree_add_95_22_pad_groupi_n_1158);
  nor csa_tree_add_95_22_pad_groupi_g4471(csa_tree_add_95_22_pad_groupi_n_1248 ,csa_tree_add_95_22_pad_groupi_n_1042 ,csa_tree_add_95_22_pad_groupi_n_1153);
  nor csa_tree_add_95_22_pad_groupi_g4472(csa_tree_add_95_22_pad_groupi_n_1247 ,csa_tree_add_95_22_pad_groupi_n_1099 ,csa_tree_add_95_22_pad_groupi_n_1169);
  and csa_tree_add_95_22_pad_groupi_g4473(csa_tree_add_95_22_pad_groupi_n_1246 ,csa_tree_add_95_22_pad_groupi_n_1164 ,csa_tree_add_95_22_pad_groupi_n_1167);
  nor csa_tree_add_95_22_pad_groupi_g4474(csa_tree_add_95_22_pad_groupi_n_1245 ,csa_tree_add_95_22_pad_groupi_n_1164 ,csa_tree_add_95_22_pad_groupi_n_1167);
  nor csa_tree_add_95_22_pad_groupi_g4475(csa_tree_add_95_22_pad_groupi_n_1244 ,csa_tree_add_95_22_pad_groupi_n_1039 ,csa_tree_add_95_22_pad_groupi_n_1148);
  or csa_tree_add_95_22_pad_groupi_g4476(csa_tree_add_95_22_pad_groupi_n_1243 ,csa_tree_add_95_22_pad_groupi_n_1205 ,csa_tree_add_95_22_pad_groupi_n_1170);
  and csa_tree_add_95_22_pad_groupi_g4477(csa_tree_add_95_22_pad_groupi_n_1242 ,csa_tree_add_95_22_pad_groupi_n_1099 ,csa_tree_add_95_22_pad_groupi_n_1169);
  or csa_tree_add_95_22_pad_groupi_g4478(csa_tree_add_95_22_pad_groupi_n_1241 ,csa_tree_add_95_22_pad_groupi_n_1207 ,csa_tree_add_95_22_pad_groupi_n_1098);
  and csa_tree_add_95_22_pad_groupi_g4479(csa_tree_add_95_22_pad_groupi_n_1240 ,csa_tree_add_95_22_pad_groupi_n_1207 ,csa_tree_add_95_22_pad_groupi_n_1098);
  or csa_tree_add_95_22_pad_groupi_g4480(csa_tree_add_95_22_pad_groupi_n_1265 ,csa_tree_add_95_22_pad_groupi_n_1051 ,csa_tree_add_95_22_pad_groupi_n_1180);
  and csa_tree_add_95_22_pad_groupi_g4481(csa_tree_add_95_22_pad_groupi_n_1264 ,csa_tree_add_95_22_pad_groupi_n_1115 ,csa_tree_add_95_22_pad_groupi_n_1199);
  or csa_tree_add_95_22_pad_groupi_g4482(csa_tree_add_95_22_pad_groupi_n_1263 ,csa_tree_add_95_22_pad_groupi_n_1123 ,csa_tree_add_95_22_pad_groupi_n_1182);
  and csa_tree_add_95_22_pad_groupi_g4483(csa_tree_add_95_22_pad_groupi_n_1262 ,csa_tree_add_95_22_pad_groupi_n_1114 ,csa_tree_add_95_22_pad_groupi_n_1149);
  or csa_tree_add_95_22_pad_groupi_g4484(csa_tree_add_95_22_pad_groupi_n_1261 ,csa_tree_add_95_22_pad_groupi_n_1124 ,csa_tree_add_95_22_pad_groupi_n_1196);
  not csa_tree_add_95_22_pad_groupi_g4485(csa_tree_add_95_22_pad_groupi_n_1239 ,csa_tree_add_95_22_pad_groupi_n_1238);
  not csa_tree_add_95_22_pad_groupi_g4486(csa_tree_add_95_22_pad_groupi_n_1237 ,csa_tree_add_95_22_pad_groupi_n_1236);
  not csa_tree_add_95_22_pad_groupi_g4487(csa_tree_add_95_22_pad_groupi_n_1234 ,csa_tree_add_95_22_pad_groupi_n_1233);
  and csa_tree_add_95_22_pad_groupi_g4488(csa_tree_add_95_22_pad_groupi_n_1232 ,csa_tree_add_95_22_pad_groupi_n_1208 ,csa_tree_add_95_22_pad_groupi_n_1174);
  or csa_tree_add_95_22_pad_groupi_g4489(csa_tree_add_95_22_pad_groupi_n_1231 ,csa_tree_add_95_22_pad_groupi_n_1208 ,csa_tree_add_95_22_pad_groupi_n_1174);
  and csa_tree_add_95_22_pad_groupi_g4490(csa_tree_add_95_22_pad_groupi_n_1230 ,csa_tree_add_95_22_pad_groupi_n_1173 ,csa_tree_add_95_22_pad_groupi_n_1172);
  nor csa_tree_add_95_22_pad_groupi_g4491(csa_tree_add_95_22_pad_groupi_n_1229 ,csa_tree_add_95_22_pad_groupi_n_1152 ,csa_tree_add_95_22_pad_groupi_n_1175);
  or csa_tree_add_95_22_pad_groupi_g4492(csa_tree_add_95_22_pad_groupi_n_1228 ,csa_tree_add_95_22_pad_groupi_n_1173 ,csa_tree_add_95_22_pad_groupi_n_1172);
  and csa_tree_add_95_22_pad_groupi_g4493(csa_tree_add_95_22_pad_groupi_n_1227 ,csa_tree_add_95_22_pad_groupi_n_1161 ,csa_tree_add_95_22_pad_groupi_n_1168);
  or csa_tree_add_95_22_pad_groupi_g4494(csa_tree_add_95_22_pad_groupi_n_1226 ,csa_tree_add_95_22_pad_groupi_n_1161 ,csa_tree_add_95_22_pad_groupi_n_1168);
  or csa_tree_add_95_22_pad_groupi_g4495(csa_tree_add_95_22_pad_groupi_n_1225 ,csa_tree_add_95_22_pad_groupi_n_1162 ,csa_tree_add_95_22_pad_groupi_n_1165);
  nor csa_tree_add_95_22_pad_groupi_g4496(csa_tree_add_95_22_pad_groupi_n_1224 ,csa_tree_add_95_22_pad_groupi_n_1204 ,csa_tree_add_95_22_pad_groupi_n_1160);
  nor csa_tree_add_95_22_pad_groupi_g4497(csa_tree_add_95_22_pad_groupi_n_1223 ,csa_tree_add_95_22_pad_groupi_n_1163 ,csa_tree_add_95_22_pad_groupi_n_1166);
  xnor csa_tree_add_95_22_pad_groupi_g4498(csa_tree_add_95_22_pad_groupi_n_1222 ,csa_tree_add_95_22_pad_groupi_n_1035 ,csa_tree_add_95_22_pad_groupi_n_1094);
  xnor csa_tree_add_95_22_pad_groupi_g4499(csa_tree_add_95_22_pad_groupi_n_1221 ,csa_tree_add_95_22_pad_groupi_n_1100 ,csa_tree_add_95_22_pad_groupi_n_1074);
  xnor csa_tree_add_95_22_pad_groupi_g4500(csa_tree_add_95_22_pad_groupi_n_1220 ,csa_tree_add_95_22_pad_groupi_n_1072 ,csa_tree_add_95_22_pad_groupi_n_1090);
  xnor csa_tree_add_95_22_pad_groupi_g4501(csa_tree_add_95_22_pad_groupi_n_1219 ,csa_tree_add_95_22_pad_groupi_n_1016 ,csa_tree_add_95_22_pad_groupi_n_1097);
  xnor csa_tree_add_95_22_pad_groupi_g4502(csa_tree_add_95_22_pad_groupi_n_1218 ,csa_tree_add_95_22_pad_groupi_n_1056 ,csa_tree_add_95_22_pad_groupi_n_3);
  xnor csa_tree_add_95_22_pad_groupi_g4503(csa_tree_add_95_22_pad_groupi_n_1238 ,csa_tree_add_95_22_pad_groupi_n_1140 ,csa_tree_add_95_22_pad_groupi_n_1076);
  xnor csa_tree_add_95_22_pad_groupi_g4504(csa_tree_add_95_22_pad_groupi_n_1217 ,csa_tree_add_95_22_pad_groupi_n_1055 ,csa_tree_add_95_22_pad_groupi_n_1095);
  xnor csa_tree_add_95_22_pad_groupi_g4505(csa_tree_add_95_22_pad_groupi_n_1216 ,csa_tree_add_95_22_pad_groupi_n_1036 ,csa_tree_add_95_22_pad_groupi_n_1087);
  xnor csa_tree_add_95_22_pad_groupi_g4506(csa_tree_add_95_22_pad_groupi_n_1215 ,csa_tree_add_95_22_pad_groupi_n_1137 ,csa_tree_add_95_22_pad_groupi_n_1086);
  xnor csa_tree_add_95_22_pad_groupi_g4507(csa_tree_add_95_22_pad_groupi_n_1214 ,csa_tree_add_95_22_pad_groupi_n_1042 ,csa_tree_add_95_22_pad_groupi_n_1093);
  xnor csa_tree_add_95_22_pad_groupi_g4508(csa_tree_add_95_22_pad_groupi_n_1213 ,csa_tree_add_95_22_pad_groupi_n_1034 ,csa_tree_add_95_22_pad_groupi_n_1104);
  xnor csa_tree_add_95_22_pad_groupi_g4509(csa_tree_add_95_22_pad_groupi_n_1212 ,csa_tree_add_95_22_pad_groupi_n_1131 ,csa_tree_add_95_22_pad_groupi_n_1082);
  xnor csa_tree_add_95_22_pad_groupi_g4510(csa_tree_add_95_22_pad_groupi_n_1211 ,csa_tree_add_95_22_pad_groupi_n_1134 ,csa_tree_add_95_22_pad_groupi_n_1135);
  xnor csa_tree_add_95_22_pad_groupi_g4511(csa_tree_add_95_22_pad_groupi_n_1210 ,csa_tree_add_95_22_pad_groupi_n_1062 ,csa_tree_add_95_22_pad_groupi_n_1133);
  xnor csa_tree_add_95_22_pad_groupi_g4512(csa_tree_add_95_22_pad_groupi_n_1236 ,csa_tree_add_95_22_pad_groupi_n_1043 ,csa_tree_add_95_22_pad_groupi_n_1078);
  xnor csa_tree_add_95_22_pad_groupi_g4513(csa_tree_add_95_22_pad_groupi_n_1235 ,csa_tree_add_95_22_pad_groupi_n_1070 ,csa_tree_add_95_22_pad_groupi_n_1079);
  xnor csa_tree_add_95_22_pad_groupi_g4514(csa_tree_add_95_22_pad_groupi_n_1233 ,csa_tree_add_95_22_pad_groupi_n_976 ,csa_tree_add_95_22_pad_groupi_n_1077);
  not csa_tree_add_95_22_pad_groupi_g4515(csa_tree_add_95_22_pad_groupi_n_1206 ,csa_tree_add_95_22_pad_groupi_n_1205);
  not csa_tree_add_95_22_pad_groupi_g4516(csa_tree_add_95_22_pad_groupi_n_1204 ,csa_tree_add_95_22_pad_groupi_n_1203);
  not csa_tree_add_95_22_pad_groupi_g4517(csa_tree_add_95_22_pad_groupi_n_1202 ,csa_tree_add_95_22_pad_groupi_n_1201);
  and csa_tree_add_95_22_pad_groupi_g4518(csa_tree_add_95_22_pad_groupi_n_1200 ,csa_tree_add_95_22_pad_groupi_n_1035 ,csa_tree_add_95_22_pad_groupi_n_1094);
  or csa_tree_add_95_22_pad_groupi_g4519(csa_tree_add_95_22_pad_groupi_n_1199 ,csa_tree_add_95_22_pad_groupi_n_1105 ,csa_tree_add_95_22_pad_groupi_n_1128);
  nor csa_tree_add_95_22_pad_groupi_g4520(csa_tree_add_95_22_pad_groupi_n_1198 ,csa_tree_add_95_22_pad_groupi_n_1100 ,csa_tree_add_95_22_pad_groupi_n_1139);
  or csa_tree_add_95_22_pad_groupi_g4521(csa_tree_add_95_22_pad_groupi_n_1197 ,csa_tree_add_95_22_pad_groupi_n_1136 ,csa_tree_add_95_22_pad_groupi_n_1086);
  and csa_tree_add_95_22_pad_groupi_g4522(csa_tree_add_95_22_pad_groupi_n_1196 ,csa_tree_add_95_22_pad_groupi_n_1118 ,csa_tree_add_95_22_pad_groupi_n_1103);
  and csa_tree_add_95_22_pad_groupi_g4523(csa_tree_add_95_22_pad_groupi_n_1195 ,csa_tree_add_95_22_pad_groupi_n_1100 ,csa_tree_add_95_22_pad_groupi_n_1139);
  or csa_tree_add_95_22_pad_groupi_g4524(csa_tree_add_95_22_pad_groupi_n_1194 ,csa_tree_add_95_22_pad_groupi_n_1055 ,csa_tree_add_95_22_pad_groupi_n_1095);
  nor csa_tree_add_95_22_pad_groupi_g4525(csa_tree_add_95_22_pad_groupi_n_1193 ,csa_tree_add_95_22_pad_groupi_n_1137 ,csa_tree_add_95_22_pad_groupi_n_1085);
  or csa_tree_add_95_22_pad_groupi_g4526(csa_tree_add_95_22_pad_groupi_n_1192 ,csa_tree_add_95_22_pad_groupi_n_1083 ,csa_tree_add_95_22_pad_groupi_n_1089);
  nor csa_tree_add_95_22_pad_groupi_g4527(csa_tree_add_95_22_pad_groupi_n_1191 ,csa_tree_add_95_22_pad_groupi_n_1022 ,csa_tree_add_95_22_pad_groupi_n_1109);
  nor csa_tree_add_95_22_pad_groupi_g4528(csa_tree_add_95_22_pad_groupi_n_1190 ,csa_tree_add_95_22_pad_groupi_n_1084 ,csa_tree_add_95_22_pad_groupi_n_1090);
  or csa_tree_add_95_22_pad_groupi_g4529(csa_tree_add_95_22_pad_groupi_n_1189 ,csa_tree_add_95_22_pad_groupi_n_1056 ,csa_tree_add_95_22_pad_groupi_n_3);
  nor csa_tree_add_95_22_pad_groupi_g4530(csa_tree_add_95_22_pad_groupi_n_1188 ,csa_tree_add_95_22_pad_groupi_n_1019 ,csa_tree_add_95_22_pad_groupi_n_1080);
  and csa_tree_add_95_22_pad_groupi_g4531(csa_tree_add_95_22_pad_groupi_n_1187 ,csa_tree_add_95_22_pad_groupi_n_1056 ,csa_tree_add_95_22_pad_groupi_n_3);
  and csa_tree_add_95_22_pad_groupi_g4532(csa_tree_add_95_22_pad_groupi_n_1186 ,csa_tree_add_95_22_pad_groupi_n_1019 ,csa_tree_add_95_22_pad_groupi_n_1080);
  and csa_tree_add_95_22_pad_groupi_g4533(csa_tree_add_95_22_pad_groupi_n_1185 ,csa_tree_add_95_22_pad_groupi_n_1134 ,csa_tree_add_95_22_pad_groupi_n_1135);
  nor csa_tree_add_95_22_pad_groupi_g4534(csa_tree_add_95_22_pad_groupi_n_1184 ,csa_tree_add_95_22_pad_groupi_n_1134 ,csa_tree_add_95_22_pad_groupi_n_1135);
  and csa_tree_add_95_22_pad_groupi_g4535(csa_tree_add_95_22_pad_groupi_n_1183 ,csa_tree_add_95_22_pad_groupi_n_1062 ,csa_tree_add_95_22_pad_groupi_n_1133);
  and csa_tree_add_95_22_pad_groupi_g4536(csa_tree_add_95_22_pad_groupi_n_1182 ,csa_tree_add_95_22_pad_groupi_n_1120 ,csa_tree_add_95_22_pad_groupi_n_1106);
  or csa_tree_add_95_22_pad_groupi_g4537(csa_tree_add_95_22_pad_groupi_n_1181 ,csa_tree_add_95_22_pad_groupi_n_1062 ,csa_tree_add_95_22_pad_groupi_n_1133);
  and csa_tree_add_95_22_pad_groupi_g4538(csa_tree_add_95_22_pad_groupi_n_1180 ,csa_tree_add_95_22_pad_groupi_n_1050 ,csa_tree_add_95_22_pad_groupi_n_1140);
  and csa_tree_add_95_22_pad_groupi_g4539(csa_tree_add_95_22_pad_groupi_n_1179 ,csa_tree_add_95_22_pad_groupi_n_1055 ,csa_tree_add_95_22_pad_groupi_n_1095);
  nor csa_tree_add_95_22_pad_groupi_g4540(csa_tree_add_95_22_pad_groupi_n_1178 ,csa_tree_add_95_22_pad_groupi_n_1023 ,csa_tree_add_95_22_pad_groupi_n_1108);
  nor csa_tree_add_95_22_pad_groupi_g4541(csa_tree_add_95_22_pad_groupi_n_1177 ,csa_tree_add_95_22_pad_groupi_n_1031 ,csa_tree_add_95_22_pad_groupi_n_1119);
  and csa_tree_add_95_22_pad_groupi_g4542(csa_tree_add_95_22_pad_groupi_n_1209 ,csa_tree_add_95_22_pad_groupi_n_1054 ,csa_tree_add_95_22_pad_groupi_n_1127);
  or csa_tree_add_95_22_pad_groupi_g4543(csa_tree_add_95_22_pad_groupi_n_1208 ,csa_tree_add_95_22_pad_groupi_n_901 ,csa_tree_add_95_22_pad_groupi_n_1122);
  or csa_tree_add_95_22_pad_groupi_g4544(csa_tree_add_95_22_pad_groupi_n_1207 ,csa_tree_add_95_22_pad_groupi_n_914 ,csa_tree_add_95_22_pad_groupi_n_1125);
  and csa_tree_add_95_22_pad_groupi_g4545(csa_tree_add_95_22_pad_groupi_n_1205 ,csa_tree_add_95_22_pad_groupi_n_884 ,csa_tree_add_95_22_pad_groupi_n_1116);
  and csa_tree_add_95_22_pad_groupi_g4546(csa_tree_add_95_22_pad_groupi_n_1203 ,csa_tree_add_95_22_pad_groupi_n_921 ,csa_tree_add_95_22_pad_groupi_n_1126);
  or csa_tree_add_95_22_pad_groupi_g4547(csa_tree_add_95_22_pad_groupi_n_1201 ,csa_tree_add_95_22_pad_groupi_n_1049 ,csa_tree_add_95_22_pad_groupi_n_1117);
  not csa_tree_add_95_22_pad_groupi_g4548(csa_tree_add_95_22_pad_groupi_n_1170 ,csa_tree_add_95_22_pad_groupi_n_1171);
  not csa_tree_add_95_22_pad_groupi_g4549(csa_tree_add_95_22_pad_groupi_n_1166 ,csa_tree_add_95_22_pad_groupi_n_1165);
  not csa_tree_add_95_22_pad_groupi_g4550(csa_tree_add_95_22_pad_groupi_n_1163 ,csa_tree_add_95_22_pad_groupi_n_1162);
  not csa_tree_add_95_22_pad_groupi_g4551(csa_tree_add_95_22_pad_groupi_n_1160 ,csa_tree_add_95_22_pad_groupi_n_1159);
  or csa_tree_add_95_22_pad_groupi_g4552(csa_tree_add_95_22_pad_groupi_n_1158 ,csa_tree_add_95_22_pad_groupi_n_1035 ,csa_tree_add_95_22_pad_groupi_n_1094);
  and csa_tree_add_95_22_pad_groupi_g4553(csa_tree_add_95_22_pad_groupi_n_1157 ,csa_tree_add_95_22_pad_groupi_n_1015 ,csa_tree_add_95_22_pad_groupi_n_1097);
  or csa_tree_add_95_22_pad_groupi_g4554(csa_tree_add_95_22_pad_groupi_n_1156 ,csa_tree_add_95_22_pad_groupi_n_1130 ,csa_tree_add_95_22_pad_groupi_n_1081);
  or csa_tree_add_95_22_pad_groupi_g4555(csa_tree_add_95_22_pad_groupi_n_1155 ,csa_tree_add_95_22_pad_groupi_n_1033 ,csa_tree_add_95_22_pad_groupi_n_1091);
  and csa_tree_add_95_22_pad_groupi_g4556(csa_tree_add_95_22_pad_groupi_n_1154 ,csa_tree_add_95_22_pad_groupi_n_1093 ,csa_tree_add_95_22_pad_groupi_n_1088);
  nor csa_tree_add_95_22_pad_groupi_g4557(csa_tree_add_95_22_pad_groupi_n_1153 ,csa_tree_add_95_22_pad_groupi_n_1093 ,csa_tree_add_95_22_pad_groupi_n_1088);
  and csa_tree_add_95_22_pad_groupi_g4558(csa_tree_add_95_22_pad_groupi_n_1152 ,csa_tree_add_95_22_pad_groupi_n_1016 ,csa_tree_add_95_22_pad_groupi_n_1096);
  nor csa_tree_add_95_22_pad_groupi_g4559(csa_tree_add_95_22_pad_groupi_n_1151 ,csa_tree_add_95_22_pad_groupi_n_1034 ,csa_tree_add_95_22_pad_groupi_n_1092);
  nor csa_tree_add_95_22_pad_groupi_g4560(csa_tree_add_95_22_pad_groupi_n_1150 ,csa_tree_add_95_22_pad_groupi_n_1131 ,csa_tree_add_95_22_pad_groupi_n_1082);
  or csa_tree_add_95_22_pad_groupi_g4561(csa_tree_add_95_22_pad_groupi_n_1149 ,csa_tree_add_95_22_pad_groupi_n_1110 ,csa_tree_add_95_22_pad_groupi_n_1101);
  and csa_tree_add_95_22_pad_groupi_g4562(csa_tree_add_95_22_pad_groupi_n_1148 ,csa_tree_add_95_22_pad_groupi_n_1037 ,csa_tree_add_95_22_pad_groupi_n_1087);
  nor csa_tree_add_95_22_pad_groupi_g4563(csa_tree_add_95_22_pad_groupi_n_1147 ,csa_tree_add_95_22_pad_groupi_n_1037 ,csa_tree_add_95_22_pad_groupi_n_1087);
  xnor csa_tree_add_95_22_pad_groupi_g4564(csa_tree_add_95_22_pad_groupi_n_1146 ,csa_tree_add_95_22_pad_groupi_n_1010 ,csa_tree_add_95_22_pad_groupi_n_1064);
  xnor csa_tree_add_95_22_pad_groupi_g4565(csa_tree_add_95_22_pad_groupi_n_1145 ,csa_tree_add_95_22_pad_groupi_n_1067 ,csa_tree_add_95_22_pad_groupi_n_1019);
  xnor csa_tree_add_95_22_pad_groupi_g4566(csa_tree_add_95_22_pad_groupi_n_1144 ,csa_tree_add_95_22_pad_groupi_n_1058 ,csa_tree_add_95_22_pad_groupi_n_1061);
  xnor csa_tree_add_95_22_pad_groupi_g4567(csa_tree_add_95_22_pad_groupi_n_1143 ,csa_tree_add_95_22_pad_groupi_n_1011 ,csa_tree_add_95_22_pad_groupi_n_1059);
  xnor csa_tree_add_95_22_pad_groupi_g4568(csa_tree_add_95_22_pad_groupi_n_1142 ,csa_tree_add_95_22_pad_groupi_n_1018 ,csa_tree_add_95_22_pad_groupi_n_1066);
  xnor csa_tree_add_95_22_pad_groupi_g4569(csa_tree_add_95_22_pad_groupi_n_1176 ,csa_tree_add_95_22_pad_groupi_n_1020 ,csa_tree_add_95_22_pad_groupi_n_1025);
  and csa_tree_add_95_22_pad_groupi_g4570(csa_tree_add_95_22_pad_groupi_n_1175 ,csa_tree_add_95_22_pad_groupi_n_1030 ,csa_tree_add_95_22_pad_groupi_n_1111);
  xnor csa_tree_add_95_22_pad_groupi_g4571(csa_tree_add_95_22_pad_groupi_n_1174 ,csa_tree_add_95_22_pad_groupi_n_1068 ,csa_tree_add_95_22_pad_groupi_n_950);
  or csa_tree_add_95_22_pad_groupi_g4572(csa_tree_add_95_22_pad_groupi_n_1173 ,csa_tree_add_95_22_pad_groupi_n_908 ,csa_tree_add_95_22_pad_groupi_n_1121);
  xnor csa_tree_add_95_22_pad_groupi_g4573(csa_tree_add_95_22_pad_groupi_n_1172 ,csa_tree_add_95_22_pad_groupi_n_1045 ,csa_tree_add_95_22_pad_groupi_n_944);
  xnor csa_tree_add_95_22_pad_groupi_g4574(csa_tree_add_95_22_pad_groupi_n_1171 ,csa_tree_add_95_22_pad_groupi_n_1073 ,csa_tree_add_95_22_pad_groupi_n_941);
  xnor csa_tree_add_95_22_pad_groupi_g4575(csa_tree_add_95_22_pad_groupi_n_1169 ,csa_tree_add_95_22_pad_groupi_n_1041 ,csa_tree_add_95_22_pad_groupi_n_974);
  xnor csa_tree_add_95_22_pad_groupi_g4576(csa_tree_add_95_22_pad_groupi_n_1168 ,csa_tree_add_95_22_pad_groupi_n_1044 ,csa_tree_add_95_22_pad_groupi_n_939);
  xnor csa_tree_add_95_22_pad_groupi_g4577(csa_tree_add_95_22_pad_groupi_n_1167 ,csa_tree_add_95_22_pad_groupi_n_1040 ,csa_tree_add_95_22_pad_groupi_n_969);
  xnor csa_tree_add_95_22_pad_groupi_g4578(csa_tree_add_95_22_pad_groupi_n_1165 ,csa_tree_add_95_22_pad_groupi_n_1038 ,csa_tree_add_95_22_pad_groupi_n_970);
  or csa_tree_add_95_22_pad_groupi_g4579(csa_tree_add_95_22_pad_groupi_n_1164 ,csa_tree_add_95_22_pad_groupi_n_858 ,csa_tree_add_95_22_pad_groupi_n_1113);
  and csa_tree_add_95_22_pad_groupi_g4580(csa_tree_add_95_22_pad_groupi_n_1162 ,csa_tree_add_95_22_pad_groupi_n_857 ,csa_tree_add_95_22_pad_groupi_n_1112);
  or csa_tree_add_95_22_pad_groupi_g4581(csa_tree_add_95_22_pad_groupi_n_1161 ,csa_tree_add_95_22_pad_groupi_n_873 ,csa_tree_add_95_22_pad_groupi_n_1129);
  xnor csa_tree_add_95_22_pad_groupi_g4582(csa_tree_add_95_22_pad_groupi_n_1159 ,csa_tree_add_95_22_pad_groupi_n_1046 ,csa_tree_add_95_22_pad_groupi_n_955);
  not csa_tree_add_95_22_pad_groupi_g4583(csa_tree_add_95_22_pad_groupi_n_1139 ,csa_tree_add_95_22_pad_groupi_n_1138);
  not csa_tree_add_95_22_pad_groupi_g4584(csa_tree_add_95_22_pad_groupi_n_1136 ,csa_tree_add_95_22_pad_groupi_n_1137);
  not csa_tree_add_95_22_pad_groupi_g4585(csa_tree_add_95_22_pad_groupi_n_1130 ,csa_tree_add_95_22_pad_groupi_n_1131);
  and csa_tree_add_95_22_pad_groupi_g4586(csa_tree_add_95_22_pad_groupi_n_1129 ,csa_tree_add_95_22_pad_groupi_n_871 ,csa_tree_add_95_22_pad_groupi_n_1040);
  nor csa_tree_add_95_22_pad_groupi_g4587(csa_tree_add_95_22_pad_groupi_n_1128 ,csa_tree_add_95_22_pad_groupi_n_1058 ,csa_tree_add_95_22_pad_groupi_n_1061);
  or csa_tree_add_95_22_pad_groupi_g4588(csa_tree_add_95_22_pad_groupi_n_1127 ,csa_tree_add_95_22_pad_groupi_n_1053 ,csa_tree_add_95_22_pad_groupi_n_1071);
  or csa_tree_add_95_22_pad_groupi_g4589(csa_tree_add_95_22_pad_groupi_n_1126 ,csa_tree_add_95_22_pad_groupi_n_918 ,csa_tree_add_95_22_pad_groupi_n_1069);
  and csa_tree_add_95_22_pad_groupi_g4590(csa_tree_add_95_22_pad_groupi_n_1125 ,csa_tree_add_95_22_pad_groupi_n_932 ,csa_tree_add_95_22_pad_groupi_n_1073);
  nor csa_tree_add_95_22_pad_groupi_g4591(csa_tree_add_95_22_pad_groupi_n_1124 ,csa_tree_add_95_22_pad_groupi_n_1010 ,csa_tree_add_95_22_pad_groupi_n_1063);
  and csa_tree_add_95_22_pad_groupi_g4592(csa_tree_add_95_22_pad_groupi_n_1123 ,csa_tree_add_95_22_pad_groupi_n_1011 ,csa_tree_add_95_22_pad_groupi_n_1059);
  and csa_tree_add_95_22_pad_groupi_g4593(csa_tree_add_95_22_pad_groupi_n_1122 ,csa_tree_add_95_22_pad_groupi_n_880 ,csa_tree_add_95_22_pad_groupi_n_1045);
  and csa_tree_add_95_22_pad_groupi_g4594(csa_tree_add_95_22_pad_groupi_n_1121 ,csa_tree_add_95_22_pad_groupi_n_867 ,csa_tree_add_95_22_pad_groupi_n_1044);
  or csa_tree_add_95_22_pad_groupi_g4595(csa_tree_add_95_22_pad_groupi_n_1120 ,csa_tree_add_95_22_pad_groupi_n_1011 ,csa_tree_add_95_22_pad_groupi_n_1059);
  nor csa_tree_add_95_22_pad_groupi_g4596(csa_tree_add_95_22_pad_groupi_n_1119 ,csa_tree_add_95_22_pad_groupi_n_1026 ,csa_tree_add_95_22_pad_groupi_n_980);
  or csa_tree_add_95_22_pad_groupi_g4597(csa_tree_add_95_22_pad_groupi_n_1118 ,csa_tree_add_95_22_pad_groupi_n_1009 ,csa_tree_add_95_22_pad_groupi_n_1064);
  and csa_tree_add_95_22_pad_groupi_g4598(csa_tree_add_95_22_pad_groupi_n_1117 ,csa_tree_add_95_22_pad_groupi_n_1029 ,csa_tree_add_95_22_pad_groupi_n_1043);
  or csa_tree_add_95_22_pad_groupi_g4599(csa_tree_add_95_22_pad_groupi_n_1116 ,csa_tree_add_95_22_pad_groupi_n_882 ,csa_tree_add_95_22_pad_groupi_n_1038);
  or csa_tree_add_95_22_pad_groupi_g4600(csa_tree_add_95_22_pad_groupi_n_1115 ,csa_tree_add_95_22_pad_groupi_n_1057 ,csa_tree_add_95_22_pad_groupi_n_1060);
  or csa_tree_add_95_22_pad_groupi_g4601(csa_tree_add_95_22_pad_groupi_n_1114 ,csa_tree_add_95_22_pad_groupi_n_1017 ,csa_tree_add_95_22_pad_groupi_n_1065);
  and csa_tree_add_95_22_pad_groupi_g4602(csa_tree_add_95_22_pad_groupi_n_1113 ,csa_tree_add_95_22_pad_groupi_n_860 ,csa_tree_add_95_22_pad_groupi_n_1041);
  or csa_tree_add_95_22_pad_groupi_g4603(csa_tree_add_95_22_pad_groupi_n_1112 ,csa_tree_add_95_22_pad_groupi_n_854 ,csa_tree_add_95_22_pad_groupi_n_1046);
  or csa_tree_add_95_22_pad_groupi_g4604(csa_tree_add_95_22_pad_groupi_n_1111 ,csa_tree_add_95_22_pad_groupi_n_1028 ,csa_tree_add_95_22_pad_groupi_n_976);
  nor csa_tree_add_95_22_pad_groupi_g4605(csa_tree_add_95_22_pad_groupi_n_1110 ,csa_tree_add_95_22_pad_groupi_n_1018 ,csa_tree_add_95_22_pad_groupi_n_1066);
  xnor csa_tree_add_95_22_pad_groupi_g4606(csa_tree_add_95_22_pad_groupi_n_1141 ,csa_tree_add_95_22_pad_groupi_n_842 ,csa_tree_add_95_22_pad_groupi_n_951);
  xnor csa_tree_add_95_22_pad_groupi_g4607(csa_tree_add_95_22_pad_groupi_n_1140 ,csa_tree_add_95_22_pad_groupi_n_803 ,csa_tree_add_95_22_pad_groupi_n_964);
  xnor csa_tree_add_95_22_pad_groupi_g4608(csa_tree_add_95_22_pad_groupi_n_1138 ,csa_tree_add_95_22_pad_groupi_n_773 ,csa_tree_add_95_22_pad_groupi_n_962);
  xnor csa_tree_add_95_22_pad_groupi_g4609(csa_tree_add_95_22_pad_groupi_n_1137 ,csa_tree_add_95_22_pad_groupi_n_783 ,csa_tree_add_95_22_pad_groupi_n_960);
  xnor csa_tree_add_95_22_pad_groupi_g4610(csa_tree_add_95_22_pad_groupi_n_1135 ,csa_tree_add_95_22_pad_groupi_n_840 ,csa_tree_add_95_22_pad_groupi_n_965);
  or csa_tree_add_95_22_pad_groupi_g4611(csa_tree_add_95_22_pad_groupi_n_1134 ,csa_tree_add_95_22_pad_groupi_n_1000 ,csa_tree_add_95_22_pad_groupi_n_1052);
  xnor csa_tree_add_95_22_pad_groupi_g4612(csa_tree_add_95_22_pad_groupi_n_1133 ,csa_tree_add_95_22_pad_groupi_n_778 ,csa_tree_add_95_22_pad_groupi_n_949);
  and csa_tree_add_95_22_pad_groupi_g4613(csa_tree_add_95_22_pad_groupi_n_1132 ,csa_tree_add_95_22_pad_groupi_n_888 ,csa_tree_add_95_22_pad_groupi_n_1032);
  or csa_tree_add_95_22_pad_groupi_g4614(csa_tree_add_95_22_pad_groupi_n_1131 ,csa_tree_add_95_22_pad_groupi_n_868 ,csa_tree_add_95_22_pad_groupi_n_1027);
  not csa_tree_add_95_22_pad_groupi_g4615(csa_tree_add_95_22_pad_groupi_n_1109 ,csa_tree_add_95_22_pad_groupi_n_1108);
  not csa_tree_add_95_22_pad_groupi_g4616(csa_tree_add_95_22_pad_groupi_n_1097 ,csa_tree_add_95_22_pad_groupi_n_1096);
  not csa_tree_add_95_22_pad_groupi_g4617(csa_tree_add_95_22_pad_groupi_n_1091 ,csa_tree_add_95_22_pad_groupi_n_1092);
  not csa_tree_add_95_22_pad_groupi_g4618(csa_tree_add_95_22_pad_groupi_n_1090 ,csa_tree_add_95_22_pad_groupi_n_1089);
  not csa_tree_add_95_22_pad_groupi_g4619(csa_tree_add_95_22_pad_groupi_n_1085 ,csa_tree_add_95_22_pad_groupi_n_1086);
  not csa_tree_add_95_22_pad_groupi_g4620(csa_tree_add_95_22_pad_groupi_n_1083 ,csa_tree_add_95_22_pad_groupi_n_1084);
  not csa_tree_add_95_22_pad_groupi_g4621(csa_tree_add_95_22_pad_groupi_n_1081 ,csa_tree_add_95_22_pad_groupi_n_1082);
  xnor csa_tree_add_95_22_pad_groupi_g4622(csa_tree_add_95_22_pad_groupi_n_1079 ,csa_tree_add_95_22_pad_groupi_n_975 ,csa_tree_add_95_22_pad_groupi_n_934);
  xnor csa_tree_add_95_22_pad_groupi_g4623(csa_tree_add_95_22_pad_groupi_n_1108 ,csa_tree_add_95_22_pad_groupi_n_892 ,csa_tree_add_95_22_pad_groupi_n_961);
  xnor csa_tree_add_95_22_pad_groupi_g4624(csa_tree_add_95_22_pad_groupi_n_1078 ,csa_tree_add_95_22_pad_groupi_n_797 ,csa_tree_add_95_22_pad_groupi_n_4);
  xnor csa_tree_add_95_22_pad_groupi_g4625(csa_tree_add_95_22_pad_groupi_n_1077 ,csa_tree_add_95_22_pad_groupi_n_746 ,csa_tree_add_95_22_pad_groupi_n_1014);
  xnor csa_tree_add_95_22_pad_groupi_g4626(csa_tree_add_95_22_pad_groupi_n_1076 ,csa_tree_add_95_22_pad_groupi_n_1012 ,csa_tree_add_95_22_pad_groupi_n_933);
  xnor csa_tree_add_95_22_pad_groupi_g4628(csa_tree_add_95_22_pad_groupi_n_1107 ,csa_tree_add_95_22_pad_groupi_n_768 ,csa_tree_add_95_22_pad_groupi_n_942);
  xnor csa_tree_add_95_22_pad_groupi_g4629(csa_tree_add_95_22_pad_groupi_n_1106 ,csa_tree_add_95_22_pad_groupi_n_764 ,csa_tree_add_95_22_pad_groupi_n_968);
  xnor csa_tree_add_95_22_pad_groupi_g4630(csa_tree_add_95_22_pad_groupi_n_1105 ,csa_tree_add_95_22_pad_groupi_n_740 ,csa_tree_add_95_22_pad_groupi_n_963);
  xnor csa_tree_add_95_22_pad_groupi_g4631(csa_tree_add_95_22_pad_groupi_n_1104 ,csa_tree_add_95_22_pad_groupi_n_782 ,csa_tree_add_95_22_pad_groupi_n_967);
  xnor csa_tree_add_95_22_pad_groupi_g4632(csa_tree_add_95_22_pad_groupi_n_1103 ,csa_tree_add_95_22_pad_groupi_n_1021 ,csa_tree_add_95_22_pad_groupi_n_957);
  xnor csa_tree_add_95_22_pad_groupi_g4633(csa_tree_add_95_22_pad_groupi_n_1102 ,csa_tree_add_95_22_pad_groupi_n_769 ,csa_tree_add_95_22_pad_groupi_n_945);
  xnor csa_tree_add_95_22_pad_groupi_g4634(csa_tree_add_95_22_pad_groupi_n_1101 ,csa_tree_add_95_22_pad_groupi_n_977 ,csa_tree_add_95_22_pad_groupi_n_966);
  xnor csa_tree_add_95_22_pad_groupi_g4635(csa_tree_add_95_22_pad_groupi_n_1100 ,csa_tree_add_95_22_pad_groupi_n_838 ,csa_tree_add_95_22_pad_groupi_n_946);
  xnor csa_tree_add_95_22_pad_groupi_g4637(csa_tree_add_95_22_pad_groupi_n_1099 ,csa_tree_add_95_22_pad_groupi_n_750 ,csa_tree_add_95_22_pad_groupi_n_952);
  xnor csa_tree_add_95_22_pad_groupi_g4638(csa_tree_add_95_22_pad_groupi_n_1098 ,csa_tree_add_95_22_pad_groupi_n_743 ,csa_tree_add_95_22_pad_groupi_n_972);
  xnor csa_tree_add_95_22_pad_groupi_g4639(csa_tree_add_95_22_pad_groupi_n_1096 ,csa_tree_add_95_22_pad_groupi_n_971 ,csa_tree_add_95_22_pad_groupi_n_578);
  xnor csa_tree_add_95_22_pad_groupi_g4640(csa_tree_add_95_22_pad_groupi_n_1095 ,csa_tree_add_95_22_pad_groupi_n_770 ,csa_tree_add_95_22_pad_groupi_n_947);
  xnor csa_tree_add_95_22_pad_groupi_g4641(csa_tree_add_95_22_pad_groupi_n_1094 ,csa_tree_add_95_22_pad_groupi_n_830 ,csa_tree_add_95_22_pad_groupi_n_943);
  xnor csa_tree_add_95_22_pad_groupi_g4642(csa_tree_add_95_22_pad_groupi_n_1093 ,csa_tree_add_95_22_pad_groupi_n_780 ,csa_tree_add_95_22_pad_groupi_n_938);
  xnor csa_tree_add_95_22_pad_groupi_g4643(csa_tree_add_95_22_pad_groupi_n_1092 ,csa_tree_add_95_22_pad_groupi_n_775 ,csa_tree_add_95_22_pad_groupi_n_937);
  xnor csa_tree_add_95_22_pad_groupi_g4644(csa_tree_add_95_22_pad_groupi_n_1089 ,csa_tree_add_95_22_pad_groupi_n_827 ,csa_tree_add_95_22_pad_groupi_n_973);
  xnor csa_tree_add_95_22_pad_groupi_g4645(csa_tree_add_95_22_pad_groupi_n_1088 ,csa_tree_add_95_22_pad_groupi_n_777 ,csa_tree_add_95_22_pad_groupi_n_940);
  xnor csa_tree_add_95_22_pad_groupi_g4646(csa_tree_add_95_22_pad_groupi_n_1087 ,csa_tree_add_95_22_pad_groupi_n_774 ,csa_tree_add_95_22_pad_groupi_n_954);
  xnor csa_tree_add_95_22_pad_groupi_g4647(csa_tree_add_95_22_pad_groupi_n_1086 ,csa_tree_add_95_22_pad_groupi_n_893 ,csa_tree_add_95_22_pad_groupi_n_959);
  xnor csa_tree_add_95_22_pad_groupi_g4648(csa_tree_add_95_22_pad_groupi_n_1084 ,csa_tree_add_95_22_pad_groupi_n_785 ,csa_tree_add_95_22_pad_groupi_n_956);
  xnor csa_tree_add_95_22_pad_groupi_g4649(csa_tree_add_95_22_pad_groupi_n_1082 ,csa_tree_add_95_22_pad_groupi_n_839 ,csa_tree_add_95_22_pad_groupi_n_958);
  xnor csa_tree_add_95_22_pad_groupi_g4650(csa_tree_add_95_22_pad_groupi_n_1080 ,csa_tree_add_95_22_pad_groupi_n_936 ,csa_tree_add_95_22_pad_groupi_n_953);
  not csa_tree_add_95_22_pad_groupi_g4651(csa_tree_add_95_22_pad_groupi_n_1071 ,csa_tree_add_95_22_pad_groupi_n_1070);
  not csa_tree_add_95_22_pad_groupi_g4652(csa_tree_add_95_22_pad_groupi_n_1069 ,csa_tree_add_95_22_pad_groupi_n_1068);
  not csa_tree_add_95_22_pad_groupi_g4653(csa_tree_add_95_22_pad_groupi_n_1065 ,csa_tree_add_95_22_pad_groupi_n_1066);
  not csa_tree_add_95_22_pad_groupi_g4654(csa_tree_add_95_22_pad_groupi_n_1063 ,csa_tree_add_95_22_pad_groupi_n_1064);
  not csa_tree_add_95_22_pad_groupi_g4655(csa_tree_add_95_22_pad_groupi_n_1060 ,csa_tree_add_95_22_pad_groupi_n_1061);
  not csa_tree_add_95_22_pad_groupi_g4656(csa_tree_add_95_22_pad_groupi_n_1057 ,csa_tree_add_95_22_pad_groupi_n_1058);
  or csa_tree_add_95_22_pad_groupi_g4657(csa_tree_add_95_22_pad_groupi_n_1054 ,csa_tree_add_95_22_pad_groupi_n_276 ,csa_tree_add_95_22_pad_groupi_n_975);
  and csa_tree_add_95_22_pad_groupi_g4658(csa_tree_add_95_22_pad_groupi_n_1053 ,csa_tree_add_95_22_pad_groupi_n_934 ,csa_tree_add_95_22_pad_groupi_n_975);
  and csa_tree_add_95_22_pad_groupi_g4659(csa_tree_add_95_22_pad_groupi_n_1052 ,csa_tree_add_95_22_pad_groupi_n_998 ,csa_tree_add_95_22_pad_groupi_n_1020);
  and csa_tree_add_95_22_pad_groupi_g4660(csa_tree_add_95_22_pad_groupi_n_1051 ,csa_tree_add_95_22_pad_groupi_n_933 ,csa_tree_add_95_22_pad_groupi_n_1012);
  or csa_tree_add_95_22_pad_groupi_g4661(csa_tree_add_95_22_pad_groupi_n_1050 ,csa_tree_add_95_22_pad_groupi_n_933 ,csa_tree_add_95_22_pad_groupi_n_1012);
  and csa_tree_add_95_22_pad_groupi_g4662(csa_tree_add_95_22_pad_groupi_n_1049 ,csa_tree_add_95_22_pad_groupi_n_797 ,csa_tree_add_95_22_pad_groupi_n_4);
  and csa_tree_add_95_22_pad_groupi_g4663(csa_tree_add_95_22_pad_groupi_n_1074 ,csa_tree_add_95_22_pad_groupi_n_913 ,csa_tree_add_95_22_pad_groupi_n_1007);
  or csa_tree_add_95_22_pad_groupi_g4664(csa_tree_add_95_22_pad_groupi_n_1073 ,csa_tree_add_95_22_pad_groupi_n_910 ,csa_tree_add_95_22_pad_groupi_n_999);
  and csa_tree_add_95_22_pad_groupi_g4665(csa_tree_add_95_22_pad_groupi_n_1072 ,csa_tree_add_95_22_pad_groupi_n_915 ,csa_tree_add_95_22_pad_groupi_n_996);
  or csa_tree_add_95_22_pad_groupi_g4666(csa_tree_add_95_22_pad_groupi_n_1070 ,csa_tree_add_95_22_pad_groupi_n_890 ,csa_tree_add_95_22_pad_groupi_n_1005);
  or csa_tree_add_95_22_pad_groupi_g4667(csa_tree_add_95_22_pad_groupi_n_1068 ,csa_tree_add_95_22_pad_groupi_n_905 ,csa_tree_add_95_22_pad_groupi_n_1003);
  and csa_tree_add_95_22_pad_groupi_g4668(csa_tree_add_95_22_pad_groupi_n_1067 ,csa_tree_add_95_22_pad_groupi_n_912 ,csa_tree_add_95_22_pad_groupi_n_1002);
  or csa_tree_add_95_22_pad_groupi_g4669(csa_tree_add_95_22_pad_groupi_n_1066 ,csa_tree_add_95_22_pad_groupi_n_903 ,csa_tree_add_95_22_pad_groupi_n_1004);
  or csa_tree_add_95_22_pad_groupi_g4670(csa_tree_add_95_22_pad_groupi_n_1064 ,csa_tree_add_95_22_pad_groupi_n_925 ,csa_tree_add_95_22_pad_groupi_n_1006);
  or csa_tree_add_95_22_pad_groupi_g4671(csa_tree_add_95_22_pad_groupi_n_1062 ,csa_tree_add_95_22_pad_groupi_n_874 ,csa_tree_add_95_22_pad_groupi_n_987);
  or csa_tree_add_95_22_pad_groupi_g4672(csa_tree_add_95_22_pad_groupi_n_1061 ,csa_tree_add_95_22_pad_groupi_n_929 ,csa_tree_add_95_22_pad_groupi_n_979);
  or csa_tree_add_95_22_pad_groupi_g4673(csa_tree_add_95_22_pad_groupi_n_1059 ,csa_tree_add_95_22_pad_groupi_n_889 ,csa_tree_add_95_22_pad_groupi_n_995);
  or csa_tree_add_95_22_pad_groupi_g4674(csa_tree_add_95_22_pad_groupi_n_1058 ,csa_tree_add_95_22_pad_groupi_n_911 ,csa_tree_add_95_22_pad_groupi_n_1008);
  or csa_tree_add_95_22_pad_groupi_g4675(csa_tree_add_95_22_pad_groupi_n_1056 ,csa_tree_add_95_22_pad_groupi_n_869 ,csa_tree_add_95_22_pad_groupi_n_1001);
  or csa_tree_add_95_22_pad_groupi_g4676(csa_tree_add_95_22_pad_groupi_n_1055 ,csa_tree_add_95_22_pad_groupi_n_886 ,csa_tree_add_95_22_pad_groupi_n_993);
  not csa_tree_add_95_22_pad_groupi_g4677(csa_tree_add_95_22_pad_groupi_n_1048 ,csa_tree_add_95_22_pad_groupi_n_1047);
  not csa_tree_add_95_22_pad_groupi_g4678(csa_tree_add_95_22_pad_groupi_n_1037 ,csa_tree_add_95_22_pad_groupi_n_1036);
  not csa_tree_add_95_22_pad_groupi_g4679(csa_tree_add_95_22_pad_groupi_n_1033 ,csa_tree_add_95_22_pad_groupi_n_1034);
  or csa_tree_add_95_22_pad_groupi_g4680(csa_tree_add_95_22_pad_groupi_n_1032 ,csa_tree_add_95_22_pad_groupi_n_876 ,csa_tree_add_95_22_pad_groupi_n_977);
  nor csa_tree_add_95_22_pad_groupi_g4681(csa_tree_add_95_22_pad_groupi_n_1031 ,csa_tree_add_95_22_pad_groupi_n_646 ,csa_tree_add_95_22_pad_groupi_n_1024);
  or csa_tree_add_95_22_pad_groupi_g4682(csa_tree_add_95_22_pad_groupi_n_1030 ,csa_tree_add_95_22_pad_groupi_n_745 ,csa_tree_add_95_22_pad_groupi_n_1014);
  or csa_tree_add_95_22_pad_groupi_g4683(csa_tree_add_95_22_pad_groupi_n_1029 ,csa_tree_add_95_22_pad_groupi_n_797 ,csa_tree_add_95_22_pad_groupi_n_4);
  nor csa_tree_add_95_22_pad_groupi_g4684(csa_tree_add_95_22_pad_groupi_n_1028 ,csa_tree_add_95_22_pad_groupi_n_746 ,csa_tree_add_95_22_pad_groupi_n_1013);
  and csa_tree_add_95_22_pad_groupi_g4685(csa_tree_add_95_22_pad_groupi_n_1027 ,csa_tree_add_95_22_pad_groupi_n_865 ,csa_tree_add_95_22_pad_groupi_n_1021);
  and csa_tree_add_95_22_pad_groupi_g4686(csa_tree_add_95_22_pad_groupi_n_1026 ,csa_tree_add_95_22_pad_groupi_n_646 ,csa_tree_add_95_22_pad_groupi_n_1024);
  and csa_tree_add_95_22_pad_groupi_g4687(csa_tree_add_95_22_pad_groupi_n_1047 ,csa_tree_add_95_22_pad_groupi_n_895 ,csa_tree_add_95_22_pad_groupi_n_994);
  xnor csa_tree_add_95_22_pad_groupi_g4688(csa_tree_add_95_22_pad_groupi_n_1025 ,csa_tree_add_95_22_pad_groupi_n_935 ,csa_tree_add_95_22_pad_groupi_n_820);
  and csa_tree_add_95_22_pad_groupi_g4689(csa_tree_add_95_22_pad_groupi_n_1046 ,csa_tree_add_95_22_pad_groupi_n_853 ,csa_tree_add_95_22_pad_groupi_n_982);
  or csa_tree_add_95_22_pad_groupi_g4690(csa_tree_add_95_22_pad_groupi_n_1045 ,csa_tree_add_95_22_pad_groupi_n_906 ,csa_tree_add_95_22_pad_groupi_n_997);
  or csa_tree_add_95_22_pad_groupi_g4691(csa_tree_add_95_22_pad_groupi_n_1044 ,csa_tree_add_95_22_pad_groupi_n_887 ,csa_tree_add_95_22_pad_groupi_n_992);
  or csa_tree_add_95_22_pad_groupi_g4692(csa_tree_add_95_22_pad_groupi_n_1043 ,csa_tree_add_95_22_pad_groupi_n_926 ,csa_tree_add_95_22_pad_groupi_n_991);
  and csa_tree_add_95_22_pad_groupi_g4693(csa_tree_add_95_22_pad_groupi_n_1042 ,csa_tree_add_95_22_pad_groupi_n_864 ,csa_tree_add_95_22_pad_groupi_n_985);
  or csa_tree_add_95_22_pad_groupi_g4694(csa_tree_add_95_22_pad_groupi_n_1041 ,csa_tree_add_95_22_pad_groupi_n_879 ,csa_tree_add_95_22_pad_groupi_n_984);
  or csa_tree_add_95_22_pad_groupi_g4695(csa_tree_add_95_22_pad_groupi_n_1040 ,csa_tree_add_95_22_pad_groupi_n_870 ,csa_tree_add_95_22_pad_groupi_n_988);
  and csa_tree_add_95_22_pad_groupi_g4696(csa_tree_add_95_22_pad_groupi_n_1039 ,csa_tree_add_95_22_pad_groupi_n_852 ,csa_tree_add_95_22_pad_groupi_n_981);
  and csa_tree_add_95_22_pad_groupi_g4697(csa_tree_add_95_22_pad_groupi_n_1038 ,csa_tree_add_95_22_pad_groupi_n_878 ,csa_tree_add_95_22_pad_groupi_n_989);
  or csa_tree_add_95_22_pad_groupi_g4698(csa_tree_add_95_22_pad_groupi_n_1036 ,csa_tree_add_95_22_pad_groupi_n_897 ,csa_tree_add_95_22_pad_groupi_n_983);
  or csa_tree_add_95_22_pad_groupi_g4699(csa_tree_add_95_22_pad_groupi_n_1035 ,csa_tree_add_95_22_pad_groupi_n_907 ,csa_tree_add_95_22_pad_groupi_n_990);
  or csa_tree_add_95_22_pad_groupi_g4700(csa_tree_add_95_22_pad_groupi_n_1034 ,csa_tree_add_95_22_pad_groupi_n_866 ,csa_tree_add_95_22_pad_groupi_n_986);
  not csa_tree_add_95_22_pad_groupi_g4701(csa_tree_add_95_22_pad_groupi_n_1023 ,csa_tree_add_95_22_pad_groupi_n_1022);
  not csa_tree_add_95_22_pad_groupi_g4702(csa_tree_add_95_22_pad_groupi_n_1018 ,csa_tree_add_95_22_pad_groupi_n_1017);
  not csa_tree_add_95_22_pad_groupi_g4703(csa_tree_add_95_22_pad_groupi_n_1016 ,csa_tree_add_95_22_pad_groupi_n_1015);
  not csa_tree_add_95_22_pad_groupi_g4704(csa_tree_add_95_22_pad_groupi_n_1014 ,csa_tree_add_95_22_pad_groupi_n_1013);
  not csa_tree_add_95_22_pad_groupi_g4705(csa_tree_add_95_22_pad_groupi_n_1010 ,csa_tree_add_95_22_pad_groupi_n_1009);
  nor csa_tree_add_95_22_pad_groupi_g4706(csa_tree_add_95_22_pad_groupi_n_1008 ,csa_tree_add_95_22_pad_groupi_n_841 ,csa_tree_add_95_22_pad_groupi_n_930);
  or csa_tree_add_95_22_pad_groupi_g4707(csa_tree_add_95_22_pad_groupi_n_1007 ,csa_tree_add_95_22_pad_groupi_n_843 ,csa_tree_add_95_22_pad_groupi_n_917);
  nor csa_tree_add_95_22_pad_groupi_g4708(csa_tree_add_95_22_pad_groupi_n_1006 ,csa_tree_add_95_22_pad_groupi_n_824 ,csa_tree_add_95_22_pad_groupi_n_872);
  and csa_tree_add_95_22_pad_groupi_g4709(csa_tree_add_95_22_pad_groupi_n_1005 ,csa_tree_add_95_22_pad_groupi_n_840 ,csa_tree_add_95_22_pad_groupi_n_922);
  and csa_tree_add_95_22_pad_groupi_g4710(csa_tree_add_95_22_pad_groupi_n_1004 ,csa_tree_add_95_22_pad_groupi_n_839 ,csa_tree_add_95_22_pad_groupi_n_909);
  and csa_tree_add_95_22_pad_groupi_g4711(csa_tree_add_95_22_pad_groupi_n_1003 ,csa_tree_add_95_22_pad_groupi_n_770 ,csa_tree_add_95_22_pad_groupi_n_916);
  or csa_tree_add_95_22_pad_groupi_g4712(csa_tree_add_95_22_pad_groupi_n_1002 ,csa_tree_add_95_22_pad_groupi_n_779 ,csa_tree_add_95_22_pad_groupi_n_902);
  and csa_tree_add_95_22_pad_groupi_g4713(csa_tree_add_95_22_pad_groupi_n_1001 ,csa_tree_add_95_22_pad_groupi_n_769 ,csa_tree_add_95_22_pad_groupi_n_904);
  and csa_tree_add_95_22_pad_groupi_g4714(csa_tree_add_95_22_pad_groupi_n_1000 ,csa_tree_add_95_22_pad_groupi_n_820 ,csa_tree_add_95_22_pad_groupi_n_935);
  nor csa_tree_add_95_22_pad_groupi_g4715(csa_tree_add_95_22_pad_groupi_n_999 ,csa_tree_add_95_22_pad_groupi_n_834 ,csa_tree_add_95_22_pad_groupi_n_896);
  or csa_tree_add_95_22_pad_groupi_g4716(csa_tree_add_95_22_pad_groupi_n_998 ,csa_tree_add_95_22_pad_groupi_n_820 ,csa_tree_add_95_22_pad_groupi_n_935);
  and csa_tree_add_95_22_pad_groupi_g4717(csa_tree_add_95_22_pad_groupi_n_997 ,csa_tree_add_95_22_pad_groupi_n_830 ,csa_tree_add_95_22_pad_groupi_n_856);
  or csa_tree_add_95_22_pad_groupi_g4718(csa_tree_add_95_22_pad_groupi_n_996 ,csa_tree_add_95_22_pad_groupi_n_936 ,csa_tree_add_95_22_pad_groupi_n_919);
  and csa_tree_add_95_22_pad_groupi_g4719(csa_tree_add_95_22_pad_groupi_n_995 ,csa_tree_add_95_22_pad_groupi_n_775 ,csa_tree_add_95_22_pad_groupi_n_891);
  or csa_tree_add_95_22_pad_groupi_g4720(csa_tree_add_95_22_pad_groupi_n_994 ,csa_tree_add_95_22_pad_groupi_n_892 ,csa_tree_add_95_22_pad_groupi_n_894);
  and csa_tree_add_95_22_pad_groupi_g4721(csa_tree_add_95_22_pad_groupi_n_993 ,csa_tree_add_95_22_pad_groupi_n_768 ,csa_tree_add_95_22_pad_groupi_n_924);
  and csa_tree_add_95_22_pad_groupi_g4722(csa_tree_add_95_22_pad_groupi_n_992 ,csa_tree_add_95_22_pad_groupi_n_780 ,csa_tree_add_95_22_pad_groupi_n_885);
  nor csa_tree_add_95_22_pad_groupi_g4723(csa_tree_add_95_22_pad_groupi_n_991 ,csa_tree_add_95_22_pad_groupi_n_837 ,csa_tree_add_95_22_pad_groupi_n_877);
  and csa_tree_add_95_22_pad_groupi_g4724(csa_tree_add_95_22_pad_groupi_n_990 ,csa_tree_add_95_22_pad_groupi_n_777 ,csa_tree_add_95_22_pad_groupi_n_928);
  or csa_tree_add_95_22_pad_groupi_g4725(csa_tree_add_95_22_pad_groupi_n_989 ,csa_tree_add_95_22_pad_groupi_n_838 ,csa_tree_add_95_22_pad_groupi_n_875);
  nor csa_tree_add_95_22_pad_groupi_g4726(csa_tree_add_95_22_pad_groupi_n_988 ,csa_tree_add_95_22_pad_groupi_n_774 ,csa_tree_add_95_22_pad_groupi_n_855);
  nor csa_tree_add_95_22_pad_groupi_g4727(csa_tree_add_95_22_pad_groupi_n_987 ,csa_tree_add_95_22_pad_groupi_n_776 ,csa_tree_add_95_22_pad_groupi_n_883);
  and csa_tree_add_95_22_pad_groupi_g4728(csa_tree_add_95_22_pad_groupi_n_986 ,csa_tree_add_95_22_pad_groupi_n_773 ,csa_tree_add_95_22_pad_groupi_n_863);
  or csa_tree_add_95_22_pad_groupi_g4729(csa_tree_add_95_22_pad_groupi_n_985 ,csa_tree_add_95_22_pad_groupi_n_823 ,csa_tree_add_95_22_pad_groupi_n_862);
  nor csa_tree_add_95_22_pad_groupi_g4730(csa_tree_add_95_22_pad_groupi_n_984 ,csa_tree_add_95_22_pad_groupi_n_772 ,csa_tree_add_95_22_pad_groupi_n_859);
  nor csa_tree_add_95_22_pad_groupi_g4731(csa_tree_add_95_22_pad_groupi_n_983 ,csa_tree_add_95_22_pad_groupi_n_771 ,csa_tree_add_95_22_pad_groupi_n_900);
  or csa_tree_add_95_22_pad_groupi_g4732(csa_tree_add_95_22_pad_groupi_n_982 ,csa_tree_add_95_22_pad_groupi_n_835 ,csa_tree_add_95_22_pad_groupi_n_851);
  or csa_tree_add_95_22_pad_groupi_g4733(csa_tree_add_95_22_pad_groupi_n_981 ,csa_tree_add_95_22_pad_groupi_n_893 ,csa_tree_add_95_22_pad_groupi_n_920);
  xnor csa_tree_add_95_22_pad_groupi_g4734(csa_tree_add_95_22_pad_groupi_n_980 ,csa_tree_add_95_22_pad_groupi_n_846 ,csa_tree_add_95_22_pad_groupi_n_848);
  and csa_tree_add_95_22_pad_groupi_g4735(csa_tree_add_95_22_pad_groupi_n_979 ,csa_tree_add_95_22_pad_groupi_n_827 ,csa_tree_add_95_22_pad_groupi_n_927);
  or csa_tree_add_95_22_pad_groupi_g4736(csa_tree_add_95_22_pad_groupi_n_1024 ,csa_tree_add_95_22_pad_groupi_n_19 ,csa_tree_add_95_22_pad_groupi_n_898);
  xnor csa_tree_add_95_22_pad_groupi_g4737(csa_tree_add_95_22_pad_groupi_n_1022 ,csa_tree_add_95_22_pad_groupi_n_706 ,csa_tree_add_95_22_pad_groupi_n_844);
  xnor csa_tree_add_95_22_pad_groupi_g4739(csa_tree_add_95_22_pad_groupi_n_1021 ,csa_tree_add_95_22_pad_groupi_n_711 ,in17[9]);
  xnor csa_tree_add_95_22_pad_groupi_g4740(csa_tree_add_95_22_pad_groupi_n_1020 ,csa_tree_add_95_22_pad_groupi_n_645 ,csa_tree_add_95_22_pad_groupi_n_832);
  and csa_tree_add_95_22_pad_groupi_g4741(csa_tree_add_95_22_pad_groupi_n_1019 ,csa_tree_add_95_22_pad_groupi_n_899 ,csa_tree_add_95_22_pad_groupi_n_359);
  and csa_tree_add_95_22_pad_groupi_g4742(csa_tree_add_95_22_pad_groupi_n_1017 ,csa_tree_add_95_22_pad_groupi_n_656 ,csa_tree_add_95_22_pad_groupi_n_923);
  or csa_tree_add_95_22_pad_groupi_g4743(csa_tree_add_95_22_pad_groupi_n_1015 ,csa_tree_add_95_22_pad_groupi_n_682 ,csa_tree_add_95_22_pad_groupi_n_881);
  or csa_tree_add_95_22_pad_groupi_g4744(csa_tree_add_95_22_pad_groupi_n_1013 ,csa_tree_add_95_22_pad_groupi_n_666 ,csa_tree_add_95_22_pad_groupi_n_861);
  xnor csa_tree_add_95_22_pad_groupi_g4745(csa_tree_add_95_22_pad_groupi_n_1012 ,csa_tree_add_95_22_pad_groupi_n_704 ,csa_tree_add_95_22_pad_groupi_n_767);
  xnor csa_tree_add_95_22_pad_groupi_g4746(csa_tree_add_95_22_pad_groupi_n_1011 ,csa_tree_add_95_22_pad_groupi_n_831 ,csa_tree_add_95_22_pad_groupi_n_1);
  or csa_tree_add_95_22_pad_groupi_g4747(csa_tree_add_95_22_pad_groupi_n_1009 ,csa_tree_add_95_22_pad_groupi_n_702 ,csa_tree_add_95_22_pad_groupi_n_931);
  xnor csa_tree_add_95_22_pad_groupi_g4748(csa_tree_add_95_22_pad_groupi_n_974 ,csa_tree_add_95_22_pad_groupi_n_726 ,csa_tree_add_95_22_pad_groupi_n_821);
  xnor csa_tree_add_95_22_pad_groupi_g4749(csa_tree_add_95_22_pad_groupi_n_973 ,csa_tree_add_95_22_pad_groupi_n_802 ,csa_tree_add_95_22_pad_groupi_n_795);
  xnor csa_tree_add_95_22_pad_groupi_g4750(csa_tree_add_95_22_pad_groupi_n_972 ,csa_tree_add_95_22_pad_groupi_n_837 ,csa_tree_add_95_22_pad_groupi_n_766);
  xnor csa_tree_add_95_22_pad_groupi_g4751(csa_tree_add_95_22_pad_groupi_n_971 ,csa_tree_add_95_22_pad_groupi_n_829 ,in17[12]);
  xnor csa_tree_add_95_22_pad_groupi_g4752(csa_tree_add_95_22_pad_groupi_n_970 ,csa_tree_add_95_22_pad_groupi_n_739 ,csa_tree_add_95_22_pad_groupi_n_728);
  xnor csa_tree_add_95_22_pad_groupi_g4753(csa_tree_add_95_22_pad_groupi_n_969 ,csa_tree_add_95_22_pad_groupi_n_758 ,csa_tree_add_95_22_pad_groupi_n_757);
  xor csa_tree_add_95_22_pad_groupi_g4754(csa_tree_add_95_22_pad_groupi_n_968 ,csa_tree_add_95_22_pad_groupi_n_824 ,csa_tree_add_95_22_pad_groupi_n_809);
  xor csa_tree_add_95_22_pad_groupi_g4755(csa_tree_add_95_22_pad_groupi_n_967 ,csa_tree_add_95_22_pad_groupi_n_834 ,in17[8]);
  xnor csa_tree_add_95_22_pad_groupi_g4756(csa_tree_add_95_22_pad_groupi_n_966 ,csa_tree_add_95_22_pad_groupi_n_733 ,csa_tree_add_95_22_pad_groupi_n_755);
  xnor csa_tree_add_95_22_pad_groupi_g4757(csa_tree_add_95_22_pad_groupi_n_965 ,csa_tree_add_95_22_pad_groupi_n_800 ,csa_tree_add_95_22_pad_groupi_n_799);
  xor csa_tree_add_95_22_pad_groupi_g4758(csa_tree_add_95_22_pad_groupi_n_964 ,csa_tree_add_95_22_pad_groupi_n_776 ,csa_tree_add_95_22_pad_groupi_n_721);
  xor csa_tree_add_95_22_pad_groupi_g4759(csa_tree_add_95_22_pad_groupi_n_963 ,csa_tree_add_95_22_pad_groupi_n_772 ,in17[1]);
  xnor csa_tree_add_95_22_pad_groupi_g4760(csa_tree_add_95_22_pad_groupi_n_962 ,csa_tree_add_95_22_pad_groupi_n_765 ,csa_tree_add_95_22_pad_groupi_n_751);
  xnor csa_tree_add_95_22_pad_groupi_g4761(csa_tree_add_95_22_pad_groupi_n_961 ,csa_tree_add_95_22_pad_groupi_n_735 ,csa_tree_add_95_22_pad_groupi_n_792);
  xor csa_tree_add_95_22_pad_groupi_g4762(csa_tree_add_95_22_pad_groupi_n_960 ,csa_tree_add_95_22_pad_groupi_n_771 ,csa_tree_add_95_22_pad_groupi_n_729);
  xnor csa_tree_add_95_22_pad_groupi_g4763(csa_tree_add_95_22_pad_groupi_n_959 ,csa_tree_add_95_22_pad_groupi_n_725 ,csa_tree_add_95_22_pad_groupi_n_723);
  xnor csa_tree_add_95_22_pad_groupi_g4764(csa_tree_add_95_22_pad_groupi_n_958 ,csa_tree_add_95_22_pad_groupi_n_814 ,csa_tree_add_95_22_pad_groupi_n_796);
  xnor csa_tree_add_95_22_pad_groupi_g4765(csa_tree_add_95_22_pad_groupi_n_957 ,csa_tree_add_95_22_pad_groupi_n_784 ,csa_tree_add_95_22_pad_groupi_n_747);
  xor csa_tree_add_95_22_pad_groupi_g4766(csa_tree_add_95_22_pad_groupi_n_956 ,csa_tree_add_95_22_pad_groupi_n_841 ,csa_tree_add_95_22_pad_groupi_n_748);
  xnor csa_tree_add_95_22_pad_groupi_g4767(csa_tree_add_95_22_pad_groupi_n_955 ,csa_tree_add_95_22_pad_groupi_n_760 ,csa_tree_add_95_22_pad_groupi_n_737);
  xnor csa_tree_add_95_22_pad_groupi_g4768(csa_tree_add_95_22_pad_groupi_n_954 ,csa_tree_add_95_22_pad_groupi_n_756 ,in17[2]);
  xnor csa_tree_add_95_22_pad_groupi_g4769(csa_tree_add_95_22_pad_groupi_n_953 ,csa_tree_add_95_22_pad_groupi_n_763 ,csa_tree_add_95_22_pad_groupi_n_817);
  xor csa_tree_add_95_22_pad_groupi_g4770(csa_tree_add_95_22_pad_groupi_n_952 ,csa_tree_add_95_22_pad_groupi_n_823 ,csa_tree_add_95_22_pad_groupi_n_742);
  xnor csa_tree_add_95_22_pad_groupi_g4771(csa_tree_add_95_22_pad_groupi_n_951 ,csa_tree_add_95_22_pad_groupi_n_806 ,csa_tree_add_95_22_pad_groupi_n_753);
  xnor csa_tree_add_95_22_pad_groupi_g4772(csa_tree_add_95_22_pad_groupi_n_950 ,csa_tree_add_95_22_pad_groupi_n_790 ,csa_tree_add_95_22_pad_groupi_n_819);
  xnor csa_tree_add_95_22_pad_groupi_g4773(csa_tree_add_95_22_pad_groupi_n_949 ,csa_tree_add_95_22_pad_groupi_n_813 ,csa_tree_add_95_22_pad_groupi_n_716);
  xnor csa_tree_add_95_22_pad_groupi_g4774(csa_tree_add_95_22_pad_groupi_n_948 ,csa_tree_add_95_22_pad_groupi_n_731 ,in17[6]);
  xnor csa_tree_add_95_22_pad_groupi_g4775(csa_tree_add_95_22_pad_groupi_n_947 ,csa_tree_add_95_22_pad_groupi_n_787 ,in17[5]);
  xnor csa_tree_add_95_22_pad_groupi_g4776(csa_tree_add_95_22_pad_groupi_n_946 ,csa_tree_add_95_22_pad_groupi_n_713 ,in17[7]);
  xnor csa_tree_add_95_22_pad_groupi_g4777(csa_tree_add_95_22_pad_groupi_n_945 ,csa_tree_add_95_22_pad_groupi_n_808 ,csa_tree_add_95_22_pad_groupi_n_788);
  xnor csa_tree_add_95_22_pad_groupi_g4778(csa_tree_add_95_22_pad_groupi_n_944 ,csa_tree_add_95_22_pad_groupi_n_761 ,csa_tree_add_95_22_pad_groupi_n_786);
  xnor csa_tree_add_95_22_pad_groupi_g4779(csa_tree_add_95_22_pad_groupi_n_943 ,csa_tree_add_95_22_pad_groupi_n_798 ,in17[4]);
  xnor csa_tree_add_95_22_pad_groupi_g4780(csa_tree_add_95_22_pad_groupi_n_942 ,csa_tree_add_95_22_pad_groupi_n_719 ,csa_tree_add_95_22_pad_groupi_n_720);
  xnor csa_tree_add_95_22_pad_groupi_g4781(csa_tree_add_95_22_pad_groupi_n_941 ,csa_tree_add_95_22_pad_groupi_n_815 ,csa_tree_add_95_22_pad_groupi_n_717);
  xnor csa_tree_add_95_22_pad_groupi_g4782(csa_tree_add_95_22_pad_groupi_n_940 ,csa_tree_add_95_22_pad_groupi_n_807 ,csa_tree_add_95_22_pad_groupi_n_714);
  xnor csa_tree_add_95_22_pad_groupi_g4783(csa_tree_add_95_22_pad_groupi_n_939 ,csa_tree_add_95_22_pad_groupi_n_810 ,csa_tree_add_95_22_pad_groupi_n_811);
  xnor csa_tree_add_95_22_pad_groupi_g4784(csa_tree_add_95_22_pad_groupi_n_938 ,csa_tree_add_95_22_pad_groupi_n_804 ,in17[3]);
  xnor csa_tree_add_95_22_pad_groupi_g4785(csa_tree_add_95_22_pad_groupi_n_937 ,csa_tree_add_95_22_pad_groupi_n_718 ,csa_tree_add_95_22_pad_groupi_n_793);
  xnor csa_tree_add_95_22_pad_groupi_g4786(csa_tree_add_95_22_pad_groupi_n_977 ,csa_tree_add_95_22_pad_groupi_n_822 ,csa_tree_add_95_22_pad_groupi_n_709);
  xnor csa_tree_add_95_22_pad_groupi_g4787(csa_tree_add_95_22_pad_groupi_n_976 ,csa_tree_add_95_22_pad_groupi_n_828 ,csa_tree_add_95_22_pad_groupi_n_710);
  xnor csa_tree_add_95_22_pad_groupi_g4788(csa_tree_add_95_22_pad_groupi_n_975 ,csa_tree_add_95_22_pad_groupi_n_825 ,in17[0]);
  or csa_tree_add_95_22_pad_groupi_g4791(csa_tree_add_95_22_pad_groupi_n_932 ,csa_tree_add_95_22_pad_groupi_n_815 ,csa_tree_add_95_22_pad_groupi_n_717);
  nor csa_tree_add_95_22_pad_groupi_g4792(csa_tree_add_95_22_pad_groupi_n_931 ,csa_tree_add_95_22_pad_groupi_n_673 ,csa_tree_add_95_22_pad_groupi_n_831);
  nor csa_tree_add_95_22_pad_groupi_g4793(csa_tree_add_95_22_pad_groupi_n_930 ,csa_tree_add_95_22_pad_groupi_n_748 ,csa_tree_add_95_22_pad_groupi_n_785);
  nor csa_tree_add_95_22_pad_groupi_g4794(csa_tree_add_95_22_pad_groupi_n_929 ,csa_tree_add_95_22_pad_groupi_n_802 ,csa_tree_add_95_22_pad_groupi_n_794);
  or csa_tree_add_95_22_pad_groupi_g4795(csa_tree_add_95_22_pad_groupi_n_928 ,csa_tree_add_95_22_pad_groupi_n_807 ,csa_tree_add_95_22_pad_groupi_n_714);
  or csa_tree_add_95_22_pad_groupi_g4796(csa_tree_add_95_22_pad_groupi_n_927 ,csa_tree_add_95_22_pad_groupi_n_801 ,csa_tree_add_95_22_pad_groupi_n_795);
  nor csa_tree_add_95_22_pad_groupi_g4797(csa_tree_add_95_22_pad_groupi_n_926 ,csa_tree_add_95_22_pad_groupi_n_766 ,csa_tree_add_95_22_pad_groupi_n_744);
  and csa_tree_add_95_22_pad_groupi_g4798(csa_tree_add_95_22_pad_groupi_n_925 ,csa_tree_add_95_22_pad_groupi_n_764 ,csa_tree_add_95_22_pad_groupi_n_809);
  or csa_tree_add_95_22_pad_groupi_g4799(csa_tree_add_95_22_pad_groupi_n_924 ,csa_tree_add_95_22_pad_groupi_n_719 ,csa_tree_add_95_22_pad_groupi_n_720);
  or csa_tree_add_95_22_pad_groupi_g4800(csa_tree_add_95_22_pad_groupi_n_923 ,csa_tree_add_95_22_pad_groupi_n_593 ,csa_tree_add_95_22_pad_groupi_n_836);
  or csa_tree_add_95_22_pad_groupi_g4801(csa_tree_add_95_22_pad_groupi_n_922 ,csa_tree_add_95_22_pad_groupi_n_800 ,csa_tree_add_95_22_pad_groupi_n_799);
  or csa_tree_add_95_22_pad_groupi_g4802(csa_tree_add_95_22_pad_groupi_n_921 ,csa_tree_add_95_22_pad_groupi_n_789 ,csa_tree_add_95_22_pad_groupi_n_818);
  nor csa_tree_add_95_22_pad_groupi_g4803(csa_tree_add_95_22_pad_groupi_n_920 ,csa_tree_add_95_22_pad_groupi_n_725 ,csa_tree_add_95_22_pad_groupi_n_723);
  nor csa_tree_add_95_22_pad_groupi_g4804(csa_tree_add_95_22_pad_groupi_n_919 ,csa_tree_add_95_22_pad_groupi_n_763 ,csa_tree_add_95_22_pad_groupi_n_817);
  nor csa_tree_add_95_22_pad_groupi_g4805(csa_tree_add_95_22_pad_groupi_n_918 ,csa_tree_add_95_22_pad_groupi_n_790 ,csa_tree_add_95_22_pad_groupi_n_819);
  nor csa_tree_add_95_22_pad_groupi_g4806(csa_tree_add_95_22_pad_groupi_n_917 ,csa_tree_add_95_22_pad_groupi_n_806 ,csa_tree_add_95_22_pad_groupi_n_753);
  or csa_tree_add_95_22_pad_groupi_g4807(csa_tree_add_95_22_pad_groupi_n_916 ,in17[5] ,csa_tree_add_95_22_pad_groupi_n_787);
  or csa_tree_add_95_22_pad_groupi_g4808(csa_tree_add_95_22_pad_groupi_n_915 ,csa_tree_add_95_22_pad_groupi_n_762 ,csa_tree_add_95_22_pad_groupi_n_816);
  and csa_tree_add_95_22_pad_groupi_g4809(csa_tree_add_95_22_pad_groupi_n_914 ,csa_tree_add_95_22_pad_groupi_n_815 ,csa_tree_add_95_22_pad_groupi_n_717);
  or csa_tree_add_95_22_pad_groupi_g4810(csa_tree_add_95_22_pad_groupi_n_913 ,csa_tree_add_95_22_pad_groupi_n_805 ,csa_tree_add_95_22_pad_groupi_n_752);
  or csa_tree_add_95_22_pad_groupi_g4811(csa_tree_add_95_22_pad_groupi_n_912 ,csa_tree_add_95_22_pad_groupi_n_812 ,csa_tree_add_95_22_pad_groupi_n_715);
  and csa_tree_add_95_22_pad_groupi_g4812(csa_tree_add_95_22_pad_groupi_n_911 ,csa_tree_add_95_22_pad_groupi_n_748 ,csa_tree_add_95_22_pad_groupi_n_785);
  nor csa_tree_add_95_22_pad_groupi_g4813(csa_tree_add_95_22_pad_groupi_n_910 ,csa_tree_add_95_22_pad_groupi_n_372 ,csa_tree_add_95_22_pad_groupi_n_782);
  or csa_tree_add_95_22_pad_groupi_g4814(csa_tree_add_95_22_pad_groupi_n_909 ,csa_tree_add_95_22_pad_groupi_n_814 ,csa_tree_add_95_22_pad_groupi_n_796);
  and csa_tree_add_95_22_pad_groupi_g4815(csa_tree_add_95_22_pad_groupi_n_908 ,csa_tree_add_95_22_pad_groupi_n_810 ,csa_tree_add_95_22_pad_groupi_n_811);
  and csa_tree_add_95_22_pad_groupi_g4816(csa_tree_add_95_22_pad_groupi_n_907 ,csa_tree_add_95_22_pad_groupi_n_807 ,csa_tree_add_95_22_pad_groupi_n_714);
  and csa_tree_add_95_22_pad_groupi_g4817(csa_tree_add_95_22_pad_groupi_n_906 ,in17[4] ,csa_tree_add_95_22_pad_groupi_n_798);
  and csa_tree_add_95_22_pad_groupi_g4818(csa_tree_add_95_22_pad_groupi_n_905 ,in17[5] ,csa_tree_add_95_22_pad_groupi_n_787);
  or csa_tree_add_95_22_pad_groupi_g4819(csa_tree_add_95_22_pad_groupi_n_904 ,csa_tree_add_95_22_pad_groupi_n_808 ,csa_tree_add_95_22_pad_groupi_n_788);
  and csa_tree_add_95_22_pad_groupi_g4820(csa_tree_add_95_22_pad_groupi_n_903 ,csa_tree_add_95_22_pad_groupi_n_814 ,csa_tree_add_95_22_pad_groupi_n_796);
  nor csa_tree_add_95_22_pad_groupi_g4821(csa_tree_add_95_22_pad_groupi_n_902 ,csa_tree_add_95_22_pad_groupi_n_813 ,csa_tree_add_95_22_pad_groupi_n_716);
  and csa_tree_add_95_22_pad_groupi_g4822(csa_tree_add_95_22_pad_groupi_n_901 ,csa_tree_add_95_22_pad_groupi_n_761 ,csa_tree_add_95_22_pad_groupi_n_786);
  nor csa_tree_add_95_22_pad_groupi_g4823(csa_tree_add_95_22_pad_groupi_n_900 ,csa_tree_add_95_22_pad_groupi_n_783 ,csa_tree_add_95_22_pad_groupi_n_729);
  or csa_tree_add_95_22_pad_groupi_g4824(csa_tree_add_95_22_pad_groupi_n_899 ,csa_tree_add_95_22_pad_groupi_n_708 ,csa_tree_add_95_22_pad_groupi_n_845);
  or csa_tree_add_95_22_pad_groupi_g4825(csa_tree_add_95_22_pad_groupi_n_898 ,csa_tree_add_95_22_pad_groupi_n_112 ,csa_tree_add_95_22_pad_groupi_n_781);
  and csa_tree_add_95_22_pad_groupi_g4826(csa_tree_add_95_22_pad_groupi_n_897 ,csa_tree_add_95_22_pad_groupi_n_783 ,csa_tree_add_95_22_pad_groupi_n_729);
  and csa_tree_add_95_22_pad_groupi_g4827(csa_tree_add_95_22_pad_groupi_n_896 ,csa_tree_add_95_22_pad_groupi_n_372 ,csa_tree_add_95_22_pad_groupi_n_782);
  or csa_tree_add_95_22_pad_groupi_g4828(csa_tree_add_95_22_pad_groupi_n_895 ,csa_tree_add_95_22_pad_groupi_n_734 ,csa_tree_add_95_22_pad_groupi_n_791);
  nor csa_tree_add_95_22_pad_groupi_g4829(csa_tree_add_95_22_pad_groupi_n_894 ,csa_tree_add_95_22_pad_groupi_n_735 ,csa_tree_add_95_22_pad_groupi_n_792);
  or csa_tree_add_95_22_pad_groupi_g4830(csa_tree_add_95_22_pad_groupi_n_936 ,csa_tree_add_95_22_pad_groupi_n_645 ,csa_tree_add_95_22_pad_groupi_n_833);
  and csa_tree_add_95_22_pad_groupi_g4831(csa_tree_add_95_22_pad_groupi_n_935 ,csa_tree_add_95_22_pad_groupi_n_705 ,csa_tree_add_95_22_pad_groupi_n_767);
  and csa_tree_add_95_22_pad_groupi_g4832(csa_tree_add_95_22_pad_groupi_n_934 ,csa_tree_add_95_22_pad_groupi_n_708 ,csa_tree_add_95_22_pad_groupi_n_845);
  and csa_tree_add_95_22_pad_groupi_g4833(csa_tree_add_95_22_pad_groupi_n_933 ,csa_tree_add_95_22_pad_groupi_n_707 ,csa_tree_add_95_22_pad_groupi_n_844);
  or csa_tree_add_95_22_pad_groupi_g4834(csa_tree_add_95_22_pad_groupi_n_891 ,csa_tree_add_95_22_pad_groupi_n_718 ,csa_tree_add_95_22_pad_groupi_n_793);
  and csa_tree_add_95_22_pad_groupi_g4835(csa_tree_add_95_22_pad_groupi_n_890 ,csa_tree_add_95_22_pad_groupi_n_800 ,csa_tree_add_95_22_pad_groupi_n_799);
  and csa_tree_add_95_22_pad_groupi_g4836(csa_tree_add_95_22_pad_groupi_n_889 ,csa_tree_add_95_22_pad_groupi_n_718 ,csa_tree_add_95_22_pad_groupi_n_793);
  or csa_tree_add_95_22_pad_groupi_g4837(csa_tree_add_95_22_pad_groupi_n_888 ,csa_tree_add_95_22_pad_groupi_n_732 ,csa_tree_add_95_22_pad_groupi_n_754);
  and csa_tree_add_95_22_pad_groupi_g4838(csa_tree_add_95_22_pad_groupi_n_887 ,in17[3] ,csa_tree_add_95_22_pad_groupi_n_804);
  and csa_tree_add_95_22_pad_groupi_g4839(csa_tree_add_95_22_pad_groupi_n_886 ,csa_tree_add_95_22_pad_groupi_n_719 ,csa_tree_add_95_22_pad_groupi_n_720);
  or csa_tree_add_95_22_pad_groupi_g4840(csa_tree_add_95_22_pad_groupi_n_885 ,in17[3] ,csa_tree_add_95_22_pad_groupi_n_804);
  or csa_tree_add_95_22_pad_groupi_g4841(csa_tree_add_95_22_pad_groupi_n_884 ,csa_tree_add_95_22_pad_groupi_n_738 ,csa_tree_add_95_22_pad_groupi_n_727);
  nor csa_tree_add_95_22_pad_groupi_g4842(csa_tree_add_95_22_pad_groupi_n_883 ,csa_tree_add_95_22_pad_groupi_n_803 ,csa_tree_add_95_22_pad_groupi_n_721);
  nor csa_tree_add_95_22_pad_groupi_g4843(csa_tree_add_95_22_pad_groupi_n_882 ,csa_tree_add_95_22_pad_groupi_n_739 ,csa_tree_add_95_22_pad_groupi_n_728);
  nor csa_tree_add_95_22_pad_groupi_g4844(csa_tree_add_95_22_pad_groupi_n_881 ,csa_tree_add_95_22_pad_groupi_n_700 ,csa_tree_add_95_22_pad_groupi_n_828);
  or csa_tree_add_95_22_pad_groupi_g4845(csa_tree_add_95_22_pad_groupi_n_880 ,csa_tree_add_95_22_pad_groupi_n_761 ,csa_tree_add_95_22_pad_groupi_n_786);
  nor csa_tree_add_95_22_pad_groupi_g4846(csa_tree_add_95_22_pad_groupi_n_879 ,csa_tree_add_95_22_pad_groupi_n_371 ,csa_tree_add_95_22_pad_groupi_n_740);
  or csa_tree_add_95_22_pad_groupi_g4847(csa_tree_add_95_22_pad_groupi_n_878 ,csa_tree_add_95_22_pad_groupi_n_387 ,csa_tree_add_95_22_pad_groupi_n_712);
  and csa_tree_add_95_22_pad_groupi_g4848(csa_tree_add_95_22_pad_groupi_n_877 ,csa_tree_add_95_22_pad_groupi_n_766 ,csa_tree_add_95_22_pad_groupi_n_744);
  nor csa_tree_add_95_22_pad_groupi_g4849(csa_tree_add_95_22_pad_groupi_n_876 ,csa_tree_add_95_22_pad_groupi_n_733 ,csa_tree_add_95_22_pad_groupi_n_755);
  nor csa_tree_add_95_22_pad_groupi_g4850(csa_tree_add_95_22_pad_groupi_n_875 ,in17[7] ,csa_tree_add_95_22_pad_groupi_n_713);
  and csa_tree_add_95_22_pad_groupi_g4851(csa_tree_add_95_22_pad_groupi_n_874 ,csa_tree_add_95_22_pad_groupi_n_803 ,csa_tree_add_95_22_pad_groupi_n_721);
  and csa_tree_add_95_22_pad_groupi_g4852(csa_tree_add_95_22_pad_groupi_n_873 ,csa_tree_add_95_22_pad_groupi_n_758 ,csa_tree_add_95_22_pad_groupi_n_757);
  nor csa_tree_add_95_22_pad_groupi_g4853(csa_tree_add_95_22_pad_groupi_n_872 ,csa_tree_add_95_22_pad_groupi_n_764 ,csa_tree_add_95_22_pad_groupi_n_809);
  or csa_tree_add_95_22_pad_groupi_g4854(csa_tree_add_95_22_pad_groupi_n_871 ,csa_tree_add_95_22_pad_groupi_n_758 ,csa_tree_add_95_22_pad_groupi_n_757);
  and csa_tree_add_95_22_pad_groupi_g4855(csa_tree_add_95_22_pad_groupi_n_870 ,in17[2] ,csa_tree_add_95_22_pad_groupi_n_756);
  and csa_tree_add_95_22_pad_groupi_g4856(csa_tree_add_95_22_pad_groupi_n_869 ,csa_tree_add_95_22_pad_groupi_n_808 ,csa_tree_add_95_22_pad_groupi_n_788);
  and csa_tree_add_95_22_pad_groupi_g4857(csa_tree_add_95_22_pad_groupi_n_868 ,csa_tree_add_95_22_pad_groupi_n_784 ,csa_tree_add_95_22_pad_groupi_n_747);
  or csa_tree_add_95_22_pad_groupi_g4858(csa_tree_add_95_22_pad_groupi_n_867 ,csa_tree_add_95_22_pad_groupi_n_810 ,csa_tree_add_95_22_pad_groupi_n_811);
  and csa_tree_add_95_22_pad_groupi_g4859(csa_tree_add_95_22_pad_groupi_n_866 ,csa_tree_add_95_22_pad_groupi_n_765 ,csa_tree_add_95_22_pad_groupi_n_751);
  or csa_tree_add_95_22_pad_groupi_g4860(csa_tree_add_95_22_pad_groupi_n_865 ,csa_tree_add_95_22_pad_groupi_n_784 ,csa_tree_add_95_22_pad_groupi_n_747);
  or csa_tree_add_95_22_pad_groupi_g4861(csa_tree_add_95_22_pad_groupi_n_864 ,csa_tree_add_95_22_pad_groupi_n_749 ,csa_tree_add_95_22_pad_groupi_n_741);
  or csa_tree_add_95_22_pad_groupi_g4862(csa_tree_add_95_22_pad_groupi_n_863 ,csa_tree_add_95_22_pad_groupi_n_765 ,csa_tree_add_95_22_pad_groupi_n_751);
  nor csa_tree_add_95_22_pad_groupi_g4863(csa_tree_add_95_22_pad_groupi_n_862 ,csa_tree_add_95_22_pad_groupi_n_750 ,csa_tree_add_95_22_pad_groupi_n_742);
  nor csa_tree_add_95_22_pad_groupi_g4864(csa_tree_add_95_22_pad_groupi_n_861 ,csa_tree_add_95_22_pad_groupi_n_600 ,csa_tree_add_95_22_pad_groupi_n_822);
  or csa_tree_add_95_22_pad_groupi_g4865(csa_tree_add_95_22_pad_groupi_n_860 ,csa_tree_add_95_22_pad_groupi_n_726 ,csa_tree_add_95_22_pad_groupi_n_821);
  and csa_tree_add_95_22_pad_groupi_g4866(csa_tree_add_95_22_pad_groupi_n_859 ,csa_tree_add_95_22_pad_groupi_n_371 ,csa_tree_add_95_22_pad_groupi_n_740);
  and csa_tree_add_95_22_pad_groupi_g4867(csa_tree_add_95_22_pad_groupi_n_858 ,csa_tree_add_95_22_pad_groupi_n_726 ,csa_tree_add_95_22_pad_groupi_n_821);
  or csa_tree_add_95_22_pad_groupi_g4868(csa_tree_add_95_22_pad_groupi_n_857 ,csa_tree_add_95_22_pad_groupi_n_759 ,csa_tree_add_95_22_pad_groupi_n_736);
  or csa_tree_add_95_22_pad_groupi_g4869(csa_tree_add_95_22_pad_groupi_n_856 ,in17[4] ,csa_tree_add_95_22_pad_groupi_n_798);
  nor csa_tree_add_95_22_pad_groupi_g4870(csa_tree_add_95_22_pad_groupi_n_855 ,in17[2] ,csa_tree_add_95_22_pad_groupi_n_756);
  nor csa_tree_add_95_22_pad_groupi_g4871(csa_tree_add_95_22_pad_groupi_n_854 ,csa_tree_add_95_22_pad_groupi_n_760 ,csa_tree_add_95_22_pad_groupi_n_737);
  or csa_tree_add_95_22_pad_groupi_g4872(csa_tree_add_95_22_pad_groupi_n_853 ,csa_tree_add_95_22_pad_groupi_n_370 ,csa_tree_add_95_22_pad_groupi_n_730);
  or csa_tree_add_95_22_pad_groupi_g4873(csa_tree_add_95_22_pad_groupi_n_852 ,csa_tree_add_95_22_pad_groupi_n_724 ,csa_tree_add_95_22_pad_groupi_n_722);
  nor csa_tree_add_95_22_pad_groupi_g4874(csa_tree_add_95_22_pad_groupi_n_851 ,in17[6] ,csa_tree_add_95_22_pad_groupi_n_731);
  or csa_tree_add_95_22_pad_groupi_g4876(csa_tree_add_95_22_pad_groupi_n_893 ,csa_tree_add_95_22_pad_groupi_n_374 ,csa_tree_add_95_22_pad_groupi_n_826);
  or csa_tree_add_95_22_pad_groupi_g4877(csa_tree_add_95_22_pad_groupi_n_892 ,csa_tree_add_95_22_pad_groupi_n_847 ,csa_tree_add_95_22_pad_groupi_n_849);
  not csa_tree_add_95_22_pad_groupi_g4878(csa_tree_add_95_22_pad_groupi_n_849 ,csa_tree_add_95_22_pad_groupi_n_848);
  not csa_tree_add_95_22_pad_groupi_g4879(csa_tree_add_95_22_pad_groupi_n_847 ,csa_tree_add_95_22_pad_groupi_n_846);
  not csa_tree_add_95_22_pad_groupi_g4880(csa_tree_add_95_22_pad_groupi_n_843 ,csa_tree_add_95_22_pad_groupi_n_842);
  not csa_tree_add_95_22_pad_groupi_g4883(csa_tree_add_95_22_pad_groupi_n_833 ,csa_tree_add_95_22_pad_groupi_n_832);
  not csa_tree_add_95_22_pad_groupi_g4884(csa_tree_add_95_22_pad_groupi_n_826 ,csa_tree_add_95_22_pad_groupi_n_825);
  not csa_tree_add_95_22_pad_groupi_g4885(csa_tree_add_95_22_pad_groupi_n_818 ,csa_tree_add_95_22_pad_groupi_n_819);
  not csa_tree_add_95_22_pad_groupi_g4886(csa_tree_add_95_22_pad_groupi_n_816 ,csa_tree_add_95_22_pad_groupi_n_817);
  not csa_tree_add_95_22_pad_groupi_g4887(csa_tree_add_95_22_pad_groupi_n_812 ,csa_tree_add_95_22_pad_groupi_n_813);
  not csa_tree_add_95_22_pad_groupi_g4888(csa_tree_add_95_22_pad_groupi_n_805 ,csa_tree_add_95_22_pad_groupi_n_806);
  not csa_tree_add_95_22_pad_groupi_g4889(csa_tree_add_95_22_pad_groupi_n_801 ,csa_tree_add_95_22_pad_groupi_n_802);
  not csa_tree_add_95_22_pad_groupi_g4890(csa_tree_add_95_22_pad_groupi_n_794 ,csa_tree_add_95_22_pad_groupi_n_795);
  not csa_tree_add_95_22_pad_groupi_g4891(csa_tree_add_95_22_pad_groupi_n_791 ,csa_tree_add_95_22_pad_groupi_n_792);
  not csa_tree_add_95_22_pad_groupi_g4892(csa_tree_add_95_22_pad_groupi_n_789 ,csa_tree_add_95_22_pad_groupi_n_790);
  and csa_tree_add_95_22_pad_groupi_g4893(csa_tree_add_95_22_pad_groupi_n_781 ,csa_tree_add_95_22_pad_groupi_n_459 ,csa_tree_add_95_22_pad_groupi_n_612);
  or csa_tree_add_95_22_pad_groupi_g4894(csa_tree_add_95_22_pad_groupi_n_848 ,csa_tree_add_95_22_pad_groupi_n_466 ,csa_tree_add_95_22_pad_groupi_n_621);
  or csa_tree_add_95_22_pad_groupi_g4895(csa_tree_add_95_22_pad_groupi_n_846 ,csa_tree_add_95_22_pad_groupi_n_576 ,csa_tree_add_95_22_pad_groupi_n_703);
  and csa_tree_add_95_22_pad_groupi_g4896(csa_tree_add_95_22_pad_groupi_n_845 ,csa_tree_add_95_22_pad_groupi_n_531 ,csa_tree_add_95_22_pad_groupi_n_685);
  or csa_tree_add_95_22_pad_groupi_g4897(csa_tree_add_95_22_pad_groupi_n_844 ,csa_tree_add_95_22_pad_groupi_n_526 ,csa_tree_add_95_22_pad_groupi_n_652);
  or csa_tree_add_95_22_pad_groupi_g4898(csa_tree_add_95_22_pad_groupi_n_842 ,csa_tree_add_95_22_pad_groupi_n_533 ,csa_tree_add_95_22_pad_groupi_n_618);
  and csa_tree_add_95_22_pad_groupi_g4899(csa_tree_add_95_22_pad_groupi_n_841 ,csa_tree_add_95_22_pad_groupi_n_472 ,csa_tree_add_95_22_pad_groupi_n_642);
  or csa_tree_add_95_22_pad_groupi_g4900(csa_tree_add_95_22_pad_groupi_n_840 ,csa_tree_add_95_22_pad_groupi_n_557 ,csa_tree_add_95_22_pad_groupi_n_598);
  or csa_tree_add_95_22_pad_groupi_g4901(csa_tree_add_95_22_pad_groupi_n_839 ,csa_tree_add_95_22_pad_groupi_n_574 ,csa_tree_add_95_22_pad_groupi_n_588);
  and csa_tree_add_95_22_pad_groupi_g4903(csa_tree_add_95_22_pad_groupi_n_837 ,csa_tree_add_95_22_pad_groupi_n_483 ,csa_tree_add_95_22_pad_groupi_n_587);
  and csa_tree_add_95_22_pad_groupi_g4906(csa_tree_add_95_22_pad_groupi_n_834 ,csa_tree_add_95_22_pad_groupi_n_460 ,csa_tree_add_95_22_pad_groupi_n_586);
  or csa_tree_add_95_22_pad_groupi_g4907(csa_tree_add_95_22_pad_groupi_n_832 ,csa_tree_add_95_22_pad_groupi_n_548 ,csa_tree_add_95_22_pad_groupi_n_699);
  or csa_tree_add_95_22_pad_groupi_g4912(csa_tree_add_95_22_pad_groupi_n_827 ,csa_tree_add_95_22_pad_groupi_n_487 ,csa_tree_add_95_22_pad_groupi_n_647);
  or csa_tree_add_95_22_pad_groupi_g4913(csa_tree_add_95_22_pad_groupi_n_825 ,csa_tree_add_95_22_pad_groupi_n_462 ,csa_tree_add_95_22_pad_groupi_n_662);
  and csa_tree_add_95_22_pad_groupi_g4914(csa_tree_add_95_22_pad_groupi_n_824 ,csa_tree_add_95_22_pad_groupi_n_485 ,csa_tree_add_95_22_pad_groupi_n_683);
  and csa_tree_add_95_22_pad_groupi_g4915(csa_tree_add_95_22_pad_groupi_n_823 ,csa_tree_add_95_22_pad_groupi_n_518 ,csa_tree_add_95_22_pad_groupi_n_595);
  or csa_tree_add_95_22_pad_groupi_g4917(csa_tree_add_95_22_pad_groupi_n_821 ,csa_tree_add_95_22_pad_groupi_n_551 ,csa_tree_add_95_22_pad_groupi_n_665);
  or csa_tree_add_95_22_pad_groupi_g4918(csa_tree_add_95_22_pad_groupi_n_820 ,csa_tree_add_95_22_pad_groupi_n_556 ,csa_tree_add_95_22_pad_groupi_n_677);
  or csa_tree_add_95_22_pad_groupi_g4919(csa_tree_add_95_22_pad_groupi_n_819 ,csa_tree_add_95_22_pad_groupi_n_516 ,csa_tree_add_95_22_pad_groupi_n_681);
  or csa_tree_add_95_22_pad_groupi_g4920(csa_tree_add_95_22_pad_groupi_n_817 ,csa_tree_add_95_22_pad_groupi_n_527 ,csa_tree_add_95_22_pad_groupi_n_674);
  or csa_tree_add_95_22_pad_groupi_g4921(csa_tree_add_95_22_pad_groupi_n_815 ,csa_tree_add_95_22_pad_groupi_n_491 ,csa_tree_add_95_22_pad_groupi_n_649);
  or csa_tree_add_95_22_pad_groupi_g4922(csa_tree_add_95_22_pad_groupi_n_814 ,csa_tree_add_95_22_pad_groupi_n_475 ,csa_tree_add_95_22_pad_groupi_n_633);
  or csa_tree_add_95_22_pad_groupi_g4923(csa_tree_add_95_22_pad_groupi_n_813 ,csa_tree_add_95_22_pad_groupi_n_525 ,csa_tree_add_95_22_pad_groupi_n_695);
  or csa_tree_add_95_22_pad_groupi_g4924(csa_tree_add_95_22_pad_groupi_n_811 ,csa_tree_add_95_22_pad_groupi_n_476 ,csa_tree_add_95_22_pad_groupi_n_599);
  or csa_tree_add_95_22_pad_groupi_g4925(csa_tree_add_95_22_pad_groupi_n_810 ,csa_tree_add_95_22_pad_groupi_n_470 ,csa_tree_add_95_22_pad_groupi_n_627);
  or csa_tree_add_95_22_pad_groupi_g4926(csa_tree_add_95_22_pad_groupi_n_809 ,csa_tree_add_95_22_pad_groupi_n_528 ,csa_tree_add_95_22_pad_groupi_n_651);
  or csa_tree_add_95_22_pad_groupi_g4927(csa_tree_add_95_22_pad_groupi_n_808 ,csa_tree_add_95_22_pad_groupi_n_541 ,csa_tree_add_95_22_pad_groupi_n_635);
  or csa_tree_add_95_22_pad_groupi_g4928(csa_tree_add_95_22_pad_groupi_n_807 ,csa_tree_add_95_22_pad_groupi_n_512 ,csa_tree_add_95_22_pad_groupi_n_625);
  or csa_tree_add_95_22_pad_groupi_g4929(csa_tree_add_95_22_pad_groupi_n_806 ,csa_tree_add_95_22_pad_groupi_n_523 ,csa_tree_add_95_22_pad_groupi_n_623);
  or csa_tree_add_95_22_pad_groupi_g4930(csa_tree_add_95_22_pad_groupi_n_804 ,csa_tree_add_95_22_pad_groupi_n_461 ,csa_tree_add_95_22_pad_groupi_n_694);
  or csa_tree_add_95_22_pad_groupi_g4931(csa_tree_add_95_22_pad_groupi_n_803 ,csa_tree_add_95_22_pad_groupi_n_529 ,csa_tree_add_95_22_pad_groupi_n_653);
  or csa_tree_add_95_22_pad_groupi_g4933(csa_tree_add_95_22_pad_groupi_n_800 ,csa_tree_add_95_22_pad_groupi_n_477 ,csa_tree_add_95_22_pad_groupi_n_658);
  or csa_tree_add_95_22_pad_groupi_g4934(csa_tree_add_95_22_pad_groupi_n_799 ,csa_tree_add_95_22_pad_groupi_n_467 ,csa_tree_add_95_22_pad_groupi_n_680);
  or csa_tree_add_95_22_pad_groupi_g4935(csa_tree_add_95_22_pad_groupi_n_798 ,csa_tree_add_95_22_pad_groupi_n_468 ,csa_tree_add_95_22_pad_groupi_n_607);
  or csa_tree_add_95_22_pad_groupi_g4936(csa_tree_add_95_22_pad_groupi_n_797 ,csa_tree_add_95_22_pad_groupi_n_394 ,csa_tree_add_95_22_pad_groupi_n_663);
  or csa_tree_add_95_22_pad_groupi_g4937(csa_tree_add_95_22_pad_groupi_n_796 ,csa_tree_add_95_22_pad_groupi_n_555 ,csa_tree_add_95_22_pad_groupi_n_669);
  or csa_tree_add_95_22_pad_groupi_g4938(csa_tree_add_95_22_pad_groupi_n_795 ,csa_tree_add_95_22_pad_groupi_n_547 ,csa_tree_add_95_22_pad_groupi_n_696);
  or csa_tree_add_95_22_pad_groupi_g4939(csa_tree_add_95_22_pad_groupi_n_793 ,csa_tree_add_95_22_pad_groupi_n_540 ,csa_tree_add_95_22_pad_groupi_n_697);
  or csa_tree_add_95_22_pad_groupi_g4940(csa_tree_add_95_22_pad_groupi_n_792 ,csa_tree_add_95_22_pad_groupi_n_456 ,csa_tree_add_95_22_pad_groupi_n_638);
  or csa_tree_add_95_22_pad_groupi_g4941(csa_tree_add_95_22_pad_groupi_n_790 ,csa_tree_add_95_22_pad_groupi_n_524 ,csa_tree_add_95_22_pad_groupi_n_661);
  or csa_tree_add_95_22_pad_groupi_g4942(csa_tree_add_95_22_pad_groupi_n_788 ,csa_tree_add_95_22_pad_groupi_n_537 ,csa_tree_add_95_22_pad_groupi_n_616);
  or csa_tree_add_95_22_pad_groupi_g4943(csa_tree_add_95_22_pad_groupi_n_787 ,csa_tree_add_95_22_pad_groupi_n_469 ,csa_tree_add_95_22_pad_groupi_n_672);
  or csa_tree_add_95_22_pad_groupi_g4944(csa_tree_add_95_22_pad_groupi_n_786 ,csa_tree_add_95_22_pad_groupi_n_473 ,csa_tree_add_95_22_pad_groupi_n_589);
  or csa_tree_add_95_22_pad_groupi_g4945(csa_tree_add_95_22_pad_groupi_n_785 ,csa_tree_add_95_22_pad_groupi_n_484 ,csa_tree_add_95_22_pad_groupi_n_698);
  or csa_tree_add_95_22_pad_groupi_g4946(csa_tree_add_95_22_pad_groupi_n_784 ,csa_tree_add_95_22_pad_groupi_n_488 ,csa_tree_add_95_22_pad_groupi_n_608);
  or csa_tree_add_95_22_pad_groupi_g4947(csa_tree_add_95_22_pad_groupi_n_783 ,csa_tree_add_95_22_pad_groupi_n_546 ,csa_tree_add_95_22_pad_groupi_n_648);
  not csa_tree_add_95_22_pad_groupi_g4949(csa_tree_add_95_22_pad_groupi_n_779 ,csa_tree_add_95_22_pad_groupi_n_778);
  not csa_tree_add_95_22_pad_groupi_g4950(csa_tree_add_95_22_pad_groupi_n_762 ,csa_tree_add_95_22_pad_groupi_n_763);
  not csa_tree_add_95_22_pad_groupi_g4951(csa_tree_add_95_22_pad_groupi_n_759 ,csa_tree_add_95_22_pad_groupi_n_760);
  not csa_tree_add_95_22_pad_groupi_g4952(csa_tree_add_95_22_pad_groupi_n_754 ,csa_tree_add_95_22_pad_groupi_n_755);
  not csa_tree_add_95_22_pad_groupi_g4953(csa_tree_add_95_22_pad_groupi_n_752 ,csa_tree_add_95_22_pad_groupi_n_753);
  not csa_tree_add_95_22_pad_groupi_g4954(csa_tree_add_95_22_pad_groupi_n_749 ,csa_tree_add_95_22_pad_groupi_n_750);
  not csa_tree_add_95_22_pad_groupi_g4955(csa_tree_add_95_22_pad_groupi_n_745 ,csa_tree_add_95_22_pad_groupi_n_746);
  not csa_tree_add_95_22_pad_groupi_g4956(csa_tree_add_95_22_pad_groupi_n_744 ,csa_tree_add_95_22_pad_groupi_n_743);
  not csa_tree_add_95_22_pad_groupi_g4957(csa_tree_add_95_22_pad_groupi_n_741 ,csa_tree_add_95_22_pad_groupi_n_742);
  not csa_tree_add_95_22_pad_groupi_g4958(csa_tree_add_95_22_pad_groupi_n_738 ,csa_tree_add_95_22_pad_groupi_n_739);
  not csa_tree_add_95_22_pad_groupi_g4959(csa_tree_add_95_22_pad_groupi_n_736 ,csa_tree_add_95_22_pad_groupi_n_737);
  not csa_tree_add_95_22_pad_groupi_g4960(csa_tree_add_95_22_pad_groupi_n_734 ,csa_tree_add_95_22_pad_groupi_n_735);
  not csa_tree_add_95_22_pad_groupi_g4961(csa_tree_add_95_22_pad_groupi_n_732 ,csa_tree_add_95_22_pad_groupi_n_733);
  not csa_tree_add_95_22_pad_groupi_g4962(csa_tree_add_95_22_pad_groupi_n_730 ,csa_tree_add_95_22_pad_groupi_n_731);
  not csa_tree_add_95_22_pad_groupi_g4963(csa_tree_add_95_22_pad_groupi_n_727 ,csa_tree_add_95_22_pad_groupi_n_728);
  not csa_tree_add_95_22_pad_groupi_g4964(csa_tree_add_95_22_pad_groupi_n_724 ,csa_tree_add_95_22_pad_groupi_n_725);
  not csa_tree_add_95_22_pad_groupi_g4965(csa_tree_add_95_22_pad_groupi_n_722 ,csa_tree_add_95_22_pad_groupi_n_723);
  not csa_tree_add_95_22_pad_groupi_g4966(csa_tree_add_95_22_pad_groupi_n_715 ,csa_tree_add_95_22_pad_groupi_n_716);
  not csa_tree_add_95_22_pad_groupi_g4967(csa_tree_add_95_22_pad_groupi_n_712 ,csa_tree_add_95_22_pad_groupi_n_713);
  xnor csa_tree_add_95_22_pad_groupi_g4968(csa_tree_add_95_22_pad_groupi_n_711 ,csa_tree_add_95_22_pad_groupi_n_583 ,in17[10]);
  xnor csa_tree_add_95_22_pad_groupi_g4970(csa_tree_add_95_22_pad_groupi_n_710 ,csa_tree_add_95_22_pad_groupi_n_282 ,in17[12]);
  xnor csa_tree_add_95_22_pad_groupi_g4972(csa_tree_add_95_22_pad_groupi_n_709 ,csa_tree_add_95_22_pad_groupi_n_582 ,in17[12]);
  or csa_tree_add_95_22_pad_groupi_g4975(csa_tree_add_95_22_pad_groupi_n_778 ,csa_tree_add_95_22_pad_groupi_n_539 ,csa_tree_add_95_22_pad_groupi_n_626);
  or csa_tree_add_95_22_pad_groupi_g4976(csa_tree_add_95_22_pad_groupi_n_777 ,csa_tree_add_95_22_pad_groupi_n_550 ,csa_tree_add_95_22_pad_groupi_n_624);
  and csa_tree_add_95_22_pad_groupi_g4977(csa_tree_add_95_22_pad_groupi_n_776 ,csa_tree_add_95_22_pad_groupi_n_464 ,csa_tree_add_95_22_pad_groupi_n_655);
  or csa_tree_add_95_22_pad_groupi_g4978(csa_tree_add_95_22_pad_groupi_n_775 ,csa_tree_add_95_22_pad_groupi_n_482 ,csa_tree_add_95_22_pad_groupi_n_637);
  or csa_tree_add_95_22_pad_groupi_g4980(csa_tree_add_95_22_pad_groupi_n_773 ,csa_tree_add_95_22_pad_groupi_n_519 ,csa_tree_add_95_22_pad_groupi_n_605);
  and csa_tree_add_95_22_pad_groupi_g4981(csa_tree_add_95_22_pad_groupi_n_772 ,csa_tree_add_95_22_pad_groupi_n_457 ,csa_tree_add_95_22_pad_groupi_n_594);
  and csa_tree_add_95_22_pad_groupi_g4982(csa_tree_add_95_22_pad_groupi_n_771 ,csa_tree_add_95_22_pad_groupi_n_492 ,csa_tree_add_95_22_pad_groupi_n_606);
  or csa_tree_add_95_22_pad_groupi_g4984(csa_tree_add_95_22_pad_groupi_n_769 ,csa_tree_add_95_22_pad_groupi_n_490 ,csa_tree_add_95_22_pad_groupi_n_689);
  or csa_tree_add_95_22_pad_groupi_g4985(csa_tree_add_95_22_pad_groupi_n_768 ,csa_tree_add_95_22_pad_groupi_n_545 ,csa_tree_add_95_22_pad_groupi_n_640);
  or csa_tree_add_95_22_pad_groupi_g4986(csa_tree_add_95_22_pad_groupi_n_767 ,csa_tree_add_95_22_pad_groupi_n_552 ,csa_tree_add_95_22_pad_groupi_n_659);
  or csa_tree_add_95_22_pad_groupi_g4988(csa_tree_add_95_22_pad_groupi_n_765 ,csa_tree_add_95_22_pad_groupi_n_517 ,csa_tree_add_95_22_pad_groupi_n_688);
  or csa_tree_add_95_22_pad_groupi_g4989(csa_tree_add_95_22_pad_groupi_n_764 ,csa_tree_add_95_22_pad_groupi_n_554 ,csa_tree_add_95_22_pad_groupi_n_654);
  or csa_tree_add_95_22_pad_groupi_g4990(csa_tree_add_95_22_pad_groupi_n_763 ,csa_tree_add_95_22_pad_groupi_n_480 ,csa_tree_add_95_22_pad_groupi_n_602);
  or csa_tree_add_95_22_pad_groupi_g4991(csa_tree_add_95_22_pad_groupi_n_761 ,csa_tree_add_95_22_pad_groupi_n_577 ,csa_tree_add_95_22_pad_groupi_n_693);
  or csa_tree_add_95_22_pad_groupi_g4992(csa_tree_add_95_22_pad_groupi_n_760 ,csa_tree_add_95_22_pad_groupi_n_478 ,csa_tree_add_95_22_pad_groupi_n_591);
  or csa_tree_add_95_22_pad_groupi_g4993(csa_tree_add_95_22_pad_groupi_n_758 ,csa_tree_add_95_22_pad_groupi_n_514 ,csa_tree_add_95_22_pad_groupi_n_604);
  or csa_tree_add_95_22_pad_groupi_g4994(csa_tree_add_95_22_pad_groupi_n_757 ,csa_tree_add_95_22_pad_groupi_n_532 ,csa_tree_add_95_22_pad_groupi_n_617);
  or csa_tree_add_95_22_pad_groupi_g4995(csa_tree_add_95_22_pad_groupi_n_756 ,csa_tree_add_95_22_pad_groupi_n_455 ,csa_tree_add_95_22_pad_groupi_n_670);
  or csa_tree_add_95_22_pad_groupi_g4996(csa_tree_add_95_22_pad_groupi_n_755 ,csa_tree_add_95_22_pad_groupi_n_544 ,csa_tree_add_95_22_pad_groupi_n_660);
  or csa_tree_add_95_22_pad_groupi_g4997(csa_tree_add_95_22_pad_groupi_n_753 ,csa_tree_add_95_22_pad_groupi_n_486 ,csa_tree_add_95_22_pad_groupi_n_679);
  or csa_tree_add_95_22_pad_groupi_g4998(csa_tree_add_95_22_pad_groupi_n_751 ,csa_tree_add_95_22_pad_groupi_n_575 ,csa_tree_add_95_22_pad_groupi_n_619);
  or csa_tree_add_95_22_pad_groupi_g4999(csa_tree_add_95_22_pad_groupi_n_750 ,csa_tree_add_95_22_pad_groupi_n_522 ,csa_tree_add_95_22_pad_groupi_n_671);
  or csa_tree_add_95_22_pad_groupi_g5000(csa_tree_add_95_22_pad_groupi_n_748 ,csa_tree_add_95_22_pad_groupi_n_515 ,csa_tree_add_95_22_pad_groupi_n_631);
  or csa_tree_add_95_22_pad_groupi_g5001(csa_tree_add_95_22_pad_groupi_n_747 ,csa_tree_add_95_22_pad_groupi_n_573 ,csa_tree_add_95_22_pad_groupi_n_620);
  or csa_tree_add_95_22_pad_groupi_g5002(csa_tree_add_95_22_pad_groupi_n_746 ,csa_tree_add_95_22_pad_groupi_n_534 ,csa_tree_add_95_22_pad_groupi_n_643);
  or csa_tree_add_95_22_pad_groupi_g5003(csa_tree_add_95_22_pad_groupi_n_743 ,csa_tree_add_95_22_pad_groupi_n_481 ,csa_tree_add_95_22_pad_groupi_n_629);
  or csa_tree_add_95_22_pad_groupi_g5004(csa_tree_add_95_22_pad_groupi_n_742 ,csa_tree_add_95_22_pad_groupi_n_536 ,csa_tree_add_95_22_pad_groupi_n_650);
  or csa_tree_add_95_22_pad_groupi_g5006(csa_tree_add_95_22_pad_groupi_n_739 ,csa_tree_add_95_22_pad_groupi_n_564 ,csa_tree_add_95_22_pad_groupi_n_628);
  or csa_tree_add_95_22_pad_groupi_g5007(csa_tree_add_95_22_pad_groupi_n_737 ,csa_tree_add_95_22_pad_groupi_n_513 ,csa_tree_add_95_22_pad_groupi_n_603);
  or csa_tree_add_95_22_pad_groupi_g5008(csa_tree_add_95_22_pad_groupi_n_735 ,csa_tree_add_95_22_pad_groupi_n_553 ,csa_tree_add_95_22_pad_groupi_n_691);
  or csa_tree_add_95_22_pad_groupi_g5009(csa_tree_add_95_22_pad_groupi_n_733 ,csa_tree_add_95_22_pad_groupi_n_530 ,csa_tree_add_95_22_pad_groupi_n_622);
  or csa_tree_add_95_22_pad_groupi_g5010(csa_tree_add_95_22_pad_groupi_n_731 ,csa_tree_add_95_22_pad_groupi_n_463 ,csa_tree_add_95_22_pad_groupi_n_590);
  or csa_tree_add_95_22_pad_groupi_g5011(csa_tree_add_95_22_pad_groupi_n_729 ,csa_tree_add_95_22_pad_groupi_n_471 ,csa_tree_add_95_22_pad_groupi_n_610);
  or csa_tree_add_95_22_pad_groupi_g5012(csa_tree_add_95_22_pad_groupi_n_728 ,csa_tree_add_95_22_pad_groupi_n_520 ,csa_tree_add_95_22_pad_groupi_n_639);
  or csa_tree_add_95_22_pad_groupi_g5013(csa_tree_add_95_22_pad_groupi_n_726 ,csa_tree_add_95_22_pad_groupi_n_535 ,csa_tree_add_95_22_pad_groupi_n_690);
  or csa_tree_add_95_22_pad_groupi_g5014(csa_tree_add_95_22_pad_groupi_n_725 ,csa_tree_add_95_22_pad_groupi_n_538 ,csa_tree_add_95_22_pad_groupi_n_675);
  or csa_tree_add_95_22_pad_groupi_g5015(csa_tree_add_95_22_pad_groupi_n_723 ,csa_tree_add_95_22_pad_groupi_n_543 ,csa_tree_add_95_22_pad_groupi_n_676);
  or csa_tree_add_95_22_pad_groupi_g5016(csa_tree_add_95_22_pad_groupi_n_721 ,csa_tree_add_95_22_pad_groupi_n_542 ,csa_tree_add_95_22_pad_groupi_n_634);
  or csa_tree_add_95_22_pad_groupi_g5017(csa_tree_add_95_22_pad_groupi_n_720 ,csa_tree_add_95_22_pad_groupi_n_479 ,csa_tree_add_95_22_pad_groupi_n_644);
  or csa_tree_add_95_22_pad_groupi_g5018(csa_tree_add_95_22_pad_groupi_n_719 ,csa_tree_add_95_22_pad_groupi_n_521 ,csa_tree_add_95_22_pad_groupi_n_611);
  or csa_tree_add_95_22_pad_groupi_g5019(csa_tree_add_95_22_pad_groupi_n_718 ,csa_tree_add_95_22_pad_groupi_n_489 ,csa_tree_add_95_22_pad_groupi_n_609);
  or csa_tree_add_95_22_pad_groupi_g5020(csa_tree_add_95_22_pad_groupi_n_717 ,csa_tree_add_95_22_pad_groupi_n_549 ,csa_tree_add_95_22_pad_groupi_n_692);
  or csa_tree_add_95_22_pad_groupi_g5021(csa_tree_add_95_22_pad_groupi_n_716 ,csa_tree_add_95_22_pad_groupi_n_465 ,csa_tree_add_95_22_pad_groupi_n_613);
  or csa_tree_add_95_22_pad_groupi_g5022(csa_tree_add_95_22_pad_groupi_n_714 ,csa_tree_add_95_22_pad_groupi_n_474 ,csa_tree_add_95_22_pad_groupi_n_657);
  or csa_tree_add_95_22_pad_groupi_g5023(csa_tree_add_95_22_pad_groupi_n_713 ,csa_tree_add_95_22_pad_groupi_n_458 ,csa_tree_add_95_22_pad_groupi_n_667);
  not csa_tree_add_95_22_pad_groupi_g5024(csa_tree_add_95_22_pad_groupi_n_707 ,csa_tree_add_95_22_pad_groupi_n_706);
  not csa_tree_add_95_22_pad_groupi_g5025(csa_tree_add_95_22_pad_groupi_n_705 ,csa_tree_add_95_22_pad_groupi_n_704);
  nor csa_tree_add_95_22_pad_groupi_g5026(csa_tree_add_95_22_pad_groupi_n_703 ,csa_tree_add_95_22_pad_groupi_n_113 ,csa_tree_add_95_22_pad_groupi_n_218);
  nor csa_tree_add_95_22_pad_groupi_g5027(csa_tree_add_95_22_pad_groupi_n_702 ,in17[9] ,csa_tree_add_95_22_pad_groupi_n_358);
  nor csa_tree_add_95_22_pad_groupi_g5029(csa_tree_add_95_22_pad_groupi_n_700 ,in17[12] ,csa_tree_add_95_22_pad_groupi_n_579);
  nor csa_tree_add_95_22_pad_groupi_g5030(csa_tree_add_95_22_pad_groupi_n_699 ,csa_tree_add_95_22_pad_groupi_n_115 ,csa_tree_add_95_22_pad_groupi_n_189);
  and csa_tree_add_95_22_pad_groupi_g5031(csa_tree_add_95_22_pad_groupi_n_698 ,in9[5] ,csa_tree_add_95_22_pad_groupi_n_172);
  nor csa_tree_add_95_22_pad_groupi_g5032(csa_tree_add_95_22_pad_groupi_n_697 ,csa_tree_add_95_22_pad_groupi_n_119 ,csa_tree_add_95_22_pad_groupi_n_38);
  nor csa_tree_add_95_22_pad_groupi_g5033(csa_tree_add_95_22_pad_groupi_n_696 ,csa_tree_add_95_22_pad_groupi_n_93 ,csa_tree_add_95_22_pad_groupi_n_66);
  and csa_tree_add_95_22_pad_groupi_g5034(csa_tree_add_95_22_pad_groupi_n_695 ,in9[2] ,csa_tree_add_95_22_pad_groupi_n_133);
  and csa_tree_add_95_22_pad_groupi_g5035(csa_tree_add_95_22_pad_groupi_n_694 ,in9[10] ,csa_tree_add_95_22_pad_groupi_n_433);
  and csa_tree_add_95_22_pad_groupi_g5036(csa_tree_add_95_22_pad_groupi_n_693 ,in9[8] ,csa_tree_add_95_22_pad_groupi_n_287);
  and csa_tree_add_95_22_pad_groupi_g5037(csa_tree_add_95_22_pad_groupi_n_692 ,in9[14] ,csa_tree_add_95_22_pad_groupi_n_169);
  and csa_tree_add_95_22_pad_groupi_g5038(csa_tree_add_95_22_pad_groupi_n_691 ,in9[1] ,csa_tree_add_95_22_pad_groupi_n_168);
  and csa_tree_add_95_22_pad_groupi_g5039(csa_tree_add_95_22_pad_groupi_n_690 ,in9[5] ,csa_tree_add_95_22_pad_groupi_n_142);
  and csa_tree_add_95_22_pad_groupi_g5040(csa_tree_add_95_22_pad_groupi_n_689 ,in9[7] ,csa_tree_add_95_22_pad_groupi_n_126);
  and csa_tree_add_95_22_pad_groupi_g5041(csa_tree_add_95_22_pad_groupi_n_688 ,in9[11] ,csa_tree_add_95_22_pad_groupi_n_285);
  or csa_tree_add_95_22_pad_groupi_g5044(csa_tree_add_95_22_pad_groupi_n_685 ,csa_tree_add_95_22_pad_groupi_n_17 ,csa_tree_add_95_22_pad_groupi_n_118);
  or csa_tree_add_95_22_pad_groupi_g5046(csa_tree_add_95_22_pad_groupi_n_683 ,csa_tree_add_95_22_pad_groupi_n_149 ,csa_tree_add_95_22_pad_groupi_n_583);
  and csa_tree_add_95_22_pad_groupi_g5047(csa_tree_add_95_22_pad_groupi_n_682 ,in17[12] ,csa_tree_add_95_22_pad_groupi_n_579);
  and csa_tree_add_95_22_pad_groupi_g5048(csa_tree_add_95_22_pad_groupi_n_681 ,in9[11] ,csa_tree_add_95_22_pad_groupi_n_135);
  and csa_tree_add_95_22_pad_groupi_g5049(csa_tree_add_95_22_pad_groupi_n_680 ,in9[6] ,csa_tree_add_95_22_pad_groupi_n_445);
  nor csa_tree_add_95_22_pad_groupi_g5050(csa_tree_add_95_22_pad_groupi_n_679 ,csa_tree_add_95_22_pad_groupi_n_252 ,csa_tree_add_95_22_pad_groupi_n_223);
  and csa_tree_add_95_22_pad_groupi_g5052(csa_tree_add_95_22_pad_groupi_n_677 ,in9[3] ,csa_tree_add_95_22_pad_groupi_n_139);
  and csa_tree_add_95_22_pad_groupi_g5053(csa_tree_add_95_22_pad_groupi_n_676 ,in9[6] ,csa_tree_add_95_22_pad_groupi_n_136);
  and csa_tree_add_95_22_pad_groupi_g5054(csa_tree_add_95_22_pad_groupi_n_675 ,in9[4] ,csa_tree_add_95_22_pad_groupi_n_144);
  and csa_tree_add_95_22_pad_groupi_g5055(csa_tree_add_95_22_pad_groupi_n_674 ,in9[4] ,csa_tree_add_95_22_pad_groupi_n_138);
  nor csa_tree_add_95_22_pad_groupi_g5056(csa_tree_add_95_22_pad_groupi_n_673 ,csa_tree_add_95_22_pad_groupi_n_369 ,csa_tree_add_95_22_pad_groupi_n_581);
  and csa_tree_add_95_22_pad_groupi_g5057(csa_tree_add_95_22_pad_groupi_n_672 ,in9[12] ,csa_tree_add_95_22_pad_groupi_n_428);
  and csa_tree_add_95_22_pad_groupi_g5058(csa_tree_add_95_22_pad_groupi_n_671 ,in9[4] ,csa_tree_add_95_22_pad_groupi_n_124);
  and csa_tree_add_95_22_pad_groupi_g5059(csa_tree_add_95_22_pad_groupi_n_670 ,in9[9] ,csa_tree_add_95_22_pad_groupi_n_439);
  and csa_tree_add_95_22_pad_groupi_g5060(csa_tree_add_95_22_pad_groupi_n_669 ,in9[14] ,csa_tree_add_95_22_pad_groupi_n_288);
  and csa_tree_add_95_22_pad_groupi_g5062(csa_tree_add_95_22_pad_groupi_n_667 ,in9[14] ,csa_tree_add_95_22_pad_groupi_n_425);
  and csa_tree_add_95_22_pad_groupi_g5063(csa_tree_add_95_22_pad_groupi_n_666 ,in17[12] ,csa_tree_add_95_22_pad_groupi_n_280);
  and csa_tree_add_95_22_pad_groupi_g5064(csa_tree_add_95_22_pad_groupi_n_665 ,in9[7] ,csa_tree_add_95_22_pad_groupi_n_171);
  and csa_tree_add_95_22_pad_groupi_g5066(csa_tree_add_95_22_pad_groupi_n_663 ,csa_tree_add_95_22_pad_groupi_n_406 ,csa_tree_add_95_22_pad_groupi_n_583);
  and csa_tree_add_95_22_pad_groupi_g5067(csa_tree_add_95_22_pad_groupi_n_662 ,in9[7] ,csa_tree_add_95_22_pad_groupi_n_429);
  and csa_tree_add_95_22_pad_groupi_g5068(csa_tree_add_95_22_pad_groupi_n_661 ,in9[9] ,csa_tree_add_95_22_pad_groupi_n_145);
  and csa_tree_add_95_22_pad_groupi_g5069(csa_tree_add_95_22_pad_groupi_n_660 ,in9[14] ,csa_tree_add_95_22_pad_groupi_n_127);
  nor csa_tree_add_95_22_pad_groupi_g5070(csa_tree_add_95_22_pad_groupi_n_659 ,csa_tree_add_95_22_pad_groupi_n_112 ,csa_tree_add_95_22_pad_groupi_n_202);
  and csa_tree_add_95_22_pad_groupi_g5071(csa_tree_add_95_22_pad_groupi_n_658 ,in9[3] ,csa_tree_add_95_22_pad_groupi_n_133);
  nor csa_tree_add_95_22_pad_groupi_g5072(csa_tree_add_95_22_pad_groupi_n_657 ,csa_tree_add_95_22_pad_groupi_n_118 ,csa_tree_add_95_22_pad_groupi_n_215);
  or csa_tree_add_95_22_pad_groupi_g5073(csa_tree_add_95_22_pad_groupi_n_656 ,csa_tree_add_95_22_pad_groupi_n_373 ,csa_tree_add_95_22_pad_groupi_n_357);
  or csa_tree_add_95_22_pad_groupi_g5074(csa_tree_add_95_22_pad_groupi_n_655 ,csa_tree_add_95_22_pad_groupi_n_27 ,csa_tree_add_95_22_pad_groupi_n_427);
  and csa_tree_add_95_22_pad_groupi_g5075(csa_tree_add_95_22_pad_groupi_n_654 ,in9[11] ,csa_tree_add_95_22_pad_groupi_n_130);
  and csa_tree_add_95_22_pad_groupi_g5076(csa_tree_add_95_22_pad_groupi_n_653 ,in9[1] ,csa_tree_add_95_22_pad_groupi_n_147);
  nor csa_tree_add_95_22_pad_groupi_g5077(csa_tree_add_95_22_pad_groupi_n_652 ,csa_tree_add_95_22_pad_groupi_n_93 ,csa_tree_add_95_22_pad_groupi_n_74);
  and csa_tree_add_95_22_pad_groupi_g5078(csa_tree_add_95_22_pad_groupi_n_651 ,in9[13] ,csa_tree_add_95_22_pad_groupi_n_148);
  and csa_tree_add_95_22_pad_groupi_g5079(csa_tree_add_95_22_pad_groupi_n_650 ,in9[6] ,csa_tree_add_95_22_pad_groupi_n_148);
  and csa_tree_add_95_22_pad_groupi_g5080(csa_tree_add_95_22_pad_groupi_n_649 ,in9[12] ,csa_tree_add_95_22_pad_groupi_n_142);
  and csa_tree_add_95_22_pad_groupi_g5081(csa_tree_add_95_22_pad_groupi_n_648 ,in9[3] ,csa_tree_add_95_22_pad_groupi_n_129);
  and csa_tree_add_95_22_pad_groupi_g5082(csa_tree_add_95_22_pad_groupi_n_647 ,in9[4] ,csa_tree_add_95_22_pad_groupi_n_284);
  or csa_tree_add_95_22_pad_groupi_g5084(csa_tree_add_95_22_pad_groupi_n_706 ,csa_tree_add_95_22_pad_groupi_n_24 ,csa_tree_add_95_22_pad_groupi_n_502);
  or csa_tree_add_95_22_pad_groupi_g5085(csa_tree_add_95_22_pad_groupi_n_704 ,csa_tree_add_95_22_pad_groupi_n_24 ,csa_tree_add_95_22_pad_groupi_n_257);
  nor csa_tree_add_95_22_pad_groupi_g5086(csa_tree_add_95_22_pad_groupi_n_644 ,csa_tree_add_95_22_pad_groupi_n_113 ,csa_tree_add_95_22_pad_groupi_n_178);
  nor csa_tree_add_95_22_pad_groupi_g5087(csa_tree_add_95_22_pad_groupi_n_643 ,csa_tree_add_95_22_pad_groupi_n_160 ,csa_tree_add_95_22_pad_groupi_n_578);
  or csa_tree_add_95_22_pad_groupi_g5088(csa_tree_add_95_22_pad_groupi_n_642 ,csa_tree_add_95_22_pad_groupi_n_47 ,csa_tree_add_95_22_pad_groupi_n_497);
  and csa_tree_add_95_22_pad_groupi_g5090(csa_tree_add_95_22_pad_groupi_n_640 ,in9[6] ,csa_tree_add_95_22_pad_groupi_n_130);
  and csa_tree_add_95_22_pad_groupi_g5091(csa_tree_add_95_22_pad_groupi_n_639 ,in9[13] ,csa_tree_add_95_22_pad_groupi_n_171);
  nor csa_tree_add_95_22_pad_groupi_g5092(csa_tree_add_95_22_pad_groupi_n_638 ,csa_tree_add_95_22_pad_groupi_n_87 ,csa_tree_add_95_22_pad_groupi_n_434);
  and csa_tree_add_95_22_pad_groupi_g5093(csa_tree_add_95_22_pad_groupi_n_637 ,in9[10] ,csa_tree_add_95_22_pad_groupi_n_166);
  nor csa_tree_add_95_22_pad_groupi_g5095(csa_tree_add_95_22_pad_groupi_n_635 ,csa_tree_add_95_22_pad_groupi_n_96 ,csa_tree_add_95_22_pad_groupi_n_255);
  and csa_tree_add_95_22_pad_groupi_g5096(csa_tree_add_95_22_pad_groupi_n_634 ,in9[2] ,csa_tree_add_95_22_pad_groupi_n_168);
  and csa_tree_add_95_22_pad_groupi_g5097(csa_tree_add_95_22_pad_groupi_n_633 ,in9[13] ,csa_tree_add_95_22_pad_groupi_n_124);
  nor csa_tree_add_95_22_pad_groupi_g5099(csa_tree_add_95_22_pad_groupi_n_631 ,csa_tree_add_95_22_pad_groupi_n_231 ,csa_tree_add_95_22_pad_groupi_n_257);
  and csa_tree_add_95_22_pad_groupi_g5101(csa_tree_add_95_22_pad_groupi_n_629 ,in9[13] ,csa_tree_add_95_22_pad_groupi_n_287);
  and csa_tree_add_95_22_pad_groupi_g5102(csa_tree_add_95_22_pad_groupi_n_628 ,in9[11] ,csa_tree_add_95_22_pad_groupi_n_145);
  and csa_tree_add_95_22_pad_groupi_g5103(csa_tree_add_95_22_pad_groupi_n_627 ,in9[7] ,csa_tree_add_95_22_pad_groupi_n_141);
  nor csa_tree_add_95_22_pad_groupi_g5104(csa_tree_add_95_22_pad_groupi_n_626 ,csa_tree_add_95_22_pad_groupi_n_71 ,csa_tree_add_95_22_pad_groupi_n_507);
  and csa_tree_add_95_22_pad_groupi_g5105(csa_tree_add_95_22_pad_groupi_n_625 ,in9[7] ,csa_tree_add_95_22_pad_groupi_n_285);
  and csa_tree_add_95_22_pad_groupi_g5106(csa_tree_add_95_22_pad_groupi_n_624 ,in9[5] ,csa_tree_add_95_22_pad_groupi_n_165);
  and csa_tree_add_95_22_pad_groupi_g5107(csa_tree_add_95_22_pad_groupi_n_623 ,in9[10] ,csa_tree_add_95_22_pad_groupi_n_132);
  nor csa_tree_add_95_22_pad_groupi_g5108(csa_tree_add_95_22_pad_groupi_n_622 ,csa_tree_add_95_22_pad_groupi_n_159 ,csa_tree_add_95_22_pad_groupi_n_282);
  nor csa_tree_add_95_22_pad_groupi_g5109(csa_tree_add_95_22_pad_groupi_n_621 ,csa_tree_add_95_22_pad_groupi_n_98 ,csa_tree_add_95_22_pad_groupi_n_430);
  nor csa_tree_add_95_22_pad_groupi_g5110(csa_tree_add_95_22_pad_groupi_n_620 ,csa_tree_add_95_22_pad_groupi_n_194 ,csa_tree_add_95_22_pad_groupi_n_502);
  nor csa_tree_add_95_22_pad_groupi_g5111(csa_tree_add_95_22_pad_groupi_n_619 ,csa_tree_add_95_22_pad_groupi_n_116 ,csa_tree_add_95_22_pad_groupi_n_187);
  and csa_tree_add_95_22_pad_groupi_g5112(csa_tree_add_95_22_pad_groupi_n_618 ,in9[8] ,csa_tree_add_95_22_pad_groupi_n_165);
  and csa_tree_add_95_22_pad_groupi_g5113(csa_tree_add_95_22_pad_groupi_n_617 ,in9[8] ,csa_tree_add_95_22_pad_groupi_n_136);
  nor csa_tree_add_95_22_pad_groupi_g5114(csa_tree_add_95_22_pad_groupi_n_616 ,csa_tree_add_95_22_pad_groupi_n_119 ,csa_tree_add_95_22_pad_groupi_n_181);
  nor csa_tree_add_95_22_pad_groupi_g5117(csa_tree_add_95_22_pad_groupi_n_613 ,csa_tree_add_95_22_pad_groupi_n_204 ,csa_tree_add_95_22_pad_groupi_n_432);
  or csa_tree_add_95_22_pad_groupi_g5118(csa_tree_add_95_22_pad_groupi_n_612 ,csa_tree_add_95_22_pad_groupi_n_64 ,csa_tree_add_95_22_pad_groupi_n_438);
  and csa_tree_add_95_22_pad_groupi_g5119(csa_tree_add_95_22_pad_groupi_n_611 ,in9[8] ,csa_tree_add_95_22_pad_groupi_n_284);
  nor csa_tree_add_95_22_pad_groupi_g5120(csa_tree_add_95_22_pad_groupi_n_610 ,csa_tree_add_95_22_pad_groupi_n_116 ,csa_tree_add_95_22_pad_groupi_n_184);
  nor csa_tree_add_95_22_pad_groupi_g5121(csa_tree_add_95_22_pad_groupi_n_609 ,csa_tree_add_95_22_pad_groupi_n_91 ,csa_tree_add_95_22_pad_groupi_n_501);
  and csa_tree_add_95_22_pad_groupi_g5122(csa_tree_add_95_22_pad_groupi_n_608 ,in9[12] ,csa_tree_add_95_22_pad_groupi_n_166);
  and csa_tree_add_95_22_pad_groupi_g5123(csa_tree_add_95_22_pad_groupi_n_607 ,in9[11] ,csa_tree_add_95_22_pad_groupi_n_431);
  or csa_tree_add_95_22_pad_groupi_g5124(csa_tree_add_95_22_pad_groupi_n_606 ,csa_tree_add_95_22_pad_groupi_n_17 ,csa_tree_add_95_22_pad_groupi_n_255);
  and csa_tree_add_95_22_pad_groupi_g5125(csa_tree_add_95_22_pad_groupi_n_605 ,in9[9] ,csa_tree_add_95_22_pad_groupi_n_127);
  nor csa_tree_add_95_22_pad_groupi_g5126(csa_tree_add_95_22_pad_groupi_n_604 ,csa_tree_add_95_22_pad_groupi_n_211 ,csa_tree_add_95_22_pad_groupi_n_508);
  and csa_tree_add_95_22_pad_groupi_g5127(csa_tree_add_95_22_pad_groupi_n_603 ,in9[12] ,csa_tree_add_95_22_pad_groupi_n_169);
  and csa_tree_add_95_22_pad_groupi_g5128(csa_tree_add_95_22_pad_groupi_n_602 ,in9[1] ,csa_tree_add_95_22_pad_groupi_n_123);
  nor csa_tree_add_95_22_pad_groupi_g5130(csa_tree_add_95_22_pad_groupi_n_600 ,in17[12] ,csa_tree_add_95_22_pad_groupi_n_582);
  and csa_tree_add_95_22_pad_groupi_g5131(csa_tree_add_95_22_pad_groupi_n_599 ,in9[9] ,csa_tree_add_95_22_pad_groupi_n_139);
  nor csa_tree_add_95_22_pad_groupi_g5132(csa_tree_add_95_22_pad_groupi_n_598 ,csa_tree_add_95_22_pad_groupi_n_101 ,csa_tree_add_95_22_pad_groupi_n_508);
  or csa_tree_add_95_22_pad_groupi_g5135(csa_tree_add_95_22_pad_groupi_n_595 ,csa_tree_add_95_22_pad_groupi_n_55 ,csa_tree_add_95_22_pad_groupi_n_115);
  or csa_tree_add_95_22_pad_groupi_g5136(csa_tree_add_95_22_pad_groupi_n_594 ,csa_tree_add_95_22_pad_groupi_n_50 ,csa_tree_add_95_22_pad_groupi_n_426);
  nor csa_tree_add_95_22_pad_groupi_g5137(csa_tree_add_95_22_pad_groupi_n_593 ,in17[11] ,csa_tree_add_95_22_pad_groupi_n_580);
  and csa_tree_add_95_22_pad_groupi_g5139(csa_tree_add_95_22_pad_groupi_n_591 ,in9[10] ,csa_tree_add_95_22_pad_groupi_n_288);
  and csa_tree_add_95_22_pad_groupi_g5140(csa_tree_add_95_22_pad_groupi_n_590 ,in9[13] ,csa_tree_add_95_22_pad_groupi_n_435);
  and csa_tree_add_95_22_pad_groupi_g5141(csa_tree_add_95_22_pad_groupi_n_589 ,in9[10] ,csa_tree_add_95_22_pad_groupi_n_172);
  nor csa_tree_add_95_22_pad_groupi_g5142(csa_tree_add_95_22_pad_groupi_n_588 ,csa_tree_add_95_22_pad_groupi_n_158 ,csa_tree_add_95_22_pad_groupi_n_280);
  or csa_tree_add_95_22_pad_groupi_g5143(csa_tree_add_95_22_pad_groupi_n_587 ,csa_tree_add_95_22_pad_groupi_n_151 ,csa_tree_add_95_22_pad_groupi_n_580);
  or csa_tree_add_95_22_pad_groupi_g5144(csa_tree_add_95_22_pad_groupi_n_586 ,csa_tree_add_95_22_pad_groupi_n_15 ,csa_tree_add_95_22_pad_groupi_n_581);
  or csa_tree_add_95_22_pad_groupi_g5145(csa_tree_add_95_22_pad_groupi_n_646 ,csa_tree_add_95_22_pad_groupi_n_57 ,csa_tree_add_95_22_pad_groupi_n_493);
  or csa_tree_add_95_22_pad_groupi_g5146(csa_tree_add_95_22_pad_groupi_n_645 ,csa_tree_add_95_22_pad_groupi_n_42 ,csa_tree_add_95_22_pad_groupi_n_278);
  nor csa_tree_add_95_22_pad_groupi_g5150(csa_tree_add_95_22_pad_groupi_n_577 ,csa_tree_add_95_22_pad_groupi_n_183 ,csa_tree_add_95_22_pad_groupi_n_332);
  nor csa_tree_add_95_22_pad_groupi_g5151(csa_tree_add_95_22_pad_groupi_n_576 ,csa_tree_add_95_22_pad_groupi_n_42 ,csa_tree_add_95_22_pad_groupi_n_302);
  nor csa_tree_add_95_22_pad_groupi_g5152(csa_tree_add_95_22_pad_groupi_n_575 ,csa_tree_add_95_22_pad_groupi_n_233 ,csa_tree_add_95_22_pad_groupi_n_306);
  nor csa_tree_add_95_22_pad_groupi_g5153(csa_tree_add_95_22_pad_groupi_n_574 ,csa_tree_add_95_22_pad_groupi_n_193 ,csa_tree_add_95_22_pad_groupi_n_341);
  nor csa_tree_add_95_22_pad_groupi_g5154(csa_tree_add_95_22_pad_groupi_n_573 ,csa_tree_add_95_22_pad_groupi_n_84 ,csa_tree_add_95_22_pad_groupi_n_312);
  nor csa_tree_add_95_22_pad_groupi_g5163(csa_tree_add_95_22_pad_groupi_n_564 ,csa_tree_add_95_22_pad_groupi_n_78 ,csa_tree_add_95_22_pad_groupi_n_330);
  nor csa_tree_add_95_22_pad_groupi_g5170(csa_tree_add_95_22_pad_groupi_n_557 ,csa_tree_add_95_22_pad_groupi_n_71 ,csa_tree_add_95_22_pad_groupi_n_335);
  nor csa_tree_add_95_22_pad_groupi_g5171(csa_tree_add_95_22_pad_groupi_n_556 ,csa_tree_add_95_22_pad_groupi_n_101 ,csa_tree_add_95_22_pad_groupi_n_315);
  nor csa_tree_add_95_22_pad_groupi_g5172(csa_tree_add_95_22_pad_groupi_n_555 ,csa_tree_add_95_22_pad_groupi_n_186 ,csa_tree_add_95_22_pad_groupi_n_336);
  nor csa_tree_add_95_22_pad_groupi_g5173(csa_tree_add_95_22_pad_groupi_n_554 ,csa_tree_add_95_22_pad_groupi_n_177 ,csa_tree_add_95_22_pad_groupi_n_309);
  nor csa_tree_add_95_22_pad_groupi_g5174(csa_tree_add_95_22_pad_groupi_n_553 ,csa_tree_add_95_22_pad_groupi_n_244 ,csa_tree_add_95_22_pad_groupi_n_320);
  nor csa_tree_add_95_22_pad_groupi_g5175(csa_tree_add_95_22_pad_groupi_n_552 ,csa_tree_add_95_22_pad_groupi_n_247 ,csa_tree_add_95_22_pad_groupi_n_323);
  nor csa_tree_add_95_22_pad_groupi_g5176(csa_tree_add_95_22_pad_groupi_n_551 ,csa_tree_add_95_22_pad_groupi_n_67 ,csa_tree_add_95_22_pad_groupi_n_317);
  nor csa_tree_add_95_22_pad_groupi_g5177(csa_tree_add_95_22_pad_groupi_n_550 ,csa_tree_add_95_22_pad_groupi_n_175 ,csa_tree_add_95_22_pad_groupi_n_339);
  nor csa_tree_add_95_22_pad_groupi_g5178(csa_tree_add_95_22_pad_groupi_n_549 ,csa_tree_add_95_22_pad_groupi_n_85 ,csa_tree_add_95_22_pad_groupi_n_321);
  nor csa_tree_add_95_22_pad_groupi_g5179(csa_tree_add_95_22_pad_groupi_n_548 ,csa_tree_add_95_22_pad_groupi_n_88 ,csa_tree_add_95_22_pad_groupi_n_305);
  nor csa_tree_add_95_22_pad_groupi_g5180(csa_tree_add_95_22_pad_groupi_n_547 ,csa_tree_add_95_22_pad_groupi_n_197 ,csa_tree_add_95_22_pad_groupi_n_323);
  nor csa_tree_add_95_22_pad_groupi_g5181(csa_tree_add_95_22_pad_groupi_n_546 ,csa_tree_add_95_22_pad_groupi_n_100 ,csa_tree_add_95_22_pad_groupi_n_326);
  nor csa_tree_add_95_22_pad_groupi_g5182(csa_tree_add_95_22_pad_groupi_n_545 ,csa_tree_add_95_22_pad_groupi_n_53 ,csa_tree_add_95_22_pad_groupi_n_327);
  nor csa_tree_add_95_22_pad_groupi_g5183(csa_tree_add_95_22_pad_groupi_n_544 ,csa_tree_add_95_22_pad_groupi_n_187 ,csa_tree_add_95_22_pad_groupi_n_326);
  nor csa_tree_add_95_22_pad_groupi_g5184(csa_tree_add_95_22_pad_groupi_n_543 ,csa_tree_add_95_22_pad_groupi_n_196 ,csa_tree_add_95_22_pad_groupi_n_317);
  nor csa_tree_add_95_22_pad_groupi_g5185(csa_tree_add_95_22_pad_groupi_n_542 ,csa_tree_add_95_22_pad_groupi_n_217 ,csa_tree_add_95_22_pad_groupi_n_318);
  nor csa_tree_add_95_22_pad_groupi_g5186(csa_tree_add_95_22_pad_groupi_n_541 ,csa_tree_add_95_22_pad_groupi_n_209 ,csa_tree_add_95_22_pad_groupi_n_344);
  nor csa_tree_add_95_22_pad_groupi_g5187(csa_tree_add_95_22_pad_groupi_n_540 ,csa_tree_add_95_22_pad_groupi_n_229 ,csa_tree_add_95_22_pad_groupi_n_324);
  nor csa_tree_add_95_22_pad_groupi_g5188(csa_tree_add_95_22_pad_groupi_n_539 ,csa_tree_add_95_22_pad_groupi_n_41 ,csa_tree_add_95_22_pad_groupi_n_335);
  nor csa_tree_add_95_22_pad_groupi_g5189(csa_tree_add_95_22_pad_groupi_n_538 ,csa_tree_add_95_22_pad_groupi_n_36 ,csa_tree_add_95_22_pad_groupi_n_336);
  nor csa_tree_add_95_22_pad_groupi_g5190(csa_tree_add_95_22_pad_groupi_n_537 ,csa_tree_add_95_22_pad_groupi_n_79 ,csa_tree_add_95_22_pad_groupi_n_324);
  nor csa_tree_add_95_22_pad_groupi_g5191(csa_tree_add_95_22_pad_groupi_n_536 ,csa_tree_add_95_22_pad_groupi_n_204 ,csa_tree_add_95_22_pad_groupi_n_345);
  nor csa_tree_add_95_22_pad_groupi_g5192(csa_tree_add_95_22_pad_groupi_n_535 ,csa_tree_add_95_22_pad_groupi_n_28 ,csa_tree_add_95_22_pad_groupi_n_329);
  nor csa_tree_add_95_22_pad_groupi_g5193(csa_tree_add_95_22_pad_groupi_n_534 ,csa_tree_add_95_22_pad_groupi_n_194 ,csa_tree_add_95_22_pad_groupi_n_327);
  nor csa_tree_add_95_22_pad_groupi_g5194(csa_tree_add_95_22_pad_groupi_n_533 ,csa_tree_add_95_22_pad_groupi_n_191 ,csa_tree_add_95_22_pad_groupi_n_338);
  nor csa_tree_add_95_22_pad_groupi_g5195(csa_tree_add_95_22_pad_groupi_n_532 ,csa_tree_add_95_22_pad_groupi_n_184 ,csa_tree_add_95_22_pad_groupi_n_318);
  or csa_tree_add_95_22_pad_groupi_g5196(csa_tree_add_95_22_pad_groupi_n_531 ,csa_tree_add_95_22_pad_groupi_n_174 ,csa_tree_add_95_22_pad_groupi_n_305);
  nor csa_tree_add_95_22_pad_groupi_g5197(csa_tree_add_95_22_pad_groupi_n_530 ,csa_tree_add_95_22_pad_groupi_n_39 ,csa_tree_add_95_22_pad_groupi_n_330);
  nor csa_tree_add_95_22_pad_groupi_g5198(csa_tree_add_95_22_pad_groupi_n_529 ,csa_tree_add_95_22_pad_groupi_n_243 ,csa_tree_add_95_22_pad_groupi_n_344);
  nor csa_tree_add_95_22_pad_groupi_g5199(csa_tree_add_95_22_pad_groupi_n_528 ,csa_tree_add_95_22_pad_groupi_n_91 ,csa_tree_add_95_22_pad_groupi_n_345);
  nor csa_tree_add_95_22_pad_groupi_g5200(csa_tree_add_95_22_pad_groupi_n_527 ,csa_tree_add_95_22_pad_groupi_n_231 ,csa_tree_add_95_22_pad_groupi_n_321);
  nor csa_tree_add_95_22_pad_groupi_g5201(csa_tree_add_95_22_pad_groupi_n_526 ,csa_tree_add_95_22_pad_groupi_n_217 ,csa_tree_add_95_22_pad_groupi_n_265);
  nor csa_tree_add_95_22_pad_groupi_g5202(csa_tree_add_95_22_pad_groupi_n_525 ,csa_tree_add_95_22_pad_groupi_n_64 ,csa_tree_add_95_22_pad_groupi_n_311);
  nor csa_tree_add_95_22_pad_groupi_g5203(csa_tree_add_95_22_pad_groupi_n_524 ,csa_tree_add_95_22_pad_groupi_n_55 ,csa_tree_add_95_22_pad_groupi_n_269);
  nor csa_tree_add_95_22_pad_groupi_g5204(csa_tree_add_95_22_pad_groupi_n_523 ,csa_tree_add_95_22_pad_groupi_n_76 ,csa_tree_add_95_22_pad_groupi_n_312);
  nor csa_tree_add_95_22_pad_groupi_g5205(csa_tree_add_95_22_pad_groupi_n_522 ,csa_tree_add_95_22_pad_groupi_n_201 ,csa_tree_add_95_22_pad_groupi_n_339);
  nor csa_tree_add_95_22_pad_groupi_g5206(csa_tree_add_95_22_pad_groupi_n_521 ,csa_tree_add_95_22_pad_groupi_n_22 ,csa_tree_add_95_22_pad_groupi_n_275);
  nor csa_tree_add_95_22_pad_groupi_g5207(csa_tree_add_95_22_pad_groupi_n_520 ,csa_tree_add_95_22_pad_groupi_n_222 ,csa_tree_add_95_22_pad_groupi_n_262);
  nor csa_tree_add_95_22_pad_groupi_g5208(csa_tree_add_95_22_pad_groupi_n_519 ,csa_tree_add_95_22_pad_groupi_n_50 ,csa_tree_add_95_22_pad_groupi_n_272);
  or csa_tree_add_95_22_pad_groupi_g5209(csa_tree_add_95_22_pad_groupi_n_518 ,csa_tree_add_95_22_pad_groupi_n_21 ,csa_tree_add_95_22_pad_groupi_n_266);
  nor csa_tree_add_95_22_pad_groupi_g5210(csa_tree_add_95_22_pad_groupi_n_517 ,csa_tree_add_95_22_pad_groupi_n_178 ,csa_tree_add_95_22_pad_groupi_n_274);
  nor csa_tree_add_95_22_pad_groupi_g5211(csa_tree_add_95_22_pad_groupi_n_516 ,csa_tree_add_95_22_pad_groupi_n_225 ,csa_tree_add_95_22_pad_groupi_n_263);
  nor csa_tree_add_95_22_pad_groupi_g5212(csa_tree_add_95_22_pad_groupi_n_515 ,csa_tree_add_95_22_pad_groupi_n_47 ,csa_tree_add_95_22_pad_groupi_n_268);
  nor csa_tree_add_95_22_pad_groupi_g5213(csa_tree_add_95_22_pad_groupi_n_514 ,csa_tree_add_95_22_pad_groupi_n_197 ,csa_tree_add_95_22_pad_groupi_n_333);
  nor csa_tree_add_95_22_pad_groupi_g5214(csa_tree_add_95_22_pad_groupi_n_513 ,csa_tree_add_95_22_pad_groupi_n_227 ,csa_tree_add_95_22_pad_groupi_n_320);
  nor csa_tree_add_95_22_pad_groupi_g5215(csa_tree_add_95_22_pad_groupi_n_512 ,csa_tree_add_95_22_pad_groupi_n_59 ,csa_tree_add_95_22_pad_groupi_n_342);
  or csa_tree_add_95_22_pad_groupi_g5217(csa_tree_add_95_22_pad_groupi_n_583 ,csa_tree_add_95_22_pad_groupi_n_121 ,csa_tree_add_95_22_pad_groupi_n_424);
  or csa_tree_add_95_22_pad_groupi_g5218(csa_tree_add_95_22_pad_groupi_n_582 ,csa_tree_add_95_22_pad_groupi_n_162 ,csa_tree_add_95_22_pad_groupi_n_402);
  or csa_tree_add_95_22_pad_groupi_g5219(csa_tree_add_95_22_pad_groupi_n_581 ,csa_tree_add_95_22_pad_groupi_n_121 ,csa_tree_add_95_22_pad_groupi_n_109);
  or csa_tree_add_95_22_pad_groupi_g5220(csa_tree_add_95_22_pad_groupi_n_580 ,csa_tree_add_95_22_pad_groupi_n_162 ,csa_tree_add_95_22_pad_groupi_n_404);
  or csa_tree_add_95_22_pad_groupi_g5221(csa_tree_add_95_22_pad_groupi_n_579 ,csa_tree_add_95_22_pad_groupi_n_163 ,csa_tree_add_95_22_pad_groupi_n_403);
  not csa_tree_add_95_22_pad_groupi_g5223(csa_tree_add_95_22_pad_groupi_n_510 ,csa_tree_add_95_22_pad_groupi_n_505);
  not csa_tree_add_95_22_pad_groupi_g5224(csa_tree_add_95_22_pad_groupi_n_509 ,csa_tree_add_95_22_pad_groupi_n_505);
  not csa_tree_add_95_22_pad_groupi_g5225(csa_tree_add_95_22_pad_groupi_n_508 ,csa_tree_add_95_22_pad_groupi_n_506);
  not csa_tree_add_95_22_pad_groupi_g5226(csa_tree_add_95_22_pad_groupi_n_507 ,csa_tree_add_95_22_pad_groupi_n_506);
  not csa_tree_add_95_22_pad_groupi_g5227(csa_tree_add_95_22_pad_groupi_n_506 ,csa_tree_add_95_22_pad_groupi_n_505);
  not csa_tree_add_95_22_pad_groupi_g5228(csa_tree_add_95_22_pad_groupi_n_504 ,csa_tree_add_95_22_pad_groupi_n_499);
  not csa_tree_add_95_22_pad_groupi_g5229(csa_tree_add_95_22_pad_groupi_n_503 ,csa_tree_add_95_22_pad_groupi_n_499);
  not csa_tree_add_95_22_pad_groupi_g5230(csa_tree_add_95_22_pad_groupi_n_502 ,csa_tree_add_95_22_pad_groupi_n_500);
  not csa_tree_add_95_22_pad_groupi_g5231(csa_tree_add_95_22_pad_groupi_n_501 ,csa_tree_add_95_22_pad_groupi_n_500);
  not csa_tree_add_95_22_pad_groupi_g5232(csa_tree_add_95_22_pad_groupi_n_500 ,csa_tree_add_95_22_pad_groupi_n_499);
  not csa_tree_add_95_22_pad_groupi_g5233(csa_tree_add_95_22_pad_groupi_n_498 ,csa_tree_add_95_22_pad_groupi_n_278);
  not csa_tree_add_95_22_pad_groupi_g5234(csa_tree_add_95_22_pad_groupi_n_496 ,csa_tree_add_95_22_pad_groupi_n_497);
  not csa_tree_add_95_22_pad_groupi_g5235(csa_tree_add_95_22_pad_groupi_n_495 ,csa_tree_add_95_22_pad_groupi_n_493);
  not csa_tree_add_95_22_pad_groupi_g5236(csa_tree_add_95_22_pad_groupi_n_494 ,csa_tree_add_95_22_pad_groupi_n_493);
  or csa_tree_add_95_22_pad_groupi_g5237(csa_tree_add_95_22_pad_groupi_n_492 ,csa_tree_add_95_22_pad_groupi_n_27 ,csa_tree_add_95_22_pad_groupi_n_311);
  nor csa_tree_add_95_22_pad_groupi_g5238(csa_tree_add_95_22_pad_groupi_n_491 ,csa_tree_add_95_22_pad_groupi_n_180 ,csa_tree_add_95_22_pad_groupi_n_329);
  nor csa_tree_add_95_22_pad_groupi_g5239(csa_tree_add_95_22_pad_groupi_n_490 ,csa_tree_add_95_22_pad_groupi_n_220 ,csa_tree_add_95_22_pad_groupi_n_271);
  nor csa_tree_add_95_22_pad_groupi_g5240(csa_tree_add_95_22_pad_groupi_n_489 ,csa_tree_add_95_22_pad_groupi_n_82 ,csa_tree_add_95_22_pad_groupi_n_275);
  nor csa_tree_add_95_22_pad_groupi_g5241(csa_tree_add_95_22_pad_groupi_n_488 ,csa_tree_add_95_22_pad_groupi_n_181 ,csa_tree_add_95_22_pad_groupi_n_309);
  nor csa_tree_add_95_22_pad_groupi_g5242(csa_tree_add_95_22_pad_groupi_n_487 ,csa_tree_add_95_22_pad_groupi_n_88 ,csa_tree_add_95_22_pad_groupi_n_341);
  nor csa_tree_add_95_22_pad_groupi_g5243(csa_tree_add_95_22_pad_groupi_n_486 ,csa_tree_add_95_22_pad_groupi_n_227 ,csa_tree_add_95_22_pad_groupi_n_306);
  or csa_tree_add_95_22_pad_groupi_g5244(csa_tree_add_95_22_pad_groupi_n_485 ,csa_tree_add_95_22_pad_groupi_n_30 ,csa_tree_add_95_22_pad_groupi_n_302);
  nor csa_tree_add_95_22_pad_groupi_g5245(csa_tree_add_95_22_pad_groupi_n_484 ,csa_tree_add_95_22_pad_groupi_n_174 ,csa_tree_add_95_22_pad_groupi_n_315);
  or csa_tree_add_95_22_pad_groupi_g5246(csa_tree_add_95_22_pad_groupi_n_483 ,csa_tree_add_95_22_pad_groupi_n_30 ,csa_tree_add_95_22_pad_groupi_n_263);
  nor csa_tree_add_95_22_pad_groupi_g5247(csa_tree_add_95_22_pad_groupi_n_482 ,csa_tree_add_95_22_pad_groupi_n_96 ,csa_tree_add_95_22_pad_groupi_n_338);
  nor csa_tree_add_95_22_pad_groupi_g5248(csa_tree_add_95_22_pad_groupi_n_481 ,csa_tree_add_95_22_pad_groupi_n_233 ,csa_tree_add_95_22_pad_groupi_n_269);
  nor csa_tree_add_95_22_pad_groupi_g5249(csa_tree_add_95_22_pad_groupi_n_480 ,csa_tree_add_95_22_pad_groupi_n_25 ,csa_tree_add_95_22_pad_groupi_n_272);
  nor csa_tree_add_95_22_pad_groupi_g5250(csa_tree_add_95_22_pad_groupi_n_479 ,csa_tree_add_95_22_pad_groupi_n_214 ,csa_tree_add_95_22_pad_groupi_n_266);
  nor csa_tree_add_95_22_pad_groupi_g5251(csa_tree_add_95_22_pad_groupi_n_478 ,csa_tree_add_95_22_pad_groupi_n_235 ,csa_tree_add_95_22_pad_groupi_n_332);
  nor csa_tree_add_95_22_pad_groupi_g5252(csa_tree_add_95_22_pad_groupi_n_477 ,csa_tree_add_95_22_pad_groupi_n_73 ,csa_tree_add_95_22_pad_groupi_n_342);
  nor csa_tree_add_95_22_pad_groupi_g5253(csa_tree_add_95_22_pad_groupi_n_476 ,csa_tree_add_95_22_pad_groupi_n_206 ,csa_tree_add_95_22_pad_groupi_n_314);
  nor csa_tree_add_95_22_pad_groupi_g5254(csa_tree_add_95_22_pad_groupi_n_475 ,csa_tree_add_95_22_pad_groupi_n_69 ,csa_tree_add_95_22_pad_groupi_n_308);
  nor csa_tree_add_95_22_pad_groupi_g5255(csa_tree_add_95_22_pad_groupi_n_474 ,csa_tree_add_95_22_pad_groupi_n_209 ,csa_tree_add_95_22_pad_groupi_n_303);
  nor csa_tree_add_95_22_pad_groupi_g5256(csa_tree_add_95_22_pad_groupi_n_473 ,csa_tree_add_95_22_pad_groupi_n_76 ,csa_tree_add_95_22_pad_groupi_n_314);
  or csa_tree_add_95_22_pad_groupi_g5257(csa_tree_add_95_22_pad_groupi_n_472 ,csa_tree_add_95_22_pad_groupi_n_45 ,csa_tree_add_95_22_pad_groupi_n_308);
  nor csa_tree_add_95_22_pad_groupi_g5258(csa_tree_add_95_22_pad_groupi_n_471 ,csa_tree_add_95_22_pad_groupi_n_211 ,csa_tree_add_95_22_pad_groupi_n_303);
  nor csa_tree_add_95_22_pad_groupi_g5259(csa_tree_add_95_22_pad_groupi_n_470 ,csa_tree_add_95_22_pad_groupi_n_67 ,csa_tree_add_95_22_pad_groupi_n_333);
  nor csa_tree_add_95_22_pad_groupi_g5260(csa_tree_add_95_22_pad_groupi_n_469 ,csa_tree_add_95_22_pad_groupi_n_180 ,csa_tree_add_95_22_pad_groupi_n_300);
  nor csa_tree_add_95_22_pad_groupi_g5261(csa_tree_add_95_22_pad_groupi_n_468 ,csa_tree_add_95_22_pad_groupi_n_177 ,csa_tree_add_95_22_pad_groupi_n_399);
  nor csa_tree_add_95_22_pad_groupi_g5262(csa_tree_add_95_22_pad_groupi_n_467 ,csa_tree_add_95_22_pad_groupi_n_52 ,csa_tree_add_95_22_pad_groupi_n_291);
  nor csa_tree_add_95_22_pad_groupi_g5263(csa_tree_add_95_22_pad_groupi_n_466 ,csa_tree_add_95_22_pad_groupi_n_45 ,csa_tree_add_95_22_pad_groupi_n_290);
  nor csa_tree_add_95_22_pad_groupi_g5264(csa_tree_add_95_22_pad_groupi_n_465 ,csa_tree_add_95_22_pad_groupi_n_175 ,csa_tree_add_95_22_pad_groupi_n_297);
  or csa_tree_add_95_22_pad_groupi_g5265(csa_tree_add_95_22_pad_groupi_n_464 ,csa_tree_add_95_22_pad_groupi_n_36 ,csa_tree_add_95_22_pad_groupi_n_296);
  nor csa_tree_add_95_22_pad_groupi_g5266(csa_tree_add_95_22_pad_groupi_n_463 ,csa_tree_add_95_22_pad_groupi_n_90 ,csa_tree_add_95_22_pad_groupi_n_260);
  nor csa_tree_add_95_22_pad_groupi_g5267(csa_tree_add_95_22_pad_groupi_n_462 ,csa_tree_add_95_22_pad_groupi_n_212 ,csa_tree_add_95_22_pad_groupi_n_299);
  nor csa_tree_add_95_22_pad_groupi_g5268(csa_tree_add_95_22_pad_groupi_n_461 ,csa_tree_add_95_22_pad_groupi_n_95 ,csa_tree_add_95_22_pad_groupi_n_299);
  or csa_tree_add_95_22_pad_groupi_g5269(csa_tree_add_95_22_pad_groupi_n_460 ,csa_tree_add_95_22_pad_groupi_n_39 ,csa_tree_add_95_22_pad_groupi_n_290);
  nor csa_tree_add_95_22_pad_groupi_g5271(csa_tree_add_95_22_pad_groupi_n_458 ,csa_tree_add_95_22_pad_groupi_n_186 ,csa_tree_add_95_22_pad_groupi_n_300);
  or csa_tree_add_95_22_pad_groupi_g5272(csa_tree_add_95_22_pad_groupi_n_457 ,csa_tree_add_95_22_pad_groupi_n_21 ,csa_tree_add_95_22_pad_groupi_n_291);
  nor csa_tree_add_95_22_pad_groupi_g5273(csa_tree_add_95_22_pad_groupi_n_456 ,csa_tree_add_95_22_pad_groupi_n_98 ,csa_tree_add_95_22_pad_groupi_n_296);
  nor csa_tree_add_95_22_pad_groupi_g5274(csa_tree_add_95_22_pad_groupi_n_455 ,csa_tree_add_95_22_pad_groupi_n_207 ,csa_tree_add_95_22_pad_groupi_n_297);
  nor csa_tree_add_95_22_pad_groupi_g5284(csa_tree_add_95_22_pad_groupi_n_445 ,csa_tree_add_95_22_pad_groupi_n_106 ,csa_tree_add_95_22_pad_groupi_n_294);
  nor csa_tree_add_95_22_pad_groupi_g5290(csa_tree_add_95_22_pad_groupi_n_439 ,csa_tree_add_95_22_pad_groupi_n_109 ,csa_tree_add_95_22_pad_groupi_n_241);
  or csa_tree_add_95_22_pad_groupi_g5291(csa_tree_add_95_22_pad_groupi_n_438 ,csa_tree_add_95_22_pad_groupi_n_32 ,csa_tree_add_95_22_pad_groupi_n_103);
  nor csa_tree_add_95_22_pad_groupi_g5294(csa_tree_add_95_22_pad_groupi_n_435 ,csa_tree_add_95_22_pad_groupi_n_107 ,csa_tree_add_95_22_pad_groupi_n_240);
  or csa_tree_add_95_22_pad_groupi_g5295(csa_tree_add_95_22_pad_groupi_n_434 ,csa_tree_add_95_22_pad_groupi_n_293 ,csa_tree_add_95_22_pad_groupi_n_110);
  nor csa_tree_add_95_22_pad_groupi_g5296(csa_tree_add_95_22_pad_groupi_n_433 ,csa_tree_add_95_22_pad_groupi_n_103 ,csa_tree_add_95_22_pad_groupi_n_294);
  or csa_tree_add_95_22_pad_groupi_g5297(csa_tree_add_95_22_pad_groupi_n_432 ,csa_tree_add_95_22_pad_groupi_n_13 ,csa_tree_add_95_22_pad_groupi_n_61);
  nor csa_tree_add_95_22_pad_groupi_g5298(csa_tree_add_95_22_pad_groupi_n_431 ,csa_tree_add_95_22_pad_groupi_n_110 ,csa_tree_add_95_22_pad_groupi_n_238);
  or csa_tree_add_95_22_pad_groupi_g5299(csa_tree_add_95_22_pad_groupi_n_430 ,csa_tree_add_95_22_pad_groupi_n_13 ,csa_tree_add_95_22_pad_groupi_n_104);
  nor csa_tree_add_95_22_pad_groupi_g5300(csa_tree_add_95_22_pad_groupi_n_429 ,csa_tree_add_95_22_pad_groupi_n_61 ,csa_tree_add_95_22_pad_groupi_n_32);
  nor csa_tree_add_95_22_pad_groupi_g5301(csa_tree_add_95_22_pad_groupi_n_428 ,csa_tree_add_95_22_pad_groupi_n_249 ,csa_tree_add_95_22_pad_groupi_n_34);
  or csa_tree_add_95_22_pad_groupi_g5302(csa_tree_add_95_22_pad_groupi_n_427 ,csa_tree_add_95_22_pad_groupi_n_15 ,csa_tree_add_95_22_pad_groupi_n_106);
  or csa_tree_add_95_22_pad_groupi_g5303(csa_tree_add_95_22_pad_groupi_n_426 ,csa_tree_add_95_22_pad_groupi_n_34 ,csa_tree_add_95_22_pad_groupi_n_107);
  nor csa_tree_add_95_22_pad_groupi_g5304(csa_tree_add_95_22_pad_groupi_n_425 ,csa_tree_add_95_22_pad_groupi_n_104 ,csa_tree_add_95_22_pad_groupi_n_237);
  or csa_tree_add_95_22_pad_groupi_g5305(csa_tree_add_95_22_pad_groupi_n_511 ,csa_tree_add_95_22_pad_groupi_n_154 ,csa_tree_add_95_22_pad_groupi_n_424);
  or csa_tree_add_95_22_pad_groupi_g5306(csa_tree_add_95_22_pad_groupi_n_505 ,csa_tree_add_95_22_pad_groupi_n_150 ,csa_tree_add_95_22_pad_groupi_n_403);
  or csa_tree_add_95_22_pad_groupi_g5307(csa_tree_add_95_22_pad_groupi_n_499 ,csa_tree_add_95_22_pad_groupi_n_155 ,csa_tree_add_95_22_pad_groupi_n_402);
  or csa_tree_add_95_22_pad_groupi_g5309(csa_tree_add_95_22_pad_groupi_n_493 ,csa_tree_add_95_22_pad_groupi_n_152 ,csa_tree_add_95_22_pad_groupi_n_404);
  not csa_tree_add_95_22_pad_groupi_g5311(csa_tree_add_95_22_pad_groupi_n_423 ,csa_tree_add_95_22_pad_groupi_n_158);
  not csa_tree_add_95_22_pad_groupi_g5312(csa_tree_add_95_22_pad_groupi_n_422 ,csa_tree_add_95_22_pad_groupi_n_155);
  not csa_tree_add_95_22_pad_groupi_g5315(csa_tree_add_95_22_pad_groupi_n_419 ,csa_tree_add_95_22_pad_groupi_n_154);
  not csa_tree_add_95_22_pad_groupi_g5317(csa_tree_add_95_22_pad_groupi_n_418 ,csa_tree_add_95_22_pad_groupi_n_149);
  not csa_tree_add_95_22_pad_groupi_g5319(csa_tree_add_95_22_pad_groupi_n_416 ,csa_tree_add_95_22_pad_groupi_n_152);
  not csa_tree_add_95_22_pad_groupi_g5321(csa_tree_add_95_22_pad_groupi_n_415 ,csa_tree_add_95_22_pad_groupi_n_151);
  not csa_tree_add_95_22_pad_groupi_g5323(csa_tree_add_95_22_pad_groupi_n_414 ,csa_tree_add_95_22_pad_groupi_n_160);
  not csa_tree_add_95_22_pad_groupi_g5324(csa_tree_add_95_22_pad_groupi_n_413 ,csa_tree_add_95_22_pad_groupi_n_153);
  not csa_tree_add_95_22_pad_groupi_g5327(csa_tree_add_95_22_pad_groupi_n_411 ,csa_tree_add_95_22_pad_groupi_n_159);
  not csa_tree_add_95_22_pad_groupi_g5328(csa_tree_add_95_22_pad_groupi_n_410 ,csa_tree_add_95_22_pad_groupi_n_150);
  or csa_tree_add_95_22_pad_groupi_g5331(csa_tree_add_95_22_pad_groupi_n_406 ,in17[10] ,in17[9]);
  and csa_tree_add_95_22_pad_groupi_g5332(csa_tree_add_95_22_pad_groupi_n_424 ,csa_tree_add_95_22_pad_groupi_n_375 ,csa_tree_add_95_22_pad_groupi_n_388);
  and csa_tree_add_95_22_pad_groupi_g5333(csa_tree_add_95_22_pad_groupi_n_421 ,n_551 ,n_558);
  and csa_tree_add_95_22_pad_groupi_g5334(csa_tree_add_95_22_pad_groupi_n_420 ,in18[0] ,n_560);
  and csa_tree_add_95_22_pad_groupi_g5335(csa_tree_add_95_22_pad_groupi_n_417 ,n_552 ,n_559);
  and csa_tree_add_95_22_pad_groupi_g5337(csa_tree_add_95_22_pad_groupi_n_409 ,n_550 ,n_557);
  not csa_tree_add_95_22_pad_groupi_g5339(csa_tree_add_95_22_pad_groupi_n_399 ,csa_tree_add_95_22_pad_groupi_n_293);
  not csa_tree_add_95_22_pad_groupi_g5340(csa_tree_add_95_22_pad_groupi_n_398 ,csa_tree_add_95_22_pad_groupi_n_395);
  not csa_tree_add_95_22_pad_groupi_g5341(csa_tree_add_95_22_pad_groupi_n_397 ,csa_tree_add_95_22_pad_groupi_n_258);
  not csa_tree_add_95_22_pad_groupi_g5345(csa_tree_add_95_22_pad_groupi_n_396 ,csa_tree_add_95_22_pad_groupi_n_395);
  and csa_tree_add_95_22_pad_groupi_g5346(csa_tree_add_95_22_pad_groupi_n_394 ,in17[10] ,in17[9]);
  and csa_tree_add_95_22_pad_groupi_g5348(csa_tree_add_95_22_pad_groupi_n_404 ,csa_tree_add_95_22_pad_groupi_n_391 ,csa_tree_add_95_22_pad_groupi_n_393);
  and csa_tree_add_95_22_pad_groupi_g5349(csa_tree_add_95_22_pad_groupi_n_403 ,csa_tree_add_95_22_pad_groupi_n_378 ,csa_tree_add_95_22_pad_groupi_n_377);
  and csa_tree_add_95_22_pad_groupi_g5350(csa_tree_add_95_22_pad_groupi_n_402 ,csa_tree_add_95_22_pad_groupi_n_392 ,csa_tree_add_95_22_pad_groupi_n_376);
  and csa_tree_add_95_22_pad_groupi_g5351(csa_tree_add_95_22_pad_groupi_n_401 ,csa_tree_add_95_22_pad_groupi_n_390 ,csa_tree_add_95_22_pad_groupi_n_389);
  or csa_tree_add_95_22_pad_groupi_g5353(csa_tree_add_95_22_pad_groupi_n_395 ,csa_tree_add_95_22_pad_groupi_n_390 ,csa_tree_add_95_22_pad_groupi_n_389);
  not csa_tree_add_95_22_pad_groupi_g5354(csa_tree_add_95_22_pad_groupi_n_393 ,n_559);
  not csa_tree_add_95_22_pad_groupi_g5355(csa_tree_add_95_22_pad_groupi_n_392 ,n_551);
  not csa_tree_add_95_22_pad_groupi_g5356(csa_tree_add_95_22_pad_groupi_n_391 ,n_552);
  not csa_tree_add_95_22_pad_groupi_g5357(csa_tree_add_95_22_pad_groupi_n_390 ,n_554);
  not csa_tree_add_95_22_pad_groupi_g5358(csa_tree_add_95_22_pad_groupi_n_389 ,n_561);
  not csa_tree_add_95_22_pad_groupi_g5359(csa_tree_add_95_22_pad_groupi_n_388 ,n_560);
  not csa_tree_add_95_22_pad_groupi_g5360(csa_tree_add_95_22_pad_groupi_n_387 ,in17[7]);
  not csa_tree_add_95_22_pad_groupi_g5361(csa_tree_add_95_22_pad_groupi_n_386 ,in9[15]);
  not csa_tree_add_95_22_pad_groupi_g5362(csa_tree_add_95_22_pad_groupi_n_385 ,in9[2]);
  not csa_tree_add_95_22_pad_groupi_g5363(csa_tree_add_95_22_pad_groupi_n_384 ,in9[5]);
  not csa_tree_add_95_22_pad_groupi_g5364(csa_tree_add_95_22_pad_groupi_n_383 ,in9[13]);
  not csa_tree_add_95_22_pad_groupi_g5365(csa_tree_add_95_22_pad_groupi_n_382 ,in9[3]);
  not csa_tree_add_95_22_pad_groupi_g5366(csa_tree_add_95_22_pad_groupi_n_381 ,in9[9]);
  not csa_tree_add_95_22_pad_groupi_g5367(csa_tree_add_95_22_pad_groupi_n_380 ,in9[1]);
  not csa_tree_add_95_22_pad_groupi_g5368(csa_tree_add_95_22_pad_groupi_n_379 ,in9[8]);
  not csa_tree_add_95_22_pad_groupi_g5369(csa_tree_add_95_22_pad_groupi_n_378 ,n_550);
  not csa_tree_add_95_22_pad_groupi_g5370(csa_tree_add_95_22_pad_groupi_n_377 ,n_557);
  not csa_tree_add_95_22_pad_groupi_g5371(csa_tree_add_95_22_pad_groupi_n_376 ,n_558);
  not csa_tree_add_95_22_pad_groupi_g5372(csa_tree_add_95_22_pad_groupi_n_375 ,in18[0]);
  not csa_tree_add_95_22_pad_groupi_g5373(csa_tree_add_95_22_pad_groupi_n_374 ,in17[0]);
  not csa_tree_add_95_22_pad_groupi_g5374(csa_tree_add_95_22_pad_groupi_n_373 ,in17[11]);
  not csa_tree_add_95_22_pad_groupi_g5375(csa_tree_add_95_22_pad_groupi_n_372 ,in17[8]);
  not csa_tree_add_95_22_pad_groupi_g5376(csa_tree_add_95_22_pad_groupi_n_371 ,in17[1]);
  not csa_tree_add_95_22_pad_groupi_g5377(csa_tree_add_95_22_pad_groupi_n_370 ,in17[6]);
  not csa_tree_add_95_22_pad_groupi_g5378(csa_tree_add_95_22_pad_groupi_n_369 ,in17[9]);
  not csa_tree_add_95_22_pad_groupi_g5379(csa_tree_add_95_22_pad_groupi_n_368 ,in9[0]);
  not csa_tree_add_95_22_pad_groupi_g5380(csa_tree_add_95_22_pad_groupi_n_367 ,in9[4]);
  not csa_tree_add_95_22_pad_groupi_g5381(csa_tree_add_95_22_pad_groupi_n_366 ,in9[12]);
  not csa_tree_add_95_22_pad_groupi_g5382(csa_tree_add_95_22_pad_groupi_n_365 ,in9[11]);
  not csa_tree_add_95_22_pad_groupi_g5383(csa_tree_add_95_22_pad_groupi_n_364 ,in9[7]);
  not csa_tree_add_95_22_pad_groupi_g5384(csa_tree_add_95_22_pad_groupi_n_363 ,in9[10]);
  not csa_tree_add_95_22_pad_groupi_g5385(csa_tree_add_95_22_pad_groupi_n_362 ,in9[6]);
  not csa_tree_add_95_22_pad_groupi_g5386(csa_tree_add_95_22_pad_groupi_n_361 ,in9[14]);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5534(csa_tree_add_95_22_pad_groupi_n_345 ,csa_tree_add_95_22_pad_groupi_n_343);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5535(csa_tree_add_95_22_pad_groupi_n_344 ,csa_tree_add_95_22_pad_groupi_n_343);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5536(csa_tree_add_95_22_pad_groupi_n_343 ,csa_tree_add_95_22_pad_groupi_n_356);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5538(csa_tree_add_95_22_pad_groupi_n_342 ,csa_tree_add_95_22_pad_groupi_n_340);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5539(csa_tree_add_95_22_pad_groupi_n_341 ,csa_tree_add_95_22_pad_groupi_n_340);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5540(csa_tree_add_95_22_pad_groupi_n_340 ,csa_tree_add_95_22_pad_groupi_n_422);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5542(csa_tree_add_95_22_pad_groupi_n_339 ,csa_tree_add_95_22_pad_groupi_n_337);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5543(csa_tree_add_95_22_pad_groupi_n_338 ,csa_tree_add_95_22_pad_groupi_n_337);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5544(csa_tree_add_95_22_pad_groupi_n_337 ,csa_tree_add_95_22_pad_groupi_n_413);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5546(csa_tree_add_95_22_pad_groupi_n_336 ,csa_tree_add_95_22_pad_groupi_n_334);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5547(csa_tree_add_95_22_pad_groupi_n_335 ,csa_tree_add_95_22_pad_groupi_n_334);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5548(csa_tree_add_95_22_pad_groupi_n_334 ,csa_tree_add_95_22_pad_groupi_n_348);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5550(csa_tree_add_95_22_pad_groupi_n_333 ,csa_tree_add_95_22_pad_groupi_n_331);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5551(csa_tree_add_95_22_pad_groupi_n_332 ,csa_tree_add_95_22_pad_groupi_n_331);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5552(csa_tree_add_95_22_pad_groupi_n_331 ,csa_tree_add_95_22_pad_groupi_n_411);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5554(csa_tree_add_95_22_pad_groupi_n_330 ,csa_tree_add_95_22_pad_groupi_n_328);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5555(csa_tree_add_95_22_pad_groupi_n_329 ,csa_tree_add_95_22_pad_groupi_n_328);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5556(csa_tree_add_95_22_pad_groupi_n_328 ,csa_tree_add_95_22_pad_groupi_n_410);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5558(csa_tree_add_95_22_pad_groupi_n_327 ,csa_tree_add_95_22_pad_groupi_n_325);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5559(csa_tree_add_95_22_pad_groupi_n_326 ,csa_tree_add_95_22_pad_groupi_n_325);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5560(csa_tree_add_95_22_pad_groupi_n_325 ,csa_tree_add_95_22_pad_groupi_n_350);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5562(csa_tree_add_95_22_pad_groupi_n_324 ,csa_tree_add_95_22_pad_groupi_n_322);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5563(csa_tree_add_95_22_pad_groupi_n_323 ,csa_tree_add_95_22_pad_groupi_n_322);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5564(csa_tree_add_95_22_pad_groupi_n_322 ,csa_tree_add_95_22_pad_groupi_n_419);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5566(csa_tree_add_95_22_pad_groupi_n_321 ,csa_tree_add_95_22_pad_groupi_n_319);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5567(csa_tree_add_95_22_pad_groupi_n_320 ,csa_tree_add_95_22_pad_groupi_n_319);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5568(csa_tree_add_95_22_pad_groupi_n_319 ,csa_tree_add_95_22_pad_groupi_n_416);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5570(csa_tree_add_95_22_pad_groupi_n_318 ,csa_tree_add_95_22_pad_groupi_n_316);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5571(csa_tree_add_95_22_pad_groupi_n_317 ,csa_tree_add_95_22_pad_groupi_n_316);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5572(csa_tree_add_95_22_pad_groupi_n_316 ,csa_tree_add_95_22_pad_groupi_n_351);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5574(csa_tree_add_95_22_pad_groupi_n_315 ,csa_tree_add_95_22_pad_groupi_n_313);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5575(csa_tree_add_95_22_pad_groupi_n_314 ,csa_tree_add_95_22_pad_groupi_n_313);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5576(csa_tree_add_95_22_pad_groupi_n_313 ,csa_tree_add_95_22_pad_groupi_n_415);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5578(csa_tree_add_95_22_pad_groupi_n_312 ,csa_tree_add_95_22_pad_groupi_n_310);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5579(csa_tree_add_95_22_pad_groupi_n_311 ,csa_tree_add_95_22_pad_groupi_n_310);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5580(csa_tree_add_95_22_pad_groupi_n_310 ,csa_tree_add_95_22_pad_groupi_n_423);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5582(csa_tree_add_95_22_pad_groupi_n_309 ,csa_tree_add_95_22_pad_groupi_n_307);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5583(csa_tree_add_95_22_pad_groupi_n_308 ,csa_tree_add_95_22_pad_groupi_n_307);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5584(csa_tree_add_95_22_pad_groupi_n_307 ,csa_tree_add_95_22_pad_groupi_n_414);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5586(csa_tree_add_95_22_pad_groupi_n_306 ,csa_tree_add_95_22_pad_groupi_n_304);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5587(csa_tree_add_95_22_pad_groupi_n_305 ,csa_tree_add_95_22_pad_groupi_n_304);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5588(csa_tree_add_95_22_pad_groupi_n_304 ,csa_tree_add_95_22_pad_groupi_n_353);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5590(csa_tree_add_95_22_pad_groupi_n_303 ,csa_tree_add_95_22_pad_groupi_n_301);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5591(csa_tree_add_95_22_pad_groupi_n_302 ,csa_tree_add_95_22_pad_groupi_n_301);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5592(csa_tree_add_95_22_pad_groupi_n_301 ,csa_tree_add_95_22_pad_groupi_n_418);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5594(csa_tree_add_95_22_pad_groupi_n_300 ,csa_tree_add_95_22_pad_groupi_n_298);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5595(csa_tree_add_95_22_pad_groupi_n_299 ,csa_tree_add_95_22_pad_groupi_n_298);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5596(csa_tree_add_95_22_pad_groupi_n_298 ,csa_tree_add_95_22_pad_groupi_n_397);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5598(csa_tree_add_95_22_pad_groupi_n_297 ,csa_tree_add_95_22_pad_groupi_n_295);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5599(csa_tree_add_95_22_pad_groupi_n_296 ,csa_tree_add_95_22_pad_groupi_n_295);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5600(csa_tree_add_95_22_pad_groupi_n_295 ,csa_tree_add_95_22_pad_groupi_n_346);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5602(csa_tree_add_95_22_pad_groupi_n_294 ,csa_tree_add_95_22_pad_groupi_n_292);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5603(csa_tree_add_95_22_pad_groupi_n_293 ,csa_tree_add_95_22_pad_groupi_n_292);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5604(csa_tree_add_95_22_pad_groupi_n_292 ,csa_tree_add_95_22_pad_groupi_n_398);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5606(csa_tree_add_95_22_pad_groupi_n_291 ,csa_tree_add_95_22_pad_groupi_n_289);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5607(csa_tree_add_95_22_pad_groupi_n_290 ,csa_tree_add_95_22_pad_groupi_n_289);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5608(csa_tree_add_95_22_pad_groupi_n_289 ,csa_tree_add_95_22_pad_groupi_n_397);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5610(csa_tree_add_95_22_pad_groupi_n_288 ,csa_tree_add_95_22_pad_groupi_n_286);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5611(csa_tree_add_95_22_pad_groupi_n_287 ,csa_tree_add_95_22_pad_groupi_n_286);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5612(csa_tree_add_95_22_pad_groupi_n_286 ,csa_tree_add_95_22_pad_groupi_n_509);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5614(csa_tree_add_95_22_pad_groupi_n_285 ,csa_tree_add_95_22_pad_groupi_n_283);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5615(csa_tree_add_95_22_pad_groupi_n_284 ,csa_tree_add_95_22_pad_groupi_n_283);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5616(csa_tree_add_95_22_pad_groupi_n_283 ,csa_tree_add_95_22_pad_groupi_n_503);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5620(csa_tree_add_95_22_pad_groupi_n_358 ,csa_tree_add_95_22_pad_groupi_n_581);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5623(csa_tree_add_95_22_pad_groupi_n_282 ,csa_tree_add_95_22_pad_groupi_n_281);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5624(csa_tree_add_95_22_pad_groupi_n_281 ,csa_tree_add_95_22_pad_groupi_n_579);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5627(csa_tree_add_95_22_pad_groupi_n_280 ,csa_tree_add_95_22_pad_groupi_n_279);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5628(csa_tree_add_95_22_pad_groupi_n_279 ,csa_tree_add_95_22_pad_groupi_n_582);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5632(csa_tree_add_95_22_pad_groupi_n_357 ,csa_tree_add_95_22_pad_groupi_n_580);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5635(csa_tree_add_95_22_pad_groupi_n_278 ,csa_tree_add_95_22_pad_groupi_n_277);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5636(csa_tree_add_95_22_pad_groupi_n_277 ,csa_tree_add_95_22_pad_groupi_n_497);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5639(csa_tree_add_95_22_pad_groupi_n_276 ,csa_tree_add_95_22_pad_groupi_n_359);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5640(csa_tree_add_95_22_pad_groupi_n_359 ,csa_tree_add_95_22_pad_groupi_n_934);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5642(csa_tree_add_95_22_pad_groupi_n_275 ,csa_tree_add_95_22_pad_groupi_n_273);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5643(csa_tree_add_95_22_pad_groupi_n_274 ,csa_tree_add_95_22_pad_groupi_n_273);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5644(csa_tree_add_95_22_pad_groupi_n_273 ,csa_tree_add_95_22_pad_groupi_n_355);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5646(csa_tree_add_95_22_pad_groupi_n_272 ,csa_tree_add_95_22_pad_groupi_n_270);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5647(csa_tree_add_95_22_pad_groupi_n_271 ,csa_tree_add_95_22_pad_groupi_n_270);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5648(csa_tree_add_95_22_pad_groupi_n_270 ,csa_tree_add_95_22_pad_groupi_n_349);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5650(csa_tree_add_95_22_pad_groupi_n_269 ,csa_tree_add_95_22_pad_groupi_n_267);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5651(csa_tree_add_95_22_pad_groupi_n_268 ,csa_tree_add_95_22_pad_groupi_n_267);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5652(csa_tree_add_95_22_pad_groupi_n_267 ,csa_tree_add_95_22_pad_groupi_n_347);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5654(csa_tree_add_95_22_pad_groupi_n_266 ,csa_tree_add_95_22_pad_groupi_n_264);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5655(csa_tree_add_95_22_pad_groupi_n_265 ,csa_tree_add_95_22_pad_groupi_n_264);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5656(csa_tree_add_95_22_pad_groupi_n_264 ,csa_tree_add_95_22_pad_groupi_n_354);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5658(csa_tree_add_95_22_pad_groupi_n_263 ,csa_tree_add_95_22_pad_groupi_n_261);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5659(csa_tree_add_95_22_pad_groupi_n_262 ,csa_tree_add_95_22_pad_groupi_n_261);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5660(csa_tree_add_95_22_pad_groupi_n_261 ,csa_tree_add_95_22_pad_groupi_n_352);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5662(csa_tree_add_95_22_pad_groupi_n_260 ,csa_tree_add_95_22_pad_groupi_n_259);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5664(csa_tree_add_95_22_pad_groupi_n_259 ,csa_tree_add_95_22_pad_groupi_n_399);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5686(csa_tree_add_95_22_pad_groupi_n_258 ,csa_tree_add_95_22_pad_groupi_n_346);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5688(csa_tree_add_95_22_pad_groupi_n_346 ,csa_tree_add_95_22_pad_groupi_n_398);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5690(csa_tree_add_95_22_pad_groupi_n_257 ,csa_tree_add_95_22_pad_groupi_n_256);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5692(csa_tree_add_95_22_pad_groupi_n_256 ,csa_tree_add_95_22_pad_groupi_n_507);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5694(csa_tree_add_95_22_pad_groupi_n_255 ,csa_tree_add_95_22_pad_groupi_n_254);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5696(csa_tree_add_95_22_pad_groupi_n_254 ,csa_tree_add_95_22_pad_groupi_n_501);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5709(csa_tree_add_95_22_pad_groupi_n_253 ,csa_tree_add_95_22_pad_groupi_n_251);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5710(csa_tree_add_95_22_pad_groupi_n_252 ,csa_tree_add_95_22_pad_groupi_n_251);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5711(csa_tree_add_95_22_pad_groupi_n_251 ,csa_tree_add_95_22_pad_groupi_n_511);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5713(csa_tree_add_95_22_pad_groupi_n_250 ,csa_tree_add_95_22_pad_groupi_n_248);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5714(csa_tree_add_95_22_pad_groupi_n_249 ,csa_tree_add_95_22_pad_groupi_n_248);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5715(csa_tree_add_95_22_pad_groupi_n_248 ,csa_tree_add_95_22_pad_groupi_n_401);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5721(csa_tree_add_95_22_pad_groupi_n_247 ,csa_tree_add_95_22_pad_groupi_n_245);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5722(csa_tree_add_95_22_pad_groupi_n_246 ,csa_tree_add_95_22_pad_groupi_n_245);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5723(csa_tree_add_95_22_pad_groupi_n_245 ,csa_tree_add_95_22_pad_groupi_n_385);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5733(csa_tree_add_95_22_pad_groupi_n_244 ,csa_tree_add_95_22_pad_groupi_n_242);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5734(csa_tree_add_95_22_pad_groupi_n_243 ,csa_tree_add_95_22_pad_groupi_n_242);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5735(csa_tree_add_95_22_pad_groupi_n_242 ,csa_tree_add_95_22_pad_groupi_n_368);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5737(csa_tree_add_95_22_pad_groupi_n_241 ,csa_tree_add_95_22_pad_groupi_n_239);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5738(csa_tree_add_95_22_pad_groupi_n_240 ,csa_tree_add_95_22_pad_groupi_n_239);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5739(csa_tree_add_95_22_pad_groupi_n_239 ,csa_tree_add_95_22_pad_groupi_n_396);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5741(csa_tree_add_95_22_pad_groupi_n_238 ,csa_tree_add_95_22_pad_groupi_n_236);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5742(csa_tree_add_95_22_pad_groupi_n_237 ,csa_tree_add_95_22_pad_groupi_n_236);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5743(csa_tree_add_95_22_pad_groupi_n_236 ,csa_tree_add_95_22_pad_groupi_n_396);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5746(csa_tree_add_95_22_pad_groupi_n_235 ,csa_tree_add_95_22_pad_groupi_n_234);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5747(csa_tree_add_95_22_pad_groupi_n_234 ,csa_tree_add_95_22_pad_groupi_n_381);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5750(csa_tree_add_95_22_pad_groupi_n_233 ,csa_tree_add_95_22_pad_groupi_n_232);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5751(csa_tree_add_95_22_pad_groupi_n_232 ,csa_tree_add_95_22_pad_groupi_n_366);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5754(csa_tree_add_95_22_pad_groupi_n_231 ,csa_tree_add_95_22_pad_groupi_n_230);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5755(csa_tree_add_95_22_pad_groupi_n_230 ,csa_tree_add_95_22_pad_groupi_n_382);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5758(csa_tree_add_95_22_pad_groupi_n_229 ,csa_tree_add_95_22_pad_groupi_n_228);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5759(csa_tree_add_95_22_pad_groupi_n_228 ,csa_tree_add_95_22_pad_groupi_n_383);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5762(csa_tree_add_95_22_pad_groupi_n_227 ,csa_tree_add_95_22_pad_groupi_n_226);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5763(csa_tree_add_95_22_pad_groupi_n_226 ,csa_tree_add_95_22_pad_groupi_n_365);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5766(csa_tree_add_95_22_pad_groupi_n_225 ,csa_tree_add_95_22_pad_groupi_n_224);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5767(csa_tree_add_95_22_pad_groupi_n_224 ,csa_tree_add_95_22_pad_groupi_n_363);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5769(csa_tree_add_95_22_pad_groupi_n_223 ,csa_tree_add_95_22_pad_groupi_n_221);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5770(csa_tree_add_95_22_pad_groupi_n_222 ,csa_tree_add_95_22_pad_groupi_n_221);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5771(csa_tree_add_95_22_pad_groupi_n_221 ,csa_tree_add_95_22_pad_groupi_n_366);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5774(csa_tree_add_95_22_pad_groupi_n_220 ,csa_tree_add_95_22_pad_groupi_n_219);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5775(csa_tree_add_95_22_pad_groupi_n_219 ,csa_tree_add_95_22_pad_groupi_n_362);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5777(csa_tree_add_95_22_pad_groupi_n_218 ,csa_tree_add_95_22_pad_groupi_n_216);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5778(csa_tree_add_95_22_pad_groupi_n_217 ,csa_tree_add_95_22_pad_groupi_n_216);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5779(csa_tree_add_95_22_pad_groupi_n_216 ,csa_tree_add_95_22_pad_groupi_n_380);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5781(csa_tree_add_95_22_pad_groupi_n_215 ,csa_tree_add_95_22_pad_groupi_n_213);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5782(csa_tree_add_95_22_pad_groupi_n_214 ,csa_tree_add_95_22_pad_groupi_n_213);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5783(csa_tree_add_95_22_pad_groupi_n_213 ,csa_tree_add_95_22_pad_groupi_n_381);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5785(csa_tree_add_95_22_pad_groupi_n_212 ,csa_tree_add_95_22_pad_groupi_n_210);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5786(csa_tree_add_95_22_pad_groupi_n_211 ,csa_tree_add_95_22_pad_groupi_n_210);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5787(csa_tree_add_95_22_pad_groupi_n_210 ,csa_tree_add_95_22_pad_groupi_n_362);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5790(csa_tree_add_95_22_pad_groupi_n_209 ,csa_tree_add_95_22_pad_groupi_n_208);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5791(csa_tree_add_95_22_pad_groupi_n_208 ,csa_tree_add_95_22_pad_groupi_n_379);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5793(csa_tree_add_95_22_pad_groupi_n_207 ,csa_tree_add_95_22_pad_groupi_n_205);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5794(csa_tree_add_95_22_pad_groupi_n_206 ,csa_tree_add_95_22_pad_groupi_n_205);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5795(csa_tree_add_95_22_pad_groupi_n_205 ,csa_tree_add_95_22_pad_groupi_n_379);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5798(csa_tree_add_95_22_pad_groupi_n_204 ,csa_tree_add_95_22_pad_groupi_n_203);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5799(csa_tree_add_95_22_pad_groupi_n_203 ,csa_tree_add_95_22_pad_groupi_n_384);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5801(csa_tree_add_95_22_pad_groupi_n_202 ,csa_tree_add_95_22_pad_groupi_n_200);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5802(csa_tree_add_95_22_pad_groupi_n_201 ,csa_tree_add_95_22_pad_groupi_n_200);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5803(csa_tree_add_95_22_pad_groupi_n_200 ,csa_tree_add_95_22_pad_groupi_n_382);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5807(csa_tree_add_95_22_pad_groupi_n_198 ,csa_tree_add_95_22_pad_groupi_n_361);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5809(csa_tree_add_95_22_pad_groupi_n_197 ,csa_tree_add_95_22_pad_groupi_n_195);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5810(csa_tree_add_95_22_pad_groupi_n_196 ,csa_tree_add_95_22_pad_groupi_n_195);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5811(csa_tree_add_95_22_pad_groupi_n_195 ,csa_tree_add_95_22_pad_groupi_n_384);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5813(csa_tree_add_95_22_pad_groupi_n_194 ,csa_tree_add_95_22_pad_groupi_n_192);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5814(csa_tree_add_95_22_pad_groupi_n_193 ,csa_tree_add_95_22_pad_groupi_n_192);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5815(csa_tree_add_95_22_pad_groupi_n_192 ,csa_tree_add_95_22_pad_groupi_n_361);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5817(csa_tree_add_95_22_pad_groupi_n_191 ,csa_tree_add_95_22_pad_groupi_n_190);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5819(csa_tree_add_95_22_pad_groupi_n_190 ,csa_tree_add_95_22_pad_groupi_n_364);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5822(csa_tree_add_95_22_pad_groupi_n_189 ,csa_tree_add_95_22_pad_groupi_n_188);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5823(csa_tree_add_95_22_pad_groupi_n_188 ,csa_tree_add_95_22_pad_groupi_n_367);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5825(csa_tree_add_95_22_pad_groupi_n_187 ,csa_tree_add_95_22_pad_groupi_n_185);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5826(csa_tree_add_95_22_pad_groupi_n_186 ,csa_tree_add_95_22_pad_groupi_n_185);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5827(csa_tree_add_95_22_pad_groupi_n_185 ,csa_tree_add_95_22_pad_groupi_n_383);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5829(csa_tree_add_95_22_pad_groupi_n_184 ,csa_tree_add_95_22_pad_groupi_n_182);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5830(csa_tree_add_95_22_pad_groupi_n_183 ,csa_tree_add_95_22_pad_groupi_n_182);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5831(csa_tree_add_95_22_pad_groupi_n_182 ,csa_tree_add_95_22_pad_groupi_n_364);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5833(csa_tree_add_95_22_pad_groupi_n_181 ,csa_tree_add_95_22_pad_groupi_n_179);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5834(csa_tree_add_95_22_pad_groupi_n_180 ,csa_tree_add_95_22_pad_groupi_n_179);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5835(csa_tree_add_95_22_pad_groupi_n_179 ,csa_tree_add_95_22_pad_groupi_n_365);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5837(csa_tree_add_95_22_pad_groupi_n_178 ,csa_tree_add_95_22_pad_groupi_n_176);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5838(csa_tree_add_95_22_pad_groupi_n_177 ,csa_tree_add_95_22_pad_groupi_n_176);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5839(csa_tree_add_95_22_pad_groupi_n_176 ,csa_tree_add_95_22_pad_groupi_n_363);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5841(csa_tree_add_95_22_pad_groupi_n_175 ,csa_tree_add_95_22_pad_groupi_n_173);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5842(csa_tree_add_95_22_pad_groupi_n_174 ,csa_tree_add_95_22_pad_groupi_n_173);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5843(csa_tree_add_95_22_pad_groupi_n_173 ,csa_tree_add_95_22_pad_groupi_n_367);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5845(csa_tree_add_95_22_pad_groupi_n_172 ,csa_tree_add_95_22_pad_groupi_n_170);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5846(csa_tree_add_95_22_pad_groupi_n_171 ,csa_tree_add_95_22_pad_groupi_n_170);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5847(csa_tree_add_95_22_pad_groupi_n_170 ,csa_tree_add_95_22_pad_groupi_n_495);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5849(csa_tree_add_95_22_pad_groupi_n_169 ,csa_tree_add_95_22_pad_groupi_n_167);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5850(csa_tree_add_95_22_pad_groupi_n_168 ,csa_tree_add_95_22_pad_groupi_n_167);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5851(csa_tree_add_95_22_pad_groupi_n_167 ,csa_tree_add_95_22_pad_groupi_n_495);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5853(csa_tree_add_95_22_pad_groupi_n_166 ,csa_tree_add_95_22_pad_groupi_n_164);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5854(csa_tree_add_95_22_pad_groupi_n_165 ,csa_tree_add_95_22_pad_groupi_n_164);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5855(csa_tree_add_95_22_pad_groupi_n_164 ,csa_tree_add_95_22_pad_groupi_n_498);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5857(csa_tree_add_95_22_pad_groupi_n_163 ,csa_tree_add_95_22_pad_groupi_n_161);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5858(csa_tree_add_95_22_pad_groupi_n_162 ,csa_tree_add_95_22_pad_groupi_n_161);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5859(csa_tree_add_95_22_pad_groupi_n_161 ,csa_tree_add_95_22_pad_groupi_n_386);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5861(csa_tree_add_95_22_pad_groupi_n_160 ,csa_tree_add_95_22_pad_groupi_n_350);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5863(csa_tree_add_95_22_pad_groupi_n_350 ,csa_tree_add_95_22_pad_groupi_n_412);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5865(csa_tree_add_95_22_pad_groupi_n_159 ,csa_tree_add_95_22_pad_groupi_n_348);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5867(csa_tree_add_95_22_pad_groupi_n_348 ,csa_tree_add_95_22_pad_groupi_n_409);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5869(csa_tree_add_95_22_pad_groupi_n_158 ,csa_tree_add_95_22_pad_groupi_n_356);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5871(csa_tree_add_95_22_pad_groupi_n_356 ,csa_tree_add_95_22_pad_groupi_n_421);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5877(csa_tree_add_95_22_pad_groupi_n_155 ,csa_tree_add_95_22_pad_groupi_n_355);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5879(csa_tree_add_95_22_pad_groupi_n_355 ,csa_tree_add_95_22_pad_groupi_n_421);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5881(csa_tree_add_95_22_pad_groupi_n_154 ,csa_tree_add_95_22_pad_groupi_n_353);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5883(csa_tree_add_95_22_pad_groupi_n_353 ,csa_tree_add_95_22_pad_groupi_n_420);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5885(csa_tree_add_95_22_pad_groupi_n_153 ,csa_tree_add_95_22_pad_groupi_n_349);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5887(csa_tree_add_95_22_pad_groupi_n_349 ,csa_tree_add_95_22_pad_groupi_n_412);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5889(csa_tree_add_95_22_pad_groupi_n_152 ,csa_tree_add_95_22_pad_groupi_n_351);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5891(csa_tree_add_95_22_pad_groupi_n_351 ,csa_tree_add_95_22_pad_groupi_n_417);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5893(csa_tree_add_95_22_pad_groupi_n_151 ,csa_tree_add_95_22_pad_groupi_n_352);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5895(csa_tree_add_95_22_pad_groupi_n_352 ,csa_tree_add_95_22_pad_groupi_n_417);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5897(csa_tree_add_95_22_pad_groupi_n_150 ,csa_tree_add_95_22_pad_groupi_n_347);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5899(csa_tree_add_95_22_pad_groupi_n_347 ,csa_tree_add_95_22_pad_groupi_n_409);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5901(csa_tree_add_95_22_pad_groupi_n_149 ,csa_tree_add_95_22_pad_groupi_n_354);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5903(csa_tree_add_95_22_pad_groupi_n_354 ,csa_tree_add_95_22_pad_groupi_n_420);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5905(csa_tree_add_95_22_pad_groupi_n_148 ,csa_tree_add_95_22_pad_groupi_n_146);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5906(csa_tree_add_95_22_pad_groupi_n_147 ,csa_tree_add_95_22_pad_groupi_n_146);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5907(csa_tree_add_95_22_pad_groupi_n_146 ,csa_tree_add_95_22_pad_groupi_n_504);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5909(csa_tree_add_95_22_pad_groupi_n_145 ,csa_tree_add_95_22_pad_groupi_n_143);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5910(csa_tree_add_95_22_pad_groupi_n_144 ,csa_tree_add_95_22_pad_groupi_n_143);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5911(csa_tree_add_95_22_pad_groupi_n_143 ,csa_tree_add_95_22_pad_groupi_n_510);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5913(csa_tree_add_95_22_pad_groupi_n_142 ,csa_tree_add_95_22_pad_groupi_n_140);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5914(csa_tree_add_95_22_pad_groupi_n_141 ,csa_tree_add_95_22_pad_groupi_n_140);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5915(csa_tree_add_95_22_pad_groupi_n_140 ,csa_tree_add_95_22_pad_groupi_n_510);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5917(csa_tree_add_95_22_pad_groupi_n_139 ,csa_tree_add_95_22_pad_groupi_n_137);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5918(csa_tree_add_95_22_pad_groupi_n_138 ,csa_tree_add_95_22_pad_groupi_n_137);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5919(csa_tree_add_95_22_pad_groupi_n_137 ,csa_tree_add_95_22_pad_groupi_n_494);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5921(csa_tree_add_95_22_pad_groupi_n_136 ,csa_tree_add_95_22_pad_groupi_n_134);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5922(csa_tree_add_95_22_pad_groupi_n_135 ,csa_tree_add_95_22_pad_groupi_n_134);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5923(csa_tree_add_95_22_pad_groupi_n_134 ,csa_tree_add_95_22_pad_groupi_n_494);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5925(csa_tree_add_95_22_pad_groupi_n_133 ,csa_tree_add_95_22_pad_groupi_n_131);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5926(csa_tree_add_95_22_pad_groupi_n_132 ,csa_tree_add_95_22_pad_groupi_n_131);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5927(csa_tree_add_95_22_pad_groupi_n_131 ,csa_tree_add_95_22_pad_groupi_n_504);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5929(csa_tree_add_95_22_pad_groupi_n_130 ,csa_tree_add_95_22_pad_groupi_n_128);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5930(csa_tree_add_95_22_pad_groupi_n_129 ,csa_tree_add_95_22_pad_groupi_n_128);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5931(csa_tree_add_95_22_pad_groupi_n_128 ,csa_tree_add_95_22_pad_groupi_n_498);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5933(csa_tree_add_95_22_pad_groupi_n_127 ,csa_tree_add_95_22_pad_groupi_n_125);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5934(csa_tree_add_95_22_pad_groupi_n_126 ,csa_tree_add_95_22_pad_groupi_n_125);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5935(csa_tree_add_95_22_pad_groupi_n_125 ,csa_tree_add_95_22_pad_groupi_n_496);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5937(csa_tree_add_95_22_pad_groupi_n_124 ,csa_tree_add_95_22_pad_groupi_n_122);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5938(csa_tree_add_95_22_pad_groupi_n_123 ,csa_tree_add_95_22_pad_groupi_n_122);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5939(csa_tree_add_95_22_pad_groupi_n_122 ,csa_tree_add_95_22_pad_groupi_n_496);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5941(csa_tree_add_95_22_pad_groupi_n_121 ,csa_tree_add_95_22_pad_groupi_n_120);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5943(csa_tree_add_95_22_pad_groupi_n_120 ,csa_tree_add_95_22_pad_groupi_n_386);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5945(csa_tree_add_95_22_pad_groupi_n_119 ,csa_tree_add_95_22_pad_groupi_n_117);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5946(csa_tree_add_95_22_pad_groupi_n_118 ,csa_tree_add_95_22_pad_groupi_n_117);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5947(csa_tree_add_95_22_pad_groupi_n_117 ,csa_tree_add_95_22_pad_groupi_n_511);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5949(csa_tree_add_95_22_pad_groupi_n_116 ,csa_tree_add_95_22_pad_groupi_n_114);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5950(csa_tree_add_95_22_pad_groupi_n_115 ,csa_tree_add_95_22_pad_groupi_n_114);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5951(csa_tree_add_95_22_pad_groupi_n_114 ,csa_tree_add_95_22_pad_groupi_n_511);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5953(csa_tree_add_95_22_pad_groupi_n_113 ,csa_tree_add_95_22_pad_groupi_n_111);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5954(csa_tree_add_95_22_pad_groupi_n_112 ,csa_tree_add_95_22_pad_groupi_n_111);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5955(csa_tree_add_95_22_pad_groupi_n_111 ,csa_tree_add_95_22_pad_groupi_n_253);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5957(csa_tree_add_95_22_pad_groupi_n_110 ,csa_tree_add_95_22_pad_groupi_n_108);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5958(csa_tree_add_95_22_pad_groupi_n_109 ,csa_tree_add_95_22_pad_groupi_n_108);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5959(csa_tree_add_95_22_pad_groupi_n_108 ,csa_tree_add_95_22_pad_groupi_n_401);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5961(csa_tree_add_95_22_pad_groupi_n_107 ,csa_tree_add_95_22_pad_groupi_n_105);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5962(csa_tree_add_95_22_pad_groupi_n_106 ,csa_tree_add_95_22_pad_groupi_n_105);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5963(csa_tree_add_95_22_pad_groupi_n_105 ,csa_tree_add_95_22_pad_groupi_n_401);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5965(csa_tree_add_95_22_pad_groupi_n_104 ,csa_tree_add_95_22_pad_groupi_n_102);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5966(csa_tree_add_95_22_pad_groupi_n_103 ,csa_tree_add_95_22_pad_groupi_n_102);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5967(csa_tree_add_95_22_pad_groupi_n_102 ,csa_tree_add_95_22_pad_groupi_n_250);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5969(csa_tree_add_95_22_pad_groupi_n_101 ,csa_tree_add_95_22_pad_groupi_n_99);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5970(csa_tree_add_95_22_pad_groupi_n_100 ,csa_tree_add_95_22_pad_groupi_n_99);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5971(csa_tree_add_95_22_pad_groupi_n_99 ,csa_tree_add_95_22_pad_groupi_n_385);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5973(csa_tree_add_95_22_pad_groupi_n_98 ,csa_tree_add_95_22_pad_groupi_n_97);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5975(csa_tree_add_95_22_pad_groupi_n_97 ,csa_tree_add_95_22_pad_groupi_n_247);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5977(csa_tree_add_95_22_pad_groupi_n_96 ,csa_tree_add_95_22_pad_groupi_n_94);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5978(csa_tree_add_95_22_pad_groupi_n_95 ,csa_tree_add_95_22_pad_groupi_n_94);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5979(csa_tree_add_95_22_pad_groupi_n_94 ,csa_tree_add_95_22_pad_groupi_n_381);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5981(csa_tree_add_95_22_pad_groupi_n_93 ,csa_tree_add_95_22_pad_groupi_n_92);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5983(csa_tree_add_95_22_pad_groupi_n_92 ,csa_tree_add_95_22_pad_groupi_n_252);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5985(csa_tree_add_95_22_pad_groupi_n_91 ,csa_tree_add_95_22_pad_groupi_n_89);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5986(csa_tree_add_95_22_pad_groupi_n_90 ,csa_tree_add_95_22_pad_groupi_n_89);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5987(csa_tree_add_95_22_pad_groupi_n_89 ,csa_tree_add_95_22_pad_groupi_n_366);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5989(csa_tree_add_95_22_pad_groupi_n_88 ,csa_tree_add_95_22_pad_groupi_n_86);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5990(csa_tree_add_95_22_pad_groupi_n_87 ,csa_tree_add_95_22_pad_groupi_n_86);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5991(csa_tree_add_95_22_pad_groupi_n_86 ,csa_tree_add_95_22_pad_groupi_n_382);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5993(csa_tree_add_95_22_pad_groupi_n_85 ,csa_tree_add_95_22_pad_groupi_n_83);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5994(csa_tree_add_95_22_pad_groupi_n_84 ,csa_tree_add_95_22_pad_groupi_n_83);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5995(csa_tree_add_95_22_pad_groupi_n_83 ,csa_tree_add_95_22_pad_groupi_n_383);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5997(csa_tree_add_95_22_pad_groupi_n_82 ,csa_tree_add_95_22_pad_groupi_n_80);
  not csa_tree_add_95_22_pad_groupi_drc_bufs5999(csa_tree_add_95_22_pad_groupi_n_80 ,csa_tree_add_95_22_pad_groupi_n_365);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6001(csa_tree_add_95_22_pad_groupi_n_79 ,csa_tree_add_95_22_pad_groupi_n_77);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6002(csa_tree_add_95_22_pad_groupi_n_78 ,csa_tree_add_95_22_pad_groupi_n_77);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6003(csa_tree_add_95_22_pad_groupi_n_77 ,csa_tree_add_95_22_pad_groupi_n_363);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6005(csa_tree_add_95_22_pad_groupi_n_76 ,csa_tree_add_95_22_pad_groupi_n_75);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6007(csa_tree_add_95_22_pad_groupi_n_75 ,csa_tree_add_95_22_pad_groupi_n_215);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6009(csa_tree_add_95_22_pad_groupi_n_74 ,csa_tree_add_95_22_pad_groupi_n_72);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6010(csa_tree_add_95_22_pad_groupi_n_73 ,csa_tree_add_95_22_pad_groupi_n_72);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6011(csa_tree_add_95_22_pad_groupi_n_72 ,csa_tree_add_95_22_pad_groupi_n_385);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6013(csa_tree_add_95_22_pad_groupi_n_71 ,csa_tree_add_95_22_pad_groupi_n_70);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6015(csa_tree_add_95_22_pad_groupi_n_70 ,csa_tree_add_95_22_pad_groupi_n_218);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6017(csa_tree_add_95_22_pad_groupi_n_69 ,csa_tree_add_95_22_pad_groupi_n_68);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6019(csa_tree_add_95_22_pad_groupi_n_68 ,csa_tree_add_95_22_pad_groupi_n_223);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6021(csa_tree_add_95_22_pad_groupi_n_67 ,csa_tree_add_95_22_pad_groupi_n_65);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6022(csa_tree_add_95_22_pad_groupi_n_66 ,csa_tree_add_95_22_pad_groupi_n_65);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6023(csa_tree_add_95_22_pad_groupi_n_65 ,csa_tree_add_95_22_pad_groupi_n_362);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6025(csa_tree_add_95_22_pad_groupi_n_64 ,csa_tree_add_95_22_pad_groupi_n_62);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6027(csa_tree_add_95_22_pad_groupi_n_62 ,csa_tree_add_95_22_pad_groupi_n_380);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6029(csa_tree_add_95_22_pad_groupi_n_61 ,csa_tree_add_95_22_pad_groupi_n_60);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6031(csa_tree_add_95_22_pad_groupi_n_60 ,csa_tree_add_95_22_pad_groupi_n_249);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6033(csa_tree_add_95_22_pad_groupi_n_59 ,csa_tree_add_95_22_pad_groupi_n_58);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6035(csa_tree_add_95_22_pad_groupi_n_58 ,csa_tree_add_95_22_pad_groupi_n_212);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6037(csa_tree_add_95_22_pad_groupi_n_57 ,csa_tree_add_95_22_pad_groupi_n_56);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6039(csa_tree_add_95_22_pad_groupi_n_56 ,csa_tree_add_95_22_pad_groupi_n_244);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6041(csa_tree_add_95_22_pad_groupi_n_55 ,csa_tree_add_95_22_pad_groupi_n_54);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6043(csa_tree_add_95_22_pad_groupi_n_54 ,csa_tree_add_95_22_pad_groupi_n_207);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6045(csa_tree_add_95_22_pad_groupi_n_53 ,csa_tree_add_95_22_pad_groupi_n_51);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6046(csa_tree_add_95_22_pad_groupi_n_52 ,csa_tree_add_95_22_pad_groupi_n_51);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6047(csa_tree_add_95_22_pad_groupi_n_51 ,csa_tree_add_95_22_pad_groupi_n_384);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6049(csa_tree_add_95_22_pad_groupi_n_50 ,csa_tree_add_95_22_pad_groupi_n_48);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6051(csa_tree_add_95_22_pad_groupi_n_48 ,csa_tree_add_95_22_pad_groupi_n_379);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6053(csa_tree_add_95_22_pad_groupi_n_47 ,csa_tree_add_95_22_pad_groupi_n_46);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6055(csa_tree_add_95_22_pad_groupi_n_46 ,csa_tree_add_95_22_pad_groupi_n_246);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6057(csa_tree_add_95_22_pad_groupi_n_45 ,csa_tree_add_95_22_pad_groupi_n_43);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6059(csa_tree_add_95_22_pad_groupi_n_43 ,csa_tree_add_95_22_pad_groupi_n_380);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6061(csa_tree_add_95_22_pad_groupi_n_42 ,csa_tree_add_95_22_pad_groupi_n_40);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6062(csa_tree_add_95_22_pad_groupi_n_41 ,csa_tree_add_95_22_pad_groupi_n_40);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6063(csa_tree_add_95_22_pad_groupi_n_40 ,csa_tree_add_95_22_pad_groupi_n_368);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6065(csa_tree_add_95_22_pad_groupi_n_39 ,csa_tree_add_95_22_pad_groupi_n_37);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6066(csa_tree_add_95_22_pad_groupi_n_38 ,csa_tree_add_95_22_pad_groupi_n_37);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6067(csa_tree_add_95_22_pad_groupi_n_37 ,csa_tree_add_95_22_pad_groupi_n_361);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6069(csa_tree_add_95_22_pad_groupi_n_36 ,csa_tree_add_95_22_pad_groupi_n_35);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6071(csa_tree_add_95_22_pad_groupi_n_35 ,csa_tree_add_95_22_pad_groupi_n_202);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6073(csa_tree_add_95_22_pad_groupi_n_34 ,csa_tree_add_95_22_pad_groupi_n_33);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6075(csa_tree_add_95_22_pad_groupi_n_33 ,csa_tree_add_95_22_pad_groupi_n_238);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6077(csa_tree_add_95_22_pad_groupi_n_32 ,csa_tree_add_95_22_pad_groupi_n_31);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6079(csa_tree_add_95_22_pad_groupi_n_31 ,csa_tree_add_95_22_pad_groupi_n_241);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6082(csa_tree_add_95_22_pad_groupi_n_30 ,csa_tree_add_95_22_pad_groupi_n_29);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6083(csa_tree_add_95_22_pad_groupi_n_29 ,csa_tree_add_95_22_pad_groupi_n_193);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6085(csa_tree_add_95_22_pad_groupi_n_28 ,csa_tree_add_95_22_pad_groupi_n_26);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6086(csa_tree_add_95_22_pad_groupi_n_27 ,csa_tree_add_95_22_pad_groupi_n_26);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6087(csa_tree_add_95_22_pad_groupi_n_26 ,csa_tree_add_95_22_pad_groupi_n_367);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6089(csa_tree_add_95_22_pad_groupi_n_25 ,csa_tree_add_95_22_pad_groupi_n_23);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6090(csa_tree_add_95_22_pad_groupi_n_24 ,csa_tree_add_95_22_pad_groupi_n_23);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6091(csa_tree_add_95_22_pad_groupi_n_23 ,csa_tree_add_95_22_pad_groupi_n_368);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6093(csa_tree_add_95_22_pad_groupi_n_22 ,csa_tree_add_95_22_pad_groupi_n_20);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6094(csa_tree_add_95_22_pad_groupi_n_21 ,csa_tree_add_95_22_pad_groupi_n_20);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6095(csa_tree_add_95_22_pad_groupi_n_20 ,csa_tree_add_95_22_pad_groupi_n_364);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6098(csa_tree_add_95_22_pad_groupi_n_19 ,csa_tree_add_95_22_pad_groupi_n_18);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6099(csa_tree_add_95_22_pad_groupi_n_18 ,csa_tree_add_95_22_pad_groupi_n_243);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6102(csa_tree_add_95_22_pad_groupi_n_17 ,csa_tree_add_95_22_pad_groupi_n_16);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6103(csa_tree_add_95_22_pad_groupi_n_16 ,csa_tree_add_95_22_pad_groupi_n_196);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6106(csa_tree_add_95_22_pad_groupi_n_15 ,csa_tree_add_95_22_pad_groupi_n_14);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6107(csa_tree_add_95_22_pad_groupi_n_14 ,csa_tree_add_95_22_pad_groupi_n_237);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6110(csa_tree_add_95_22_pad_groupi_n_13 ,csa_tree_add_95_22_pad_groupi_n_12);
  not csa_tree_add_95_22_pad_groupi_drc_bufs6111(csa_tree_add_95_22_pad_groupi_n_12 ,csa_tree_add_95_22_pad_groupi_n_240);
  xor csa_tree_add_95_22_pad_groupi_g2(n_279 ,csa_tree_add_95_22_pad_groupi_n_1537 ,csa_tree_add_95_22_pad_groupi_n_1520);
  xor csa_tree_add_95_22_pad_groupi_g6113(n_277 ,csa_tree_add_95_22_pad_groupi_n_1532 ,csa_tree_add_95_22_pad_groupi_n_1518);
  xor csa_tree_add_95_22_pad_groupi_g6114(n_274 ,csa_tree_add_95_22_pad_groupi_n_1524 ,csa_tree_add_95_22_pad_groupi_n_1482);
  xor csa_tree_add_95_22_pad_groupi_g6115(n_273 ,csa_tree_add_95_22_pad_groupi_n_1522 ,csa_tree_add_95_22_pad_groupi_n_1502);
  xor csa_tree_add_95_22_pad_groupi_g6116(n_272 ,csa_tree_add_95_22_pad_groupi_n_1515 ,csa_tree_add_95_22_pad_groupi_n_1461);
  xor csa_tree_add_95_22_pad_groupi_g6117(csa_tree_add_95_22_pad_groupi_n_6 ,csa_tree_add_95_22_pad_groupi_n_1368 ,csa_tree_add_95_22_pad_groupi_n_1406);
  xor csa_tree_add_95_22_pad_groupi_g6118(csa_tree_add_95_22_pad_groupi_n_5 ,csa_tree_add_95_22_pad_groupi_n_1332 ,csa_tree_add_95_22_pad_groupi_n_1350);
  xor csa_tree_add_95_22_pad_groupi_g6119(csa_tree_add_95_22_pad_groupi_n_4 ,csa_tree_add_95_22_pad_groupi_n_836 ,csa_tree_add_95_22_pad_groupi_n_0);
  xor csa_tree_add_95_22_pad_groupi_g6120(csa_tree_add_95_22_pad_groupi_n_3 ,csa_tree_add_95_22_pad_groupi_n_835 ,csa_tree_add_95_22_pad_groupi_n_948);
  xor csa_tree_add_95_22_pad_groupi_g6122(csa_tree_add_95_22_pad_groupi_n_1 ,csa_tree_add_95_22_pad_groupi_n_358 ,in17[9]);
  xor csa_tree_add_95_22_pad_groupi_g6123(csa_tree_add_95_22_pad_groupi_n_0 ,csa_tree_add_95_22_pad_groupi_n_357 ,in17[11]);
  xnor csa_tree_add_101_22_pad_groupi_g4151(n_238 ,csa_tree_add_101_22_pad_groupi_n_1336 ,csa_tree_add_101_22_pad_groupi_n_1558);
  or csa_tree_add_101_22_pad_groupi_g4152(csa_tree_add_101_22_pad_groupi_n_1558 ,csa_tree_add_101_22_pad_groupi_n_1393 ,csa_tree_add_101_22_pad_groupi_n_1556);
  xnor csa_tree_add_101_22_pad_groupi_g4153(n_237 ,csa_tree_add_101_22_pad_groupi_n_1555 ,csa_tree_add_101_22_pad_groupi_n_1404);
  and csa_tree_add_101_22_pad_groupi_g4154(csa_tree_add_101_22_pad_groupi_n_1556 ,csa_tree_add_101_22_pad_groupi_n_1389 ,csa_tree_add_101_22_pad_groupi_n_1555);
  or csa_tree_add_101_22_pad_groupi_g4155(csa_tree_add_101_22_pad_groupi_n_1555 ,csa_tree_add_101_22_pad_groupi_n_1407 ,csa_tree_add_101_22_pad_groupi_n_1553);
  xnor csa_tree_add_101_22_pad_groupi_g4156(n_236 ,csa_tree_add_101_22_pad_groupi_n_1552 ,csa_tree_add_101_22_pad_groupi_n_1434);
  and csa_tree_add_101_22_pad_groupi_g4157(csa_tree_add_101_22_pad_groupi_n_1553 ,csa_tree_add_101_22_pad_groupi_n_1410 ,csa_tree_add_101_22_pad_groupi_n_1552);
  or csa_tree_add_101_22_pad_groupi_g4158(csa_tree_add_101_22_pad_groupi_n_1552 ,csa_tree_add_101_22_pad_groupi_n_1453 ,csa_tree_add_101_22_pad_groupi_n_1550);
  xnor csa_tree_add_101_22_pad_groupi_g4159(n_235 ,csa_tree_add_101_22_pad_groupi_n_1549 ,csa_tree_add_101_22_pad_groupi_n_1462);
  and csa_tree_add_101_22_pad_groupi_g4160(csa_tree_add_101_22_pad_groupi_n_1550 ,csa_tree_add_101_22_pad_groupi_n_1459 ,csa_tree_add_101_22_pad_groupi_n_1549);
  or csa_tree_add_101_22_pad_groupi_g4161(csa_tree_add_101_22_pad_groupi_n_1549 ,csa_tree_add_101_22_pad_groupi_n_1463 ,csa_tree_add_101_22_pad_groupi_n_1547);
  xnor csa_tree_add_101_22_pad_groupi_g4162(n_234 ,csa_tree_add_101_22_pad_groupi_n_1546 ,csa_tree_add_101_22_pad_groupi_n_1483);
  nor csa_tree_add_101_22_pad_groupi_g4163(csa_tree_add_101_22_pad_groupi_n_1547 ,csa_tree_add_101_22_pad_groupi_n_1546 ,csa_tree_add_101_22_pad_groupi_n_1464);
  and csa_tree_add_101_22_pad_groupi_g4164(csa_tree_add_101_22_pad_groupi_n_1546 ,csa_tree_add_101_22_pad_groupi_n_1500 ,csa_tree_add_101_22_pad_groupi_n_1544);
  xnor csa_tree_add_101_22_pad_groupi_g4165(n_233 ,csa_tree_add_101_22_pad_groupi_n_1542 ,csa_tree_add_101_22_pad_groupi_n_1501);
  or csa_tree_add_101_22_pad_groupi_g4166(csa_tree_add_101_22_pad_groupi_n_1544 ,csa_tree_add_101_22_pad_groupi_n_1494 ,csa_tree_add_101_22_pad_groupi_n_1543);
  not csa_tree_add_101_22_pad_groupi_g4167(csa_tree_add_101_22_pad_groupi_n_1543 ,csa_tree_add_101_22_pad_groupi_n_1542);
  or csa_tree_add_101_22_pad_groupi_g4168(csa_tree_add_101_22_pad_groupi_n_1542 ,csa_tree_add_101_22_pad_groupi_n_1499 ,csa_tree_add_101_22_pad_groupi_n_1540);
  xnor csa_tree_add_101_22_pad_groupi_g4169(n_232 ,csa_tree_add_101_22_pad_groupi_n_1539 ,csa_tree_add_101_22_pad_groupi_n_1503);
  nor csa_tree_add_101_22_pad_groupi_g4170(csa_tree_add_101_22_pad_groupi_n_1540 ,csa_tree_add_101_22_pad_groupi_n_1496 ,csa_tree_add_101_22_pad_groupi_n_1539);
  and csa_tree_add_101_22_pad_groupi_g4171(csa_tree_add_101_22_pad_groupi_n_1539 ,csa_tree_add_101_22_pad_groupi_n_1538 ,csa_tree_add_101_22_pad_groupi_n_1510);
  or csa_tree_add_101_22_pad_groupi_g4173(csa_tree_add_101_22_pad_groupi_n_1538 ,csa_tree_add_101_22_pad_groupi_n_1513 ,csa_tree_add_101_22_pad_groupi_n_1537);
  and csa_tree_add_101_22_pad_groupi_g4175(csa_tree_add_101_22_pad_groupi_n_1537 ,csa_tree_add_101_22_pad_groupi_n_1512 ,csa_tree_add_101_22_pad_groupi_n_1535);
  xnor csa_tree_add_101_22_pad_groupi_g4176(n_230 ,csa_tree_add_101_22_pad_groupi_n_1534 ,csa_tree_add_101_22_pad_groupi_n_1519);
  or csa_tree_add_101_22_pad_groupi_g4177(csa_tree_add_101_22_pad_groupi_n_1535 ,csa_tree_add_101_22_pad_groupi_n_1514 ,csa_tree_add_101_22_pad_groupi_n_1534);
  and csa_tree_add_101_22_pad_groupi_g4178(csa_tree_add_101_22_pad_groupi_n_1534 ,csa_tree_add_101_22_pad_groupi_n_1533 ,csa_tree_add_101_22_pad_groupi_n_1511);
  or csa_tree_add_101_22_pad_groupi_g4180(csa_tree_add_101_22_pad_groupi_n_1533 ,csa_tree_add_101_22_pad_groupi_n_1505 ,csa_tree_add_101_22_pad_groupi_n_1532);
  and csa_tree_add_101_22_pad_groupi_g4182(csa_tree_add_101_22_pad_groupi_n_1532 ,csa_tree_add_101_22_pad_groupi_n_1506 ,csa_tree_add_101_22_pad_groupi_n_1530);
  xnor csa_tree_add_101_22_pad_groupi_g4183(n_228 ,csa_tree_add_101_22_pad_groupi_n_1529 ,csa_tree_add_101_22_pad_groupi_n_1517);
  or csa_tree_add_101_22_pad_groupi_g4184(csa_tree_add_101_22_pad_groupi_n_1530 ,csa_tree_add_101_22_pad_groupi_n_1507 ,csa_tree_add_101_22_pad_groupi_n_1529);
  and csa_tree_add_101_22_pad_groupi_g4185(csa_tree_add_101_22_pad_groupi_n_1529 ,csa_tree_add_101_22_pad_groupi_n_1508 ,csa_tree_add_101_22_pad_groupi_n_1527);
  xnor csa_tree_add_101_22_pad_groupi_g4186(n_227 ,csa_tree_add_101_22_pad_groupi_n_1526 ,csa_tree_add_101_22_pad_groupi_n_1516);
  or csa_tree_add_101_22_pad_groupi_g4187(csa_tree_add_101_22_pad_groupi_n_1527 ,csa_tree_add_101_22_pad_groupi_n_1526 ,csa_tree_add_101_22_pad_groupi_n_1509);
  and csa_tree_add_101_22_pad_groupi_g4188(csa_tree_add_101_22_pad_groupi_n_1526 ,csa_tree_add_101_22_pad_groupi_n_1471 ,csa_tree_add_101_22_pad_groupi_n_1525);
  or csa_tree_add_101_22_pad_groupi_g4190(csa_tree_add_101_22_pad_groupi_n_1525 ,csa_tree_add_101_22_pad_groupi_n_1470 ,csa_tree_add_101_22_pad_groupi_n_1524);
  and csa_tree_add_101_22_pad_groupi_g4192(csa_tree_add_101_22_pad_groupi_n_1524 ,csa_tree_add_101_22_pad_groupi_n_1498 ,csa_tree_add_101_22_pad_groupi_n_1523);
  or csa_tree_add_101_22_pad_groupi_g4194(csa_tree_add_101_22_pad_groupi_n_1523 ,csa_tree_add_101_22_pad_groupi_n_1497 ,csa_tree_add_101_22_pad_groupi_n_1522);
  and csa_tree_add_101_22_pad_groupi_g4196(csa_tree_add_101_22_pad_groupi_n_1522 ,csa_tree_add_101_22_pad_groupi_n_1452 ,csa_tree_add_101_22_pad_groupi_n_1521);
  or csa_tree_add_101_22_pad_groupi_g4198(csa_tree_add_101_22_pad_groupi_n_1521 ,csa_tree_add_101_22_pad_groupi_n_1451 ,csa_tree_add_101_22_pad_groupi_n_1515);
  xnor csa_tree_add_101_22_pad_groupi_g4199(csa_tree_add_101_22_pad_groupi_n_1520 ,csa_tree_add_101_22_pad_groupi_n_1475 ,csa_tree_add_101_22_pad_groupi_n_1491);
  xnor csa_tree_add_101_22_pad_groupi_g4200(csa_tree_add_101_22_pad_groupi_n_1519 ,csa_tree_add_101_22_pad_groupi_n_1473 ,csa_tree_add_101_22_pad_groupi_n_1489);
  xnor csa_tree_add_101_22_pad_groupi_g4201(csa_tree_add_101_22_pad_groupi_n_1518 ,csa_tree_add_101_22_pad_groupi_n_1480 ,csa_tree_add_101_22_pad_groupi_n_1487);
  xnor csa_tree_add_101_22_pad_groupi_g4202(csa_tree_add_101_22_pad_groupi_n_1517 ,csa_tree_add_101_22_pad_groupi_n_1477 ,csa_tree_add_101_22_pad_groupi_n_1493);
  xnor csa_tree_add_101_22_pad_groupi_g4203(csa_tree_add_101_22_pad_groupi_n_1516 ,csa_tree_add_101_22_pad_groupi_n_1448 ,csa_tree_add_101_22_pad_groupi_n_1485);
  nor csa_tree_add_101_22_pad_groupi_g4205(csa_tree_add_101_22_pad_groupi_n_1514 ,csa_tree_add_101_22_pad_groupi_n_1472 ,csa_tree_add_101_22_pad_groupi_n_1489);
  nor csa_tree_add_101_22_pad_groupi_g4206(csa_tree_add_101_22_pad_groupi_n_1513 ,csa_tree_add_101_22_pad_groupi_n_1475 ,csa_tree_add_101_22_pad_groupi_n_1491);
  or csa_tree_add_101_22_pad_groupi_g4207(csa_tree_add_101_22_pad_groupi_n_1512 ,csa_tree_add_101_22_pad_groupi_n_1473 ,csa_tree_add_101_22_pad_groupi_n_1488);
  or csa_tree_add_101_22_pad_groupi_g4208(csa_tree_add_101_22_pad_groupi_n_1511 ,csa_tree_add_101_22_pad_groupi_n_1479 ,csa_tree_add_101_22_pad_groupi_n_1486);
  or csa_tree_add_101_22_pad_groupi_g4209(csa_tree_add_101_22_pad_groupi_n_1510 ,csa_tree_add_101_22_pad_groupi_n_1474 ,csa_tree_add_101_22_pad_groupi_n_1490);
  nor csa_tree_add_101_22_pad_groupi_g4210(csa_tree_add_101_22_pad_groupi_n_1509 ,csa_tree_add_101_22_pad_groupi_n_1447 ,csa_tree_add_101_22_pad_groupi_n_1485);
  and csa_tree_add_101_22_pad_groupi_g4211(csa_tree_add_101_22_pad_groupi_n_1515 ,csa_tree_add_101_22_pad_groupi_n_1450 ,csa_tree_add_101_22_pad_groupi_n_1495);
  or csa_tree_add_101_22_pad_groupi_g4212(csa_tree_add_101_22_pad_groupi_n_1508 ,csa_tree_add_101_22_pad_groupi_n_1448 ,csa_tree_add_101_22_pad_groupi_n_1484);
  nor csa_tree_add_101_22_pad_groupi_g4213(csa_tree_add_101_22_pad_groupi_n_1507 ,csa_tree_add_101_22_pad_groupi_n_1476 ,csa_tree_add_101_22_pad_groupi_n_1493);
  or csa_tree_add_101_22_pad_groupi_g4214(csa_tree_add_101_22_pad_groupi_n_1506 ,csa_tree_add_101_22_pad_groupi_n_1477 ,csa_tree_add_101_22_pad_groupi_n_1492);
  nor csa_tree_add_101_22_pad_groupi_g4215(csa_tree_add_101_22_pad_groupi_n_1505 ,csa_tree_add_101_22_pad_groupi_n_1480 ,csa_tree_add_101_22_pad_groupi_n_1487);
  xnor csa_tree_add_101_22_pad_groupi_g4216(n_223 ,csa_tree_add_101_22_pad_groupi_n_1481 ,csa_tree_add_101_22_pad_groupi_n_1460);
  xnor csa_tree_add_101_22_pad_groupi_g4217(csa_tree_add_101_22_pad_groupi_n_1503 ,csa_tree_add_101_22_pad_groupi_n_1478 ,csa_tree_add_101_22_pad_groupi_n_1467);
  xnor csa_tree_add_101_22_pad_groupi_g4218(csa_tree_add_101_22_pad_groupi_n_1502 ,csa_tree_add_101_22_pad_groupi_n_1412 ,csa_tree_add_101_22_pad_groupi_n_1466);
  xnor csa_tree_add_101_22_pad_groupi_g4219(csa_tree_add_101_22_pad_groupi_n_1501 ,csa_tree_add_101_22_pad_groupi_n_1442 ,csa_tree_add_101_22_pad_groupi_n_1469);
  or csa_tree_add_101_22_pad_groupi_g4220(csa_tree_add_101_22_pad_groupi_n_1500 ,csa_tree_add_101_22_pad_groupi_n_1441 ,csa_tree_add_101_22_pad_groupi_n_6);
  nor csa_tree_add_101_22_pad_groupi_g4221(csa_tree_add_101_22_pad_groupi_n_1499 ,csa_tree_add_101_22_pad_groupi_n_1478 ,csa_tree_add_101_22_pad_groupi_n_1468);
  or csa_tree_add_101_22_pad_groupi_g4222(csa_tree_add_101_22_pad_groupi_n_1498 ,csa_tree_add_101_22_pad_groupi_n_1411 ,csa_tree_add_101_22_pad_groupi_n_1465);
  nor csa_tree_add_101_22_pad_groupi_g4223(csa_tree_add_101_22_pad_groupi_n_1497 ,csa_tree_add_101_22_pad_groupi_n_1412 ,csa_tree_add_101_22_pad_groupi_n_1466);
  and csa_tree_add_101_22_pad_groupi_g4224(csa_tree_add_101_22_pad_groupi_n_1496 ,csa_tree_add_101_22_pad_groupi_n_1478 ,csa_tree_add_101_22_pad_groupi_n_1468);
  or csa_tree_add_101_22_pad_groupi_g4225(csa_tree_add_101_22_pad_groupi_n_1495 ,csa_tree_add_101_22_pad_groupi_n_1449 ,csa_tree_add_101_22_pad_groupi_n_1481);
  nor csa_tree_add_101_22_pad_groupi_g4226(csa_tree_add_101_22_pad_groupi_n_1494 ,csa_tree_add_101_22_pad_groupi_n_1442 ,csa_tree_add_101_22_pad_groupi_n_1469);
  not csa_tree_add_101_22_pad_groupi_g4227(csa_tree_add_101_22_pad_groupi_n_1493 ,csa_tree_add_101_22_pad_groupi_n_1492);
  not csa_tree_add_101_22_pad_groupi_g4228(csa_tree_add_101_22_pad_groupi_n_1491 ,csa_tree_add_101_22_pad_groupi_n_1490);
  not csa_tree_add_101_22_pad_groupi_g4229(csa_tree_add_101_22_pad_groupi_n_1489 ,csa_tree_add_101_22_pad_groupi_n_1488);
  not csa_tree_add_101_22_pad_groupi_g4230(csa_tree_add_101_22_pad_groupi_n_1487 ,csa_tree_add_101_22_pad_groupi_n_1486);
  not csa_tree_add_101_22_pad_groupi_g4231(csa_tree_add_101_22_pad_groupi_n_1485 ,csa_tree_add_101_22_pad_groupi_n_1484);
  xnor csa_tree_add_101_22_pad_groupi_g4232(csa_tree_add_101_22_pad_groupi_n_1483 ,csa_tree_add_101_22_pad_groupi_n_1440 ,csa_tree_add_101_22_pad_groupi_n_1445);
  xnor csa_tree_add_101_22_pad_groupi_g4233(csa_tree_add_101_22_pad_groupi_n_1482 ,csa_tree_add_101_22_pad_groupi_n_1419 ,csa_tree_add_101_22_pad_groupi_n_1444);
  xnor csa_tree_add_101_22_pad_groupi_g4234(csa_tree_add_101_22_pad_groupi_n_1492 ,csa_tree_add_101_22_pad_groupi_n_1387 ,csa_tree_add_101_22_pad_groupi_n_1438);
  xnor csa_tree_add_101_22_pad_groupi_g4235(csa_tree_add_101_22_pad_groupi_n_1490 ,csa_tree_add_101_22_pad_groupi_n_1400 ,csa_tree_add_101_22_pad_groupi_n_1433);
  xnor csa_tree_add_101_22_pad_groupi_g4236(csa_tree_add_101_22_pad_groupi_n_1488 ,csa_tree_add_101_22_pad_groupi_n_1401 ,csa_tree_add_101_22_pad_groupi_n_1436);
  xnor csa_tree_add_101_22_pad_groupi_g4237(csa_tree_add_101_22_pad_groupi_n_1486 ,csa_tree_add_101_22_pad_groupi_n_1402 ,csa_tree_add_101_22_pad_groupi_n_1437);
  xnor csa_tree_add_101_22_pad_groupi_g4238(csa_tree_add_101_22_pad_groupi_n_1484 ,csa_tree_add_101_22_pad_groupi_n_1403 ,csa_tree_add_101_22_pad_groupi_n_1435);
  not csa_tree_add_101_22_pad_groupi_g4239(csa_tree_add_101_22_pad_groupi_n_1479 ,csa_tree_add_101_22_pad_groupi_n_1480);
  not csa_tree_add_101_22_pad_groupi_g4240(csa_tree_add_101_22_pad_groupi_n_1477 ,csa_tree_add_101_22_pad_groupi_n_1476);
  not csa_tree_add_101_22_pad_groupi_g4241(csa_tree_add_101_22_pad_groupi_n_1474 ,csa_tree_add_101_22_pad_groupi_n_1475);
  not csa_tree_add_101_22_pad_groupi_g4242(csa_tree_add_101_22_pad_groupi_n_1473 ,csa_tree_add_101_22_pad_groupi_n_1472);
  or csa_tree_add_101_22_pad_groupi_g4243(csa_tree_add_101_22_pad_groupi_n_1471 ,csa_tree_add_101_22_pad_groupi_n_1418 ,csa_tree_add_101_22_pad_groupi_n_1443);
  nor csa_tree_add_101_22_pad_groupi_g4244(csa_tree_add_101_22_pad_groupi_n_1470 ,csa_tree_add_101_22_pad_groupi_n_1419 ,csa_tree_add_101_22_pad_groupi_n_1444);
  and csa_tree_add_101_22_pad_groupi_g4245(csa_tree_add_101_22_pad_groupi_n_1481 ,csa_tree_add_101_22_pad_groupi_n_1371 ,csa_tree_add_101_22_pad_groupi_n_1439);
  or csa_tree_add_101_22_pad_groupi_g4246(csa_tree_add_101_22_pad_groupi_n_1480 ,csa_tree_add_101_22_pad_groupi_n_1424 ,csa_tree_add_101_22_pad_groupi_n_1456);
  and csa_tree_add_101_22_pad_groupi_g4247(csa_tree_add_101_22_pad_groupi_n_1478 ,csa_tree_add_101_22_pad_groupi_n_1431 ,csa_tree_add_101_22_pad_groupi_n_1454);
  or csa_tree_add_101_22_pad_groupi_g4248(csa_tree_add_101_22_pad_groupi_n_1476 ,csa_tree_add_101_22_pad_groupi_n_1422 ,csa_tree_add_101_22_pad_groupi_n_1455);
  or csa_tree_add_101_22_pad_groupi_g4249(csa_tree_add_101_22_pad_groupi_n_1475 ,csa_tree_add_101_22_pad_groupi_n_1429 ,csa_tree_add_101_22_pad_groupi_n_1458);
  or csa_tree_add_101_22_pad_groupi_g4250(csa_tree_add_101_22_pad_groupi_n_1472 ,csa_tree_add_101_22_pad_groupi_n_1426 ,csa_tree_add_101_22_pad_groupi_n_1457);
  not csa_tree_add_101_22_pad_groupi_g4251(csa_tree_add_101_22_pad_groupi_n_1469 ,csa_tree_add_101_22_pad_groupi_n_6);
  not csa_tree_add_101_22_pad_groupi_g4252(csa_tree_add_101_22_pad_groupi_n_1468 ,csa_tree_add_101_22_pad_groupi_n_1467);
  not csa_tree_add_101_22_pad_groupi_g4253(csa_tree_add_101_22_pad_groupi_n_1466 ,csa_tree_add_101_22_pad_groupi_n_1465);
  and csa_tree_add_101_22_pad_groupi_g4254(csa_tree_add_101_22_pad_groupi_n_1464 ,csa_tree_add_101_22_pad_groupi_n_1440 ,csa_tree_add_101_22_pad_groupi_n_1446);
  nor csa_tree_add_101_22_pad_groupi_g4255(csa_tree_add_101_22_pad_groupi_n_1463 ,csa_tree_add_101_22_pad_groupi_n_1440 ,csa_tree_add_101_22_pad_groupi_n_1446);
  xnor csa_tree_add_101_22_pad_groupi_g4256(csa_tree_add_101_22_pad_groupi_n_1462 ,csa_tree_add_101_22_pad_groupi_n_1432 ,csa_tree_add_101_22_pad_groupi_n_1413);
  xnor csa_tree_add_101_22_pad_groupi_g4257(csa_tree_add_101_22_pad_groupi_n_1461 ,csa_tree_add_101_22_pad_groupi_n_1397 ,csa_tree_add_101_22_pad_groupi_n_1417);
  xnor csa_tree_add_101_22_pad_groupi_g4258(csa_tree_add_101_22_pad_groupi_n_1460 ,csa_tree_add_101_22_pad_groupi_n_1367 ,csa_tree_add_101_22_pad_groupi_n_1415);
  xnor csa_tree_add_101_22_pad_groupi_g4260(csa_tree_add_101_22_pad_groupi_n_1467 ,csa_tree_add_101_22_pad_groupi_n_1384 ,csa_tree_add_101_22_pad_groupi_n_1405);
  xnor csa_tree_add_101_22_pad_groupi_g4261(csa_tree_add_101_22_pad_groupi_n_1465 ,csa_tree_add_101_22_pad_groupi_n_1295 ,csa_tree_add_101_22_pad_groupi_n_5);
  or csa_tree_add_101_22_pad_groupi_g4262(csa_tree_add_101_22_pad_groupi_n_1459 ,csa_tree_add_101_22_pad_groupi_n_1432 ,csa_tree_add_101_22_pad_groupi_n_1413);
  and csa_tree_add_101_22_pad_groupi_g4263(csa_tree_add_101_22_pad_groupi_n_1458 ,csa_tree_add_101_22_pad_groupi_n_1401 ,csa_tree_add_101_22_pad_groupi_n_1427);
  and csa_tree_add_101_22_pad_groupi_g4264(csa_tree_add_101_22_pad_groupi_n_1457 ,csa_tree_add_101_22_pad_groupi_n_1402 ,csa_tree_add_101_22_pad_groupi_n_1425);
  and csa_tree_add_101_22_pad_groupi_g4265(csa_tree_add_101_22_pad_groupi_n_1456 ,csa_tree_add_101_22_pad_groupi_n_1387 ,csa_tree_add_101_22_pad_groupi_n_1423);
  and csa_tree_add_101_22_pad_groupi_g4266(csa_tree_add_101_22_pad_groupi_n_1455 ,csa_tree_add_101_22_pad_groupi_n_1403 ,csa_tree_add_101_22_pad_groupi_n_1421);
  or csa_tree_add_101_22_pad_groupi_g4267(csa_tree_add_101_22_pad_groupi_n_1454 ,csa_tree_add_101_22_pad_groupi_n_1430 ,csa_tree_add_101_22_pad_groupi_n_1386);
  and csa_tree_add_101_22_pad_groupi_g4268(csa_tree_add_101_22_pad_groupi_n_1453 ,csa_tree_add_101_22_pad_groupi_n_1432 ,csa_tree_add_101_22_pad_groupi_n_1413);
  or csa_tree_add_101_22_pad_groupi_g4269(csa_tree_add_101_22_pad_groupi_n_1452 ,csa_tree_add_101_22_pad_groupi_n_1396 ,csa_tree_add_101_22_pad_groupi_n_1416);
  nor csa_tree_add_101_22_pad_groupi_g4270(csa_tree_add_101_22_pad_groupi_n_1451 ,csa_tree_add_101_22_pad_groupi_n_1397 ,csa_tree_add_101_22_pad_groupi_n_1417);
  or csa_tree_add_101_22_pad_groupi_g4271(csa_tree_add_101_22_pad_groupi_n_1450 ,csa_tree_add_101_22_pad_groupi_n_1367 ,csa_tree_add_101_22_pad_groupi_n_1414);
  nor csa_tree_add_101_22_pad_groupi_g4272(csa_tree_add_101_22_pad_groupi_n_1449 ,csa_tree_add_101_22_pad_groupi_n_1366 ,csa_tree_add_101_22_pad_groupi_n_1415);
  not csa_tree_add_101_22_pad_groupi_g4273(csa_tree_add_101_22_pad_groupi_n_1448 ,csa_tree_add_101_22_pad_groupi_n_1447);
  not csa_tree_add_101_22_pad_groupi_g4274(csa_tree_add_101_22_pad_groupi_n_1446 ,csa_tree_add_101_22_pad_groupi_n_1445);
  not csa_tree_add_101_22_pad_groupi_g4275(csa_tree_add_101_22_pad_groupi_n_1444 ,csa_tree_add_101_22_pad_groupi_n_1443);
  not csa_tree_add_101_22_pad_groupi_g4276(csa_tree_add_101_22_pad_groupi_n_1441 ,csa_tree_add_101_22_pad_groupi_n_1442);
  or csa_tree_add_101_22_pad_groupi_g4277(csa_tree_add_101_22_pad_groupi_n_1439 ,csa_tree_add_101_22_pad_groupi_n_1372 ,csa_tree_add_101_22_pad_groupi_n_1428);
  xnor csa_tree_add_101_22_pad_groupi_g4278(csa_tree_add_101_22_pad_groupi_n_1438 ,csa_tree_add_101_22_pad_groupi_n_1291 ,csa_tree_add_101_22_pad_groupi_n_1379);
  xnor csa_tree_add_101_22_pad_groupi_g4279(csa_tree_add_101_22_pad_groupi_n_1437 ,csa_tree_add_101_22_pad_groupi_n_1293 ,csa_tree_add_101_22_pad_groupi_n_1381);
  xnor csa_tree_add_101_22_pad_groupi_g4280(csa_tree_add_101_22_pad_groupi_n_1436 ,csa_tree_add_101_22_pad_groupi_n_1301 ,csa_tree_add_101_22_pad_groupi_n_1376);
  xnor csa_tree_add_101_22_pad_groupi_g4281(csa_tree_add_101_22_pad_groupi_n_1435 ,csa_tree_add_101_22_pad_groupi_n_1303 ,csa_tree_add_101_22_pad_groupi_n_1383);
  xnor csa_tree_add_101_22_pad_groupi_g4282(csa_tree_add_101_22_pad_groupi_n_1434 ,csa_tree_add_101_22_pad_groupi_n_1377 ,csa_tree_add_101_22_pad_groupi_n_1398);
  xnor csa_tree_add_101_22_pad_groupi_g4283(csa_tree_add_101_22_pad_groupi_n_1433 ,csa_tree_add_101_22_pad_groupi_n_1298 ,csa_tree_add_101_22_pad_groupi_n_1386);
  or csa_tree_add_101_22_pad_groupi_g4284(csa_tree_add_101_22_pad_groupi_n_1447 ,csa_tree_add_101_22_pad_groupi_n_1340 ,csa_tree_add_101_22_pad_groupi_n_1420);
  xnor csa_tree_add_101_22_pad_groupi_g4285(csa_tree_add_101_22_pad_groupi_n_1445 ,csa_tree_add_101_22_pad_groupi_n_1334 ,csa_tree_add_101_22_pad_groupi_n_1370);
  xnor csa_tree_add_101_22_pad_groupi_g4286(csa_tree_add_101_22_pad_groupi_n_1443 ,csa_tree_add_101_22_pad_groupi_n_1385 ,csa_tree_add_101_22_pad_groupi_n_1369);
  or csa_tree_add_101_22_pad_groupi_g4287(csa_tree_add_101_22_pad_groupi_n_1442 ,csa_tree_add_101_22_pad_groupi_n_1374 ,csa_tree_add_101_22_pad_groupi_n_1409);
  and csa_tree_add_101_22_pad_groupi_g4288(csa_tree_add_101_22_pad_groupi_n_1440 ,csa_tree_add_101_22_pad_groupi_n_1395 ,csa_tree_add_101_22_pad_groupi_n_1408);
  or csa_tree_add_101_22_pad_groupi_g4289(csa_tree_add_101_22_pad_groupi_n_1431 ,csa_tree_add_101_22_pad_groupi_n_1297 ,csa_tree_add_101_22_pad_groupi_n_1399);
  nor csa_tree_add_101_22_pad_groupi_g4290(csa_tree_add_101_22_pad_groupi_n_1430 ,csa_tree_add_101_22_pad_groupi_n_1298 ,csa_tree_add_101_22_pad_groupi_n_1400);
  nor csa_tree_add_101_22_pad_groupi_g4291(csa_tree_add_101_22_pad_groupi_n_1429 ,csa_tree_add_101_22_pad_groupi_n_1300 ,csa_tree_add_101_22_pad_groupi_n_1376);
  nor csa_tree_add_101_22_pad_groupi_g4292(csa_tree_add_101_22_pad_groupi_n_1428 ,csa_tree_add_101_22_pad_groupi_n_1363 ,csa_tree_add_101_22_pad_groupi_n_1394);
  or csa_tree_add_101_22_pad_groupi_g4293(csa_tree_add_101_22_pad_groupi_n_1427 ,csa_tree_add_101_22_pad_groupi_n_1301 ,csa_tree_add_101_22_pad_groupi_n_1375);
  nor csa_tree_add_101_22_pad_groupi_g4294(csa_tree_add_101_22_pad_groupi_n_1426 ,csa_tree_add_101_22_pad_groupi_n_1292 ,csa_tree_add_101_22_pad_groupi_n_1381);
  or csa_tree_add_101_22_pad_groupi_g4295(csa_tree_add_101_22_pad_groupi_n_1425 ,csa_tree_add_101_22_pad_groupi_n_1293 ,csa_tree_add_101_22_pad_groupi_n_1380);
  nor csa_tree_add_101_22_pad_groupi_g4296(csa_tree_add_101_22_pad_groupi_n_1424 ,csa_tree_add_101_22_pad_groupi_n_1290 ,csa_tree_add_101_22_pad_groupi_n_1379);
  or csa_tree_add_101_22_pad_groupi_g4297(csa_tree_add_101_22_pad_groupi_n_1423 ,csa_tree_add_101_22_pad_groupi_n_1291 ,csa_tree_add_101_22_pad_groupi_n_1378);
  nor csa_tree_add_101_22_pad_groupi_g4298(csa_tree_add_101_22_pad_groupi_n_1422 ,csa_tree_add_101_22_pad_groupi_n_1302 ,csa_tree_add_101_22_pad_groupi_n_1383);
  or csa_tree_add_101_22_pad_groupi_g4299(csa_tree_add_101_22_pad_groupi_n_1421 ,csa_tree_add_101_22_pad_groupi_n_1303 ,csa_tree_add_101_22_pad_groupi_n_1382);
  nor csa_tree_add_101_22_pad_groupi_g4300(csa_tree_add_101_22_pad_groupi_n_1420 ,csa_tree_add_101_22_pad_groupi_n_1355 ,csa_tree_add_101_22_pad_groupi_n_1385);
  or csa_tree_add_101_22_pad_groupi_g4301(csa_tree_add_101_22_pad_groupi_n_1432 ,csa_tree_add_101_22_pad_groupi_n_1365 ,csa_tree_add_101_22_pad_groupi_n_1391);
  not csa_tree_add_101_22_pad_groupi_g4302(csa_tree_add_101_22_pad_groupi_n_1419 ,csa_tree_add_101_22_pad_groupi_n_1418);
  not csa_tree_add_101_22_pad_groupi_g4303(csa_tree_add_101_22_pad_groupi_n_1417 ,csa_tree_add_101_22_pad_groupi_n_1416);
  not csa_tree_add_101_22_pad_groupi_g4304(csa_tree_add_101_22_pad_groupi_n_1415 ,csa_tree_add_101_22_pad_groupi_n_1414);
  not csa_tree_add_101_22_pad_groupi_g4305(csa_tree_add_101_22_pad_groupi_n_1412 ,csa_tree_add_101_22_pad_groupi_n_1411);
  or csa_tree_add_101_22_pad_groupi_g4306(csa_tree_add_101_22_pad_groupi_n_1410 ,csa_tree_add_101_22_pad_groupi_n_1377 ,csa_tree_add_101_22_pad_groupi_n_1398);
  nor csa_tree_add_101_22_pad_groupi_g4307(csa_tree_add_101_22_pad_groupi_n_1409 ,csa_tree_add_101_22_pad_groupi_n_1384 ,csa_tree_add_101_22_pad_groupi_n_1392);
  or csa_tree_add_101_22_pad_groupi_g4308(csa_tree_add_101_22_pad_groupi_n_1408 ,csa_tree_add_101_22_pad_groupi_n_1368 ,csa_tree_add_101_22_pad_groupi_n_1373);
  and csa_tree_add_101_22_pad_groupi_g4309(csa_tree_add_101_22_pad_groupi_n_1407 ,csa_tree_add_101_22_pad_groupi_n_1377 ,csa_tree_add_101_22_pad_groupi_n_1398);
  xnor csa_tree_add_101_22_pad_groupi_g4310(csa_tree_add_101_22_pad_groupi_n_1406 ,csa_tree_add_101_22_pad_groupi_n_1280 ,csa_tree_add_101_22_pad_groupi_n_1346);
  xnor csa_tree_add_101_22_pad_groupi_g4312(csa_tree_add_101_22_pad_groupi_n_1405 ,csa_tree_add_101_22_pad_groupi_n_1304 ,csa_tree_add_101_22_pad_groupi_n_1348);
  xnor csa_tree_add_101_22_pad_groupi_g4313(csa_tree_add_101_22_pad_groupi_n_1404 ,csa_tree_add_101_22_pad_groupi_n_1309 ,csa_tree_add_101_22_pad_groupi_n_1345);
  and csa_tree_add_101_22_pad_groupi_g4314(csa_tree_add_101_22_pad_groupi_n_1418 ,csa_tree_add_101_22_pad_groupi_n_1354 ,csa_tree_add_101_22_pad_groupi_n_1390);
  xnor csa_tree_add_101_22_pad_groupi_g4315(csa_tree_add_101_22_pad_groupi_n_1416 ,csa_tree_add_101_22_pad_groupi_n_1311 ,csa_tree_add_101_22_pad_groupi_n_1337);
  xnor csa_tree_add_101_22_pad_groupi_g4316(csa_tree_add_101_22_pad_groupi_n_1414 ,csa_tree_add_101_22_pad_groupi_n_1320 ,csa_tree_add_101_22_pad_groupi_n_1335);
  xnor csa_tree_add_101_22_pad_groupi_g4317(csa_tree_add_101_22_pad_groupi_n_1413 ,csa_tree_add_101_22_pad_groupi_n_1333 ,csa_tree_add_101_22_pad_groupi_n_1338);
  and csa_tree_add_101_22_pad_groupi_g4318(csa_tree_add_101_22_pad_groupi_n_1411 ,csa_tree_add_101_22_pad_groupi_n_1356 ,csa_tree_add_101_22_pad_groupi_n_1388);
  not csa_tree_add_101_22_pad_groupi_g4319(csa_tree_add_101_22_pad_groupi_n_1400 ,csa_tree_add_101_22_pad_groupi_n_1399);
  not csa_tree_add_101_22_pad_groupi_g4320(csa_tree_add_101_22_pad_groupi_n_1396 ,csa_tree_add_101_22_pad_groupi_n_1397);
  or csa_tree_add_101_22_pad_groupi_g4321(csa_tree_add_101_22_pad_groupi_n_1395 ,csa_tree_add_101_22_pad_groupi_n_1280 ,csa_tree_add_101_22_pad_groupi_n_1347);
  nor csa_tree_add_101_22_pad_groupi_g4322(csa_tree_add_101_22_pad_groupi_n_1394 ,csa_tree_add_101_22_pad_groupi_n_1362 ,csa_tree_add_101_22_pad_groupi_n_1361);
  and csa_tree_add_101_22_pad_groupi_g4323(csa_tree_add_101_22_pad_groupi_n_1393 ,csa_tree_add_101_22_pad_groupi_n_1309 ,csa_tree_add_101_22_pad_groupi_n_1345);
  and csa_tree_add_101_22_pad_groupi_g4324(csa_tree_add_101_22_pad_groupi_n_1392 ,csa_tree_add_101_22_pad_groupi_n_1304 ,csa_tree_add_101_22_pad_groupi_n_1349);
  and csa_tree_add_101_22_pad_groupi_g4325(csa_tree_add_101_22_pad_groupi_n_1391 ,csa_tree_add_101_22_pad_groupi_n_1334 ,csa_tree_add_101_22_pad_groupi_n_1360);
  or csa_tree_add_101_22_pad_groupi_g4326(csa_tree_add_101_22_pad_groupi_n_1390 ,csa_tree_add_101_22_pad_groupi_n_1353 ,csa_tree_add_101_22_pad_groupi_n_1350);
  or csa_tree_add_101_22_pad_groupi_g4327(csa_tree_add_101_22_pad_groupi_n_1389 ,csa_tree_add_101_22_pad_groupi_n_1309 ,csa_tree_add_101_22_pad_groupi_n_1345);
  or csa_tree_add_101_22_pad_groupi_g4328(csa_tree_add_101_22_pad_groupi_n_1388 ,csa_tree_add_101_22_pad_groupi_n_1305 ,csa_tree_add_101_22_pad_groupi_n_1342);
  or csa_tree_add_101_22_pad_groupi_g4329(csa_tree_add_101_22_pad_groupi_n_1403 ,csa_tree_add_101_22_pad_groupi_n_1246 ,csa_tree_add_101_22_pad_groupi_n_1359);
  or csa_tree_add_101_22_pad_groupi_g4330(csa_tree_add_101_22_pad_groupi_n_1402 ,csa_tree_add_101_22_pad_groupi_n_1230 ,csa_tree_add_101_22_pad_groupi_n_1343);
  or csa_tree_add_101_22_pad_groupi_g4331(csa_tree_add_101_22_pad_groupi_n_1401 ,csa_tree_add_101_22_pad_groupi_n_1232 ,csa_tree_add_101_22_pad_groupi_n_1339);
  and csa_tree_add_101_22_pad_groupi_g4332(csa_tree_add_101_22_pad_groupi_n_1399 ,csa_tree_add_101_22_pad_groupi_n_1254 ,csa_tree_add_101_22_pad_groupi_n_1364);
  or csa_tree_add_101_22_pad_groupi_g4333(csa_tree_add_101_22_pad_groupi_n_1398 ,csa_tree_add_101_22_pad_groupi_n_1329 ,csa_tree_add_101_22_pad_groupi_n_1357);
  or csa_tree_add_101_22_pad_groupi_g4334(csa_tree_add_101_22_pad_groupi_n_1397 ,csa_tree_add_101_22_pad_groupi_n_1323 ,csa_tree_add_101_22_pad_groupi_n_1358);
  not csa_tree_add_101_22_pad_groupi_g4335(csa_tree_add_101_22_pad_groupi_n_1383 ,csa_tree_add_101_22_pad_groupi_n_1382);
  not csa_tree_add_101_22_pad_groupi_g4336(csa_tree_add_101_22_pad_groupi_n_1381 ,csa_tree_add_101_22_pad_groupi_n_1380);
  not csa_tree_add_101_22_pad_groupi_g4337(csa_tree_add_101_22_pad_groupi_n_1379 ,csa_tree_add_101_22_pad_groupi_n_1378);
  not csa_tree_add_101_22_pad_groupi_g4338(csa_tree_add_101_22_pad_groupi_n_1376 ,csa_tree_add_101_22_pad_groupi_n_1375);
  nor csa_tree_add_101_22_pad_groupi_g4339(csa_tree_add_101_22_pad_groupi_n_1374 ,csa_tree_add_101_22_pad_groupi_n_1304 ,csa_tree_add_101_22_pad_groupi_n_1349);
  and csa_tree_add_101_22_pad_groupi_g4340(csa_tree_add_101_22_pad_groupi_n_1373 ,csa_tree_add_101_22_pad_groupi_n_1280 ,csa_tree_add_101_22_pad_groupi_n_1347);
  nor csa_tree_add_101_22_pad_groupi_g4341(csa_tree_add_101_22_pad_groupi_n_1372 ,csa_tree_add_101_22_pad_groupi_n_1306 ,csa_tree_add_101_22_pad_groupi_n_1352);
  or csa_tree_add_101_22_pad_groupi_g4342(csa_tree_add_101_22_pad_groupi_n_1371 ,csa_tree_add_101_22_pad_groupi_n_1307 ,csa_tree_add_101_22_pad_groupi_n_1351);
  xnor csa_tree_add_101_22_pad_groupi_g4343(csa_tree_add_101_22_pad_groupi_n_1370 ,csa_tree_add_101_22_pad_groupi_n_1261 ,csa_tree_add_101_22_pad_groupi_n_1310);
  xnor csa_tree_add_101_22_pad_groupi_g4344(csa_tree_add_101_22_pad_groupi_n_1369 ,csa_tree_add_101_22_pad_groupi_n_1299 ,csa_tree_add_101_22_pad_groupi_n_1330);
  or csa_tree_add_101_22_pad_groupi_g4345(csa_tree_add_101_22_pad_groupi_n_1387 ,csa_tree_add_101_22_pad_groupi_n_1227 ,csa_tree_add_101_22_pad_groupi_n_1341);
  xnor csa_tree_add_101_22_pad_groupi_g4346(csa_tree_add_101_22_pad_groupi_n_1386 ,csa_tree_add_101_22_pad_groupi_n_1317 ,csa_tree_add_101_22_pad_groupi_n_1273);
  xnor csa_tree_add_101_22_pad_groupi_g4347(csa_tree_add_101_22_pad_groupi_n_1385 ,csa_tree_add_101_22_pad_groupi_n_1316 ,csa_tree_add_101_22_pad_groupi_n_1268);
  and csa_tree_add_101_22_pad_groupi_g4348(csa_tree_add_101_22_pad_groupi_n_1384 ,csa_tree_add_101_22_pad_groupi_n_1225 ,csa_tree_add_101_22_pad_groupi_n_1344);
  xnor csa_tree_add_101_22_pad_groupi_g4349(csa_tree_add_101_22_pad_groupi_n_1382 ,csa_tree_add_101_22_pad_groupi_n_1313 ,csa_tree_add_101_22_pad_groupi_n_1266);
  xnor csa_tree_add_101_22_pad_groupi_g4350(csa_tree_add_101_22_pad_groupi_n_1380 ,csa_tree_add_101_22_pad_groupi_n_1315 ,csa_tree_add_101_22_pad_groupi_n_1270);
  xnor csa_tree_add_101_22_pad_groupi_g4351(csa_tree_add_101_22_pad_groupi_n_1378 ,csa_tree_add_101_22_pad_groupi_n_1314 ,csa_tree_add_101_22_pad_groupi_n_1267);
  xnor csa_tree_add_101_22_pad_groupi_g4352(csa_tree_add_101_22_pad_groupi_n_1377 ,csa_tree_add_101_22_pad_groupi_n_1262 ,csa_tree_add_101_22_pad_groupi_n_1308);
  xnor csa_tree_add_101_22_pad_groupi_g4353(csa_tree_add_101_22_pad_groupi_n_1375 ,csa_tree_add_101_22_pad_groupi_n_1318 ,csa_tree_add_101_22_pad_groupi_n_1271);
  not csa_tree_add_101_22_pad_groupi_g4355(csa_tree_add_101_22_pad_groupi_n_1367 ,csa_tree_add_101_22_pad_groupi_n_1366);
  and csa_tree_add_101_22_pad_groupi_g4356(csa_tree_add_101_22_pad_groupi_n_1365 ,csa_tree_add_101_22_pad_groupi_n_1261 ,csa_tree_add_101_22_pad_groupi_n_1310);
  or csa_tree_add_101_22_pad_groupi_g4357(csa_tree_add_101_22_pad_groupi_n_1364 ,csa_tree_add_101_22_pad_groupi_n_1224 ,csa_tree_add_101_22_pad_groupi_n_1319);
  and csa_tree_add_101_22_pad_groupi_g4358(csa_tree_add_101_22_pad_groupi_n_1363 ,csa_tree_add_101_22_pad_groupi_n_1265 ,csa_tree_add_101_22_pad_groupi_n_1321);
  nor csa_tree_add_101_22_pad_groupi_g4359(csa_tree_add_101_22_pad_groupi_n_1362 ,csa_tree_add_101_22_pad_groupi_n_1265 ,csa_tree_add_101_22_pad_groupi_n_1321);
  nor csa_tree_add_101_22_pad_groupi_g4360(csa_tree_add_101_22_pad_groupi_n_1361 ,csa_tree_add_101_22_pad_groupi_n_1285 ,csa_tree_add_101_22_pad_groupi_n_1326);
  or csa_tree_add_101_22_pad_groupi_g4361(csa_tree_add_101_22_pad_groupi_n_1360 ,csa_tree_add_101_22_pad_groupi_n_1261 ,csa_tree_add_101_22_pad_groupi_n_1310);
  nor csa_tree_add_101_22_pad_groupi_g4362(csa_tree_add_101_22_pad_groupi_n_1359 ,csa_tree_add_101_22_pad_groupi_n_1245 ,csa_tree_add_101_22_pad_groupi_n_1316);
  nor csa_tree_add_101_22_pad_groupi_g4363(csa_tree_add_101_22_pad_groupi_n_1358 ,csa_tree_add_101_22_pad_groupi_n_1328 ,csa_tree_add_101_22_pad_groupi_n_1320);
  nor csa_tree_add_101_22_pad_groupi_g4364(csa_tree_add_101_22_pad_groupi_n_1357 ,csa_tree_add_101_22_pad_groupi_n_1333 ,csa_tree_add_101_22_pad_groupi_n_1322);
  or csa_tree_add_101_22_pad_groupi_g4365(csa_tree_add_101_22_pad_groupi_n_1356 ,csa_tree_add_101_22_pad_groupi_n_1278 ,csa_tree_add_101_22_pad_groupi_n_1312);
  nor csa_tree_add_101_22_pad_groupi_g4366(csa_tree_add_101_22_pad_groupi_n_1355 ,csa_tree_add_101_22_pad_groupi_n_1299 ,csa_tree_add_101_22_pad_groupi_n_1330);
  or csa_tree_add_101_22_pad_groupi_g4367(csa_tree_add_101_22_pad_groupi_n_1354 ,csa_tree_add_101_22_pad_groupi_n_1294 ,csa_tree_add_101_22_pad_groupi_n_1332);
  nor csa_tree_add_101_22_pad_groupi_g4368(csa_tree_add_101_22_pad_groupi_n_1353 ,csa_tree_add_101_22_pad_groupi_n_1295 ,csa_tree_add_101_22_pad_groupi_n_1331);
  and csa_tree_add_101_22_pad_groupi_g4369(csa_tree_add_101_22_pad_groupi_n_1368 ,csa_tree_add_101_22_pad_groupi_n_1243 ,csa_tree_add_101_22_pad_groupi_n_1324);
  or csa_tree_add_101_22_pad_groupi_g4370(csa_tree_add_101_22_pad_groupi_n_1366 ,csa_tree_add_101_22_pad_groupi_n_1185 ,csa_tree_add_101_22_pad_groupi_n_1327);
  not csa_tree_add_101_22_pad_groupi_g4371(csa_tree_add_101_22_pad_groupi_n_1352 ,csa_tree_add_101_22_pad_groupi_n_1351);
  not csa_tree_add_101_22_pad_groupi_g4373(csa_tree_add_101_22_pad_groupi_n_1349 ,csa_tree_add_101_22_pad_groupi_n_1348);
  not csa_tree_add_101_22_pad_groupi_g4374(csa_tree_add_101_22_pad_groupi_n_1347 ,csa_tree_add_101_22_pad_groupi_n_1346);
  or csa_tree_add_101_22_pad_groupi_g4375(csa_tree_add_101_22_pad_groupi_n_1344 ,csa_tree_add_101_22_pad_groupi_n_1223 ,csa_tree_add_101_22_pad_groupi_n_1317);
  and csa_tree_add_101_22_pad_groupi_g4376(csa_tree_add_101_22_pad_groupi_n_1343 ,csa_tree_add_101_22_pad_groupi_n_1228 ,csa_tree_add_101_22_pad_groupi_n_1314);
  and csa_tree_add_101_22_pad_groupi_g4377(csa_tree_add_101_22_pad_groupi_n_1342 ,csa_tree_add_101_22_pad_groupi_n_1278 ,csa_tree_add_101_22_pad_groupi_n_1312);
  and csa_tree_add_101_22_pad_groupi_g4378(csa_tree_add_101_22_pad_groupi_n_1341 ,csa_tree_add_101_22_pad_groupi_n_1226 ,csa_tree_add_101_22_pad_groupi_n_1313);
  and csa_tree_add_101_22_pad_groupi_g4379(csa_tree_add_101_22_pad_groupi_n_1340 ,csa_tree_add_101_22_pad_groupi_n_1299 ,csa_tree_add_101_22_pad_groupi_n_1330);
  and csa_tree_add_101_22_pad_groupi_g4380(csa_tree_add_101_22_pad_groupi_n_1339 ,csa_tree_add_101_22_pad_groupi_n_1231 ,csa_tree_add_101_22_pad_groupi_n_1315);
  xnor csa_tree_add_101_22_pad_groupi_g4381(csa_tree_add_101_22_pad_groupi_n_1338 ,csa_tree_add_101_22_pad_groupi_n_1201 ,csa_tree_add_101_22_pad_groupi_n_1279);
  xnor csa_tree_add_101_22_pad_groupi_g4382(csa_tree_add_101_22_pad_groupi_n_1351 ,csa_tree_add_101_22_pad_groupi_n_1281 ,csa_tree_add_101_22_pad_groupi_n_1211);
  xor csa_tree_add_101_22_pad_groupi_g4383(csa_tree_add_101_22_pad_groupi_n_1337 ,csa_tree_add_101_22_pad_groupi_n_1278 ,csa_tree_add_101_22_pad_groupi_n_1305);
  xnor csa_tree_add_101_22_pad_groupi_g4384(csa_tree_add_101_22_pad_groupi_n_1336 ,csa_tree_add_101_22_pad_groupi_n_1075 ,csa_tree_add_101_22_pad_groupi_n_1274);
  xnor csa_tree_add_101_22_pad_groupi_g4385(csa_tree_add_101_22_pad_groupi_n_1335 ,csa_tree_add_101_22_pad_groupi_n_1235 ,csa_tree_add_101_22_pad_groupi_n_1296);
  xnor csa_tree_add_101_22_pad_groupi_g4386(csa_tree_add_101_22_pad_groupi_n_1350 ,csa_tree_add_101_22_pad_groupi_n_1264 ,csa_tree_add_101_22_pad_groupi_n_1272);
  xnor csa_tree_add_101_22_pad_groupi_g4387(csa_tree_add_101_22_pad_groupi_n_1348 ,csa_tree_add_101_22_pad_groupi_n_1282 ,csa_tree_add_101_22_pad_groupi_n_1269);
  xnor csa_tree_add_101_22_pad_groupi_g4388(csa_tree_add_101_22_pad_groupi_n_1346 ,csa_tree_add_101_22_pad_groupi_n_1263 ,csa_tree_add_101_22_pad_groupi_n_1275);
  or csa_tree_add_101_22_pad_groupi_g4389(csa_tree_add_101_22_pad_groupi_n_1345 ,csa_tree_add_101_22_pad_groupi_n_1277 ,csa_tree_add_101_22_pad_groupi_n_1325);
  not csa_tree_add_101_22_pad_groupi_g4390(csa_tree_add_101_22_pad_groupi_n_1332 ,csa_tree_add_101_22_pad_groupi_n_1331);
  nor csa_tree_add_101_22_pad_groupi_g4391(csa_tree_add_101_22_pad_groupi_n_1329 ,csa_tree_add_101_22_pad_groupi_n_1202 ,csa_tree_add_101_22_pad_groupi_n_1279);
  nor csa_tree_add_101_22_pad_groupi_g4392(csa_tree_add_101_22_pad_groupi_n_1328 ,csa_tree_add_101_22_pad_groupi_n_1235 ,csa_tree_add_101_22_pad_groupi_n_1296);
  nor csa_tree_add_101_22_pad_groupi_g4393(csa_tree_add_101_22_pad_groupi_n_1327 ,csa_tree_add_101_22_pad_groupi_n_1184 ,csa_tree_add_101_22_pad_groupi_n_1281);
  nor csa_tree_add_101_22_pad_groupi_g4394(csa_tree_add_101_22_pad_groupi_n_1326 ,csa_tree_add_101_22_pad_groupi_n_1287 ,csa_tree_add_101_22_pad_groupi_n_1288);
  nor csa_tree_add_101_22_pad_groupi_g4395(csa_tree_add_101_22_pad_groupi_n_1325 ,csa_tree_add_101_22_pad_groupi_n_1276 ,csa_tree_add_101_22_pad_groupi_n_1262);
  or csa_tree_add_101_22_pad_groupi_g4396(csa_tree_add_101_22_pad_groupi_n_1324 ,csa_tree_add_101_22_pad_groupi_n_1252 ,csa_tree_add_101_22_pad_groupi_n_1283);
  and csa_tree_add_101_22_pad_groupi_g4397(csa_tree_add_101_22_pad_groupi_n_1323 ,csa_tree_add_101_22_pad_groupi_n_1235 ,csa_tree_add_101_22_pad_groupi_n_1296);
  and csa_tree_add_101_22_pad_groupi_g4398(csa_tree_add_101_22_pad_groupi_n_1322 ,csa_tree_add_101_22_pad_groupi_n_1202 ,csa_tree_add_101_22_pad_groupi_n_1279);
  or csa_tree_add_101_22_pad_groupi_g4399(csa_tree_add_101_22_pad_groupi_n_1334 ,csa_tree_add_101_22_pad_groupi_n_1240 ,csa_tree_add_101_22_pad_groupi_n_1284);
  and csa_tree_add_101_22_pad_groupi_g4400(csa_tree_add_101_22_pad_groupi_n_1333 ,csa_tree_add_101_22_pad_groupi_n_1156 ,csa_tree_add_101_22_pad_groupi_n_1286);
  xnor csa_tree_add_101_22_pad_groupi_g4401(csa_tree_add_101_22_pad_groupi_n_1331 ,csa_tree_add_101_22_pad_groupi_n_1039 ,csa_tree_add_101_22_pad_groupi_n_1216);
  or csa_tree_add_101_22_pad_groupi_g4402(csa_tree_add_101_22_pad_groupi_n_1330 ,csa_tree_add_101_22_pad_groupi_n_1242 ,csa_tree_add_101_22_pad_groupi_n_1289);
  not csa_tree_add_101_22_pad_groupi_g4403(csa_tree_add_101_22_pad_groupi_n_1319 ,csa_tree_add_101_22_pad_groupi_n_1318);
  not csa_tree_add_101_22_pad_groupi_g4404(csa_tree_add_101_22_pad_groupi_n_1312 ,csa_tree_add_101_22_pad_groupi_n_1311);
  xnor csa_tree_add_101_22_pad_groupi_g4405(csa_tree_add_101_22_pad_groupi_n_1321 ,csa_tree_add_101_22_pad_groupi_n_1176 ,csa_tree_add_101_22_pad_groupi_n_1210);
  xnor csa_tree_add_101_22_pad_groupi_g4406(csa_tree_add_101_22_pad_groupi_n_1308 ,csa_tree_add_101_22_pad_groupi_n_1132 ,csa_tree_add_101_22_pad_groupi_n_1233);
  xnor csa_tree_add_101_22_pad_groupi_g4407(csa_tree_add_101_22_pad_groupi_n_1320 ,csa_tree_add_101_22_pad_groupi_n_1084 ,csa_tree_add_101_22_pad_groupi_n_1220);
  xnor csa_tree_add_101_22_pad_groupi_g4408(csa_tree_add_101_22_pad_groupi_n_1318 ,csa_tree_add_101_22_pad_groupi_n_1138 ,csa_tree_add_101_22_pad_groupi_n_1221);
  xnor csa_tree_add_101_22_pad_groupi_g4409(csa_tree_add_101_22_pad_groupi_n_1317 ,csa_tree_add_101_22_pad_groupi_n_1092 ,csa_tree_add_101_22_pad_groupi_n_1213);
  xnor csa_tree_add_101_22_pad_groupi_g4410(csa_tree_add_101_22_pad_groupi_n_1316 ,csa_tree_add_101_22_pad_groupi_n_1088 ,csa_tree_add_101_22_pad_groupi_n_1214);
  xnor csa_tree_add_101_22_pad_groupi_g4411(csa_tree_add_101_22_pad_groupi_n_1315 ,csa_tree_add_101_22_pad_groupi_n_1141 ,csa_tree_add_101_22_pad_groupi_n_1218);
  xnor csa_tree_add_101_22_pad_groupi_g4412(csa_tree_add_101_22_pad_groupi_n_1314 ,csa_tree_add_101_22_pad_groupi_n_1102 ,csa_tree_add_101_22_pad_groupi_n_1217);
  xnor csa_tree_add_101_22_pad_groupi_g4413(csa_tree_add_101_22_pad_groupi_n_1313 ,csa_tree_add_101_22_pad_groupi_n_1107 ,csa_tree_add_101_22_pad_groupi_n_1222);
  xnor csa_tree_add_101_22_pad_groupi_g4414(csa_tree_add_101_22_pad_groupi_n_1311 ,csa_tree_add_101_22_pad_groupi_n_1209 ,csa_tree_add_101_22_pad_groupi_n_1215);
  xnor csa_tree_add_101_22_pad_groupi_g4415(csa_tree_add_101_22_pad_groupi_n_1310 ,csa_tree_add_101_22_pad_groupi_n_1236 ,csa_tree_add_101_22_pad_groupi_n_1212);
  xnor csa_tree_add_101_22_pad_groupi_g4416(csa_tree_add_101_22_pad_groupi_n_1309 ,csa_tree_add_101_22_pad_groupi_n_1175 ,csa_tree_add_101_22_pad_groupi_n_1219);
  not csa_tree_add_101_22_pad_groupi_g4417(csa_tree_add_101_22_pad_groupi_n_1307 ,csa_tree_add_101_22_pad_groupi_n_1306);
  not csa_tree_add_101_22_pad_groupi_g4418(csa_tree_add_101_22_pad_groupi_n_1302 ,csa_tree_add_101_22_pad_groupi_n_1303);
  not csa_tree_add_101_22_pad_groupi_g4419(csa_tree_add_101_22_pad_groupi_n_1300 ,csa_tree_add_101_22_pad_groupi_n_1301);
  not csa_tree_add_101_22_pad_groupi_g4420(csa_tree_add_101_22_pad_groupi_n_1297 ,csa_tree_add_101_22_pad_groupi_n_1298);
  not csa_tree_add_101_22_pad_groupi_g4421(csa_tree_add_101_22_pad_groupi_n_1295 ,csa_tree_add_101_22_pad_groupi_n_1294);
  not csa_tree_add_101_22_pad_groupi_g4422(csa_tree_add_101_22_pad_groupi_n_1292 ,csa_tree_add_101_22_pad_groupi_n_1293);
  not csa_tree_add_101_22_pad_groupi_g4423(csa_tree_add_101_22_pad_groupi_n_1290 ,csa_tree_add_101_22_pad_groupi_n_1291);
  nor csa_tree_add_101_22_pad_groupi_g4424(csa_tree_add_101_22_pad_groupi_n_1289 ,csa_tree_add_101_22_pad_groupi_n_1247 ,csa_tree_add_101_22_pad_groupi_n_1264);
  nor csa_tree_add_101_22_pad_groupi_g4425(csa_tree_add_101_22_pad_groupi_n_1288 ,csa_tree_add_101_22_pad_groupi_n_1048 ,csa_tree_add_101_22_pad_groupi_n_1238);
  nor csa_tree_add_101_22_pad_groupi_g4426(csa_tree_add_101_22_pad_groupi_n_1287 ,csa_tree_add_101_22_pad_groupi_n_1178 ,csa_tree_add_101_22_pad_groupi_n_1251);
  or csa_tree_add_101_22_pad_groupi_g4427(csa_tree_add_101_22_pad_groupi_n_1286 ,csa_tree_add_101_22_pad_groupi_n_1150 ,csa_tree_add_101_22_pad_groupi_n_1237);
  nor csa_tree_add_101_22_pad_groupi_g4428(csa_tree_add_101_22_pad_groupi_n_1285 ,csa_tree_add_101_22_pad_groupi_n_1047 ,csa_tree_add_101_22_pad_groupi_n_1239);
  and csa_tree_add_101_22_pad_groupi_g4429(csa_tree_add_101_22_pad_groupi_n_1284 ,csa_tree_add_101_22_pad_groupi_n_1241 ,csa_tree_add_101_22_pad_groupi_n_1263);
  or csa_tree_add_101_22_pad_groupi_g4430(csa_tree_add_101_22_pad_groupi_n_1306 ,csa_tree_add_101_22_pad_groupi_n_1183 ,csa_tree_add_101_22_pad_groupi_n_1253);
  and csa_tree_add_101_22_pad_groupi_g4431(csa_tree_add_101_22_pad_groupi_n_1305 ,csa_tree_add_101_22_pad_groupi_n_1192 ,csa_tree_add_101_22_pad_groupi_n_1257);
  and csa_tree_add_101_22_pad_groupi_g4432(csa_tree_add_101_22_pad_groupi_n_1304 ,csa_tree_add_101_22_pad_groupi_n_1155 ,csa_tree_add_101_22_pad_groupi_n_1260);
  or csa_tree_add_101_22_pad_groupi_g4433(csa_tree_add_101_22_pad_groupi_n_1303 ,csa_tree_add_101_22_pad_groupi_n_1154 ,csa_tree_add_101_22_pad_groupi_n_1248);
  or csa_tree_add_101_22_pad_groupi_g4434(csa_tree_add_101_22_pad_groupi_n_1301 ,csa_tree_add_101_22_pad_groupi_n_1187 ,csa_tree_add_101_22_pad_groupi_n_1255);
  or csa_tree_add_101_22_pad_groupi_g4435(csa_tree_add_101_22_pad_groupi_n_1299 ,csa_tree_add_101_22_pad_groupi_n_1147 ,csa_tree_add_101_22_pad_groupi_n_1244);
  or csa_tree_add_101_22_pad_groupi_g4436(csa_tree_add_101_22_pad_groupi_n_1298 ,csa_tree_add_101_22_pad_groupi_n_1198 ,csa_tree_add_101_22_pad_groupi_n_1258);
  or csa_tree_add_101_22_pad_groupi_g4437(csa_tree_add_101_22_pad_groupi_n_1296 ,csa_tree_add_101_22_pad_groupi_n_1188 ,csa_tree_add_101_22_pad_groupi_n_1256);
  and csa_tree_add_101_22_pad_groupi_g4438(csa_tree_add_101_22_pad_groupi_n_1294 ,csa_tree_add_101_22_pad_groupi_n_1197 ,csa_tree_add_101_22_pad_groupi_n_1259);
  or csa_tree_add_101_22_pad_groupi_g4439(csa_tree_add_101_22_pad_groupi_n_1293 ,csa_tree_add_101_22_pad_groupi_n_1179 ,csa_tree_add_101_22_pad_groupi_n_1250);
  or csa_tree_add_101_22_pad_groupi_g4440(csa_tree_add_101_22_pad_groupi_n_1291 ,csa_tree_add_101_22_pad_groupi_n_1200 ,csa_tree_add_101_22_pad_groupi_n_1249);
  not csa_tree_add_101_22_pad_groupi_g4441(csa_tree_add_101_22_pad_groupi_n_1283 ,csa_tree_add_101_22_pad_groupi_n_1282);
  nor csa_tree_add_101_22_pad_groupi_g4442(csa_tree_add_101_22_pad_groupi_n_1277 ,csa_tree_add_101_22_pad_groupi_n_1132 ,csa_tree_add_101_22_pad_groupi_n_1234);
  and csa_tree_add_101_22_pad_groupi_g4443(csa_tree_add_101_22_pad_groupi_n_1276 ,csa_tree_add_101_22_pad_groupi_n_1132 ,csa_tree_add_101_22_pad_groupi_n_1234);
  xnor csa_tree_add_101_22_pad_groupi_g4444(csa_tree_add_101_22_pad_groupi_n_1275 ,csa_tree_add_101_22_pad_groupi_n_1207 ,csa_tree_add_101_22_pad_groupi_n_1098);
  nor csa_tree_add_101_22_pad_groupi_g4445(csa_tree_add_101_22_pad_groupi_n_1274 ,csa_tree_add_101_22_pad_groupi_n_1157 ,csa_tree_add_101_22_pad_groupi_n_1229);
  xnor csa_tree_add_101_22_pad_groupi_g4446(csa_tree_add_101_22_pad_groupi_n_1273 ,csa_tree_add_101_22_pad_groupi_n_1163 ,csa_tree_add_101_22_pad_groupi_n_1166);
  xnor csa_tree_add_101_22_pad_groupi_g4447(csa_tree_add_101_22_pad_groupi_n_1272 ,csa_tree_add_101_22_pad_groupi_n_1099 ,csa_tree_add_101_22_pad_groupi_n_1169);
  xnor csa_tree_add_101_22_pad_groupi_g4448(csa_tree_add_101_22_pad_groupi_n_1271 ,csa_tree_add_101_22_pad_groupi_n_1204 ,csa_tree_add_101_22_pad_groupi_n_1160);
  xnor csa_tree_add_101_22_pad_groupi_g4449(csa_tree_add_101_22_pad_groupi_n_1270 ,csa_tree_add_101_22_pad_groupi_n_1208 ,csa_tree_add_101_22_pad_groupi_n_1174);
  xnor csa_tree_add_101_22_pad_groupi_g4450(csa_tree_add_101_22_pad_groupi_n_1269 ,csa_tree_add_101_22_pad_groupi_n_1206 ,csa_tree_add_101_22_pad_groupi_n_1171);
  xnor csa_tree_add_101_22_pad_groupi_g4451(csa_tree_add_101_22_pad_groupi_n_1268 ,csa_tree_add_101_22_pad_groupi_n_1164 ,csa_tree_add_101_22_pad_groupi_n_1167);
  xnor csa_tree_add_101_22_pad_groupi_g4452(csa_tree_add_101_22_pad_groupi_n_1267 ,csa_tree_add_101_22_pad_groupi_n_1173 ,csa_tree_add_101_22_pad_groupi_n_1172);
  xnor csa_tree_add_101_22_pad_groupi_g4453(csa_tree_add_101_22_pad_groupi_n_1266 ,csa_tree_add_101_22_pad_groupi_n_1161 ,csa_tree_add_101_22_pad_groupi_n_1168);
  xnor csa_tree_add_101_22_pad_groupi_g4454(csa_tree_add_101_22_pad_groupi_n_1282 ,csa_tree_add_101_22_pad_groupi_n_1106 ,csa_tree_add_101_22_pad_groupi_n_1143);
  xnor csa_tree_add_101_22_pad_groupi_g4455(csa_tree_add_101_22_pad_groupi_n_1281 ,csa_tree_add_101_22_pad_groupi_n_1080 ,csa_tree_add_101_22_pad_groupi_n_1145);
  xnor csa_tree_add_101_22_pad_groupi_g4456(csa_tree_add_101_22_pad_groupi_n_1280 ,csa_tree_add_101_22_pad_groupi_n_1103 ,csa_tree_add_101_22_pad_groupi_n_1146);
  xnor csa_tree_add_101_22_pad_groupi_g4457(csa_tree_add_101_22_pad_groupi_n_1279 ,csa_tree_add_101_22_pad_groupi_n_1101 ,csa_tree_add_101_22_pad_groupi_n_1142);
  xnor csa_tree_add_101_22_pad_groupi_g4458(csa_tree_add_101_22_pad_groupi_n_1278 ,csa_tree_add_101_22_pad_groupi_n_1105 ,csa_tree_add_101_22_pad_groupi_n_1144);
  or csa_tree_add_101_22_pad_groupi_g4459(csa_tree_add_101_22_pad_groupi_n_1260 ,csa_tree_add_101_22_pad_groupi_n_1104 ,csa_tree_add_101_22_pad_groupi_n_1151);
  or csa_tree_add_101_22_pad_groupi_g4460(csa_tree_add_101_22_pad_groupi_n_1259 ,csa_tree_add_101_22_pad_groupi_n_1209 ,csa_tree_add_101_22_pad_groupi_n_1193);
  nor csa_tree_add_101_22_pad_groupi_g4461(csa_tree_add_101_22_pad_groupi_n_1258 ,csa_tree_add_101_22_pad_groupi_n_1074 ,csa_tree_add_101_22_pad_groupi_n_1195);
  or csa_tree_add_101_22_pad_groupi_g4462(csa_tree_add_101_22_pad_groupi_n_1257 ,csa_tree_add_101_22_pad_groupi_n_1072 ,csa_tree_add_101_22_pad_groupi_n_1190);
  nor csa_tree_add_101_22_pad_groupi_g4463(csa_tree_add_101_22_pad_groupi_n_1256 ,csa_tree_add_101_22_pad_groupi_n_1067 ,csa_tree_add_101_22_pad_groupi_n_1186);
  and csa_tree_add_101_22_pad_groupi_g4464(csa_tree_add_101_22_pad_groupi_n_1255 ,csa_tree_add_101_22_pad_groupi_n_1141 ,csa_tree_add_101_22_pad_groupi_n_1189);
  or csa_tree_add_101_22_pad_groupi_g4465(csa_tree_add_101_22_pad_groupi_n_1254 ,csa_tree_add_101_22_pad_groupi_n_1203 ,csa_tree_add_101_22_pad_groupi_n_1159);
  and csa_tree_add_101_22_pad_groupi_g4466(csa_tree_add_101_22_pad_groupi_n_1253 ,csa_tree_add_101_22_pad_groupi_n_1181 ,csa_tree_add_101_22_pad_groupi_n_1176);
  nor csa_tree_add_101_22_pad_groupi_g4467(csa_tree_add_101_22_pad_groupi_n_1252 ,csa_tree_add_101_22_pad_groupi_n_1206 ,csa_tree_add_101_22_pad_groupi_n_1171);
  nor csa_tree_add_101_22_pad_groupi_g4468(csa_tree_add_101_22_pad_groupi_n_1251 ,csa_tree_add_101_22_pad_groupi_n_1177 ,csa_tree_add_101_22_pad_groupi_n_1191);
  and csa_tree_add_101_22_pad_groupi_g4469(csa_tree_add_101_22_pad_groupi_n_1250 ,csa_tree_add_101_22_pad_groupi_n_1102 ,csa_tree_add_101_22_pad_groupi_n_1194);
  and csa_tree_add_101_22_pad_groupi_g4470(csa_tree_add_101_22_pad_groupi_n_1249 ,csa_tree_add_101_22_pad_groupi_n_1107 ,csa_tree_add_101_22_pad_groupi_n_1158);
  nor csa_tree_add_101_22_pad_groupi_g4471(csa_tree_add_101_22_pad_groupi_n_1248 ,csa_tree_add_101_22_pad_groupi_n_1042 ,csa_tree_add_101_22_pad_groupi_n_1153);
  nor csa_tree_add_101_22_pad_groupi_g4472(csa_tree_add_101_22_pad_groupi_n_1247 ,csa_tree_add_101_22_pad_groupi_n_1099 ,csa_tree_add_101_22_pad_groupi_n_1169);
  and csa_tree_add_101_22_pad_groupi_g4473(csa_tree_add_101_22_pad_groupi_n_1246 ,csa_tree_add_101_22_pad_groupi_n_1164 ,csa_tree_add_101_22_pad_groupi_n_1167);
  nor csa_tree_add_101_22_pad_groupi_g4474(csa_tree_add_101_22_pad_groupi_n_1245 ,csa_tree_add_101_22_pad_groupi_n_1164 ,csa_tree_add_101_22_pad_groupi_n_1167);
  nor csa_tree_add_101_22_pad_groupi_g4475(csa_tree_add_101_22_pad_groupi_n_1244 ,csa_tree_add_101_22_pad_groupi_n_1039 ,csa_tree_add_101_22_pad_groupi_n_1148);
  or csa_tree_add_101_22_pad_groupi_g4476(csa_tree_add_101_22_pad_groupi_n_1243 ,csa_tree_add_101_22_pad_groupi_n_1205 ,csa_tree_add_101_22_pad_groupi_n_1170);
  and csa_tree_add_101_22_pad_groupi_g4477(csa_tree_add_101_22_pad_groupi_n_1242 ,csa_tree_add_101_22_pad_groupi_n_1099 ,csa_tree_add_101_22_pad_groupi_n_1169);
  or csa_tree_add_101_22_pad_groupi_g4478(csa_tree_add_101_22_pad_groupi_n_1241 ,csa_tree_add_101_22_pad_groupi_n_1207 ,csa_tree_add_101_22_pad_groupi_n_1098);
  and csa_tree_add_101_22_pad_groupi_g4479(csa_tree_add_101_22_pad_groupi_n_1240 ,csa_tree_add_101_22_pad_groupi_n_1207 ,csa_tree_add_101_22_pad_groupi_n_1098);
  or csa_tree_add_101_22_pad_groupi_g4480(csa_tree_add_101_22_pad_groupi_n_1265 ,csa_tree_add_101_22_pad_groupi_n_1051 ,csa_tree_add_101_22_pad_groupi_n_1180);
  and csa_tree_add_101_22_pad_groupi_g4481(csa_tree_add_101_22_pad_groupi_n_1264 ,csa_tree_add_101_22_pad_groupi_n_1115 ,csa_tree_add_101_22_pad_groupi_n_1199);
  or csa_tree_add_101_22_pad_groupi_g4482(csa_tree_add_101_22_pad_groupi_n_1263 ,csa_tree_add_101_22_pad_groupi_n_1123 ,csa_tree_add_101_22_pad_groupi_n_1182);
  and csa_tree_add_101_22_pad_groupi_g4483(csa_tree_add_101_22_pad_groupi_n_1262 ,csa_tree_add_101_22_pad_groupi_n_1114 ,csa_tree_add_101_22_pad_groupi_n_1149);
  or csa_tree_add_101_22_pad_groupi_g4484(csa_tree_add_101_22_pad_groupi_n_1261 ,csa_tree_add_101_22_pad_groupi_n_1124 ,csa_tree_add_101_22_pad_groupi_n_1196);
  not csa_tree_add_101_22_pad_groupi_g4485(csa_tree_add_101_22_pad_groupi_n_1239 ,csa_tree_add_101_22_pad_groupi_n_1238);
  not csa_tree_add_101_22_pad_groupi_g4486(csa_tree_add_101_22_pad_groupi_n_1237 ,csa_tree_add_101_22_pad_groupi_n_1236);
  not csa_tree_add_101_22_pad_groupi_g4487(csa_tree_add_101_22_pad_groupi_n_1234 ,csa_tree_add_101_22_pad_groupi_n_1233);
  and csa_tree_add_101_22_pad_groupi_g4488(csa_tree_add_101_22_pad_groupi_n_1232 ,csa_tree_add_101_22_pad_groupi_n_1208 ,csa_tree_add_101_22_pad_groupi_n_1174);
  or csa_tree_add_101_22_pad_groupi_g4489(csa_tree_add_101_22_pad_groupi_n_1231 ,csa_tree_add_101_22_pad_groupi_n_1208 ,csa_tree_add_101_22_pad_groupi_n_1174);
  and csa_tree_add_101_22_pad_groupi_g4490(csa_tree_add_101_22_pad_groupi_n_1230 ,csa_tree_add_101_22_pad_groupi_n_1173 ,csa_tree_add_101_22_pad_groupi_n_1172);
  nor csa_tree_add_101_22_pad_groupi_g4491(csa_tree_add_101_22_pad_groupi_n_1229 ,csa_tree_add_101_22_pad_groupi_n_1152 ,csa_tree_add_101_22_pad_groupi_n_1175);
  or csa_tree_add_101_22_pad_groupi_g4492(csa_tree_add_101_22_pad_groupi_n_1228 ,csa_tree_add_101_22_pad_groupi_n_1173 ,csa_tree_add_101_22_pad_groupi_n_1172);
  and csa_tree_add_101_22_pad_groupi_g4493(csa_tree_add_101_22_pad_groupi_n_1227 ,csa_tree_add_101_22_pad_groupi_n_1161 ,csa_tree_add_101_22_pad_groupi_n_1168);
  or csa_tree_add_101_22_pad_groupi_g4494(csa_tree_add_101_22_pad_groupi_n_1226 ,csa_tree_add_101_22_pad_groupi_n_1161 ,csa_tree_add_101_22_pad_groupi_n_1168);
  or csa_tree_add_101_22_pad_groupi_g4495(csa_tree_add_101_22_pad_groupi_n_1225 ,csa_tree_add_101_22_pad_groupi_n_1162 ,csa_tree_add_101_22_pad_groupi_n_1165);
  nor csa_tree_add_101_22_pad_groupi_g4496(csa_tree_add_101_22_pad_groupi_n_1224 ,csa_tree_add_101_22_pad_groupi_n_1204 ,csa_tree_add_101_22_pad_groupi_n_1160);
  nor csa_tree_add_101_22_pad_groupi_g4497(csa_tree_add_101_22_pad_groupi_n_1223 ,csa_tree_add_101_22_pad_groupi_n_1163 ,csa_tree_add_101_22_pad_groupi_n_1166);
  xnor csa_tree_add_101_22_pad_groupi_g4498(csa_tree_add_101_22_pad_groupi_n_1222 ,csa_tree_add_101_22_pad_groupi_n_1035 ,csa_tree_add_101_22_pad_groupi_n_1094);
  xnor csa_tree_add_101_22_pad_groupi_g4499(csa_tree_add_101_22_pad_groupi_n_1221 ,csa_tree_add_101_22_pad_groupi_n_1100 ,csa_tree_add_101_22_pad_groupi_n_1074);
  xnor csa_tree_add_101_22_pad_groupi_g4500(csa_tree_add_101_22_pad_groupi_n_1220 ,csa_tree_add_101_22_pad_groupi_n_1072 ,csa_tree_add_101_22_pad_groupi_n_1090);
  xnor csa_tree_add_101_22_pad_groupi_g4501(csa_tree_add_101_22_pad_groupi_n_1219 ,csa_tree_add_101_22_pad_groupi_n_1016 ,csa_tree_add_101_22_pad_groupi_n_1097);
  xnor csa_tree_add_101_22_pad_groupi_g4502(csa_tree_add_101_22_pad_groupi_n_1218 ,csa_tree_add_101_22_pad_groupi_n_1056 ,csa_tree_add_101_22_pad_groupi_n_3);
  xnor csa_tree_add_101_22_pad_groupi_g4503(csa_tree_add_101_22_pad_groupi_n_1238 ,csa_tree_add_101_22_pad_groupi_n_1140 ,csa_tree_add_101_22_pad_groupi_n_1076);
  xnor csa_tree_add_101_22_pad_groupi_g4504(csa_tree_add_101_22_pad_groupi_n_1217 ,csa_tree_add_101_22_pad_groupi_n_1055 ,csa_tree_add_101_22_pad_groupi_n_1095);
  xnor csa_tree_add_101_22_pad_groupi_g4505(csa_tree_add_101_22_pad_groupi_n_1216 ,csa_tree_add_101_22_pad_groupi_n_1036 ,csa_tree_add_101_22_pad_groupi_n_1087);
  xnor csa_tree_add_101_22_pad_groupi_g4506(csa_tree_add_101_22_pad_groupi_n_1215 ,csa_tree_add_101_22_pad_groupi_n_1137 ,csa_tree_add_101_22_pad_groupi_n_1086);
  xnor csa_tree_add_101_22_pad_groupi_g4507(csa_tree_add_101_22_pad_groupi_n_1214 ,csa_tree_add_101_22_pad_groupi_n_1042 ,csa_tree_add_101_22_pad_groupi_n_1093);
  xnor csa_tree_add_101_22_pad_groupi_g4508(csa_tree_add_101_22_pad_groupi_n_1213 ,csa_tree_add_101_22_pad_groupi_n_1034 ,csa_tree_add_101_22_pad_groupi_n_1104);
  xnor csa_tree_add_101_22_pad_groupi_g4509(csa_tree_add_101_22_pad_groupi_n_1212 ,csa_tree_add_101_22_pad_groupi_n_1131 ,csa_tree_add_101_22_pad_groupi_n_1082);
  xnor csa_tree_add_101_22_pad_groupi_g4510(csa_tree_add_101_22_pad_groupi_n_1211 ,csa_tree_add_101_22_pad_groupi_n_1134 ,csa_tree_add_101_22_pad_groupi_n_1135);
  xnor csa_tree_add_101_22_pad_groupi_g4511(csa_tree_add_101_22_pad_groupi_n_1210 ,csa_tree_add_101_22_pad_groupi_n_1062 ,csa_tree_add_101_22_pad_groupi_n_1133);
  xnor csa_tree_add_101_22_pad_groupi_g4512(csa_tree_add_101_22_pad_groupi_n_1236 ,csa_tree_add_101_22_pad_groupi_n_1043 ,csa_tree_add_101_22_pad_groupi_n_1078);
  xnor csa_tree_add_101_22_pad_groupi_g4513(csa_tree_add_101_22_pad_groupi_n_1235 ,csa_tree_add_101_22_pad_groupi_n_1070 ,csa_tree_add_101_22_pad_groupi_n_1079);
  xnor csa_tree_add_101_22_pad_groupi_g4514(csa_tree_add_101_22_pad_groupi_n_1233 ,csa_tree_add_101_22_pad_groupi_n_976 ,csa_tree_add_101_22_pad_groupi_n_1077);
  not csa_tree_add_101_22_pad_groupi_g4515(csa_tree_add_101_22_pad_groupi_n_1206 ,csa_tree_add_101_22_pad_groupi_n_1205);
  not csa_tree_add_101_22_pad_groupi_g4516(csa_tree_add_101_22_pad_groupi_n_1204 ,csa_tree_add_101_22_pad_groupi_n_1203);
  not csa_tree_add_101_22_pad_groupi_g4517(csa_tree_add_101_22_pad_groupi_n_1202 ,csa_tree_add_101_22_pad_groupi_n_1201);
  and csa_tree_add_101_22_pad_groupi_g4518(csa_tree_add_101_22_pad_groupi_n_1200 ,csa_tree_add_101_22_pad_groupi_n_1035 ,csa_tree_add_101_22_pad_groupi_n_1094);
  or csa_tree_add_101_22_pad_groupi_g4519(csa_tree_add_101_22_pad_groupi_n_1199 ,csa_tree_add_101_22_pad_groupi_n_1105 ,csa_tree_add_101_22_pad_groupi_n_1128);
  nor csa_tree_add_101_22_pad_groupi_g4520(csa_tree_add_101_22_pad_groupi_n_1198 ,csa_tree_add_101_22_pad_groupi_n_1100 ,csa_tree_add_101_22_pad_groupi_n_1139);
  or csa_tree_add_101_22_pad_groupi_g4521(csa_tree_add_101_22_pad_groupi_n_1197 ,csa_tree_add_101_22_pad_groupi_n_1136 ,csa_tree_add_101_22_pad_groupi_n_1086);
  and csa_tree_add_101_22_pad_groupi_g4522(csa_tree_add_101_22_pad_groupi_n_1196 ,csa_tree_add_101_22_pad_groupi_n_1118 ,csa_tree_add_101_22_pad_groupi_n_1103);
  and csa_tree_add_101_22_pad_groupi_g4523(csa_tree_add_101_22_pad_groupi_n_1195 ,csa_tree_add_101_22_pad_groupi_n_1100 ,csa_tree_add_101_22_pad_groupi_n_1139);
  or csa_tree_add_101_22_pad_groupi_g4524(csa_tree_add_101_22_pad_groupi_n_1194 ,csa_tree_add_101_22_pad_groupi_n_1055 ,csa_tree_add_101_22_pad_groupi_n_1095);
  nor csa_tree_add_101_22_pad_groupi_g4525(csa_tree_add_101_22_pad_groupi_n_1193 ,csa_tree_add_101_22_pad_groupi_n_1137 ,csa_tree_add_101_22_pad_groupi_n_1085);
  or csa_tree_add_101_22_pad_groupi_g4526(csa_tree_add_101_22_pad_groupi_n_1192 ,csa_tree_add_101_22_pad_groupi_n_1083 ,csa_tree_add_101_22_pad_groupi_n_1089);
  nor csa_tree_add_101_22_pad_groupi_g4527(csa_tree_add_101_22_pad_groupi_n_1191 ,csa_tree_add_101_22_pad_groupi_n_1022 ,csa_tree_add_101_22_pad_groupi_n_1109);
  nor csa_tree_add_101_22_pad_groupi_g4528(csa_tree_add_101_22_pad_groupi_n_1190 ,csa_tree_add_101_22_pad_groupi_n_1084 ,csa_tree_add_101_22_pad_groupi_n_1090);
  or csa_tree_add_101_22_pad_groupi_g4529(csa_tree_add_101_22_pad_groupi_n_1189 ,csa_tree_add_101_22_pad_groupi_n_1056 ,csa_tree_add_101_22_pad_groupi_n_3);
  nor csa_tree_add_101_22_pad_groupi_g4530(csa_tree_add_101_22_pad_groupi_n_1188 ,csa_tree_add_101_22_pad_groupi_n_1019 ,csa_tree_add_101_22_pad_groupi_n_1080);
  and csa_tree_add_101_22_pad_groupi_g4531(csa_tree_add_101_22_pad_groupi_n_1187 ,csa_tree_add_101_22_pad_groupi_n_1056 ,csa_tree_add_101_22_pad_groupi_n_3);
  and csa_tree_add_101_22_pad_groupi_g4532(csa_tree_add_101_22_pad_groupi_n_1186 ,csa_tree_add_101_22_pad_groupi_n_1019 ,csa_tree_add_101_22_pad_groupi_n_1080);
  and csa_tree_add_101_22_pad_groupi_g4533(csa_tree_add_101_22_pad_groupi_n_1185 ,csa_tree_add_101_22_pad_groupi_n_1134 ,csa_tree_add_101_22_pad_groupi_n_1135);
  nor csa_tree_add_101_22_pad_groupi_g4534(csa_tree_add_101_22_pad_groupi_n_1184 ,csa_tree_add_101_22_pad_groupi_n_1134 ,csa_tree_add_101_22_pad_groupi_n_1135);
  and csa_tree_add_101_22_pad_groupi_g4535(csa_tree_add_101_22_pad_groupi_n_1183 ,csa_tree_add_101_22_pad_groupi_n_1062 ,csa_tree_add_101_22_pad_groupi_n_1133);
  and csa_tree_add_101_22_pad_groupi_g4536(csa_tree_add_101_22_pad_groupi_n_1182 ,csa_tree_add_101_22_pad_groupi_n_1120 ,csa_tree_add_101_22_pad_groupi_n_1106);
  or csa_tree_add_101_22_pad_groupi_g4537(csa_tree_add_101_22_pad_groupi_n_1181 ,csa_tree_add_101_22_pad_groupi_n_1062 ,csa_tree_add_101_22_pad_groupi_n_1133);
  and csa_tree_add_101_22_pad_groupi_g4538(csa_tree_add_101_22_pad_groupi_n_1180 ,csa_tree_add_101_22_pad_groupi_n_1050 ,csa_tree_add_101_22_pad_groupi_n_1140);
  and csa_tree_add_101_22_pad_groupi_g4539(csa_tree_add_101_22_pad_groupi_n_1179 ,csa_tree_add_101_22_pad_groupi_n_1055 ,csa_tree_add_101_22_pad_groupi_n_1095);
  nor csa_tree_add_101_22_pad_groupi_g4540(csa_tree_add_101_22_pad_groupi_n_1178 ,csa_tree_add_101_22_pad_groupi_n_1023 ,csa_tree_add_101_22_pad_groupi_n_1108);
  nor csa_tree_add_101_22_pad_groupi_g4541(csa_tree_add_101_22_pad_groupi_n_1177 ,csa_tree_add_101_22_pad_groupi_n_1031 ,csa_tree_add_101_22_pad_groupi_n_1119);
  and csa_tree_add_101_22_pad_groupi_g4542(csa_tree_add_101_22_pad_groupi_n_1209 ,csa_tree_add_101_22_pad_groupi_n_1054 ,csa_tree_add_101_22_pad_groupi_n_1127);
  or csa_tree_add_101_22_pad_groupi_g4543(csa_tree_add_101_22_pad_groupi_n_1208 ,csa_tree_add_101_22_pad_groupi_n_901 ,csa_tree_add_101_22_pad_groupi_n_1122);
  or csa_tree_add_101_22_pad_groupi_g4544(csa_tree_add_101_22_pad_groupi_n_1207 ,csa_tree_add_101_22_pad_groupi_n_914 ,csa_tree_add_101_22_pad_groupi_n_1125);
  and csa_tree_add_101_22_pad_groupi_g4545(csa_tree_add_101_22_pad_groupi_n_1205 ,csa_tree_add_101_22_pad_groupi_n_884 ,csa_tree_add_101_22_pad_groupi_n_1116);
  and csa_tree_add_101_22_pad_groupi_g4546(csa_tree_add_101_22_pad_groupi_n_1203 ,csa_tree_add_101_22_pad_groupi_n_921 ,csa_tree_add_101_22_pad_groupi_n_1126);
  or csa_tree_add_101_22_pad_groupi_g4547(csa_tree_add_101_22_pad_groupi_n_1201 ,csa_tree_add_101_22_pad_groupi_n_1049 ,csa_tree_add_101_22_pad_groupi_n_1117);
  not csa_tree_add_101_22_pad_groupi_g4548(csa_tree_add_101_22_pad_groupi_n_1170 ,csa_tree_add_101_22_pad_groupi_n_1171);
  not csa_tree_add_101_22_pad_groupi_g4549(csa_tree_add_101_22_pad_groupi_n_1166 ,csa_tree_add_101_22_pad_groupi_n_1165);
  not csa_tree_add_101_22_pad_groupi_g4550(csa_tree_add_101_22_pad_groupi_n_1163 ,csa_tree_add_101_22_pad_groupi_n_1162);
  not csa_tree_add_101_22_pad_groupi_g4551(csa_tree_add_101_22_pad_groupi_n_1160 ,csa_tree_add_101_22_pad_groupi_n_1159);
  or csa_tree_add_101_22_pad_groupi_g4552(csa_tree_add_101_22_pad_groupi_n_1158 ,csa_tree_add_101_22_pad_groupi_n_1035 ,csa_tree_add_101_22_pad_groupi_n_1094);
  and csa_tree_add_101_22_pad_groupi_g4553(csa_tree_add_101_22_pad_groupi_n_1157 ,csa_tree_add_101_22_pad_groupi_n_1015 ,csa_tree_add_101_22_pad_groupi_n_1097);
  or csa_tree_add_101_22_pad_groupi_g4554(csa_tree_add_101_22_pad_groupi_n_1156 ,csa_tree_add_101_22_pad_groupi_n_1130 ,csa_tree_add_101_22_pad_groupi_n_1081);
  or csa_tree_add_101_22_pad_groupi_g4555(csa_tree_add_101_22_pad_groupi_n_1155 ,csa_tree_add_101_22_pad_groupi_n_1033 ,csa_tree_add_101_22_pad_groupi_n_1091);
  and csa_tree_add_101_22_pad_groupi_g4556(csa_tree_add_101_22_pad_groupi_n_1154 ,csa_tree_add_101_22_pad_groupi_n_1093 ,csa_tree_add_101_22_pad_groupi_n_1088);
  nor csa_tree_add_101_22_pad_groupi_g4557(csa_tree_add_101_22_pad_groupi_n_1153 ,csa_tree_add_101_22_pad_groupi_n_1093 ,csa_tree_add_101_22_pad_groupi_n_1088);
  and csa_tree_add_101_22_pad_groupi_g4558(csa_tree_add_101_22_pad_groupi_n_1152 ,csa_tree_add_101_22_pad_groupi_n_1016 ,csa_tree_add_101_22_pad_groupi_n_1096);
  nor csa_tree_add_101_22_pad_groupi_g4559(csa_tree_add_101_22_pad_groupi_n_1151 ,csa_tree_add_101_22_pad_groupi_n_1034 ,csa_tree_add_101_22_pad_groupi_n_1092);
  nor csa_tree_add_101_22_pad_groupi_g4560(csa_tree_add_101_22_pad_groupi_n_1150 ,csa_tree_add_101_22_pad_groupi_n_1131 ,csa_tree_add_101_22_pad_groupi_n_1082);
  or csa_tree_add_101_22_pad_groupi_g4561(csa_tree_add_101_22_pad_groupi_n_1149 ,csa_tree_add_101_22_pad_groupi_n_1110 ,csa_tree_add_101_22_pad_groupi_n_1101);
  and csa_tree_add_101_22_pad_groupi_g4562(csa_tree_add_101_22_pad_groupi_n_1148 ,csa_tree_add_101_22_pad_groupi_n_1037 ,csa_tree_add_101_22_pad_groupi_n_1087);
  nor csa_tree_add_101_22_pad_groupi_g4563(csa_tree_add_101_22_pad_groupi_n_1147 ,csa_tree_add_101_22_pad_groupi_n_1037 ,csa_tree_add_101_22_pad_groupi_n_1087);
  xnor csa_tree_add_101_22_pad_groupi_g4564(csa_tree_add_101_22_pad_groupi_n_1146 ,csa_tree_add_101_22_pad_groupi_n_1010 ,csa_tree_add_101_22_pad_groupi_n_1064);
  xnor csa_tree_add_101_22_pad_groupi_g4565(csa_tree_add_101_22_pad_groupi_n_1145 ,csa_tree_add_101_22_pad_groupi_n_1067 ,csa_tree_add_101_22_pad_groupi_n_1019);
  xnor csa_tree_add_101_22_pad_groupi_g4566(csa_tree_add_101_22_pad_groupi_n_1144 ,csa_tree_add_101_22_pad_groupi_n_1058 ,csa_tree_add_101_22_pad_groupi_n_1061);
  xnor csa_tree_add_101_22_pad_groupi_g4567(csa_tree_add_101_22_pad_groupi_n_1143 ,csa_tree_add_101_22_pad_groupi_n_1011 ,csa_tree_add_101_22_pad_groupi_n_1059);
  xnor csa_tree_add_101_22_pad_groupi_g4568(csa_tree_add_101_22_pad_groupi_n_1142 ,csa_tree_add_101_22_pad_groupi_n_1018 ,csa_tree_add_101_22_pad_groupi_n_1066);
  xnor csa_tree_add_101_22_pad_groupi_g4569(csa_tree_add_101_22_pad_groupi_n_1176 ,csa_tree_add_101_22_pad_groupi_n_1020 ,csa_tree_add_101_22_pad_groupi_n_1025);
  and csa_tree_add_101_22_pad_groupi_g4570(csa_tree_add_101_22_pad_groupi_n_1175 ,csa_tree_add_101_22_pad_groupi_n_1030 ,csa_tree_add_101_22_pad_groupi_n_1111);
  xnor csa_tree_add_101_22_pad_groupi_g4571(csa_tree_add_101_22_pad_groupi_n_1174 ,csa_tree_add_101_22_pad_groupi_n_1068 ,csa_tree_add_101_22_pad_groupi_n_950);
  or csa_tree_add_101_22_pad_groupi_g4572(csa_tree_add_101_22_pad_groupi_n_1173 ,csa_tree_add_101_22_pad_groupi_n_908 ,csa_tree_add_101_22_pad_groupi_n_1121);
  xnor csa_tree_add_101_22_pad_groupi_g4573(csa_tree_add_101_22_pad_groupi_n_1172 ,csa_tree_add_101_22_pad_groupi_n_1045 ,csa_tree_add_101_22_pad_groupi_n_944);
  xnor csa_tree_add_101_22_pad_groupi_g4574(csa_tree_add_101_22_pad_groupi_n_1171 ,csa_tree_add_101_22_pad_groupi_n_1073 ,csa_tree_add_101_22_pad_groupi_n_941);
  xnor csa_tree_add_101_22_pad_groupi_g4575(csa_tree_add_101_22_pad_groupi_n_1169 ,csa_tree_add_101_22_pad_groupi_n_1041 ,csa_tree_add_101_22_pad_groupi_n_974);
  xnor csa_tree_add_101_22_pad_groupi_g4576(csa_tree_add_101_22_pad_groupi_n_1168 ,csa_tree_add_101_22_pad_groupi_n_1044 ,csa_tree_add_101_22_pad_groupi_n_939);
  xnor csa_tree_add_101_22_pad_groupi_g4577(csa_tree_add_101_22_pad_groupi_n_1167 ,csa_tree_add_101_22_pad_groupi_n_1040 ,csa_tree_add_101_22_pad_groupi_n_969);
  xnor csa_tree_add_101_22_pad_groupi_g4578(csa_tree_add_101_22_pad_groupi_n_1165 ,csa_tree_add_101_22_pad_groupi_n_1038 ,csa_tree_add_101_22_pad_groupi_n_970);
  or csa_tree_add_101_22_pad_groupi_g4579(csa_tree_add_101_22_pad_groupi_n_1164 ,csa_tree_add_101_22_pad_groupi_n_858 ,csa_tree_add_101_22_pad_groupi_n_1113);
  and csa_tree_add_101_22_pad_groupi_g4580(csa_tree_add_101_22_pad_groupi_n_1162 ,csa_tree_add_101_22_pad_groupi_n_857 ,csa_tree_add_101_22_pad_groupi_n_1112);
  or csa_tree_add_101_22_pad_groupi_g4581(csa_tree_add_101_22_pad_groupi_n_1161 ,csa_tree_add_101_22_pad_groupi_n_873 ,csa_tree_add_101_22_pad_groupi_n_1129);
  xnor csa_tree_add_101_22_pad_groupi_g4582(csa_tree_add_101_22_pad_groupi_n_1159 ,csa_tree_add_101_22_pad_groupi_n_1046 ,csa_tree_add_101_22_pad_groupi_n_955);
  not csa_tree_add_101_22_pad_groupi_g4583(csa_tree_add_101_22_pad_groupi_n_1139 ,csa_tree_add_101_22_pad_groupi_n_1138);
  not csa_tree_add_101_22_pad_groupi_g4584(csa_tree_add_101_22_pad_groupi_n_1136 ,csa_tree_add_101_22_pad_groupi_n_1137);
  not csa_tree_add_101_22_pad_groupi_g4585(csa_tree_add_101_22_pad_groupi_n_1130 ,csa_tree_add_101_22_pad_groupi_n_1131);
  and csa_tree_add_101_22_pad_groupi_g4586(csa_tree_add_101_22_pad_groupi_n_1129 ,csa_tree_add_101_22_pad_groupi_n_871 ,csa_tree_add_101_22_pad_groupi_n_1040);
  nor csa_tree_add_101_22_pad_groupi_g4587(csa_tree_add_101_22_pad_groupi_n_1128 ,csa_tree_add_101_22_pad_groupi_n_1058 ,csa_tree_add_101_22_pad_groupi_n_1061);
  or csa_tree_add_101_22_pad_groupi_g4588(csa_tree_add_101_22_pad_groupi_n_1127 ,csa_tree_add_101_22_pad_groupi_n_1053 ,csa_tree_add_101_22_pad_groupi_n_1071);
  or csa_tree_add_101_22_pad_groupi_g4589(csa_tree_add_101_22_pad_groupi_n_1126 ,csa_tree_add_101_22_pad_groupi_n_918 ,csa_tree_add_101_22_pad_groupi_n_1069);
  and csa_tree_add_101_22_pad_groupi_g4590(csa_tree_add_101_22_pad_groupi_n_1125 ,csa_tree_add_101_22_pad_groupi_n_932 ,csa_tree_add_101_22_pad_groupi_n_1073);
  nor csa_tree_add_101_22_pad_groupi_g4591(csa_tree_add_101_22_pad_groupi_n_1124 ,csa_tree_add_101_22_pad_groupi_n_1010 ,csa_tree_add_101_22_pad_groupi_n_1063);
  and csa_tree_add_101_22_pad_groupi_g4592(csa_tree_add_101_22_pad_groupi_n_1123 ,csa_tree_add_101_22_pad_groupi_n_1011 ,csa_tree_add_101_22_pad_groupi_n_1059);
  and csa_tree_add_101_22_pad_groupi_g4593(csa_tree_add_101_22_pad_groupi_n_1122 ,csa_tree_add_101_22_pad_groupi_n_880 ,csa_tree_add_101_22_pad_groupi_n_1045);
  and csa_tree_add_101_22_pad_groupi_g4594(csa_tree_add_101_22_pad_groupi_n_1121 ,csa_tree_add_101_22_pad_groupi_n_867 ,csa_tree_add_101_22_pad_groupi_n_1044);
  or csa_tree_add_101_22_pad_groupi_g4595(csa_tree_add_101_22_pad_groupi_n_1120 ,csa_tree_add_101_22_pad_groupi_n_1011 ,csa_tree_add_101_22_pad_groupi_n_1059);
  nor csa_tree_add_101_22_pad_groupi_g4596(csa_tree_add_101_22_pad_groupi_n_1119 ,csa_tree_add_101_22_pad_groupi_n_1026 ,csa_tree_add_101_22_pad_groupi_n_980);
  or csa_tree_add_101_22_pad_groupi_g4597(csa_tree_add_101_22_pad_groupi_n_1118 ,csa_tree_add_101_22_pad_groupi_n_1009 ,csa_tree_add_101_22_pad_groupi_n_1064);
  and csa_tree_add_101_22_pad_groupi_g4598(csa_tree_add_101_22_pad_groupi_n_1117 ,csa_tree_add_101_22_pad_groupi_n_1029 ,csa_tree_add_101_22_pad_groupi_n_1043);
  or csa_tree_add_101_22_pad_groupi_g4599(csa_tree_add_101_22_pad_groupi_n_1116 ,csa_tree_add_101_22_pad_groupi_n_882 ,csa_tree_add_101_22_pad_groupi_n_1038);
  or csa_tree_add_101_22_pad_groupi_g4600(csa_tree_add_101_22_pad_groupi_n_1115 ,csa_tree_add_101_22_pad_groupi_n_1057 ,csa_tree_add_101_22_pad_groupi_n_1060);
  or csa_tree_add_101_22_pad_groupi_g4601(csa_tree_add_101_22_pad_groupi_n_1114 ,csa_tree_add_101_22_pad_groupi_n_1017 ,csa_tree_add_101_22_pad_groupi_n_1065);
  and csa_tree_add_101_22_pad_groupi_g4602(csa_tree_add_101_22_pad_groupi_n_1113 ,csa_tree_add_101_22_pad_groupi_n_860 ,csa_tree_add_101_22_pad_groupi_n_1041);
  or csa_tree_add_101_22_pad_groupi_g4603(csa_tree_add_101_22_pad_groupi_n_1112 ,csa_tree_add_101_22_pad_groupi_n_854 ,csa_tree_add_101_22_pad_groupi_n_1046);
  or csa_tree_add_101_22_pad_groupi_g4604(csa_tree_add_101_22_pad_groupi_n_1111 ,csa_tree_add_101_22_pad_groupi_n_1028 ,csa_tree_add_101_22_pad_groupi_n_976);
  nor csa_tree_add_101_22_pad_groupi_g4605(csa_tree_add_101_22_pad_groupi_n_1110 ,csa_tree_add_101_22_pad_groupi_n_1018 ,csa_tree_add_101_22_pad_groupi_n_1066);
  xnor csa_tree_add_101_22_pad_groupi_g4606(csa_tree_add_101_22_pad_groupi_n_1141 ,csa_tree_add_101_22_pad_groupi_n_842 ,csa_tree_add_101_22_pad_groupi_n_951);
  xnor csa_tree_add_101_22_pad_groupi_g4607(csa_tree_add_101_22_pad_groupi_n_1140 ,csa_tree_add_101_22_pad_groupi_n_803 ,csa_tree_add_101_22_pad_groupi_n_964);
  xnor csa_tree_add_101_22_pad_groupi_g4608(csa_tree_add_101_22_pad_groupi_n_1138 ,csa_tree_add_101_22_pad_groupi_n_773 ,csa_tree_add_101_22_pad_groupi_n_962);
  xnor csa_tree_add_101_22_pad_groupi_g4609(csa_tree_add_101_22_pad_groupi_n_1137 ,csa_tree_add_101_22_pad_groupi_n_783 ,csa_tree_add_101_22_pad_groupi_n_960);
  xnor csa_tree_add_101_22_pad_groupi_g4610(csa_tree_add_101_22_pad_groupi_n_1135 ,csa_tree_add_101_22_pad_groupi_n_840 ,csa_tree_add_101_22_pad_groupi_n_965);
  or csa_tree_add_101_22_pad_groupi_g4611(csa_tree_add_101_22_pad_groupi_n_1134 ,csa_tree_add_101_22_pad_groupi_n_1000 ,csa_tree_add_101_22_pad_groupi_n_1052);
  xnor csa_tree_add_101_22_pad_groupi_g4612(csa_tree_add_101_22_pad_groupi_n_1133 ,csa_tree_add_101_22_pad_groupi_n_778 ,csa_tree_add_101_22_pad_groupi_n_949);
  and csa_tree_add_101_22_pad_groupi_g4613(csa_tree_add_101_22_pad_groupi_n_1132 ,csa_tree_add_101_22_pad_groupi_n_888 ,csa_tree_add_101_22_pad_groupi_n_1032);
  or csa_tree_add_101_22_pad_groupi_g4614(csa_tree_add_101_22_pad_groupi_n_1131 ,csa_tree_add_101_22_pad_groupi_n_868 ,csa_tree_add_101_22_pad_groupi_n_1027);
  not csa_tree_add_101_22_pad_groupi_g4615(csa_tree_add_101_22_pad_groupi_n_1109 ,csa_tree_add_101_22_pad_groupi_n_1108);
  not csa_tree_add_101_22_pad_groupi_g4616(csa_tree_add_101_22_pad_groupi_n_1097 ,csa_tree_add_101_22_pad_groupi_n_1096);
  not csa_tree_add_101_22_pad_groupi_g4617(csa_tree_add_101_22_pad_groupi_n_1091 ,csa_tree_add_101_22_pad_groupi_n_1092);
  not csa_tree_add_101_22_pad_groupi_g4618(csa_tree_add_101_22_pad_groupi_n_1090 ,csa_tree_add_101_22_pad_groupi_n_1089);
  not csa_tree_add_101_22_pad_groupi_g4619(csa_tree_add_101_22_pad_groupi_n_1085 ,csa_tree_add_101_22_pad_groupi_n_1086);
  not csa_tree_add_101_22_pad_groupi_g4620(csa_tree_add_101_22_pad_groupi_n_1083 ,csa_tree_add_101_22_pad_groupi_n_1084);
  not csa_tree_add_101_22_pad_groupi_g4621(csa_tree_add_101_22_pad_groupi_n_1081 ,csa_tree_add_101_22_pad_groupi_n_1082);
  xnor csa_tree_add_101_22_pad_groupi_g4622(csa_tree_add_101_22_pad_groupi_n_1079 ,csa_tree_add_101_22_pad_groupi_n_975 ,csa_tree_add_101_22_pad_groupi_n_934);
  xnor csa_tree_add_101_22_pad_groupi_g4623(csa_tree_add_101_22_pad_groupi_n_1108 ,csa_tree_add_101_22_pad_groupi_n_892 ,csa_tree_add_101_22_pad_groupi_n_961);
  xnor csa_tree_add_101_22_pad_groupi_g4624(csa_tree_add_101_22_pad_groupi_n_1078 ,csa_tree_add_101_22_pad_groupi_n_797 ,csa_tree_add_101_22_pad_groupi_n_4);
  xnor csa_tree_add_101_22_pad_groupi_g4625(csa_tree_add_101_22_pad_groupi_n_1077 ,csa_tree_add_101_22_pad_groupi_n_746 ,csa_tree_add_101_22_pad_groupi_n_1014);
  xnor csa_tree_add_101_22_pad_groupi_g4626(csa_tree_add_101_22_pad_groupi_n_1076 ,csa_tree_add_101_22_pad_groupi_n_1012 ,csa_tree_add_101_22_pad_groupi_n_933);
  xnor csa_tree_add_101_22_pad_groupi_g4628(csa_tree_add_101_22_pad_groupi_n_1107 ,csa_tree_add_101_22_pad_groupi_n_768 ,csa_tree_add_101_22_pad_groupi_n_942);
  xnor csa_tree_add_101_22_pad_groupi_g4629(csa_tree_add_101_22_pad_groupi_n_1106 ,csa_tree_add_101_22_pad_groupi_n_764 ,csa_tree_add_101_22_pad_groupi_n_968);
  xnor csa_tree_add_101_22_pad_groupi_g4630(csa_tree_add_101_22_pad_groupi_n_1105 ,csa_tree_add_101_22_pad_groupi_n_740 ,csa_tree_add_101_22_pad_groupi_n_963);
  xnor csa_tree_add_101_22_pad_groupi_g4631(csa_tree_add_101_22_pad_groupi_n_1104 ,csa_tree_add_101_22_pad_groupi_n_782 ,csa_tree_add_101_22_pad_groupi_n_967);
  xnor csa_tree_add_101_22_pad_groupi_g4632(csa_tree_add_101_22_pad_groupi_n_1103 ,csa_tree_add_101_22_pad_groupi_n_1021 ,csa_tree_add_101_22_pad_groupi_n_957);
  xnor csa_tree_add_101_22_pad_groupi_g4633(csa_tree_add_101_22_pad_groupi_n_1102 ,csa_tree_add_101_22_pad_groupi_n_769 ,csa_tree_add_101_22_pad_groupi_n_945);
  xnor csa_tree_add_101_22_pad_groupi_g4634(csa_tree_add_101_22_pad_groupi_n_1101 ,csa_tree_add_101_22_pad_groupi_n_977 ,csa_tree_add_101_22_pad_groupi_n_966);
  xnor csa_tree_add_101_22_pad_groupi_g4635(csa_tree_add_101_22_pad_groupi_n_1100 ,csa_tree_add_101_22_pad_groupi_n_838 ,csa_tree_add_101_22_pad_groupi_n_946);
  xnor csa_tree_add_101_22_pad_groupi_g4637(csa_tree_add_101_22_pad_groupi_n_1099 ,csa_tree_add_101_22_pad_groupi_n_750 ,csa_tree_add_101_22_pad_groupi_n_952);
  xnor csa_tree_add_101_22_pad_groupi_g4638(csa_tree_add_101_22_pad_groupi_n_1098 ,csa_tree_add_101_22_pad_groupi_n_743 ,csa_tree_add_101_22_pad_groupi_n_972);
  xnor csa_tree_add_101_22_pad_groupi_g4639(csa_tree_add_101_22_pad_groupi_n_1096 ,csa_tree_add_101_22_pad_groupi_n_971 ,csa_tree_add_101_22_pad_groupi_n_578);
  xnor csa_tree_add_101_22_pad_groupi_g4640(csa_tree_add_101_22_pad_groupi_n_1095 ,csa_tree_add_101_22_pad_groupi_n_770 ,csa_tree_add_101_22_pad_groupi_n_947);
  xnor csa_tree_add_101_22_pad_groupi_g4641(csa_tree_add_101_22_pad_groupi_n_1094 ,csa_tree_add_101_22_pad_groupi_n_830 ,csa_tree_add_101_22_pad_groupi_n_943);
  xnor csa_tree_add_101_22_pad_groupi_g4642(csa_tree_add_101_22_pad_groupi_n_1093 ,csa_tree_add_101_22_pad_groupi_n_780 ,csa_tree_add_101_22_pad_groupi_n_938);
  xnor csa_tree_add_101_22_pad_groupi_g4643(csa_tree_add_101_22_pad_groupi_n_1092 ,csa_tree_add_101_22_pad_groupi_n_775 ,csa_tree_add_101_22_pad_groupi_n_937);
  xnor csa_tree_add_101_22_pad_groupi_g4644(csa_tree_add_101_22_pad_groupi_n_1089 ,csa_tree_add_101_22_pad_groupi_n_827 ,csa_tree_add_101_22_pad_groupi_n_973);
  xnor csa_tree_add_101_22_pad_groupi_g4645(csa_tree_add_101_22_pad_groupi_n_1088 ,csa_tree_add_101_22_pad_groupi_n_777 ,csa_tree_add_101_22_pad_groupi_n_940);
  xnor csa_tree_add_101_22_pad_groupi_g4646(csa_tree_add_101_22_pad_groupi_n_1087 ,csa_tree_add_101_22_pad_groupi_n_774 ,csa_tree_add_101_22_pad_groupi_n_954);
  xnor csa_tree_add_101_22_pad_groupi_g4647(csa_tree_add_101_22_pad_groupi_n_1086 ,csa_tree_add_101_22_pad_groupi_n_893 ,csa_tree_add_101_22_pad_groupi_n_959);
  xnor csa_tree_add_101_22_pad_groupi_g4648(csa_tree_add_101_22_pad_groupi_n_1084 ,csa_tree_add_101_22_pad_groupi_n_785 ,csa_tree_add_101_22_pad_groupi_n_956);
  xnor csa_tree_add_101_22_pad_groupi_g4649(csa_tree_add_101_22_pad_groupi_n_1082 ,csa_tree_add_101_22_pad_groupi_n_839 ,csa_tree_add_101_22_pad_groupi_n_958);
  xnor csa_tree_add_101_22_pad_groupi_g4650(csa_tree_add_101_22_pad_groupi_n_1080 ,csa_tree_add_101_22_pad_groupi_n_936 ,csa_tree_add_101_22_pad_groupi_n_953);
  not csa_tree_add_101_22_pad_groupi_g4651(csa_tree_add_101_22_pad_groupi_n_1071 ,csa_tree_add_101_22_pad_groupi_n_1070);
  not csa_tree_add_101_22_pad_groupi_g4652(csa_tree_add_101_22_pad_groupi_n_1069 ,csa_tree_add_101_22_pad_groupi_n_1068);
  not csa_tree_add_101_22_pad_groupi_g4653(csa_tree_add_101_22_pad_groupi_n_1065 ,csa_tree_add_101_22_pad_groupi_n_1066);
  not csa_tree_add_101_22_pad_groupi_g4654(csa_tree_add_101_22_pad_groupi_n_1063 ,csa_tree_add_101_22_pad_groupi_n_1064);
  not csa_tree_add_101_22_pad_groupi_g4655(csa_tree_add_101_22_pad_groupi_n_1060 ,csa_tree_add_101_22_pad_groupi_n_1061);
  not csa_tree_add_101_22_pad_groupi_g4656(csa_tree_add_101_22_pad_groupi_n_1057 ,csa_tree_add_101_22_pad_groupi_n_1058);
  or csa_tree_add_101_22_pad_groupi_g4657(csa_tree_add_101_22_pad_groupi_n_1054 ,csa_tree_add_101_22_pad_groupi_n_276 ,csa_tree_add_101_22_pad_groupi_n_975);
  and csa_tree_add_101_22_pad_groupi_g4658(csa_tree_add_101_22_pad_groupi_n_1053 ,csa_tree_add_101_22_pad_groupi_n_934 ,csa_tree_add_101_22_pad_groupi_n_975);
  and csa_tree_add_101_22_pad_groupi_g4659(csa_tree_add_101_22_pad_groupi_n_1052 ,csa_tree_add_101_22_pad_groupi_n_998 ,csa_tree_add_101_22_pad_groupi_n_1020);
  and csa_tree_add_101_22_pad_groupi_g4660(csa_tree_add_101_22_pad_groupi_n_1051 ,csa_tree_add_101_22_pad_groupi_n_933 ,csa_tree_add_101_22_pad_groupi_n_1012);
  or csa_tree_add_101_22_pad_groupi_g4661(csa_tree_add_101_22_pad_groupi_n_1050 ,csa_tree_add_101_22_pad_groupi_n_933 ,csa_tree_add_101_22_pad_groupi_n_1012);
  and csa_tree_add_101_22_pad_groupi_g4662(csa_tree_add_101_22_pad_groupi_n_1049 ,csa_tree_add_101_22_pad_groupi_n_797 ,csa_tree_add_101_22_pad_groupi_n_4);
  and csa_tree_add_101_22_pad_groupi_g4663(csa_tree_add_101_22_pad_groupi_n_1074 ,csa_tree_add_101_22_pad_groupi_n_913 ,csa_tree_add_101_22_pad_groupi_n_1007);
  or csa_tree_add_101_22_pad_groupi_g4664(csa_tree_add_101_22_pad_groupi_n_1073 ,csa_tree_add_101_22_pad_groupi_n_910 ,csa_tree_add_101_22_pad_groupi_n_999);
  and csa_tree_add_101_22_pad_groupi_g4665(csa_tree_add_101_22_pad_groupi_n_1072 ,csa_tree_add_101_22_pad_groupi_n_915 ,csa_tree_add_101_22_pad_groupi_n_996);
  or csa_tree_add_101_22_pad_groupi_g4666(csa_tree_add_101_22_pad_groupi_n_1070 ,csa_tree_add_101_22_pad_groupi_n_890 ,csa_tree_add_101_22_pad_groupi_n_1005);
  or csa_tree_add_101_22_pad_groupi_g4667(csa_tree_add_101_22_pad_groupi_n_1068 ,csa_tree_add_101_22_pad_groupi_n_905 ,csa_tree_add_101_22_pad_groupi_n_1003);
  and csa_tree_add_101_22_pad_groupi_g4668(csa_tree_add_101_22_pad_groupi_n_1067 ,csa_tree_add_101_22_pad_groupi_n_912 ,csa_tree_add_101_22_pad_groupi_n_1002);
  or csa_tree_add_101_22_pad_groupi_g4669(csa_tree_add_101_22_pad_groupi_n_1066 ,csa_tree_add_101_22_pad_groupi_n_903 ,csa_tree_add_101_22_pad_groupi_n_1004);
  or csa_tree_add_101_22_pad_groupi_g4670(csa_tree_add_101_22_pad_groupi_n_1064 ,csa_tree_add_101_22_pad_groupi_n_925 ,csa_tree_add_101_22_pad_groupi_n_1006);
  or csa_tree_add_101_22_pad_groupi_g4671(csa_tree_add_101_22_pad_groupi_n_1062 ,csa_tree_add_101_22_pad_groupi_n_874 ,csa_tree_add_101_22_pad_groupi_n_987);
  or csa_tree_add_101_22_pad_groupi_g4672(csa_tree_add_101_22_pad_groupi_n_1061 ,csa_tree_add_101_22_pad_groupi_n_929 ,csa_tree_add_101_22_pad_groupi_n_979);
  or csa_tree_add_101_22_pad_groupi_g4673(csa_tree_add_101_22_pad_groupi_n_1059 ,csa_tree_add_101_22_pad_groupi_n_889 ,csa_tree_add_101_22_pad_groupi_n_995);
  or csa_tree_add_101_22_pad_groupi_g4674(csa_tree_add_101_22_pad_groupi_n_1058 ,csa_tree_add_101_22_pad_groupi_n_911 ,csa_tree_add_101_22_pad_groupi_n_1008);
  or csa_tree_add_101_22_pad_groupi_g4675(csa_tree_add_101_22_pad_groupi_n_1056 ,csa_tree_add_101_22_pad_groupi_n_869 ,csa_tree_add_101_22_pad_groupi_n_1001);
  or csa_tree_add_101_22_pad_groupi_g4676(csa_tree_add_101_22_pad_groupi_n_1055 ,csa_tree_add_101_22_pad_groupi_n_886 ,csa_tree_add_101_22_pad_groupi_n_993);
  not csa_tree_add_101_22_pad_groupi_g4677(csa_tree_add_101_22_pad_groupi_n_1048 ,csa_tree_add_101_22_pad_groupi_n_1047);
  not csa_tree_add_101_22_pad_groupi_g4678(csa_tree_add_101_22_pad_groupi_n_1037 ,csa_tree_add_101_22_pad_groupi_n_1036);
  not csa_tree_add_101_22_pad_groupi_g4679(csa_tree_add_101_22_pad_groupi_n_1033 ,csa_tree_add_101_22_pad_groupi_n_1034);
  or csa_tree_add_101_22_pad_groupi_g4680(csa_tree_add_101_22_pad_groupi_n_1032 ,csa_tree_add_101_22_pad_groupi_n_876 ,csa_tree_add_101_22_pad_groupi_n_977);
  nor csa_tree_add_101_22_pad_groupi_g4681(csa_tree_add_101_22_pad_groupi_n_1031 ,csa_tree_add_101_22_pad_groupi_n_646 ,csa_tree_add_101_22_pad_groupi_n_1024);
  or csa_tree_add_101_22_pad_groupi_g4682(csa_tree_add_101_22_pad_groupi_n_1030 ,csa_tree_add_101_22_pad_groupi_n_745 ,csa_tree_add_101_22_pad_groupi_n_1014);
  or csa_tree_add_101_22_pad_groupi_g4683(csa_tree_add_101_22_pad_groupi_n_1029 ,csa_tree_add_101_22_pad_groupi_n_797 ,csa_tree_add_101_22_pad_groupi_n_4);
  nor csa_tree_add_101_22_pad_groupi_g4684(csa_tree_add_101_22_pad_groupi_n_1028 ,csa_tree_add_101_22_pad_groupi_n_746 ,csa_tree_add_101_22_pad_groupi_n_1013);
  and csa_tree_add_101_22_pad_groupi_g4685(csa_tree_add_101_22_pad_groupi_n_1027 ,csa_tree_add_101_22_pad_groupi_n_865 ,csa_tree_add_101_22_pad_groupi_n_1021);
  and csa_tree_add_101_22_pad_groupi_g4686(csa_tree_add_101_22_pad_groupi_n_1026 ,csa_tree_add_101_22_pad_groupi_n_646 ,csa_tree_add_101_22_pad_groupi_n_1024);
  and csa_tree_add_101_22_pad_groupi_g4687(csa_tree_add_101_22_pad_groupi_n_1047 ,csa_tree_add_101_22_pad_groupi_n_895 ,csa_tree_add_101_22_pad_groupi_n_994);
  xnor csa_tree_add_101_22_pad_groupi_g4688(csa_tree_add_101_22_pad_groupi_n_1025 ,csa_tree_add_101_22_pad_groupi_n_935 ,csa_tree_add_101_22_pad_groupi_n_820);
  and csa_tree_add_101_22_pad_groupi_g4689(csa_tree_add_101_22_pad_groupi_n_1046 ,csa_tree_add_101_22_pad_groupi_n_853 ,csa_tree_add_101_22_pad_groupi_n_982);
  or csa_tree_add_101_22_pad_groupi_g4690(csa_tree_add_101_22_pad_groupi_n_1045 ,csa_tree_add_101_22_pad_groupi_n_906 ,csa_tree_add_101_22_pad_groupi_n_997);
  or csa_tree_add_101_22_pad_groupi_g4691(csa_tree_add_101_22_pad_groupi_n_1044 ,csa_tree_add_101_22_pad_groupi_n_887 ,csa_tree_add_101_22_pad_groupi_n_992);
  or csa_tree_add_101_22_pad_groupi_g4692(csa_tree_add_101_22_pad_groupi_n_1043 ,csa_tree_add_101_22_pad_groupi_n_926 ,csa_tree_add_101_22_pad_groupi_n_991);
  and csa_tree_add_101_22_pad_groupi_g4693(csa_tree_add_101_22_pad_groupi_n_1042 ,csa_tree_add_101_22_pad_groupi_n_864 ,csa_tree_add_101_22_pad_groupi_n_985);
  or csa_tree_add_101_22_pad_groupi_g4694(csa_tree_add_101_22_pad_groupi_n_1041 ,csa_tree_add_101_22_pad_groupi_n_879 ,csa_tree_add_101_22_pad_groupi_n_984);
  or csa_tree_add_101_22_pad_groupi_g4695(csa_tree_add_101_22_pad_groupi_n_1040 ,csa_tree_add_101_22_pad_groupi_n_870 ,csa_tree_add_101_22_pad_groupi_n_988);
  and csa_tree_add_101_22_pad_groupi_g4696(csa_tree_add_101_22_pad_groupi_n_1039 ,csa_tree_add_101_22_pad_groupi_n_852 ,csa_tree_add_101_22_pad_groupi_n_981);
  and csa_tree_add_101_22_pad_groupi_g4697(csa_tree_add_101_22_pad_groupi_n_1038 ,csa_tree_add_101_22_pad_groupi_n_878 ,csa_tree_add_101_22_pad_groupi_n_989);
  or csa_tree_add_101_22_pad_groupi_g4698(csa_tree_add_101_22_pad_groupi_n_1036 ,csa_tree_add_101_22_pad_groupi_n_897 ,csa_tree_add_101_22_pad_groupi_n_983);
  or csa_tree_add_101_22_pad_groupi_g4699(csa_tree_add_101_22_pad_groupi_n_1035 ,csa_tree_add_101_22_pad_groupi_n_907 ,csa_tree_add_101_22_pad_groupi_n_990);
  or csa_tree_add_101_22_pad_groupi_g4700(csa_tree_add_101_22_pad_groupi_n_1034 ,csa_tree_add_101_22_pad_groupi_n_866 ,csa_tree_add_101_22_pad_groupi_n_986);
  not csa_tree_add_101_22_pad_groupi_g4701(csa_tree_add_101_22_pad_groupi_n_1023 ,csa_tree_add_101_22_pad_groupi_n_1022);
  not csa_tree_add_101_22_pad_groupi_g4702(csa_tree_add_101_22_pad_groupi_n_1018 ,csa_tree_add_101_22_pad_groupi_n_1017);
  not csa_tree_add_101_22_pad_groupi_g4703(csa_tree_add_101_22_pad_groupi_n_1016 ,csa_tree_add_101_22_pad_groupi_n_1015);
  not csa_tree_add_101_22_pad_groupi_g4704(csa_tree_add_101_22_pad_groupi_n_1014 ,csa_tree_add_101_22_pad_groupi_n_1013);
  not csa_tree_add_101_22_pad_groupi_g4705(csa_tree_add_101_22_pad_groupi_n_1010 ,csa_tree_add_101_22_pad_groupi_n_1009);
  nor csa_tree_add_101_22_pad_groupi_g4706(csa_tree_add_101_22_pad_groupi_n_1008 ,csa_tree_add_101_22_pad_groupi_n_841 ,csa_tree_add_101_22_pad_groupi_n_930);
  or csa_tree_add_101_22_pad_groupi_g4707(csa_tree_add_101_22_pad_groupi_n_1007 ,csa_tree_add_101_22_pad_groupi_n_843 ,csa_tree_add_101_22_pad_groupi_n_917);
  nor csa_tree_add_101_22_pad_groupi_g4708(csa_tree_add_101_22_pad_groupi_n_1006 ,csa_tree_add_101_22_pad_groupi_n_824 ,csa_tree_add_101_22_pad_groupi_n_872);
  and csa_tree_add_101_22_pad_groupi_g4709(csa_tree_add_101_22_pad_groupi_n_1005 ,csa_tree_add_101_22_pad_groupi_n_840 ,csa_tree_add_101_22_pad_groupi_n_922);
  and csa_tree_add_101_22_pad_groupi_g4710(csa_tree_add_101_22_pad_groupi_n_1004 ,csa_tree_add_101_22_pad_groupi_n_839 ,csa_tree_add_101_22_pad_groupi_n_909);
  and csa_tree_add_101_22_pad_groupi_g4711(csa_tree_add_101_22_pad_groupi_n_1003 ,csa_tree_add_101_22_pad_groupi_n_770 ,csa_tree_add_101_22_pad_groupi_n_916);
  or csa_tree_add_101_22_pad_groupi_g4712(csa_tree_add_101_22_pad_groupi_n_1002 ,csa_tree_add_101_22_pad_groupi_n_779 ,csa_tree_add_101_22_pad_groupi_n_902);
  and csa_tree_add_101_22_pad_groupi_g4713(csa_tree_add_101_22_pad_groupi_n_1001 ,csa_tree_add_101_22_pad_groupi_n_769 ,csa_tree_add_101_22_pad_groupi_n_904);
  and csa_tree_add_101_22_pad_groupi_g4714(csa_tree_add_101_22_pad_groupi_n_1000 ,csa_tree_add_101_22_pad_groupi_n_820 ,csa_tree_add_101_22_pad_groupi_n_935);
  nor csa_tree_add_101_22_pad_groupi_g4715(csa_tree_add_101_22_pad_groupi_n_999 ,csa_tree_add_101_22_pad_groupi_n_834 ,csa_tree_add_101_22_pad_groupi_n_896);
  or csa_tree_add_101_22_pad_groupi_g4716(csa_tree_add_101_22_pad_groupi_n_998 ,csa_tree_add_101_22_pad_groupi_n_820 ,csa_tree_add_101_22_pad_groupi_n_935);
  and csa_tree_add_101_22_pad_groupi_g4717(csa_tree_add_101_22_pad_groupi_n_997 ,csa_tree_add_101_22_pad_groupi_n_830 ,csa_tree_add_101_22_pad_groupi_n_856);
  or csa_tree_add_101_22_pad_groupi_g4718(csa_tree_add_101_22_pad_groupi_n_996 ,csa_tree_add_101_22_pad_groupi_n_936 ,csa_tree_add_101_22_pad_groupi_n_919);
  and csa_tree_add_101_22_pad_groupi_g4719(csa_tree_add_101_22_pad_groupi_n_995 ,csa_tree_add_101_22_pad_groupi_n_775 ,csa_tree_add_101_22_pad_groupi_n_891);
  or csa_tree_add_101_22_pad_groupi_g4720(csa_tree_add_101_22_pad_groupi_n_994 ,csa_tree_add_101_22_pad_groupi_n_892 ,csa_tree_add_101_22_pad_groupi_n_894);
  and csa_tree_add_101_22_pad_groupi_g4721(csa_tree_add_101_22_pad_groupi_n_993 ,csa_tree_add_101_22_pad_groupi_n_768 ,csa_tree_add_101_22_pad_groupi_n_924);
  and csa_tree_add_101_22_pad_groupi_g4722(csa_tree_add_101_22_pad_groupi_n_992 ,csa_tree_add_101_22_pad_groupi_n_780 ,csa_tree_add_101_22_pad_groupi_n_885);
  nor csa_tree_add_101_22_pad_groupi_g4723(csa_tree_add_101_22_pad_groupi_n_991 ,csa_tree_add_101_22_pad_groupi_n_837 ,csa_tree_add_101_22_pad_groupi_n_877);
  and csa_tree_add_101_22_pad_groupi_g4724(csa_tree_add_101_22_pad_groupi_n_990 ,csa_tree_add_101_22_pad_groupi_n_777 ,csa_tree_add_101_22_pad_groupi_n_928);
  or csa_tree_add_101_22_pad_groupi_g4725(csa_tree_add_101_22_pad_groupi_n_989 ,csa_tree_add_101_22_pad_groupi_n_838 ,csa_tree_add_101_22_pad_groupi_n_875);
  nor csa_tree_add_101_22_pad_groupi_g4726(csa_tree_add_101_22_pad_groupi_n_988 ,csa_tree_add_101_22_pad_groupi_n_774 ,csa_tree_add_101_22_pad_groupi_n_855);
  nor csa_tree_add_101_22_pad_groupi_g4727(csa_tree_add_101_22_pad_groupi_n_987 ,csa_tree_add_101_22_pad_groupi_n_776 ,csa_tree_add_101_22_pad_groupi_n_883);
  and csa_tree_add_101_22_pad_groupi_g4728(csa_tree_add_101_22_pad_groupi_n_986 ,csa_tree_add_101_22_pad_groupi_n_773 ,csa_tree_add_101_22_pad_groupi_n_863);
  or csa_tree_add_101_22_pad_groupi_g4729(csa_tree_add_101_22_pad_groupi_n_985 ,csa_tree_add_101_22_pad_groupi_n_823 ,csa_tree_add_101_22_pad_groupi_n_862);
  nor csa_tree_add_101_22_pad_groupi_g4730(csa_tree_add_101_22_pad_groupi_n_984 ,csa_tree_add_101_22_pad_groupi_n_772 ,csa_tree_add_101_22_pad_groupi_n_859);
  nor csa_tree_add_101_22_pad_groupi_g4731(csa_tree_add_101_22_pad_groupi_n_983 ,csa_tree_add_101_22_pad_groupi_n_771 ,csa_tree_add_101_22_pad_groupi_n_900);
  or csa_tree_add_101_22_pad_groupi_g4732(csa_tree_add_101_22_pad_groupi_n_982 ,csa_tree_add_101_22_pad_groupi_n_835 ,csa_tree_add_101_22_pad_groupi_n_851);
  or csa_tree_add_101_22_pad_groupi_g4733(csa_tree_add_101_22_pad_groupi_n_981 ,csa_tree_add_101_22_pad_groupi_n_893 ,csa_tree_add_101_22_pad_groupi_n_920);
  xnor csa_tree_add_101_22_pad_groupi_g4734(csa_tree_add_101_22_pad_groupi_n_980 ,csa_tree_add_101_22_pad_groupi_n_846 ,csa_tree_add_101_22_pad_groupi_n_848);
  and csa_tree_add_101_22_pad_groupi_g4735(csa_tree_add_101_22_pad_groupi_n_979 ,csa_tree_add_101_22_pad_groupi_n_827 ,csa_tree_add_101_22_pad_groupi_n_927);
  or csa_tree_add_101_22_pad_groupi_g4736(csa_tree_add_101_22_pad_groupi_n_1024 ,csa_tree_add_101_22_pad_groupi_n_19 ,csa_tree_add_101_22_pad_groupi_n_898);
  xnor csa_tree_add_101_22_pad_groupi_g4737(csa_tree_add_101_22_pad_groupi_n_1022 ,csa_tree_add_101_22_pad_groupi_n_706 ,csa_tree_add_101_22_pad_groupi_n_844);
  xnor csa_tree_add_101_22_pad_groupi_g4739(csa_tree_add_101_22_pad_groupi_n_1021 ,csa_tree_add_101_22_pad_groupi_n_711 ,in21[9]);
  xnor csa_tree_add_101_22_pad_groupi_g4740(csa_tree_add_101_22_pad_groupi_n_1020 ,csa_tree_add_101_22_pad_groupi_n_645 ,csa_tree_add_101_22_pad_groupi_n_832);
  and csa_tree_add_101_22_pad_groupi_g4741(csa_tree_add_101_22_pad_groupi_n_1019 ,csa_tree_add_101_22_pad_groupi_n_899 ,csa_tree_add_101_22_pad_groupi_n_359);
  and csa_tree_add_101_22_pad_groupi_g4742(csa_tree_add_101_22_pad_groupi_n_1017 ,csa_tree_add_101_22_pad_groupi_n_656 ,csa_tree_add_101_22_pad_groupi_n_923);
  or csa_tree_add_101_22_pad_groupi_g4743(csa_tree_add_101_22_pad_groupi_n_1015 ,csa_tree_add_101_22_pad_groupi_n_682 ,csa_tree_add_101_22_pad_groupi_n_881);
  or csa_tree_add_101_22_pad_groupi_g4744(csa_tree_add_101_22_pad_groupi_n_1013 ,csa_tree_add_101_22_pad_groupi_n_666 ,csa_tree_add_101_22_pad_groupi_n_861);
  xnor csa_tree_add_101_22_pad_groupi_g4745(csa_tree_add_101_22_pad_groupi_n_1012 ,csa_tree_add_101_22_pad_groupi_n_704 ,csa_tree_add_101_22_pad_groupi_n_767);
  xnor csa_tree_add_101_22_pad_groupi_g4746(csa_tree_add_101_22_pad_groupi_n_1011 ,csa_tree_add_101_22_pad_groupi_n_831 ,csa_tree_add_101_22_pad_groupi_n_1);
  or csa_tree_add_101_22_pad_groupi_g4747(csa_tree_add_101_22_pad_groupi_n_1009 ,csa_tree_add_101_22_pad_groupi_n_702 ,csa_tree_add_101_22_pad_groupi_n_931);
  xnor csa_tree_add_101_22_pad_groupi_g4748(csa_tree_add_101_22_pad_groupi_n_974 ,csa_tree_add_101_22_pad_groupi_n_726 ,csa_tree_add_101_22_pad_groupi_n_821);
  xnor csa_tree_add_101_22_pad_groupi_g4749(csa_tree_add_101_22_pad_groupi_n_973 ,csa_tree_add_101_22_pad_groupi_n_802 ,csa_tree_add_101_22_pad_groupi_n_795);
  xnor csa_tree_add_101_22_pad_groupi_g4750(csa_tree_add_101_22_pad_groupi_n_972 ,csa_tree_add_101_22_pad_groupi_n_837 ,csa_tree_add_101_22_pad_groupi_n_766);
  xnor csa_tree_add_101_22_pad_groupi_g4751(csa_tree_add_101_22_pad_groupi_n_971 ,csa_tree_add_101_22_pad_groupi_n_829 ,in21[12]);
  xnor csa_tree_add_101_22_pad_groupi_g4752(csa_tree_add_101_22_pad_groupi_n_970 ,csa_tree_add_101_22_pad_groupi_n_739 ,csa_tree_add_101_22_pad_groupi_n_728);
  xnor csa_tree_add_101_22_pad_groupi_g4753(csa_tree_add_101_22_pad_groupi_n_969 ,csa_tree_add_101_22_pad_groupi_n_758 ,csa_tree_add_101_22_pad_groupi_n_757);
  xor csa_tree_add_101_22_pad_groupi_g4754(csa_tree_add_101_22_pad_groupi_n_968 ,csa_tree_add_101_22_pad_groupi_n_824 ,csa_tree_add_101_22_pad_groupi_n_809);
  xor csa_tree_add_101_22_pad_groupi_g4755(csa_tree_add_101_22_pad_groupi_n_967 ,csa_tree_add_101_22_pad_groupi_n_834 ,in21[8]);
  xnor csa_tree_add_101_22_pad_groupi_g4756(csa_tree_add_101_22_pad_groupi_n_966 ,csa_tree_add_101_22_pad_groupi_n_733 ,csa_tree_add_101_22_pad_groupi_n_755);
  xnor csa_tree_add_101_22_pad_groupi_g4757(csa_tree_add_101_22_pad_groupi_n_965 ,csa_tree_add_101_22_pad_groupi_n_800 ,csa_tree_add_101_22_pad_groupi_n_799);
  xor csa_tree_add_101_22_pad_groupi_g4758(csa_tree_add_101_22_pad_groupi_n_964 ,csa_tree_add_101_22_pad_groupi_n_776 ,csa_tree_add_101_22_pad_groupi_n_721);
  xor csa_tree_add_101_22_pad_groupi_g4759(csa_tree_add_101_22_pad_groupi_n_963 ,csa_tree_add_101_22_pad_groupi_n_772 ,in21[1]);
  xnor csa_tree_add_101_22_pad_groupi_g4760(csa_tree_add_101_22_pad_groupi_n_962 ,csa_tree_add_101_22_pad_groupi_n_765 ,csa_tree_add_101_22_pad_groupi_n_751);
  xnor csa_tree_add_101_22_pad_groupi_g4761(csa_tree_add_101_22_pad_groupi_n_961 ,csa_tree_add_101_22_pad_groupi_n_735 ,csa_tree_add_101_22_pad_groupi_n_792);
  xor csa_tree_add_101_22_pad_groupi_g4762(csa_tree_add_101_22_pad_groupi_n_960 ,csa_tree_add_101_22_pad_groupi_n_771 ,csa_tree_add_101_22_pad_groupi_n_729);
  xnor csa_tree_add_101_22_pad_groupi_g4763(csa_tree_add_101_22_pad_groupi_n_959 ,csa_tree_add_101_22_pad_groupi_n_725 ,csa_tree_add_101_22_pad_groupi_n_723);
  xnor csa_tree_add_101_22_pad_groupi_g4764(csa_tree_add_101_22_pad_groupi_n_958 ,csa_tree_add_101_22_pad_groupi_n_814 ,csa_tree_add_101_22_pad_groupi_n_796);
  xnor csa_tree_add_101_22_pad_groupi_g4765(csa_tree_add_101_22_pad_groupi_n_957 ,csa_tree_add_101_22_pad_groupi_n_784 ,csa_tree_add_101_22_pad_groupi_n_747);
  xor csa_tree_add_101_22_pad_groupi_g4766(csa_tree_add_101_22_pad_groupi_n_956 ,csa_tree_add_101_22_pad_groupi_n_841 ,csa_tree_add_101_22_pad_groupi_n_748);
  xnor csa_tree_add_101_22_pad_groupi_g4767(csa_tree_add_101_22_pad_groupi_n_955 ,csa_tree_add_101_22_pad_groupi_n_760 ,csa_tree_add_101_22_pad_groupi_n_737);
  xnor csa_tree_add_101_22_pad_groupi_g4768(csa_tree_add_101_22_pad_groupi_n_954 ,csa_tree_add_101_22_pad_groupi_n_756 ,in21[2]);
  xnor csa_tree_add_101_22_pad_groupi_g4769(csa_tree_add_101_22_pad_groupi_n_953 ,csa_tree_add_101_22_pad_groupi_n_763 ,csa_tree_add_101_22_pad_groupi_n_817);
  xor csa_tree_add_101_22_pad_groupi_g4770(csa_tree_add_101_22_pad_groupi_n_952 ,csa_tree_add_101_22_pad_groupi_n_823 ,csa_tree_add_101_22_pad_groupi_n_742);
  xnor csa_tree_add_101_22_pad_groupi_g4771(csa_tree_add_101_22_pad_groupi_n_951 ,csa_tree_add_101_22_pad_groupi_n_806 ,csa_tree_add_101_22_pad_groupi_n_753);
  xnor csa_tree_add_101_22_pad_groupi_g4772(csa_tree_add_101_22_pad_groupi_n_950 ,csa_tree_add_101_22_pad_groupi_n_790 ,csa_tree_add_101_22_pad_groupi_n_819);
  xnor csa_tree_add_101_22_pad_groupi_g4773(csa_tree_add_101_22_pad_groupi_n_949 ,csa_tree_add_101_22_pad_groupi_n_813 ,csa_tree_add_101_22_pad_groupi_n_716);
  xnor csa_tree_add_101_22_pad_groupi_g4774(csa_tree_add_101_22_pad_groupi_n_948 ,csa_tree_add_101_22_pad_groupi_n_731 ,in21[6]);
  xnor csa_tree_add_101_22_pad_groupi_g4775(csa_tree_add_101_22_pad_groupi_n_947 ,csa_tree_add_101_22_pad_groupi_n_787 ,in21[5]);
  xnor csa_tree_add_101_22_pad_groupi_g4776(csa_tree_add_101_22_pad_groupi_n_946 ,csa_tree_add_101_22_pad_groupi_n_713 ,in21[7]);
  xnor csa_tree_add_101_22_pad_groupi_g4777(csa_tree_add_101_22_pad_groupi_n_945 ,csa_tree_add_101_22_pad_groupi_n_808 ,csa_tree_add_101_22_pad_groupi_n_788);
  xnor csa_tree_add_101_22_pad_groupi_g4778(csa_tree_add_101_22_pad_groupi_n_944 ,csa_tree_add_101_22_pad_groupi_n_761 ,csa_tree_add_101_22_pad_groupi_n_786);
  xnor csa_tree_add_101_22_pad_groupi_g4779(csa_tree_add_101_22_pad_groupi_n_943 ,csa_tree_add_101_22_pad_groupi_n_798 ,in21[4]);
  xnor csa_tree_add_101_22_pad_groupi_g4780(csa_tree_add_101_22_pad_groupi_n_942 ,csa_tree_add_101_22_pad_groupi_n_719 ,csa_tree_add_101_22_pad_groupi_n_720);
  xnor csa_tree_add_101_22_pad_groupi_g4781(csa_tree_add_101_22_pad_groupi_n_941 ,csa_tree_add_101_22_pad_groupi_n_815 ,csa_tree_add_101_22_pad_groupi_n_717);
  xnor csa_tree_add_101_22_pad_groupi_g4782(csa_tree_add_101_22_pad_groupi_n_940 ,csa_tree_add_101_22_pad_groupi_n_807 ,csa_tree_add_101_22_pad_groupi_n_714);
  xnor csa_tree_add_101_22_pad_groupi_g4783(csa_tree_add_101_22_pad_groupi_n_939 ,csa_tree_add_101_22_pad_groupi_n_810 ,csa_tree_add_101_22_pad_groupi_n_811);
  xnor csa_tree_add_101_22_pad_groupi_g4784(csa_tree_add_101_22_pad_groupi_n_938 ,csa_tree_add_101_22_pad_groupi_n_804 ,in21[3]);
  xnor csa_tree_add_101_22_pad_groupi_g4785(csa_tree_add_101_22_pad_groupi_n_937 ,csa_tree_add_101_22_pad_groupi_n_718 ,csa_tree_add_101_22_pad_groupi_n_793);
  xnor csa_tree_add_101_22_pad_groupi_g4786(csa_tree_add_101_22_pad_groupi_n_977 ,csa_tree_add_101_22_pad_groupi_n_822 ,csa_tree_add_101_22_pad_groupi_n_709);
  xnor csa_tree_add_101_22_pad_groupi_g4787(csa_tree_add_101_22_pad_groupi_n_976 ,csa_tree_add_101_22_pad_groupi_n_828 ,csa_tree_add_101_22_pad_groupi_n_710);
  xnor csa_tree_add_101_22_pad_groupi_g4788(csa_tree_add_101_22_pad_groupi_n_975 ,csa_tree_add_101_22_pad_groupi_n_825 ,in21[0]);
  or csa_tree_add_101_22_pad_groupi_g4791(csa_tree_add_101_22_pad_groupi_n_932 ,csa_tree_add_101_22_pad_groupi_n_815 ,csa_tree_add_101_22_pad_groupi_n_717);
  nor csa_tree_add_101_22_pad_groupi_g4792(csa_tree_add_101_22_pad_groupi_n_931 ,csa_tree_add_101_22_pad_groupi_n_673 ,csa_tree_add_101_22_pad_groupi_n_831);
  nor csa_tree_add_101_22_pad_groupi_g4793(csa_tree_add_101_22_pad_groupi_n_930 ,csa_tree_add_101_22_pad_groupi_n_748 ,csa_tree_add_101_22_pad_groupi_n_785);
  nor csa_tree_add_101_22_pad_groupi_g4794(csa_tree_add_101_22_pad_groupi_n_929 ,csa_tree_add_101_22_pad_groupi_n_802 ,csa_tree_add_101_22_pad_groupi_n_794);
  or csa_tree_add_101_22_pad_groupi_g4795(csa_tree_add_101_22_pad_groupi_n_928 ,csa_tree_add_101_22_pad_groupi_n_807 ,csa_tree_add_101_22_pad_groupi_n_714);
  or csa_tree_add_101_22_pad_groupi_g4796(csa_tree_add_101_22_pad_groupi_n_927 ,csa_tree_add_101_22_pad_groupi_n_801 ,csa_tree_add_101_22_pad_groupi_n_795);
  nor csa_tree_add_101_22_pad_groupi_g4797(csa_tree_add_101_22_pad_groupi_n_926 ,csa_tree_add_101_22_pad_groupi_n_766 ,csa_tree_add_101_22_pad_groupi_n_744);
  and csa_tree_add_101_22_pad_groupi_g4798(csa_tree_add_101_22_pad_groupi_n_925 ,csa_tree_add_101_22_pad_groupi_n_764 ,csa_tree_add_101_22_pad_groupi_n_809);
  or csa_tree_add_101_22_pad_groupi_g4799(csa_tree_add_101_22_pad_groupi_n_924 ,csa_tree_add_101_22_pad_groupi_n_719 ,csa_tree_add_101_22_pad_groupi_n_720);
  or csa_tree_add_101_22_pad_groupi_g4800(csa_tree_add_101_22_pad_groupi_n_923 ,csa_tree_add_101_22_pad_groupi_n_593 ,csa_tree_add_101_22_pad_groupi_n_836);
  or csa_tree_add_101_22_pad_groupi_g4801(csa_tree_add_101_22_pad_groupi_n_922 ,csa_tree_add_101_22_pad_groupi_n_800 ,csa_tree_add_101_22_pad_groupi_n_799);
  or csa_tree_add_101_22_pad_groupi_g4802(csa_tree_add_101_22_pad_groupi_n_921 ,csa_tree_add_101_22_pad_groupi_n_789 ,csa_tree_add_101_22_pad_groupi_n_818);
  nor csa_tree_add_101_22_pad_groupi_g4803(csa_tree_add_101_22_pad_groupi_n_920 ,csa_tree_add_101_22_pad_groupi_n_725 ,csa_tree_add_101_22_pad_groupi_n_723);
  nor csa_tree_add_101_22_pad_groupi_g4804(csa_tree_add_101_22_pad_groupi_n_919 ,csa_tree_add_101_22_pad_groupi_n_763 ,csa_tree_add_101_22_pad_groupi_n_817);
  nor csa_tree_add_101_22_pad_groupi_g4805(csa_tree_add_101_22_pad_groupi_n_918 ,csa_tree_add_101_22_pad_groupi_n_790 ,csa_tree_add_101_22_pad_groupi_n_819);
  nor csa_tree_add_101_22_pad_groupi_g4806(csa_tree_add_101_22_pad_groupi_n_917 ,csa_tree_add_101_22_pad_groupi_n_806 ,csa_tree_add_101_22_pad_groupi_n_753);
  or csa_tree_add_101_22_pad_groupi_g4807(csa_tree_add_101_22_pad_groupi_n_916 ,in21[5] ,csa_tree_add_101_22_pad_groupi_n_787);
  or csa_tree_add_101_22_pad_groupi_g4808(csa_tree_add_101_22_pad_groupi_n_915 ,csa_tree_add_101_22_pad_groupi_n_762 ,csa_tree_add_101_22_pad_groupi_n_816);
  and csa_tree_add_101_22_pad_groupi_g4809(csa_tree_add_101_22_pad_groupi_n_914 ,csa_tree_add_101_22_pad_groupi_n_815 ,csa_tree_add_101_22_pad_groupi_n_717);
  or csa_tree_add_101_22_pad_groupi_g4810(csa_tree_add_101_22_pad_groupi_n_913 ,csa_tree_add_101_22_pad_groupi_n_805 ,csa_tree_add_101_22_pad_groupi_n_752);
  or csa_tree_add_101_22_pad_groupi_g4811(csa_tree_add_101_22_pad_groupi_n_912 ,csa_tree_add_101_22_pad_groupi_n_812 ,csa_tree_add_101_22_pad_groupi_n_715);
  and csa_tree_add_101_22_pad_groupi_g4812(csa_tree_add_101_22_pad_groupi_n_911 ,csa_tree_add_101_22_pad_groupi_n_748 ,csa_tree_add_101_22_pad_groupi_n_785);
  nor csa_tree_add_101_22_pad_groupi_g4813(csa_tree_add_101_22_pad_groupi_n_910 ,csa_tree_add_101_22_pad_groupi_n_372 ,csa_tree_add_101_22_pad_groupi_n_782);
  or csa_tree_add_101_22_pad_groupi_g4814(csa_tree_add_101_22_pad_groupi_n_909 ,csa_tree_add_101_22_pad_groupi_n_814 ,csa_tree_add_101_22_pad_groupi_n_796);
  and csa_tree_add_101_22_pad_groupi_g4815(csa_tree_add_101_22_pad_groupi_n_908 ,csa_tree_add_101_22_pad_groupi_n_810 ,csa_tree_add_101_22_pad_groupi_n_811);
  and csa_tree_add_101_22_pad_groupi_g4816(csa_tree_add_101_22_pad_groupi_n_907 ,csa_tree_add_101_22_pad_groupi_n_807 ,csa_tree_add_101_22_pad_groupi_n_714);
  and csa_tree_add_101_22_pad_groupi_g4817(csa_tree_add_101_22_pad_groupi_n_906 ,in21[4] ,csa_tree_add_101_22_pad_groupi_n_798);
  and csa_tree_add_101_22_pad_groupi_g4818(csa_tree_add_101_22_pad_groupi_n_905 ,in21[5] ,csa_tree_add_101_22_pad_groupi_n_787);
  or csa_tree_add_101_22_pad_groupi_g4819(csa_tree_add_101_22_pad_groupi_n_904 ,csa_tree_add_101_22_pad_groupi_n_808 ,csa_tree_add_101_22_pad_groupi_n_788);
  and csa_tree_add_101_22_pad_groupi_g4820(csa_tree_add_101_22_pad_groupi_n_903 ,csa_tree_add_101_22_pad_groupi_n_814 ,csa_tree_add_101_22_pad_groupi_n_796);
  nor csa_tree_add_101_22_pad_groupi_g4821(csa_tree_add_101_22_pad_groupi_n_902 ,csa_tree_add_101_22_pad_groupi_n_813 ,csa_tree_add_101_22_pad_groupi_n_716);
  and csa_tree_add_101_22_pad_groupi_g4822(csa_tree_add_101_22_pad_groupi_n_901 ,csa_tree_add_101_22_pad_groupi_n_761 ,csa_tree_add_101_22_pad_groupi_n_786);
  nor csa_tree_add_101_22_pad_groupi_g4823(csa_tree_add_101_22_pad_groupi_n_900 ,csa_tree_add_101_22_pad_groupi_n_783 ,csa_tree_add_101_22_pad_groupi_n_729);
  or csa_tree_add_101_22_pad_groupi_g4824(csa_tree_add_101_22_pad_groupi_n_899 ,csa_tree_add_101_22_pad_groupi_n_708 ,csa_tree_add_101_22_pad_groupi_n_845);
  or csa_tree_add_101_22_pad_groupi_g4825(csa_tree_add_101_22_pad_groupi_n_898 ,csa_tree_add_101_22_pad_groupi_n_112 ,csa_tree_add_101_22_pad_groupi_n_781);
  and csa_tree_add_101_22_pad_groupi_g4826(csa_tree_add_101_22_pad_groupi_n_897 ,csa_tree_add_101_22_pad_groupi_n_783 ,csa_tree_add_101_22_pad_groupi_n_729);
  and csa_tree_add_101_22_pad_groupi_g4827(csa_tree_add_101_22_pad_groupi_n_896 ,csa_tree_add_101_22_pad_groupi_n_372 ,csa_tree_add_101_22_pad_groupi_n_782);
  or csa_tree_add_101_22_pad_groupi_g4828(csa_tree_add_101_22_pad_groupi_n_895 ,csa_tree_add_101_22_pad_groupi_n_734 ,csa_tree_add_101_22_pad_groupi_n_791);
  nor csa_tree_add_101_22_pad_groupi_g4829(csa_tree_add_101_22_pad_groupi_n_894 ,csa_tree_add_101_22_pad_groupi_n_735 ,csa_tree_add_101_22_pad_groupi_n_792);
  or csa_tree_add_101_22_pad_groupi_g4830(csa_tree_add_101_22_pad_groupi_n_936 ,csa_tree_add_101_22_pad_groupi_n_645 ,csa_tree_add_101_22_pad_groupi_n_833);
  and csa_tree_add_101_22_pad_groupi_g4831(csa_tree_add_101_22_pad_groupi_n_935 ,csa_tree_add_101_22_pad_groupi_n_705 ,csa_tree_add_101_22_pad_groupi_n_767);
  and csa_tree_add_101_22_pad_groupi_g4832(csa_tree_add_101_22_pad_groupi_n_934 ,csa_tree_add_101_22_pad_groupi_n_708 ,csa_tree_add_101_22_pad_groupi_n_845);
  and csa_tree_add_101_22_pad_groupi_g4833(csa_tree_add_101_22_pad_groupi_n_933 ,csa_tree_add_101_22_pad_groupi_n_707 ,csa_tree_add_101_22_pad_groupi_n_844);
  or csa_tree_add_101_22_pad_groupi_g4834(csa_tree_add_101_22_pad_groupi_n_891 ,csa_tree_add_101_22_pad_groupi_n_718 ,csa_tree_add_101_22_pad_groupi_n_793);
  and csa_tree_add_101_22_pad_groupi_g4835(csa_tree_add_101_22_pad_groupi_n_890 ,csa_tree_add_101_22_pad_groupi_n_800 ,csa_tree_add_101_22_pad_groupi_n_799);
  and csa_tree_add_101_22_pad_groupi_g4836(csa_tree_add_101_22_pad_groupi_n_889 ,csa_tree_add_101_22_pad_groupi_n_718 ,csa_tree_add_101_22_pad_groupi_n_793);
  or csa_tree_add_101_22_pad_groupi_g4837(csa_tree_add_101_22_pad_groupi_n_888 ,csa_tree_add_101_22_pad_groupi_n_732 ,csa_tree_add_101_22_pad_groupi_n_754);
  and csa_tree_add_101_22_pad_groupi_g4838(csa_tree_add_101_22_pad_groupi_n_887 ,in21[3] ,csa_tree_add_101_22_pad_groupi_n_804);
  and csa_tree_add_101_22_pad_groupi_g4839(csa_tree_add_101_22_pad_groupi_n_886 ,csa_tree_add_101_22_pad_groupi_n_719 ,csa_tree_add_101_22_pad_groupi_n_720);
  or csa_tree_add_101_22_pad_groupi_g4840(csa_tree_add_101_22_pad_groupi_n_885 ,in21[3] ,csa_tree_add_101_22_pad_groupi_n_804);
  or csa_tree_add_101_22_pad_groupi_g4841(csa_tree_add_101_22_pad_groupi_n_884 ,csa_tree_add_101_22_pad_groupi_n_738 ,csa_tree_add_101_22_pad_groupi_n_727);
  nor csa_tree_add_101_22_pad_groupi_g4842(csa_tree_add_101_22_pad_groupi_n_883 ,csa_tree_add_101_22_pad_groupi_n_803 ,csa_tree_add_101_22_pad_groupi_n_721);
  nor csa_tree_add_101_22_pad_groupi_g4843(csa_tree_add_101_22_pad_groupi_n_882 ,csa_tree_add_101_22_pad_groupi_n_739 ,csa_tree_add_101_22_pad_groupi_n_728);
  nor csa_tree_add_101_22_pad_groupi_g4844(csa_tree_add_101_22_pad_groupi_n_881 ,csa_tree_add_101_22_pad_groupi_n_700 ,csa_tree_add_101_22_pad_groupi_n_828);
  or csa_tree_add_101_22_pad_groupi_g4845(csa_tree_add_101_22_pad_groupi_n_880 ,csa_tree_add_101_22_pad_groupi_n_761 ,csa_tree_add_101_22_pad_groupi_n_786);
  nor csa_tree_add_101_22_pad_groupi_g4846(csa_tree_add_101_22_pad_groupi_n_879 ,csa_tree_add_101_22_pad_groupi_n_371 ,csa_tree_add_101_22_pad_groupi_n_740);
  or csa_tree_add_101_22_pad_groupi_g4847(csa_tree_add_101_22_pad_groupi_n_878 ,csa_tree_add_101_22_pad_groupi_n_387 ,csa_tree_add_101_22_pad_groupi_n_712);
  and csa_tree_add_101_22_pad_groupi_g4848(csa_tree_add_101_22_pad_groupi_n_877 ,csa_tree_add_101_22_pad_groupi_n_766 ,csa_tree_add_101_22_pad_groupi_n_744);
  nor csa_tree_add_101_22_pad_groupi_g4849(csa_tree_add_101_22_pad_groupi_n_876 ,csa_tree_add_101_22_pad_groupi_n_733 ,csa_tree_add_101_22_pad_groupi_n_755);
  nor csa_tree_add_101_22_pad_groupi_g4850(csa_tree_add_101_22_pad_groupi_n_875 ,in21[7] ,csa_tree_add_101_22_pad_groupi_n_713);
  and csa_tree_add_101_22_pad_groupi_g4851(csa_tree_add_101_22_pad_groupi_n_874 ,csa_tree_add_101_22_pad_groupi_n_803 ,csa_tree_add_101_22_pad_groupi_n_721);
  and csa_tree_add_101_22_pad_groupi_g4852(csa_tree_add_101_22_pad_groupi_n_873 ,csa_tree_add_101_22_pad_groupi_n_758 ,csa_tree_add_101_22_pad_groupi_n_757);
  nor csa_tree_add_101_22_pad_groupi_g4853(csa_tree_add_101_22_pad_groupi_n_872 ,csa_tree_add_101_22_pad_groupi_n_764 ,csa_tree_add_101_22_pad_groupi_n_809);
  or csa_tree_add_101_22_pad_groupi_g4854(csa_tree_add_101_22_pad_groupi_n_871 ,csa_tree_add_101_22_pad_groupi_n_758 ,csa_tree_add_101_22_pad_groupi_n_757);
  and csa_tree_add_101_22_pad_groupi_g4855(csa_tree_add_101_22_pad_groupi_n_870 ,in21[2] ,csa_tree_add_101_22_pad_groupi_n_756);
  and csa_tree_add_101_22_pad_groupi_g4856(csa_tree_add_101_22_pad_groupi_n_869 ,csa_tree_add_101_22_pad_groupi_n_808 ,csa_tree_add_101_22_pad_groupi_n_788);
  and csa_tree_add_101_22_pad_groupi_g4857(csa_tree_add_101_22_pad_groupi_n_868 ,csa_tree_add_101_22_pad_groupi_n_784 ,csa_tree_add_101_22_pad_groupi_n_747);
  or csa_tree_add_101_22_pad_groupi_g4858(csa_tree_add_101_22_pad_groupi_n_867 ,csa_tree_add_101_22_pad_groupi_n_810 ,csa_tree_add_101_22_pad_groupi_n_811);
  and csa_tree_add_101_22_pad_groupi_g4859(csa_tree_add_101_22_pad_groupi_n_866 ,csa_tree_add_101_22_pad_groupi_n_765 ,csa_tree_add_101_22_pad_groupi_n_751);
  or csa_tree_add_101_22_pad_groupi_g4860(csa_tree_add_101_22_pad_groupi_n_865 ,csa_tree_add_101_22_pad_groupi_n_784 ,csa_tree_add_101_22_pad_groupi_n_747);
  or csa_tree_add_101_22_pad_groupi_g4861(csa_tree_add_101_22_pad_groupi_n_864 ,csa_tree_add_101_22_pad_groupi_n_749 ,csa_tree_add_101_22_pad_groupi_n_741);
  or csa_tree_add_101_22_pad_groupi_g4862(csa_tree_add_101_22_pad_groupi_n_863 ,csa_tree_add_101_22_pad_groupi_n_765 ,csa_tree_add_101_22_pad_groupi_n_751);
  nor csa_tree_add_101_22_pad_groupi_g4863(csa_tree_add_101_22_pad_groupi_n_862 ,csa_tree_add_101_22_pad_groupi_n_750 ,csa_tree_add_101_22_pad_groupi_n_742);
  nor csa_tree_add_101_22_pad_groupi_g4864(csa_tree_add_101_22_pad_groupi_n_861 ,csa_tree_add_101_22_pad_groupi_n_600 ,csa_tree_add_101_22_pad_groupi_n_822);
  or csa_tree_add_101_22_pad_groupi_g4865(csa_tree_add_101_22_pad_groupi_n_860 ,csa_tree_add_101_22_pad_groupi_n_726 ,csa_tree_add_101_22_pad_groupi_n_821);
  and csa_tree_add_101_22_pad_groupi_g4866(csa_tree_add_101_22_pad_groupi_n_859 ,csa_tree_add_101_22_pad_groupi_n_371 ,csa_tree_add_101_22_pad_groupi_n_740);
  and csa_tree_add_101_22_pad_groupi_g4867(csa_tree_add_101_22_pad_groupi_n_858 ,csa_tree_add_101_22_pad_groupi_n_726 ,csa_tree_add_101_22_pad_groupi_n_821);
  or csa_tree_add_101_22_pad_groupi_g4868(csa_tree_add_101_22_pad_groupi_n_857 ,csa_tree_add_101_22_pad_groupi_n_759 ,csa_tree_add_101_22_pad_groupi_n_736);
  or csa_tree_add_101_22_pad_groupi_g4869(csa_tree_add_101_22_pad_groupi_n_856 ,in21[4] ,csa_tree_add_101_22_pad_groupi_n_798);
  nor csa_tree_add_101_22_pad_groupi_g4870(csa_tree_add_101_22_pad_groupi_n_855 ,in21[2] ,csa_tree_add_101_22_pad_groupi_n_756);
  nor csa_tree_add_101_22_pad_groupi_g4871(csa_tree_add_101_22_pad_groupi_n_854 ,csa_tree_add_101_22_pad_groupi_n_760 ,csa_tree_add_101_22_pad_groupi_n_737);
  or csa_tree_add_101_22_pad_groupi_g4872(csa_tree_add_101_22_pad_groupi_n_853 ,csa_tree_add_101_22_pad_groupi_n_370 ,csa_tree_add_101_22_pad_groupi_n_730);
  or csa_tree_add_101_22_pad_groupi_g4873(csa_tree_add_101_22_pad_groupi_n_852 ,csa_tree_add_101_22_pad_groupi_n_724 ,csa_tree_add_101_22_pad_groupi_n_722);
  nor csa_tree_add_101_22_pad_groupi_g4874(csa_tree_add_101_22_pad_groupi_n_851 ,in21[6] ,csa_tree_add_101_22_pad_groupi_n_731);
  or csa_tree_add_101_22_pad_groupi_g4876(csa_tree_add_101_22_pad_groupi_n_893 ,csa_tree_add_101_22_pad_groupi_n_374 ,csa_tree_add_101_22_pad_groupi_n_826);
  or csa_tree_add_101_22_pad_groupi_g4877(csa_tree_add_101_22_pad_groupi_n_892 ,csa_tree_add_101_22_pad_groupi_n_847 ,csa_tree_add_101_22_pad_groupi_n_849);
  not csa_tree_add_101_22_pad_groupi_g4878(csa_tree_add_101_22_pad_groupi_n_849 ,csa_tree_add_101_22_pad_groupi_n_848);
  not csa_tree_add_101_22_pad_groupi_g4879(csa_tree_add_101_22_pad_groupi_n_847 ,csa_tree_add_101_22_pad_groupi_n_846);
  not csa_tree_add_101_22_pad_groupi_g4880(csa_tree_add_101_22_pad_groupi_n_843 ,csa_tree_add_101_22_pad_groupi_n_842);
  not csa_tree_add_101_22_pad_groupi_g4883(csa_tree_add_101_22_pad_groupi_n_833 ,csa_tree_add_101_22_pad_groupi_n_832);
  not csa_tree_add_101_22_pad_groupi_g4884(csa_tree_add_101_22_pad_groupi_n_826 ,csa_tree_add_101_22_pad_groupi_n_825);
  not csa_tree_add_101_22_pad_groupi_g4885(csa_tree_add_101_22_pad_groupi_n_818 ,csa_tree_add_101_22_pad_groupi_n_819);
  not csa_tree_add_101_22_pad_groupi_g4886(csa_tree_add_101_22_pad_groupi_n_816 ,csa_tree_add_101_22_pad_groupi_n_817);
  not csa_tree_add_101_22_pad_groupi_g4887(csa_tree_add_101_22_pad_groupi_n_812 ,csa_tree_add_101_22_pad_groupi_n_813);
  not csa_tree_add_101_22_pad_groupi_g4888(csa_tree_add_101_22_pad_groupi_n_805 ,csa_tree_add_101_22_pad_groupi_n_806);
  not csa_tree_add_101_22_pad_groupi_g4889(csa_tree_add_101_22_pad_groupi_n_801 ,csa_tree_add_101_22_pad_groupi_n_802);
  not csa_tree_add_101_22_pad_groupi_g4890(csa_tree_add_101_22_pad_groupi_n_794 ,csa_tree_add_101_22_pad_groupi_n_795);
  not csa_tree_add_101_22_pad_groupi_g4891(csa_tree_add_101_22_pad_groupi_n_791 ,csa_tree_add_101_22_pad_groupi_n_792);
  not csa_tree_add_101_22_pad_groupi_g4892(csa_tree_add_101_22_pad_groupi_n_789 ,csa_tree_add_101_22_pad_groupi_n_790);
  and csa_tree_add_101_22_pad_groupi_g4893(csa_tree_add_101_22_pad_groupi_n_781 ,csa_tree_add_101_22_pad_groupi_n_459 ,csa_tree_add_101_22_pad_groupi_n_612);
  or csa_tree_add_101_22_pad_groupi_g4894(csa_tree_add_101_22_pad_groupi_n_848 ,csa_tree_add_101_22_pad_groupi_n_466 ,csa_tree_add_101_22_pad_groupi_n_621);
  or csa_tree_add_101_22_pad_groupi_g4895(csa_tree_add_101_22_pad_groupi_n_846 ,csa_tree_add_101_22_pad_groupi_n_576 ,csa_tree_add_101_22_pad_groupi_n_703);
  and csa_tree_add_101_22_pad_groupi_g4896(csa_tree_add_101_22_pad_groupi_n_845 ,csa_tree_add_101_22_pad_groupi_n_531 ,csa_tree_add_101_22_pad_groupi_n_685);
  or csa_tree_add_101_22_pad_groupi_g4897(csa_tree_add_101_22_pad_groupi_n_844 ,csa_tree_add_101_22_pad_groupi_n_526 ,csa_tree_add_101_22_pad_groupi_n_652);
  or csa_tree_add_101_22_pad_groupi_g4898(csa_tree_add_101_22_pad_groupi_n_842 ,csa_tree_add_101_22_pad_groupi_n_533 ,csa_tree_add_101_22_pad_groupi_n_618);
  and csa_tree_add_101_22_pad_groupi_g4899(csa_tree_add_101_22_pad_groupi_n_841 ,csa_tree_add_101_22_pad_groupi_n_472 ,csa_tree_add_101_22_pad_groupi_n_642);
  or csa_tree_add_101_22_pad_groupi_g4900(csa_tree_add_101_22_pad_groupi_n_840 ,csa_tree_add_101_22_pad_groupi_n_557 ,csa_tree_add_101_22_pad_groupi_n_598);
  or csa_tree_add_101_22_pad_groupi_g4901(csa_tree_add_101_22_pad_groupi_n_839 ,csa_tree_add_101_22_pad_groupi_n_574 ,csa_tree_add_101_22_pad_groupi_n_588);
  and csa_tree_add_101_22_pad_groupi_g4903(csa_tree_add_101_22_pad_groupi_n_837 ,csa_tree_add_101_22_pad_groupi_n_483 ,csa_tree_add_101_22_pad_groupi_n_587);
  and csa_tree_add_101_22_pad_groupi_g4906(csa_tree_add_101_22_pad_groupi_n_834 ,csa_tree_add_101_22_pad_groupi_n_460 ,csa_tree_add_101_22_pad_groupi_n_586);
  or csa_tree_add_101_22_pad_groupi_g4907(csa_tree_add_101_22_pad_groupi_n_832 ,csa_tree_add_101_22_pad_groupi_n_548 ,csa_tree_add_101_22_pad_groupi_n_699);
  or csa_tree_add_101_22_pad_groupi_g4912(csa_tree_add_101_22_pad_groupi_n_827 ,csa_tree_add_101_22_pad_groupi_n_487 ,csa_tree_add_101_22_pad_groupi_n_647);
  or csa_tree_add_101_22_pad_groupi_g4913(csa_tree_add_101_22_pad_groupi_n_825 ,csa_tree_add_101_22_pad_groupi_n_462 ,csa_tree_add_101_22_pad_groupi_n_662);
  and csa_tree_add_101_22_pad_groupi_g4914(csa_tree_add_101_22_pad_groupi_n_824 ,csa_tree_add_101_22_pad_groupi_n_485 ,csa_tree_add_101_22_pad_groupi_n_683);
  and csa_tree_add_101_22_pad_groupi_g4915(csa_tree_add_101_22_pad_groupi_n_823 ,csa_tree_add_101_22_pad_groupi_n_518 ,csa_tree_add_101_22_pad_groupi_n_595);
  or csa_tree_add_101_22_pad_groupi_g4917(csa_tree_add_101_22_pad_groupi_n_821 ,csa_tree_add_101_22_pad_groupi_n_551 ,csa_tree_add_101_22_pad_groupi_n_665);
  or csa_tree_add_101_22_pad_groupi_g4918(csa_tree_add_101_22_pad_groupi_n_820 ,csa_tree_add_101_22_pad_groupi_n_556 ,csa_tree_add_101_22_pad_groupi_n_677);
  or csa_tree_add_101_22_pad_groupi_g4919(csa_tree_add_101_22_pad_groupi_n_819 ,csa_tree_add_101_22_pad_groupi_n_516 ,csa_tree_add_101_22_pad_groupi_n_681);
  or csa_tree_add_101_22_pad_groupi_g4920(csa_tree_add_101_22_pad_groupi_n_817 ,csa_tree_add_101_22_pad_groupi_n_527 ,csa_tree_add_101_22_pad_groupi_n_674);
  or csa_tree_add_101_22_pad_groupi_g4921(csa_tree_add_101_22_pad_groupi_n_815 ,csa_tree_add_101_22_pad_groupi_n_491 ,csa_tree_add_101_22_pad_groupi_n_649);
  or csa_tree_add_101_22_pad_groupi_g4922(csa_tree_add_101_22_pad_groupi_n_814 ,csa_tree_add_101_22_pad_groupi_n_475 ,csa_tree_add_101_22_pad_groupi_n_633);
  or csa_tree_add_101_22_pad_groupi_g4923(csa_tree_add_101_22_pad_groupi_n_813 ,csa_tree_add_101_22_pad_groupi_n_525 ,csa_tree_add_101_22_pad_groupi_n_695);
  or csa_tree_add_101_22_pad_groupi_g4924(csa_tree_add_101_22_pad_groupi_n_811 ,csa_tree_add_101_22_pad_groupi_n_476 ,csa_tree_add_101_22_pad_groupi_n_599);
  or csa_tree_add_101_22_pad_groupi_g4925(csa_tree_add_101_22_pad_groupi_n_810 ,csa_tree_add_101_22_pad_groupi_n_470 ,csa_tree_add_101_22_pad_groupi_n_627);
  or csa_tree_add_101_22_pad_groupi_g4926(csa_tree_add_101_22_pad_groupi_n_809 ,csa_tree_add_101_22_pad_groupi_n_528 ,csa_tree_add_101_22_pad_groupi_n_651);
  or csa_tree_add_101_22_pad_groupi_g4927(csa_tree_add_101_22_pad_groupi_n_808 ,csa_tree_add_101_22_pad_groupi_n_541 ,csa_tree_add_101_22_pad_groupi_n_635);
  or csa_tree_add_101_22_pad_groupi_g4928(csa_tree_add_101_22_pad_groupi_n_807 ,csa_tree_add_101_22_pad_groupi_n_512 ,csa_tree_add_101_22_pad_groupi_n_625);
  or csa_tree_add_101_22_pad_groupi_g4929(csa_tree_add_101_22_pad_groupi_n_806 ,csa_tree_add_101_22_pad_groupi_n_523 ,csa_tree_add_101_22_pad_groupi_n_623);
  or csa_tree_add_101_22_pad_groupi_g4930(csa_tree_add_101_22_pad_groupi_n_804 ,csa_tree_add_101_22_pad_groupi_n_461 ,csa_tree_add_101_22_pad_groupi_n_694);
  or csa_tree_add_101_22_pad_groupi_g4931(csa_tree_add_101_22_pad_groupi_n_803 ,csa_tree_add_101_22_pad_groupi_n_529 ,csa_tree_add_101_22_pad_groupi_n_653);
  or csa_tree_add_101_22_pad_groupi_g4933(csa_tree_add_101_22_pad_groupi_n_800 ,csa_tree_add_101_22_pad_groupi_n_477 ,csa_tree_add_101_22_pad_groupi_n_658);
  or csa_tree_add_101_22_pad_groupi_g4934(csa_tree_add_101_22_pad_groupi_n_799 ,csa_tree_add_101_22_pad_groupi_n_467 ,csa_tree_add_101_22_pad_groupi_n_680);
  or csa_tree_add_101_22_pad_groupi_g4935(csa_tree_add_101_22_pad_groupi_n_798 ,csa_tree_add_101_22_pad_groupi_n_468 ,csa_tree_add_101_22_pad_groupi_n_607);
  or csa_tree_add_101_22_pad_groupi_g4936(csa_tree_add_101_22_pad_groupi_n_797 ,csa_tree_add_101_22_pad_groupi_n_394 ,csa_tree_add_101_22_pad_groupi_n_663);
  or csa_tree_add_101_22_pad_groupi_g4937(csa_tree_add_101_22_pad_groupi_n_796 ,csa_tree_add_101_22_pad_groupi_n_555 ,csa_tree_add_101_22_pad_groupi_n_669);
  or csa_tree_add_101_22_pad_groupi_g4938(csa_tree_add_101_22_pad_groupi_n_795 ,csa_tree_add_101_22_pad_groupi_n_547 ,csa_tree_add_101_22_pad_groupi_n_696);
  or csa_tree_add_101_22_pad_groupi_g4939(csa_tree_add_101_22_pad_groupi_n_793 ,csa_tree_add_101_22_pad_groupi_n_540 ,csa_tree_add_101_22_pad_groupi_n_697);
  or csa_tree_add_101_22_pad_groupi_g4940(csa_tree_add_101_22_pad_groupi_n_792 ,csa_tree_add_101_22_pad_groupi_n_456 ,csa_tree_add_101_22_pad_groupi_n_638);
  or csa_tree_add_101_22_pad_groupi_g4941(csa_tree_add_101_22_pad_groupi_n_790 ,csa_tree_add_101_22_pad_groupi_n_524 ,csa_tree_add_101_22_pad_groupi_n_661);
  or csa_tree_add_101_22_pad_groupi_g4942(csa_tree_add_101_22_pad_groupi_n_788 ,csa_tree_add_101_22_pad_groupi_n_537 ,csa_tree_add_101_22_pad_groupi_n_616);
  or csa_tree_add_101_22_pad_groupi_g4943(csa_tree_add_101_22_pad_groupi_n_787 ,csa_tree_add_101_22_pad_groupi_n_469 ,csa_tree_add_101_22_pad_groupi_n_672);
  or csa_tree_add_101_22_pad_groupi_g4944(csa_tree_add_101_22_pad_groupi_n_786 ,csa_tree_add_101_22_pad_groupi_n_473 ,csa_tree_add_101_22_pad_groupi_n_589);
  or csa_tree_add_101_22_pad_groupi_g4945(csa_tree_add_101_22_pad_groupi_n_785 ,csa_tree_add_101_22_pad_groupi_n_484 ,csa_tree_add_101_22_pad_groupi_n_698);
  or csa_tree_add_101_22_pad_groupi_g4946(csa_tree_add_101_22_pad_groupi_n_784 ,csa_tree_add_101_22_pad_groupi_n_488 ,csa_tree_add_101_22_pad_groupi_n_608);
  or csa_tree_add_101_22_pad_groupi_g4947(csa_tree_add_101_22_pad_groupi_n_783 ,csa_tree_add_101_22_pad_groupi_n_546 ,csa_tree_add_101_22_pad_groupi_n_648);
  not csa_tree_add_101_22_pad_groupi_g4949(csa_tree_add_101_22_pad_groupi_n_779 ,csa_tree_add_101_22_pad_groupi_n_778);
  not csa_tree_add_101_22_pad_groupi_g4950(csa_tree_add_101_22_pad_groupi_n_762 ,csa_tree_add_101_22_pad_groupi_n_763);
  not csa_tree_add_101_22_pad_groupi_g4951(csa_tree_add_101_22_pad_groupi_n_759 ,csa_tree_add_101_22_pad_groupi_n_760);
  not csa_tree_add_101_22_pad_groupi_g4952(csa_tree_add_101_22_pad_groupi_n_754 ,csa_tree_add_101_22_pad_groupi_n_755);
  not csa_tree_add_101_22_pad_groupi_g4953(csa_tree_add_101_22_pad_groupi_n_752 ,csa_tree_add_101_22_pad_groupi_n_753);
  not csa_tree_add_101_22_pad_groupi_g4954(csa_tree_add_101_22_pad_groupi_n_749 ,csa_tree_add_101_22_pad_groupi_n_750);
  not csa_tree_add_101_22_pad_groupi_g4955(csa_tree_add_101_22_pad_groupi_n_745 ,csa_tree_add_101_22_pad_groupi_n_746);
  not csa_tree_add_101_22_pad_groupi_g4956(csa_tree_add_101_22_pad_groupi_n_744 ,csa_tree_add_101_22_pad_groupi_n_743);
  not csa_tree_add_101_22_pad_groupi_g4957(csa_tree_add_101_22_pad_groupi_n_741 ,csa_tree_add_101_22_pad_groupi_n_742);
  not csa_tree_add_101_22_pad_groupi_g4958(csa_tree_add_101_22_pad_groupi_n_738 ,csa_tree_add_101_22_pad_groupi_n_739);
  not csa_tree_add_101_22_pad_groupi_g4959(csa_tree_add_101_22_pad_groupi_n_736 ,csa_tree_add_101_22_pad_groupi_n_737);
  not csa_tree_add_101_22_pad_groupi_g4960(csa_tree_add_101_22_pad_groupi_n_734 ,csa_tree_add_101_22_pad_groupi_n_735);
  not csa_tree_add_101_22_pad_groupi_g4961(csa_tree_add_101_22_pad_groupi_n_732 ,csa_tree_add_101_22_pad_groupi_n_733);
  not csa_tree_add_101_22_pad_groupi_g4962(csa_tree_add_101_22_pad_groupi_n_730 ,csa_tree_add_101_22_pad_groupi_n_731);
  not csa_tree_add_101_22_pad_groupi_g4963(csa_tree_add_101_22_pad_groupi_n_727 ,csa_tree_add_101_22_pad_groupi_n_728);
  not csa_tree_add_101_22_pad_groupi_g4964(csa_tree_add_101_22_pad_groupi_n_724 ,csa_tree_add_101_22_pad_groupi_n_725);
  not csa_tree_add_101_22_pad_groupi_g4965(csa_tree_add_101_22_pad_groupi_n_722 ,csa_tree_add_101_22_pad_groupi_n_723);
  not csa_tree_add_101_22_pad_groupi_g4966(csa_tree_add_101_22_pad_groupi_n_715 ,csa_tree_add_101_22_pad_groupi_n_716);
  not csa_tree_add_101_22_pad_groupi_g4967(csa_tree_add_101_22_pad_groupi_n_712 ,csa_tree_add_101_22_pad_groupi_n_713);
  xnor csa_tree_add_101_22_pad_groupi_g4968(csa_tree_add_101_22_pad_groupi_n_711 ,csa_tree_add_101_22_pad_groupi_n_583 ,in21[10]);
  xnor csa_tree_add_101_22_pad_groupi_g4970(csa_tree_add_101_22_pad_groupi_n_710 ,csa_tree_add_101_22_pad_groupi_n_282 ,in21[12]);
  xnor csa_tree_add_101_22_pad_groupi_g4972(csa_tree_add_101_22_pad_groupi_n_709 ,csa_tree_add_101_22_pad_groupi_n_582 ,in21[12]);
  or csa_tree_add_101_22_pad_groupi_g4975(csa_tree_add_101_22_pad_groupi_n_778 ,csa_tree_add_101_22_pad_groupi_n_539 ,csa_tree_add_101_22_pad_groupi_n_626);
  or csa_tree_add_101_22_pad_groupi_g4976(csa_tree_add_101_22_pad_groupi_n_777 ,csa_tree_add_101_22_pad_groupi_n_550 ,csa_tree_add_101_22_pad_groupi_n_624);
  and csa_tree_add_101_22_pad_groupi_g4977(csa_tree_add_101_22_pad_groupi_n_776 ,csa_tree_add_101_22_pad_groupi_n_464 ,csa_tree_add_101_22_pad_groupi_n_655);
  or csa_tree_add_101_22_pad_groupi_g4978(csa_tree_add_101_22_pad_groupi_n_775 ,csa_tree_add_101_22_pad_groupi_n_482 ,csa_tree_add_101_22_pad_groupi_n_637);
  or csa_tree_add_101_22_pad_groupi_g4980(csa_tree_add_101_22_pad_groupi_n_773 ,csa_tree_add_101_22_pad_groupi_n_519 ,csa_tree_add_101_22_pad_groupi_n_605);
  and csa_tree_add_101_22_pad_groupi_g4981(csa_tree_add_101_22_pad_groupi_n_772 ,csa_tree_add_101_22_pad_groupi_n_457 ,csa_tree_add_101_22_pad_groupi_n_594);
  and csa_tree_add_101_22_pad_groupi_g4982(csa_tree_add_101_22_pad_groupi_n_771 ,csa_tree_add_101_22_pad_groupi_n_492 ,csa_tree_add_101_22_pad_groupi_n_606);
  or csa_tree_add_101_22_pad_groupi_g4984(csa_tree_add_101_22_pad_groupi_n_769 ,csa_tree_add_101_22_pad_groupi_n_490 ,csa_tree_add_101_22_pad_groupi_n_689);
  or csa_tree_add_101_22_pad_groupi_g4985(csa_tree_add_101_22_pad_groupi_n_768 ,csa_tree_add_101_22_pad_groupi_n_545 ,csa_tree_add_101_22_pad_groupi_n_640);
  or csa_tree_add_101_22_pad_groupi_g4986(csa_tree_add_101_22_pad_groupi_n_767 ,csa_tree_add_101_22_pad_groupi_n_552 ,csa_tree_add_101_22_pad_groupi_n_659);
  or csa_tree_add_101_22_pad_groupi_g4988(csa_tree_add_101_22_pad_groupi_n_765 ,csa_tree_add_101_22_pad_groupi_n_517 ,csa_tree_add_101_22_pad_groupi_n_688);
  or csa_tree_add_101_22_pad_groupi_g4989(csa_tree_add_101_22_pad_groupi_n_764 ,csa_tree_add_101_22_pad_groupi_n_554 ,csa_tree_add_101_22_pad_groupi_n_654);
  or csa_tree_add_101_22_pad_groupi_g4990(csa_tree_add_101_22_pad_groupi_n_763 ,csa_tree_add_101_22_pad_groupi_n_480 ,csa_tree_add_101_22_pad_groupi_n_602);
  or csa_tree_add_101_22_pad_groupi_g4991(csa_tree_add_101_22_pad_groupi_n_761 ,csa_tree_add_101_22_pad_groupi_n_577 ,csa_tree_add_101_22_pad_groupi_n_693);
  or csa_tree_add_101_22_pad_groupi_g4992(csa_tree_add_101_22_pad_groupi_n_760 ,csa_tree_add_101_22_pad_groupi_n_478 ,csa_tree_add_101_22_pad_groupi_n_591);
  or csa_tree_add_101_22_pad_groupi_g4993(csa_tree_add_101_22_pad_groupi_n_758 ,csa_tree_add_101_22_pad_groupi_n_514 ,csa_tree_add_101_22_pad_groupi_n_604);
  or csa_tree_add_101_22_pad_groupi_g4994(csa_tree_add_101_22_pad_groupi_n_757 ,csa_tree_add_101_22_pad_groupi_n_532 ,csa_tree_add_101_22_pad_groupi_n_617);
  or csa_tree_add_101_22_pad_groupi_g4995(csa_tree_add_101_22_pad_groupi_n_756 ,csa_tree_add_101_22_pad_groupi_n_455 ,csa_tree_add_101_22_pad_groupi_n_670);
  or csa_tree_add_101_22_pad_groupi_g4996(csa_tree_add_101_22_pad_groupi_n_755 ,csa_tree_add_101_22_pad_groupi_n_544 ,csa_tree_add_101_22_pad_groupi_n_660);
  or csa_tree_add_101_22_pad_groupi_g4997(csa_tree_add_101_22_pad_groupi_n_753 ,csa_tree_add_101_22_pad_groupi_n_486 ,csa_tree_add_101_22_pad_groupi_n_679);
  or csa_tree_add_101_22_pad_groupi_g4998(csa_tree_add_101_22_pad_groupi_n_751 ,csa_tree_add_101_22_pad_groupi_n_575 ,csa_tree_add_101_22_pad_groupi_n_619);
  or csa_tree_add_101_22_pad_groupi_g4999(csa_tree_add_101_22_pad_groupi_n_750 ,csa_tree_add_101_22_pad_groupi_n_522 ,csa_tree_add_101_22_pad_groupi_n_671);
  or csa_tree_add_101_22_pad_groupi_g5000(csa_tree_add_101_22_pad_groupi_n_748 ,csa_tree_add_101_22_pad_groupi_n_515 ,csa_tree_add_101_22_pad_groupi_n_631);
  or csa_tree_add_101_22_pad_groupi_g5001(csa_tree_add_101_22_pad_groupi_n_747 ,csa_tree_add_101_22_pad_groupi_n_573 ,csa_tree_add_101_22_pad_groupi_n_620);
  or csa_tree_add_101_22_pad_groupi_g5002(csa_tree_add_101_22_pad_groupi_n_746 ,csa_tree_add_101_22_pad_groupi_n_534 ,csa_tree_add_101_22_pad_groupi_n_643);
  or csa_tree_add_101_22_pad_groupi_g5003(csa_tree_add_101_22_pad_groupi_n_743 ,csa_tree_add_101_22_pad_groupi_n_481 ,csa_tree_add_101_22_pad_groupi_n_629);
  or csa_tree_add_101_22_pad_groupi_g5004(csa_tree_add_101_22_pad_groupi_n_742 ,csa_tree_add_101_22_pad_groupi_n_536 ,csa_tree_add_101_22_pad_groupi_n_650);
  or csa_tree_add_101_22_pad_groupi_g5006(csa_tree_add_101_22_pad_groupi_n_739 ,csa_tree_add_101_22_pad_groupi_n_564 ,csa_tree_add_101_22_pad_groupi_n_628);
  or csa_tree_add_101_22_pad_groupi_g5007(csa_tree_add_101_22_pad_groupi_n_737 ,csa_tree_add_101_22_pad_groupi_n_513 ,csa_tree_add_101_22_pad_groupi_n_603);
  or csa_tree_add_101_22_pad_groupi_g5008(csa_tree_add_101_22_pad_groupi_n_735 ,csa_tree_add_101_22_pad_groupi_n_553 ,csa_tree_add_101_22_pad_groupi_n_691);
  or csa_tree_add_101_22_pad_groupi_g5009(csa_tree_add_101_22_pad_groupi_n_733 ,csa_tree_add_101_22_pad_groupi_n_530 ,csa_tree_add_101_22_pad_groupi_n_622);
  or csa_tree_add_101_22_pad_groupi_g5010(csa_tree_add_101_22_pad_groupi_n_731 ,csa_tree_add_101_22_pad_groupi_n_463 ,csa_tree_add_101_22_pad_groupi_n_590);
  or csa_tree_add_101_22_pad_groupi_g5011(csa_tree_add_101_22_pad_groupi_n_729 ,csa_tree_add_101_22_pad_groupi_n_471 ,csa_tree_add_101_22_pad_groupi_n_610);
  or csa_tree_add_101_22_pad_groupi_g5012(csa_tree_add_101_22_pad_groupi_n_728 ,csa_tree_add_101_22_pad_groupi_n_520 ,csa_tree_add_101_22_pad_groupi_n_639);
  or csa_tree_add_101_22_pad_groupi_g5013(csa_tree_add_101_22_pad_groupi_n_726 ,csa_tree_add_101_22_pad_groupi_n_535 ,csa_tree_add_101_22_pad_groupi_n_690);
  or csa_tree_add_101_22_pad_groupi_g5014(csa_tree_add_101_22_pad_groupi_n_725 ,csa_tree_add_101_22_pad_groupi_n_538 ,csa_tree_add_101_22_pad_groupi_n_675);
  or csa_tree_add_101_22_pad_groupi_g5015(csa_tree_add_101_22_pad_groupi_n_723 ,csa_tree_add_101_22_pad_groupi_n_543 ,csa_tree_add_101_22_pad_groupi_n_676);
  or csa_tree_add_101_22_pad_groupi_g5016(csa_tree_add_101_22_pad_groupi_n_721 ,csa_tree_add_101_22_pad_groupi_n_542 ,csa_tree_add_101_22_pad_groupi_n_634);
  or csa_tree_add_101_22_pad_groupi_g5017(csa_tree_add_101_22_pad_groupi_n_720 ,csa_tree_add_101_22_pad_groupi_n_479 ,csa_tree_add_101_22_pad_groupi_n_644);
  or csa_tree_add_101_22_pad_groupi_g5018(csa_tree_add_101_22_pad_groupi_n_719 ,csa_tree_add_101_22_pad_groupi_n_521 ,csa_tree_add_101_22_pad_groupi_n_611);
  or csa_tree_add_101_22_pad_groupi_g5019(csa_tree_add_101_22_pad_groupi_n_718 ,csa_tree_add_101_22_pad_groupi_n_489 ,csa_tree_add_101_22_pad_groupi_n_609);
  or csa_tree_add_101_22_pad_groupi_g5020(csa_tree_add_101_22_pad_groupi_n_717 ,csa_tree_add_101_22_pad_groupi_n_549 ,csa_tree_add_101_22_pad_groupi_n_692);
  or csa_tree_add_101_22_pad_groupi_g5021(csa_tree_add_101_22_pad_groupi_n_716 ,csa_tree_add_101_22_pad_groupi_n_465 ,csa_tree_add_101_22_pad_groupi_n_613);
  or csa_tree_add_101_22_pad_groupi_g5022(csa_tree_add_101_22_pad_groupi_n_714 ,csa_tree_add_101_22_pad_groupi_n_474 ,csa_tree_add_101_22_pad_groupi_n_657);
  or csa_tree_add_101_22_pad_groupi_g5023(csa_tree_add_101_22_pad_groupi_n_713 ,csa_tree_add_101_22_pad_groupi_n_458 ,csa_tree_add_101_22_pad_groupi_n_667);
  not csa_tree_add_101_22_pad_groupi_g5024(csa_tree_add_101_22_pad_groupi_n_707 ,csa_tree_add_101_22_pad_groupi_n_706);
  not csa_tree_add_101_22_pad_groupi_g5025(csa_tree_add_101_22_pad_groupi_n_705 ,csa_tree_add_101_22_pad_groupi_n_704);
  nor csa_tree_add_101_22_pad_groupi_g5026(csa_tree_add_101_22_pad_groupi_n_703 ,csa_tree_add_101_22_pad_groupi_n_113 ,csa_tree_add_101_22_pad_groupi_n_218);
  nor csa_tree_add_101_22_pad_groupi_g5027(csa_tree_add_101_22_pad_groupi_n_702 ,in21[9] ,csa_tree_add_101_22_pad_groupi_n_358);
  nor csa_tree_add_101_22_pad_groupi_g5029(csa_tree_add_101_22_pad_groupi_n_700 ,in21[12] ,csa_tree_add_101_22_pad_groupi_n_579);
  nor csa_tree_add_101_22_pad_groupi_g5030(csa_tree_add_101_22_pad_groupi_n_699 ,csa_tree_add_101_22_pad_groupi_n_115 ,csa_tree_add_101_22_pad_groupi_n_189);
  and csa_tree_add_101_22_pad_groupi_g5031(csa_tree_add_101_22_pad_groupi_n_698 ,in9[5] ,csa_tree_add_101_22_pad_groupi_n_172);
  nor csa_tree_add_101_22_pad_groupi_g5032(csa_tree_add_101_22_pad_groupi_n_697 ,csa_tree_add_101_22_pad_groupi_n_119 ,csa_tree_add_101_22_pad_groupi_n_38);
  nor csa_tree_add_101_22_pad_groupi_g5033(csa_tree_add_101_22_pad_groupi_n_696 ,csa_tree_add_101_22_pad_groupi_n_93 ,csa_tree_add_101_22_pad_groupi_n_66);
  and csa_tree_add_101_22_pad_groupi_g5034(csa_tree_add_101_22_pad_groupi_n_695 ,in9[2] ,csa_tree_add_101_22_pad_groupi_n_133);
  and csa_tree_add_101_22_pad_groupi_g5035(csa_tree_add_101_22_pad_groupi_n_694 ,in9[10] ,csa_tree_add_101_22_pad_groupi_n_433);
  and csa_tree_add_101_22_pad_groupi_g5036(csa_tree_add_101_22_pad_groupi_n_693 ,in9[8] ,csa_tree_add_101_22_pad_groupi_n_287);
  and csa_tree_add_101_22_pad_groupi_g5037(csa_tree_add_101_22_pad_groupi_n_692 ,in9[14] ,csa_tree_add_101_22_pad_groupi_n_169);
  and csa_tree_add_101_22_pad_groupi_g5038(csa_tree_add_101_22_pad_groupi_n_691 ,in9[1] ,csa_tree_add_101_22_pad_groupi_n_168);
  and csa_tree_add_101_22_pad_groupi_g5039(csa_tree_add_101_22_pad_groupi_n_690 ,in9[5] ,csa_tree_add_101_22_pad_groupi_n_142);
  and csa_tree_add_101_22_pad_groupi_g5040(csa_tree_add_101_22_pad_groupi_n_689 ,in9[7] ,csa_tree_add_101_22_pad_groupi_n_126);
  and csa_tree_add_101_22_pad_groupi_g5041(csa_tree_add_101_22_pad_groupi_n_688 ,in9[11] ,csa_tree_add_101_22_pad_groupi_n_285);
  or csa_tree_add_101_22_pad_groupi_g5044(csa_tree_add_101_22_pad_groupi_n_685 ,csa_tree_add_101_22_pad_groupi_n_17 ,csa_tree_add_101_22_pad_groupi_n_118);
  or csa_tree_add_101_22_pad_groupi_g5046(csa_tree_add_101_22_pad_groupi_n_683 ,csa_tree_add_101_22_pad_groupi_n_149 ,csa_tree_add_101_22_pad_groupi_n_583);
  and csa_tree_add_101_22_pad_groupi_g5047(csa_tree_add_101_22_pad_groupi_n_682 ,in21[12] ,csa_tree_add_101_22_pad_groupi_n_579);
  and csa_tree_add_101_22_pad_groupi_g5048(csa_tree_add_101_22_pad_groupi_n_681 ,in9[11] ,csa_tree_add_101_22_pad_groupi_n_135);
  and csa_tree_add_101_22_pad_groupi_g5049(csa_tree_add_101_22_pad_groupi_n_680 ,in9[6] ,csa_tree_add_101_22_pad_groupi_n_445);
  nor csa_tree_add_101_22_pad_groupi_g5050(csa_tree_add_101_22_pad_groupi_n_679 ,csa_tree_add_101_22_pad_groupi_n_252 ,csa_tree_add_101_22_pad_groupi_n_223);
  and csa_tree_add_101_22_pad_groupi_g5052(csa_tree_add_101_22_pad_groupi_n_677 ,in9[3] ,csa_tree_add_101_22_pad_groupi_n_139);
  and csa_tree_add_101_22_pad_groupi_g5053(csa_tree_add_101_22_pad_groupi_n_676 ,in9[6] ,csa_tree_add_101_22_pad_groupi_n_136);
  and csa_tree_add_101_22_pad_groupi_g5054(csa_tree_add_101_22_pad_groupi_n_675 ,in9[4] ,csa_tree_add_101_22_pad_groupi_n_144);
  and csa_tree_add_101_22_pad_groupi_g5055(csa_tree_add_101_22_pad_groupi_n_674 ,in9[4] ,csa_tree_add_101_22_pad_groupi_n_138);
  nor csa_tree_add_101_22_pad_groupi_g5056(csa_tree_add_101_22_pad_groupi_n_673 ,csa_tree_add_101_22_pad_groupi_n_369 ,csa_tree_add_101_22_pad_groupi_n_581);
  and csa_tree_add_101_22_pad_groupi_g5057(csa_tree_add_101_22_pad_groupi_n_672 ,in9[12] ,csa_tree_add_101_22_pad_groupi_n_428);
  and csa_tree_add_101_22_pad_groupi_g5058(csa_tree_add_101_22_pad_groupi_n_671 ,in9[4] ,csa_tree_add_101_22_pad_groupi_n_124);
  and csa_tree_add_101_22_pad_groupi_g5059(csa_tree_add_101_22_pad_groupi_n_670 ,in9[9] ,csa_tree_add_101_22_pad_groupi_n_439);
  and csa_tree_add_101_22_pad_groupi_g5060(csa_tree_add_101_22_pad_groupi_n_669 ,in9[14] ,csa_tree_add_101_22_pad_groupi_n_288);
  and csa_tree_add_101_22_pad_groupi_g5062(csa_tree_add_101_22_pad_groupi_n_667 ,in9[14] ,csa_tree_add_101_22_pad_groupi_n_425);
  and csa_tree_add_101_22_pad_groupi_g5063(csa_tree_add_101_22_pad_groupi_n_666 ,in21[12] ,csa_tree_add_101_22_pad_groupi_n_280);
  and csa_tree_add_101_22_pad_groupi_g5064(csa_tree_add_101_22_pad_groupi_n_665 ,in9[7] ,csa_tree_add_101_22_pad_groupi_n_171);
  and csa_tree_add_101_22_pad_groupi_g5066(csa_tree_add_101_22_pad_groupi_n_663 ,csa_tree_add_101_22_pad_groupi_n_406 ,csa_tree_add_101_22_pad_groupi_n_583);
  and csa_tree_add_101_22_pad_groupi_g5067(csa_tree_add_101_22_pad_groupi_n_662 ,in9[7] ,csa_tree_add_101_22_pad_groupi_n_429);
  and csa_tree_add_101_22_pad_groupi_g5068(csa_tree_add_101_22_pad_groupi_n_661 ,in9[9] ,csa_tree_add_101_22_pad_groupi_n_145);
  and csa_tree_add_101_22_pad_groupi_g5069(csa_tree_add_101_22_pad_groupi_n_660 ,in9[14] ,csa_tree_add_101_22_pad_groupi_n_127);
  nor csa_tree_add_101_22_pad_groupi_g5070(csa_tree_add_101_22_pad_groupi_n_659 ,csa_tree_add_101_22_pad_groupi_n_112 ,csa_tree_add_101_22_pad_groupi_n_202);
  and csa_tree_add_101_22_pad_groupi_g5071(csa_tree_add_101_22_pad_groupi_n_658 ,in9[3] ,csa_tree_add_101_22_pad_groupi_n_133);
  nor csa_tree_add_101_22_pad_groupi_g5072(csa_tree_add_101_22_pad_groupi_n_657 ,csa_tree_add_101_22_pad_groupi_n_118 ,csa_tree_add_101_22_pad_groupi_n_215);
  or csa_tree_add_101_22_pad_groupi_g5073(csa_tree_add_101_22_pad_groupi_n_656 ,csa_tree_add_101_22_pad_groupi_n_373 ,csa_tree_add_101_22_pad_groupi_n_357);
  or csa_tree_add_101_22_pad_groupi_g5074(csa_tree_add_101_22_pad_groupi_n_655 ,csa_tree_add_101_22_pad_groupi_n_27 ,csa_tree_add_101_22_pad_groupi_n_427);
  and csa_tree_add_101_22_pad_groupi_g5075(csa_tree_add_101_22_pad_groupi_n_654 ,in9[11] ,csa_tree_add_101_22_pad_groupi_n_130);
  and csa_tree_add_101_22_pad_groupi_g5076(csa_tree_add_101_22_pad_groupi_n_653 ,in9[1] ,csa_tree_add_101_22_pad_groupi_n_147);
  nor csa_tree_add_101_22_pad_groupi_g5077(csa_tree_add_101_22_pad_groupi_n_652 ,csa_tree_add_101_22_pad_groupi_n_93 ,csa_tree_add_101_22_pad_groupi_n_74);
  and csa_tree_add_101_22_pad_groupi_g5078(csa_tree_add_101_22_pad_groupi_n_651 ,in9[13] ,csa_tree_add_101_22_pad_groupi_n_148);
  and csa_tree_add_101_22_pad_groupi_g5079(csa_tree_add_101_22_pad_groupi_n_650 ,in9[6] ,csa_tree_add_101_22_pad_groupi_n_148);
  and csa_tree_add_101_22_pad_groupi_g5080(csa_tree_add_101_22_pad_groupi_n_649 ,in9[12] ,csa_tree_add_101_22_pad_groupi_n_142);
  and csa_tree_add_101_22_pad_groupi_g5081(csa_tree_add_101_22_pad_groupi_n_648 ,in9[3] ,csa_tree_add_101_22_pad_groupi_n_129);
  and csa_tree_add_101_22_pad_groupi_g5082(csa_tree_add_101_22_pad_groupi_n_647 ,in9[4] ,csa_tree_add_101_22_pad_groupi_n_284);
  or csa_tree_add_101_22_pad_groupi_g5084(csa_tree_add_101_22_pad_groupi_n_706 ,csa_tree_add_101_22_pad_groupi_n_24 ,csa_tree_add_101_22_pad_groupi_n_502);
  or csa_tree_add_101_22_pad_groupi_g5085(csa_tree_add_101_22_pad_groupi_n_704 ,csa_tree_add_101_22_pad_groupi_n_24 ,csa_tree_add_101_22_pad_groupi_n_257);
  nor csa_tree_add_101_22_pad_groupi_g5086(csa_tree_add_101_22_pad_groupi_n_644 ,csa_tree_add_101_22_pad_groupi_n_113 ,csa_tree_add_101_22_pad_groupi_n_178);
  nor csa_tree_add_101_22_pad_groupi_g5087(csa_tree_add_101_22_pad_groupi_n_643 ,csa_tree_add_101_22_pad_groupi_n_160 ,csa_tree_add_101_22_pad_groupi_n_578);
  or csa_tree_add_101_22_pad_groupi_g5088(csa_tree_add_101_22_pad_groupi_n_642 ,csa_tree_add_101_22_pad_groupi_n_47 ,csa_tree_add_101_22_pad_groupi_n_497);
  and csa_tree_add_101_22_pad_groupi_g5090(csa_tree_add_101_22_pad_groupi_n_640 ,in9[6] ,csa_tree_add_101_22_pad_groupi_n_130);
  and csa_tree_add_101_22_pad_groupi_g5091(csa_tree_add_101_22_pad_groupi_n_639 ,in9[13] ,csa_tree_add_101_22_pad_groupi_n_171);
  nor csa_tree_add_101_22_pad_groupi_g5092(csa_tree_add_101_22_pad_groupi_n_638 ,csa_tree_add_101_22_pad_groupi_n_87 ,csa_tree_add_101_22_pad_groupi_n_434);
  and csa_tree_add_101_22_pad_groupi_g5093(csa_tree_add_101_22_pad_groupi_n_637 ,in9[10] ,csa_tree_add_101_22_pad_groupi_n_166);
  nor csa_tree_add_101_22_pad_groupi_g5095(csa_tree_add_101_22_pad_groupi_n_635 ,csa_tree_add_101_22_pad_groupi_n_96 ,csa_tree_add_101_22_pad_groupi_n_255);
  and csa_tree_add_101_22_pad_groupi_g5096(csa_tree_add_101_22_pad_groupi_n_634 ,in9[2] ,csa_tree_add_101_22_pad_groupi_n_168);
  and csa_tree_add_101_22_pad_groupi_g5097(csa_tree_add_101_22_pad_groupi_n_633 ,in9[13] ,csa_tree_add_101_22_pad_groupi_n_124);
  nor csa_tree_add_101_22_pad_groupi_g5099(csa_tree_add_101_22_pad_groupi_n_631 ,csa_tree_add_101_22_pad_groupi_n_231 ,csa_tree_add_101_22_pad_groupi_n_257);
  and csa_tree_add_101_22_pad_groupi_g5101(csa_tree_add_101_22_pad_groupi_n_629 ,in9[13] ,csa_tree_add_101_22_pad_groupi_n_287);
  and csa_tree_add_101_22_pad_groupi_g5102(csa_tree_add_101_22_pad_groupi_n_628 ,in9[11] ,csa_tree_add_101_22_pad_groupi_n_145);
  and csa_tree_add_101_22_pad_groupi_g5103(csa_tree_add_101_22_pad_groupi_n_627 ,in9[7] ,csa_tree_add_101_22_pad_groupi_n_141);
  nor csa_tree_add_101_22_pad_groupi_g5104(csa_tree_add_101_22_pad_groupi_n_626 ,csa_tree_add_101_22_pad_groupi_n_71 ,csa_tree_add_101_22_pad_groupi_n_507);
  and csa_tree_add_101_22_pad_groupi_g5105(csa_tree_add_101_22_pad_groupi_n_625 ,in9[7] ,csa_tree_add_101_22_pad_groupi_n_285);
  and csa_tree_add_101_22_pad_groupi_g5106(csa_tree_add_101_22_pad_groupi_n_624 ,in9[5] ,csa_tree_add_101_22_pad_groupi_n_165);
  and csa_tree_add_101_22_pad_groupi_g5107(csa_tree_add_101_22_pad_groupi_n_623 ,in9[10] ,csa_tree_add_101_22_pad_groupi_n_132);
  nor csa_tree_add_101_22_pad_groupi_g5108(csa_tree_add_101_22_pad_groupi_n_622 ,csa_tree_add_101_22_pad_groupi_n_159 ,csa_tree_add_101_22_pad_groupi_n_282);
  nor csa_tree_add_101_22_pad_groupi_g5109(csa_tree_add_101_22_pad_groupi_n_621 ,csa_tree_add_101_22_pad_groupi_n_98 ,csa_tree_add_101_22_pad_groupi_n_430);
  nor csa_tree_add_101_22_pad_groupi_g5110(csa_tree_add_101_22_pad_groupi_n_620 ,csa_tree_add_101_22_pad_groupi_n_194 ,csa_tree_add_101_22_pad_groupi_n_502);
  nor csa_tree_add_101_22_pad_groupi_g5111(csa_tree_add_101_22_pad_groupi_n_619 ,csa_tree_add_101_22_pad_groupi_n_116 ,csa_tree_add_101_22_pad_groupi_n_187);
  and csa_tree_add_101_22_pad_groupi_g5112(csa_tree_add_101_22_pad_groupi_n_618 ,in9[8] ,csa_tree_add_101_22_pad_groupi_n_165);
  and csa_tree_add_101_22_pad_groupi_g5113(csa_tree_add_101_22_pad_groupi_n_617 ,in9[8] ,csa_tree_add_101_22_pad_groupi_n_136);
  nor csa_tree_add_101_22_pad_groupi_g5114(csa_tree_add_101_22_pad_groupi_n_616 ,csa_tree_add_101_22_pad_groupi_n_119 ,csa_tree_add_101_22_pad_groupi_n_181);
  nor csa_tree_add_101_22_pad_groupi_g5117(csa_tree_add_101_22_pad_groupi_n_613 ,csa_tree_add_101_22_pad_groupi_n_204 ,csa_tree_add_101_22_pad_groupi_n_432);
  or csa_tree_add_101_22_pad_groupi_g5118(csa_tree_add_101_22_pad_groupi_n_612 ,csa_tree_add_101_22_pad_groupi_n_64 ,csa_tree_add_101_22_pad_groupi_n_438);
  and csa_tree_add_101_22_pad_groupi_g5119(csa_tree_add_101_22_pad_groupi_n_611 ,in9[8] ,csa_tree_add_101_22_pad_groupi_n_284);
  nor csa_tree_add_101_22_pad_groupi_g5120(csa_tree_add_101_22_pad_groupi_n_610 ,csa_tree_add_101_22_pad_groupi_n_116 ,csa_tree_add_101_22_pad_groupi_n_184);
  nor csa_tree_add_101_22_pad_groupi_g5121(csa_tree_add_101_22_pad_groupi_n_609 ,csa_tree_add_101_22_pad_groupi_n_91 ,csa_tree_add_101_22_pad_groupi_n_501);
  and csa_tree_add_101_22_pad_groupi_g5122(csa_tree_add_101_22_pad_groupi_n_608 ,in9[12] ,csa_tree_add_101_22_pad_groupi_n_166);
  and csa_tree_add_101_22_pad_groupi_g5123(csa_tree_add_101_22_pad_groupi_n_607 ,in9[11] ,csa_tree_add_101_22_pad_groupi_n_431);
  or csa_tree_add_101_22_pad_groupi_g5124(csa_tree_add_101_22_pad_groupi_n_606 ,csa_tree_add_101_22_pad_groupi_n_17 ,csa_tree_add_101_22_pad_groupi_n_255);
  and csa_tree_add_101_22_pad_groupi_g5125(csa_tree_add_101_22_pad_groupi_n_605 ,in9[9] ,csa_tree_add_101_22_pad_groupi_n_127);
  nor csa_tree_add_101_22_pad_groupi_g5126(csa_tree_add_101_22_pad_groupi_n_604 ,csa_tree_add_101_22_pad_groupi_n_211 ,csa_tree_add_101_22_pad_groupi_n_508);
  and csa_tree_add_101_22_pad_groupi_g5127(csa_tree_add_101_22_pad_groupi_n_603 ,in9[12] ,csa_tree_add_101_22_pad_groupi_n_169);
  and csa_tree_add_101_22_pad_groupi_g5128(csa_tree_add_101_22_pad_groupi_n_602 ,in9[1] ,csa_tree_add_101_22_pad_groupi_n_123);
  nor csa_tree_add_101_22_pad_groupi_g5130(csa_tree_add_101_22_pad_groupi_n_600 ,in21[12] ,csa_tree_add_101_22_pad_groupi_n_582);
  and csa_tree_add_101_22_pad_groupi_g5131(csa_tree_add_101_22_pad_groupi_n_599 ,in9[9] ,csa_tree_add_101_22_pad_groupi_n_139);
  nor csa_tree_add_101_22_pad_groupi_g5132(csa_tree_add_101_22_pad_groupi_n_598 ,csa_tree_add_101_22_pad_groupi_n_101 ,csa_tree_add_101_22_pad_groupi_n_508);
  or csa_tree_add_101_22_pad_groupi_g5135(csa_tree_add_101_22_pad_groupi_n_595 ,csa_tree_add_101_22_pad_groupi_n_55 ,csa_tree_add_101_22_pad_groupi_n_115);
  or csa_tree_add_101_22_pad_groupi_g5136(csa_tree_add_101_22_pad_groupi_n_594 ,csa_tree_add_101_22_pad_groupi_n_50 ,csa_tree_add_101_22_pad_groupi_n_426);
  nor csa_tree_add_101_22_pad_groupi_g5137(csa_tree_add_101_22_pad_groupi_n_593 ,in21[11] ,csa_tree_add_101_22_pad_groupi_n_580);
  and csa_tree_add_101_22_pad_groupi_g5139(csa_tree_add_101_22_pad_groupi_n_591 ,in9[10] ,csa_tree_add_101_22_pad_groupi_n_288);
  and csa_tree_add_101_22_pad_groupi_g5140(csa_tree_add_101_22_pad_groupi_n_590 ,in9[13] ,csa_tree_add_101_22_pad_groupi_n_435);
  and csa_tree_add_101_22_pad_groupi_g5141(csa_tree_add_101_22_pad_groupi_n_589 ,in9[10] ,csa_tree_add_101_22_pad_groupi_n_172);
  nor csa_tree_add_101_22_pad_groupi_g5142(csa_tree_add_101_22_pad_groupi_n_588 ,csa_tree_add_101_22_pad_groupi_n_158 ,csa_tree_add_101_22_pad_groupi_n_280);
  or csa_tree_add_101_22_pad_groupi_g5143(csa_tree_add_101_22_pad_groupi_n_587 ,csa_tree_add_101_22_pad_groupi_n_151 ,csa_tree_add_101_22_pad_groupi_n_580);
  or csa_tree_add_101_22_pad_groupi_g5144(csa_tree_add_101_22_pad_groupi_n_586 ,csa_tree_add_101_22_pad_groupi_n_15 ,csa_tree_add_101_22_pad_groupi_n_581);
  or csa_tree_add_101_22_pad_groupi_g5145(csa_tree_add_101_22_pad_groupi_n_646 ,csa_tree_add_101_22_pad_groupi_n_57 ,csa_tree_add_101_22_pad_groupi_n_493);
  or csa_tree_add_101_22_pad_groupi_g5146(csa_tree_add_101_22_pad_groupi_n_645 ,csa_tree_add_101_22_pad_groupi_n_42 ,csa_tree_add_101_22_pad_groupi_n_278);
  nor csa_tree_add_101_22_pad_groupi_g5150(csa_tree_add_101_22_pad_groupi_n_577 ,csa_tree_add_101_22_pad_groupi_n_183 ,csa_tree_add_101_22_pad_groupi_n_332);
  nor csa_tree_add_101_22_pad_groupi_g5151(csa_tree_add_101_22_pad_groupi_n_576 ,csa_tree_add_101_22_pad_groupi_n_42 ,csa_tree_add_101_22_pad_groupi_n_302);
  nor csa_tree_add_101_22_pad_groupi_g5152(csa_tree_add_101_22_pad_groupi_n_575 ,csa_tree_add_101_22_pad_groupi_n_233 ,csa_tree_add_101_22_pad_groupi_n_306);
  nor csa_tree_add_101_22_pad_groupi_g5153(csa_tree_add_101_22_pad_groupi_n_574 ,csa_tree_add_101_22_pad_groupi_n_193 ,csa_tree_add_101_22_pad_groupi_n_341);
  nor csa_tree_add_101_22_pad_groupi_g5154(csa_tree_add_101_22_pad_groupi_n_573 ,csa_tree_add_101_22_pad_groupi_n_84 ,csa_tree_add_101_22_pad_groupi_n_312);
  nor csa_tree_add_101_22_pad_groupi_g5163(csa_tree_add_101_22_pad_groupi_n_564 ,csa_tree_add_101_22_pad_groupi_n_78 ,csa_tree_add_101_22_pad_groupi_n_330);
  nor csa_tree_add_101_22_pad_groupi_g5170(csa_tree_add_101_22_pad_groupi_n_557 ,csa_tree_add_101_22_pad_groupi_n_71 ,csa_tree_add_101_22_pad_groupi_n_335);
  nor csa_tree_add_101_22_pad_groupi_g5171(csa_tree_add_101_22_pad_groupi_n_556 ,csa_tree_add_101_22_pad_groupi_n_101 ,csa_tree_add_101_22_pad_groupi_n_315);
  nor csa_tree_add_101_22_pad_groupi_g5172(csa_tree_add_101_22_pad_groupi_n_555 ,csa_tree_add_101_22_pad_groupi_n_186 ,csa_tree_add_101_22_pad_groupi_n_336);
  nor csa_tree_add_101_22_pad_groupi_g5173(csa_tree_add_101_22_pad_groupi_n_554 ,csa_tree_add_101_22_pad_groupi_n_177 ,csa_tree_add_101_22_pad_groupi_n_309);
  nor csa_tree_add_101_22_pad_groupi_g5174(csa_tree_add_101_22_pad_groupi_n_553 ,csa_tree_add_101_22_pad_groupi_n_244 ,csa_tree_add_101_22_pad_groupi_n_320);
  nor csa_tree_add_101_22_pad_groupi_g5175(csa_tree_add_101_22_pad_groupi_n_552 ,csa_tree_add_101_22_pad_groupi_n_247 ,csa_tree_add_101_22_pad_groupi_n_323);
  nor csa_tree_add_101_22_pad_groupi_g5176(csa_tree_add_101_22_pad_groupi_n_551 ,csa_tree_add_101_22_pad_groupi_n_67 ,csa_tree_add_101_22_pad_groupi_n_317);
  nor csa_tree_add_101_22_pad_groupi_g5177(csa_tree_add_101_22_pad_groupi_n_550 ,csa_tree_add_101_22_pad_groupi_n_175 ,csa_tree_add_101_22_pad_groupi_n_339);
  nor csa_tree_add_101_22_pad_groupi_g5178(csa_tree_add_101_22_pad_groupi_n_549 ,csa_tree_add_101_22_pad_groupi_n_85 ,csa_tree_add_101_22_pad_groupi_n_321);
  nor csa_tree_add_101_22_pad_groupi_g5179(csa_tree_add_101_22_pad_groupi_n_548 ,csa_tree_add_101_22_pad_groupi_n_88 ,csa_tree_add_101_22_pad_groupi_n_305);
  nor csa_tree_add_101_22_pad_groupi_g5180(csa_tree_add_101_22_pad_groupi_n_547 ,csa_tree_add_101_22_pad_groupi_n_197 ,csa_tree_add_101_22_pad_groupi_n_323);
  nor csa_tree_add_101_22_pad_groupi_g5181(csa_tree_add_101_22_pad_groupi_n_546 ,csa_tree_add_101_22_pad_groupi_n_100 ,csa_tree_add_101_22_pad_groupi_n_326);
  nor csa_tree_add_101_22_pad_groupi_g5182(csa_tree_add_101_22_pad_groupi_n_545 ,csa_tree_add_101_22_pad_groupi_n_53 ,csa_tree_add_101_22_pad_groupi_n_327);
  nor csa_tree_add_101_22_pad_groupi_g5183(csa_tree_add_101_22_pad_groupi_n_544 ,csa_tree_add_101_22_pad_groupi_n_187 ,csa_tree_add_101_22_pad_groupi_n_326);
  nor csa_tree_add_101_22_pad_groupi_g5184(csa_tree_add_101_22_pad_groupi_n_543 ,csa_tree_add_101_22_pad_groupi_n_196 ,csa_tree_add_101_22_pad_groupi_n_317);
  nor csa_tree_add_101_22_pad_groupi_g5185(csa_tree_add_101_22_pad_groupi_n_542 ,csa_tree_add_101_22_pad_groupi_n_217 ,csa_tree_add_101_22_pad_groupi_n_318);
  nor csa_tree_add_101_22_pad_groupi_g5186(csa_tree_add_101_22_pad_groupi_n_541 ,csa_tree_add_101_22_pad_groupi_n_209 ,csa_tree_add_101_22_pad_groupi_n_344);
  nor csa_tree_add_101_22_pad_groupi_g5187(csa_tree_add_101_22_pad_groupi_n_540 ,csa_tree_add_101_22_pad_groupi_n_229 ,csa_tree_add_101_22_pad_groupi_n_324);
  nor csa_tree_add_101_22_pad_groupi_g5188(csa_tree_add_101_22_pad_groupi_n_539 ,csa_tree_add_101_22_pad_groupi_n_41 ,csa_tree_add_101_22_pad_groupi_n_335);
  nor csa_tree_add_101_22_pad_groupi_g5189(csa_tree_add_101_22_pad_groupi_n_538 ,csa_tree_add_101_22_pad_groupi_n_36 ,csa_tree_add_101_22_pad_groupi_n_336);
  nor csa_tree_add_101_22_pad_groupi_g5190(csa_tree_add_101_22_pad_groupi_n_537 ,csa_tree_add_101_22_pad_groupi_n_79 ,csa_tree_add_101_22_pad_groupi_n_324);
  nor csa_tree_add_101_22_pad_groupi_g5191(csa_tree_add_101_22_pad_groupi_n_536 ,csa_tree_add_101_22_pad_groupi_n_204 ,csa_tree_add_101_22_pad_groupi_n_345);
  nor csa_tree_add_101_22_pad_groupi_g5192(csa_tree_add_101_22_pad_groupi_n_535 ,csa_tree_add_101_22_pad_groupi_n_28 ,csa_tree_add_101_22_pad_groupi_n_329);
  nor csa_tree_add_101_22_pad_groupi_g5193(csa_tree_add_101_22_pad_groupi_n_534 ,csa_tree_add_101_22_pad_groupi_n_194 ,csa_tree_add_101_22_pad_groupi_n_327);
  nor csa_tree_add_101_22_pad_groupi_g5194(csa_tree_add_101_22_pad_groupi_n_533 ,csa_tree_add_101_22_pad_groupi_n_191 ,csa_tree_add_101_22_pad_groupi_n_338);
  nor csa_tree_add_101_22_pad_groupi_g5195(csa_tree_add_101_22_pad_groupi_n_532 ,csa_tree_add_101_22_pad_groupi_n_184 ,csa_tree_add_101_22_pad_groupi_n_318);
  or csa_tree_add_101_22_pad_groupi_g5196(csa_tree_add_101_22_pad_groupi_n_531 ,csa_tree_add_101_22_pad_groupi_n_174 ,csa_tree_add_101_22_pad_groupi_n_305);
  nor csa_tree_add_101_22_pad_groupi_g5197(csa_tree_add_101_22_pad_groupi_n_530 ,csa_tree_add_101_22_pad_groupi_n_39 ,csa_tree_add_101_22_pad_groupi_n_330);
  nor csa_tree_add_101_22_pad_groupi_g5198(csa_tree_add_101_22_pad_groupi_n_529 ,csa_tree_add_101_22_pad_groupi_n_243 ,csa_tree_add_101_22_pad_groupi_n_344);
  nor csa_tree_add_101_22_pad_groupi_g5199(csa_tree_add_101_22_pad_groupi_n_528 ,csa_tree_add_101_22_pad_groupi_n_91 ,csa_tree_add_101_22_pad_groupi_n_345);
  nor csa_tree_add_101_22_pad_groupi_g5200(csa_tree_add_101_22_pad_groupi_n_527 ,csa_tree_add_101_22_pad_groupi_n_231 ,csa_tree_add_101_22_pad_groupi_n_321);
  nor csa_tree_add_101_22_pad_groupi_g5201(csa_tree_add_101_22_pad_groupi_n_526 ,csa_tree_add_101_22_pad_groupi_n_217 ,csa_tree_add_101_22_pad_groupi_n_265);
  nor csa_tree_add_101_22_pad_groupi_g5202(csa_tree_add_101_22_pad_groupi_n_525 ,csa_tree_add_101_22_pad_groupi_n_64 ,csa_tree_add_101_22_pad_groupi_n_311);
  nor csa_tree_add_101_22_pad_groupi_g5203(csa_tree_add_101_22_pad_groupi_n_524 ,csa_tree_add_101_22_pad_groupi_n_55 ,csa_tree_add_101_22_pad_groupi_n_269);
  nor csa_tree_add_101_22_pad_groupi_g5204(csa_tree_add_101_22_pad_groupi_n_523 ,csa_tree_add_101_22_pad_groupi_n_76 ,csa_tree_add_101_22_pad_groupi_n_312);
  nor csa_tree_add_101_22_pad_groupi_g5205(csa_tree_add_101_22_pad_groupi_n_522 ,csa_tree_add_101_22_pad_groupi_n_201 ,csa_tree_add_101_22_pad_groupi_n_339);
  nor csa_tree_add_101_22_pad_groupi_g5206(csa_tree_add_101_22_pad_groupi_n_521 ,csa_tree_add_101_22_pad_groupi_n_22 ,csa_tree_add_101_22_pad_groupi_n_275);
  nor csa_tree_add_101_22_pad_groupi_g5207(csa_tree_add_101_22_pad_groupi_n_520 ,csa_tree_add_101_22_pad_groupi_n_222 ,csa_tree_add_101_22_pad_groupi_n_262);
  nor csa_tree_add_101_22_pad_groupi_g5208(csa_tree_add_101_22_pad_groupi_n_519 ,csa_tree_add_101_22_pad_groupi_n_50 ,csa_tree_add_101_22_pad_groupi_n_272);
  or csa_tree_add_101_22_pad_groupi_g5209(csa_tree_add_101_22_pad_groupi_n_518 ,csa_tree_add_101_22_pad_groupi_n_21 ,csa_tree_add_101_22_pad_groupi_n_266);
  nor csa_tree_add_101_22_pad_groupi_g5210(csa_tree_add_101_22_pad_groupi_n_517 ,csa_tree_add_101_22_pad_groupi_n_178 ,csa_tree_add_101_22_pad_groupi_n_274);
  nor csa_tree_add_101_22_pad_groupi_g5211(csa_tree_add_101_22_pad_groupi_n_516 ,csa_tree_add_101_22_pad_groupi_n_225 ,csa_tree_add_101_22_pad_groupi_n_263);
  nor csa_tree_add_101_22_pad_groupi_g5212(csa_tree_add_101_22_pad_groupi_n_515 ,csa_tree_add_101_22_pad_groupi_n_47 ,csa_tree_add_101_22_pad_groupi_n_268);
  nor csa_tree_add_101_22_pad_groupi_g5213(csa_tree_add_101_22_pad_groupi_n_514 ,csa_tree_add_101_22_pad_groupi_n_197 ,csa_tree_add_101_22_pad_groupi_n_333);
  nor csa_tree_add_101_22_pad_groupi_g5214(csa_tree_add_101_22_pad_groupi_n_513 ,csa_tree_add_101_22_pad_groupi_n_227 ,csa_tree_add_101_22_pad_groupi_n_320);
  nor csa_tree_add_101_22_pad_groupi_g5215(csa_tree_add_101_22_pad_groupi_n_512 ,csa_tree_add_101_22_pad_groupi_n_59 ,csa_tree_add_101_22_pad_groupi_n_342);
  or csa_tree_add_101_22_pad_groupi_g5217(csa_tree_add_101_22_pad_groupi_n_583 ,csa_tree_add_101_22_pad_groupi_n_121 ,csa_tree_add_101_22_pad_groupi_n_424);
  or csa_tree_add_101_22_pad_groupi_g5218(csa_tree_add_101_22_pad_groupi_n_582 ,csa_tree_add_101_22_pad_groupi_n_162 ,csa_tree_add_101_22_pad_groupi_n_402);
  or csa_tree_add_101_22_pad_groupi_g5219(csa_tree_add_101_22_pad_groupi_n_581 ,csa_tree_add_101_22_pad_groupi_n_121 ,csa_tree_add_101_22_pad_groupi_n_109);
  or csa_tree_add_101_22_pad_groupi_g5220(csa_tree_add_101_22_pad_groupi_n_580 ,csa_tree_add_101_22_pad_groupi_n_162 ,csa_tree_add_101_22_pad_groupi_n_404);
  or csa_tree_add_101_22_pad_groupi_g5221(csa_tree_add_101_22_pad_groupi_n_579 ,csa_tree_add_101_22_pad_groupi_n_163 ,csa_tree_add_101_22_pad_groupi_n_403);
  not csa_tree_add_101_22_pad_groupi_g5223(csa_tree_add_101_22_pad_groupi_n_510 ,csa_tree_add_101_22_pad_groupi_n_505);
  not csa_tree_add_101_22_pad_groupi_g5224(csa_tree_add_101_22_pad_groupi_n_509 ,csa_tree_add_101_22_pad_groupi_n_505);
  not csa_tree_add_101_22_pad_groupi_g5225(csa_tree_add_101_22_pad_groupi_n_508 ,csa_tree_add_101_22_pad_groupi_n_506);
  not csa_tree_add_101_22_pad_groupi_g5226(csa_tree_add_101_22_pad_groupi_n_507 ,csa_tree_add_101_22_pad_groupi_n_506);
  not csa_tree_add_101_22_pad_groupi_g5227(csa_tree_add_101_22_pad_groupi_n_506 ,csa_tree_add_101_22_pad_groupi_n_505);
  not csa_tree_add_101_22_pad_groupi_g5228(csa_tree_add_101_22_pad_groupi_n_504 ,csa_tree_add_101_22_pad_groupi_n_499);
  not csa_tree_add_101_22_pad_groupi_g5229(csa_tree_add_101_22_pad_groupi_n_503 ,csa_tree_add_101_22_pad_groupi_n_499);
  not csa_tree_add_101_22_pad_groupi_g5230(csa_tree_add_101_22_pad_groupi_n_502 ,csa_tree_add_101_22_pad_groupi_n_500);
  not csa_tree_add_101_22_pad_groupi_g5231(csa_tree_add_101_22_pad_groupi_n_501 ,csa_tree_add_101_22_pad_groupi_n_500);
  not csa_tree_add_101_22_pad_groupi_g5232(csa_tree_add_101_22_pad_groupi_n_500 ,csa_tree_add_101_22_pad_groupi_n_499);
  not csa_tree_add_101_22_pad_groupi_g5233(csa_tree_add_101_22_pad_groupi_n_498 ,csa_tree_add_101_22_pad_groupi_n_278);
  not csa_tree_add_101_22_pad_groupi_g5234(csa_tree_add_101_22_pad_groupi_n_496 ,csa_tree_add_101_22_pad_groupi_n_497);
  not csa_tree_add_101_22_pad_groupi_g5235(csa_tree_add_101_22_pad_groupi_n_495 ,csa_tree_add_101_22_pad_groupi_n_493);
  not csa_tree_add_101_22_pad_groupi_g5236(csa_tree_add_101_22_pad_groupi_n_494 ,csa_tree_add_101_22_pad_groupi_n_493);
  or csa_tree_add_101_22_pad_groupi_g5237(csa_tree_add_101_22_pad_groupi_n_492 ,csa_tree_add_101_22_pad_groupi_n_27 ,csa_tree_add_101_22_pad_groupi_n_311);
  nor csa_tree_add_101_22_pad_groupi_g5238(csa_tree_add_101_22_pad_groupi_n_491 ,csa_tree_add_101_22_pad_groupi_n_180 ,csa_tree_add_101_22_pad_groupi_n_329);
  nor csa_tree_add_101_22_pad_groupi_g5239(csa_tree_add_101_22_pad_groupi_n_490 ,csa_tree_add_101_22_pad_groupi_n_220 ,csa_tree_add_101_22_pad_groupi_n_271);
  nor csa_tree_add_101_22_pad_groupi_g5240(csa_tree_add_101_22_pad_groupi_n_489 ,csa_tree_add_101_22_pad_groupi_n_82 ,csa_tree_add_101_22_pad_groupi_n_275);
  nor csa_tree_add_101_22_pad_groupi_g5241(csa_tree_add_101_22_pad_groupi_n_488 ,csa_tree_add_101_22_pad_groupi_n_181 ,csa_tree_add_101_22_pad_groupi_n_309);
  nor csa_tree_add_101_22_pad_groupi_g5242(csa_tree_add_101_22_pad_groupi_n_487 ,csa_tree_add_101_22_pad_groupi_n_88 ,csa_tree_add_101_22_pad_groupi_n_341);
  nor csa_tree_add_101_22_pad_groupi_g5243(csa_tree_add_101_22_pad_groupi_n_486 ,csa_tree_add_101_22_pad_groupi_n_227 ,csa_tree_add_101_22_pad_groupi_n_306);
  or csa_tree_add_101_22_pad_groupi_g5244(csa_tree_add_101_22_pad_groupi_n_485 ,csa_tree_add_101_22_pad_groupi_n_30 ,csa_tree_add_101_22_pad_groupi_n_302);
  nor csa_tree_add_101_22_pad_groupi_g5245(csa_tree_add_101_22_pad_groupi_n_484 ,csa_tree_add_101_22_pad_groupi_n_174 ,csa_tree_add_101_22_pad_groupi_n_315);
  or csa_tree_add_101_22_pad_groupi_g5246(csa_tree_add_101_22_pad_groupi_n_483 ,csa_tree_add_101_22_pad_groupi_n_30 ,csa_tree_add_101_22_pad_groupi_n_263);
  nor csa_tree_add_101_22_pad_groupi_g5247(csa_tree_add_101_22_pad_groupi_n_482 ,csa_tree_add_101_22_pad_groupi_n_96 ,csa_tree_add_101_22_pad_groupi_n_338);
  nor csa_tree_add_101_22_pad_groupi_g5248(csa_tree_add_101_22_pad_groupi_n_481 ,csa_tree_add_101_22_pad_groupi_n_233 ,csa_tree_add_101_22_pad_groupi_n_269);
  nor csa_tree_add_101_22_pad_groupi_g5249(csa_tree_add_101_22_pad_groupi_n_480 ,csa_tree_add_101_22_pad_groupi_n_25 ,csa_tree_add_101_22_pad_groupi_n_272);
  nor csa_tree_add_101_22_pad_groupi_g5250(csa_tree_add_101_22_pad_groupi_n_479 ,csa_tree_add_101_22_pad_groupi_n_214 ,csa_tree_add_101_22_pad_groupi_n_266);
  nor csa_tree_add_101_22_pad_groupi_g5251(csa_tree_add_101_22_pad_groupi_n_478 ,csa_tree_add_101_22_pad_groupi_n_235 ,csa_tree_add_101_22_pad_groupi_n_332);
  nor csa_tree_add_101_22_pad_groupi_g5252(csa_tree_add_101_22_pad_groupi_n_477 ,csa_tree_add_101_22_pad_groupi_n_73 ,csa_tree_add_101_22_pad_groupi_n_342);
  nor csa_tree_add_101_22_pad_groupi_g5253(csa_tree_add_101_22_pad_groupi_n_476 ,csa_tree_add_101_22_pad_groupi_n_206 ,csa_tree_add_101_22_pad_groupi_n_314);
  nor csa_tree_add_101_22_pad_groupi_g5254(csa_tree_add_101_22_pad_groupi_n_475 ,csa_tree_add_101_22_pad_groupi_n_69 ,csa_tree_add_101_22_pad_groupi_n_308);
  nor csa_tree_add_101_22_pad_groupi_g5255(csa_tree_add_101_22_pad_groupi_n_474 ,csa_tree_add_101_22_pad_groupi_n_209 ,csa_tree_add_101_22_pad_groupi_n_303);
  nor csa_tree_add_101_22_pad_groupi_g5256(csa_tree_add_101_22_pad_groupi_n_473 ,csa_tree_add_101_22_pad_groupi_n_76 ,csa_tree_add_101_22_pad_groupi_n_314);
  or csa_tree_add_101_22_pad_groupi_g5257(csa_tree_add_101_22_pad_groupi_n_472 ,csa_tree_add_101_22_pad_groupi_n_45 ,csa_tree_add_101_22_pad_groupi_n_308);
  nor csa_tree_add_101_22_pad_groupi_g5258(csa_tree_add_101_22_pad_groupi_n_471 ,csa_tree_add_101_22_pad_groupi_n_211 ,csa_tree_add_101_22_pad_groupi_n_303);
  nor csa_tree_add_101_22_pad_groupi_g5259(csa_tree_add_101_22_pad_groupi_n_470 ,csa_tree_add_101_22_pad_groupi_n_67 ,csa_tree_add_101_22_pad_groupi_n_333);
  nor csa_tree_add_101_22_pad_groupi_g5260(csa_tree_add_101_22_pad_groupi_n_469 ,csa_tree_add_101_22_pad_groupi_n_180 ,csa_tree_add_101_22_pad_groupi_n_300);
  nor csa_tree_add_101_22_pad_groupi_g5261(csa_tree_add_101_22_pad_groupi_n_468 ,csa_tree_add_101_22_pad_groupi_n_177 ,csa_tree_add_101_22_pad_groupi_n_399);
  nor csa_tree_add_101_22_pad_groupi_g5262(csa_tree_add_101_22_pad_groupi_n_467 ,csa_tree_add_101_22_pad_groupi_n_52 ,csa_tree_add_101_22_pad_groupi_n_291);
  nor csa_tree_add_101_22_pad_groupi_g5263(csa_tree_add_101_22_pad_groupi_n_466 ,csa_tree_add_101_22_pad_groupi_n_45 ,csa_tree_add_101_22_pad_groupi_n_290);
  nor csa_tree_add_101_22_pad_groupi_g5264(csa_tree_add_101_22_pad_groupi_n_465 ,csa_tree_add_101_22_pad_groupi_n_175 ,csa_tree_add_101_22_pad_groupi_n_297);
  or csa_tree_add_101_22_pad_groupi_g5265(csa_tree_add_101_22_pad_groupi_n_464 ,csa_tree_add_101_22_pad_groupi_n_36 ,csa_tree_add_101_22_pad_groupi_n_296);
  nor csa_tree_add_101_22_pad_groupi_g5266(csa_tree_add_101_22_pad_groupi_n_463 ,csa_tree_add_101_22_pad_groupi_n_90 ,csa_tree_add_101_22_pad_groupi_n_260);
  nor csa_tree_add_101_22_pad_groupi_g5267(csa_tree_add_101_22_pad_groupi_n_462 ,csa_tree_add_101_22_pad_groupi_n_212 ,csa_tree_add_101_22_pad_groupi_n_299);
  nor csa_tree_add_101_22_pad_groupi_g5268(csa_tree_add_101_22_pad_groupi_n_461 ,csa_tree_add_101_22_pad_groupi_n_95 ,csa_tree_add_101_22_pad_groupi_n_299);
  or csa_tree_add_101_22_pad_groupi_g5269(csa_tree_add_101_22_pad_groupi_n_460 ,csa_tree_add_101_22_pad_groupi_n_39 ,csa_tree_add_101_22_pad_groupi_n_290);
  nor csa_tree_add_101_22_pad_groupi_g5271(csa_tree_add_101_22_pad_groupi_n_458 ,csa_tree_add_101_22_pad_groupi_n_186 ,csa_tree_add_101_22_pad_groupi_n_300);
  or csa_tree_add_101_22_pad_groupi_g5272(csa_tree_add_101_22_pad_groupi_n_457 ,csa_tree_add_101_22_pad_groupi_n_21 ,csa_tree_add_101_22_pad_groupi_n_291);
  nor csa_tree_add_101_22_pad_groupi_g5273(csa_tree_add_101_22_pad_groupi_n_456 ,csa_tree_add_101_22_pad_groupi_n_98 ,csa_tree_add_101_22_pad_groupi_n_296);
  nor csa_tree_add_101_22_pad_groupi_g5274(csa_tree_add_101_22_pad_groupi_n_455 ,csa_tree_add_101_22_pad_groupi_n_207 ,csa_tree_add_101_22_pad_groupi_n_297);
  nor csa_tree_add_101_22_pad_groupi_g5284(csa_tree_add_101_22_pad_groupi_n_445 ,csa_tree_add_101_22_pad_groupi_n_106 ,csa_tree_add_101_22_pad_groupi_n_294);
  nor csa_tree_add_101_22_pad_groupi_g5290(csa_tree_add_101_22_pad_groupi_n_439 ,csa_tree_add_101_22_pad_groupi_n_109 ,csa_tree_add_101_22_pad_groupi_n_241);
  or csa_tree_add_101_22_pad_groupi_g5291(csa_tree_add_101_22_pad_groupi_n_438 ,csa_tree_add_101_22_pad_groupi_n_32 ,csa_tree_add_101_22_pad_groupi_n_103);
  nor csa_tree_add_101_22_pad_groupi_g5294(csa_tree_add_101_22_pad_groupi_n_435 ,csa_tree_add_101_22_pad_groupi_n_107 ,csa_tree_add_101_22_pad_groupi_n_240);
  or csa_tree_add_101_22_pad_groupi_g5295(csa_tree_add_101_22_pad_groupi_n_434 ,csa_tree_add_101_22_pad_groupi_n_293 ,csa_tree_add_101_22_pad_groupi_n_110);
  nor csa_tree_add_101_22_pad_groupi_g5296(csa_tree_add_101_22_pad_groupi_n_433 ,csa_tree_add_101_22_pad_groupi_n_103 ,csa_tree_add_101_22_pad_groupi_n_294);
  or csa_tree_add_101_22_pad_groupi_g5297(csa_tree_add_101_22_pad_groupi_n_432 ,csa_tree_add_101_22_pad_groupi_n_13 ,csa_tree_add_101_22_pad_groupi_n_61);
  nor csa_tree_add_101_22_pad_groupi_g5298(csa_tree_add_101_22_pad_groupi_n_431 ,csa_tree_add_101_22_pad_groupi_n_110 ,csa_tree_add_101_22_pad_groupi_n_238);
  or csa_tree_add_101_22_pad_groupi_g5299(csa_tree_add_101_22_pad_groupi_n_430 ,csa_tree_add_101_22_pad_groupi_n_13 ,csa_tree_add_101_22_pad_groupi_n_104);
  nor csa_tree_add_101_22_pad_groupi_g5300(csa_tree_add_101_22_pad_groupi_n_429 ,csa_tree_add_101_22_pad_groupi_n_61 ,csa_tree_add_101_22_pad_groupi_n_32);
  nor csa_tree_add_101_22_pad_groupi_g5301(csa_tree_add_101_22_pad_groupi_n_428 ,csa_tree_add_101_22_pad_groupi_n_249 ,csa_tree_add_101_22_pad_groupi_n_34);
  or csa_tree_add_101_22_pad_groupi_g5302(csa_tree_add_101_22_pad_groupi_n_427 ,csa_tree_add_101_22_pad_groupi_n_15 ,csa_tree_add_101_22_pad_groupi_n_106);
  or csa_tree_add_101_22_pad_groupi_g5303(csa_tree_add_101_22_pad_groupi_n_426 ,csa_tree_add_101_22_pad_groupi_n_34 ,csa_tree_add_101_22_pad_groupi_n_107);
  nor csa_tree_add_101_22_pad_groupi_g5304(csa_tree_add_101_22_pad_groupi_n_425 ,csa_tree_add_101_22_pad_groupi_n_104 ,csa_tree_add_101_22_pad_groupi_n_237);
  or csa_tree_add_101_22_pad_groupi_g5305(csa_tree_add_101_22_pad_groupi_n_511 ,csa_tree_add_101_22_pad_groupi_n_154 ,csa_tree_add_101_22_pad_groupi_n_424);
  or csa_tree_add_101_22_pad_groupi_g5306(csa_tree_add_101_22_pad_groupi_n_505 ,csa_tree_add_101_22_pad_groupi_n_150 ,csa_tree_add_101_22_pad_groupi_n_403);
  or csa_tree_add_101_22_pad_groupi_g5307(csa_tree_add_101_22_pad_groupi_n_499 ,csa_tree_add_101_22_pad_groupi_n_155 ,csa_tree_add_101_22_pad_groupi_n_402);
  or csa_tree_add_101_22_pad_groupi_g5309(csa_tree_add_101_22_pad_groupi_n_493 ,csa_tree_add_101_22_pad_groupi_n_152 ,csa_tree_add_101_22_pad_groupi_n_404);
  not csa_tree_add_101_22_pad_groupi_g5311(csa_tree_add_101_22_pad_groupi_n_423 ,csa_tree_add_101_22_pad_groupi_n_158);
  not csa_tree_add_101_22_pad_groupi_g5312(csa_tree_add_101_22_pad_groupi_n_422 ,csa_tree_add_101_22_pad_groupi_n_155);
  not csa_tree_add_101_22_pad_groupi_g5315(csa_tree_add_101_22_pad_groupi_n_419 ,csa_tree_add_101_22_pad_groupi_n_154);
  not csa_tree_add_101_22_pad_groupi_g5317(csa_tree_add_101_22_pad_groupi_n_418 ,csa_tree_add_101_22_pad_groupi_n_149);
  not csa_tree_add_101_22_pad_groupi_g5319(csa_tree_add_101_22_pad_groupi_n_416 ,csa_tree_add_101_22_pad_groupi_n_152);
  not csa_tree_add_101_22_pad_groupi_g5321(csa_tree_add_101_22_pad_groupi_n_415 ,csa_tree_add_101_22_pad_groupi_n_151);
  not csa_tree_add_101_22_pad_groupi_g5323(csa_tree_add_101_22_pad_groupi_n_414 ,csa_tree_add_101_22_pad_groupi_n_160);
  not csa_tree_add_101_22_pad_groupi_g5324(csa_tree_add_101_22_pad_groupi_n_413 ,csa_tree_add_101_22_pad_groupi_n_153);
  not csa_tree_add_101_22_pad_groupi_g5327(csa_tree_add_101_22_pad_groupi_n_411 ,csa_tree_add_101_22_pad_groupi_n_159);
  not csa_tree_add_101_22_pad_groupi_g5328(csa_tree_add_101_22_pad_groupi_n_410 ,csa_tree_add_101_22_pad_groupi_n_150);
  or csa_tree_add_101_22_pad_groupi_g5331(csa_tree_add_101_22_pad_groupi_n_406 ,in21[10] ,in21[9]);
  and csa_tree_add_101_22_pad_groupi_g5332(csa_tree_add_101_22_pad_groupi_n_424 ,csa_tree_add_101_22_pad_groupi_n_375 ,csa_tree_add_101_22_pad_groupi_n_388);
  and csa_tree_add_101_22_pad_groupi_g5333(csa_tree_add_101_22_pad_groupi_n_421 ,n_627 ,n_634);
  and csa_tree_add_101_22_pad_groupi_g5334(csa_tree_add_101_22_pad_groupi_n_420 ,in22[0] ,n_636);
  and csa_tree_add_101_22_pad_groupi_g5335(csa_tree_add_101_22_pad_groupi_n_417 ,n_628 ,n_635);
  and csa_tree_add_101_22_pad_groupi_g5337(csa_tree_add_101_22_pad_groupi_n_409 ,n_626 ,n_633);
  not csa_tree_add_101_22_pad_groupi_g5339(csa_tree_add_101_22_pad_groupi_n_399 ,csa_tree_add_101_22_pad_groupi_n_293);
  not csa_tree_add_101_22_pad_groupi_g5340(csa_tree_add_101_22_pad_groupi_n_398 ,csa_tree_add_101_22_pad_groupi_n_395);
  not csa_tree_add_101_22_pad_groupi_g5341(csa_tree_add_101_22_pad_groupi_n_397 ,csa_tree_add_101_22_pad_groupi_n_258);
  not csa_tree_add_101_22_pad_groupi_g5345(csa_tree_add_101_22_pad_groupi_n_396 ,csa_tree_add_101_22_pad_groupi_n_395);
  and csa_tree_add_101_22_pad_groupi_g5346(csa_tree_add_101_22_pad_groupi_n_394 ,in21[10] ,in21[9]);
  and csa_tree_add_101_22_pad_groupi_g5348(csa_tree_add_101_22_pad_groupi_n_404 ,csa_tree_add_101_22_pad_groupi_n_391 ,csa_tree_add_101_22_pad_groupi_n_393);
  and csa_tree_add_101_22_pad_groupi_g5349(csa_tree_add_101_22_pad_groupi_n_403 ,csa_tree_add_101_22_pad_groupi_n_378 ,csa_tree_add_101_22_pad_groupi_n_377);
  and csa_tree_add_101_22_pad_groupi_g5350(csa_tree_add_101_22_pad_groupi_n_402 ,csa_tree_add_101_22_pad_groupi_n_392 ,csa_tree_add_101_22_pad_groupi_n_376);
  and csa_tree_add_101_22_pad_groupi_g5351(csa_tree_add_101_22_pad_groupi_n_401 ,csa_tree_add_101_22_pad_groupi_n_390 ,csa_tree_add_101_22_pad_groupi_n_389);
  or csa_tree_add_101_22_pad_groupi_g5353(csa_tree_add_101_22_pad_groupi_n_395 ,csa_tree_add_101_22_pad_groupi_n_390 ,csa_tree_add_101_22_pad_groupi_n_389);
  not csa_tree_add_101_22_pad_groupi_g5354(csa_tree_add_101_22_pad_groupi_n_393 ,n_635);
  not csa_tree_add_101_22_pad_groupi_g5355(csa_tree_add_101_22_pad_groupi_n_392 ,n_627);
  not csa_tree_add_101_22_pad_groupi_g5356(csa_tree_add_101_22_pad_groupi_n_391 ,n_628);
  not csa_tree_add_101_22_pad_groupi_g5357(csa_tree_add_101_22_pad_groupi_n_390 ,n_630);
  not csa_tree_add_101_22_pad_groupi_g5358(csa_tree_add_101_22_pad_groupi_n_389 ,n_637);
  not csa_tree_add_101_22_pad_groupi_g5359(csa_tree_add_101_22_pad_groupi_n_388 ,n_636);
  not csa_tree_add_101_22_pad_groupi_g5360(csa_tree_add_101_22_pad_groupi_n_387 ,in21[7]);
  not csa_tree_add_101_22_pad_groupi_g5361(csa_tree_add_101_22_pad_groupi_n_386 ,in9[15]);
  not csa_tree_add_101_22_pad_groupi_g5362(csa_tree_add_101_22_pad_groupi_n_385 ,in9[2]);
  not csa_tree_add_101_22_pad_groupi_g5363(csa_tree_add_101_22_pad_groupi_n_384 ,in9[5]);
  not csa_tree_add_101_22_pad_groupi_g5364(csa_tree_add_101_22_pad_groupi_n_383 ,in9[13]);
  not csa_tree_add_101_22_pad_groupi_g5365(csa_tree_add_101_22_pad_groupi_n_382 ,in9[3]);
  not csa_tree_add_101_22_pad_groupi_g5366(csa_tree_add_101_22_pad_groupi_n_381 ,in9[9]);
  not csa_tree_add_101_22_pad_groupi_g5367(csa_tree_add_101_22_pad_groupi_n_380 ,in9[1]);
  not csa_tree_add_101_22_pad_groupi_g5368(csa_tree_add_101_22_pad_groupi_n_379 ,in9[8]);
  not csa_tree_add_101_22_pad_groupi_g5369(csa_tree_add_101_22_pad_groupi_n_378 ,n_626);
  not csa_tree_add_101_22_pad_groupi_g5370(csa_tree_add_101_22_pad_groupi_n_377 ,n_633);
  not csa_tree_add_101_22_pad_groupi_g5371(csa_tree_add_101_22_pad_groupi_n_376 ,n_634);
  not csa_tree_add_101_22_pad_groupi_g5372(csa_tree_add_101_22_pad_groupi_n_375 ,in22[0]);
  not csa_tree_add_101_22_pad_groupi_g5373(csa_tree_add_101_22_pad_groupi_n_374 ,in21[0]);
  not csa_tree_add_101_22_pad_groupi_g5374(csa_tree_add_101_22_pad_groupi_n_373 ,in21[11]);
  not csa_tree_add_101_22_pad_groupi_g5375(csa_tree_add_101_22_pad_groupi_n_372 ,in21[8]);
  not csa_tree_add_101_22_pad_groupi_g5376(csa_tree_add_101_22_pad_groupi_n_371 ,in21[1]);
  not csa_tree_add_101_22_pad_groupi_g5377(csa_tree_add_101_22_pad_groupi_n_370 ,in21[6]);
  not csa_tree_add_101_22_pad_groupi_g5378(csa_tree_add_101_22_pad_groupi_n_369 ,in21[9]);
  not csa_tree_add_101_22_pad_groupi_g5379(csa_tree_add_101_22_pad_groupi_n_368 ,in9[0]);
  not csa_tree_add_101_22_pad_groupi_g5380(csa_tree_add_101_22_pad_groupi_n_367 ,in9[4]);
  not csa_tree_add_101_22_pad_groupi_g5381(csa_tree_add_101_22_pad_groupi_n_366 ,in9[12]);
  not csa_tree_add_101_22_pad_groupi_g5382(csa_tree_add_101_22_pad_groupi_n_365 ,in9[11]);
  not csa_tree_add_101_22_pad_groupi_g5383(csa_tree_add_101_22_pad_groupi_n_364 ,in9[7]);
  not csa_tree_add_101_22_pad_groupi_g5384(csa_tree_add_101_22_pad_groupi_n_363 ,in9[10]);
  not csa_tree_add_101_22_pad_groupi_g5385(csa_tree_add_101_22_pad_groupi_n_362 ,in9[6]);
  not csa_tree_add_101_22_pad_groupi_g5386(csa_tree_add_101_22_pad_groupi_n_361 ,in9[14]);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5534(csa_tree_add_101_22_pad_groupi_n_345 ,csa_tree_add_101_22_pad_groupi_n_343);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5535(csa_tree_add_101_22_pad_groupi_n_344 ,csa_tree_add_101_22_pad_groupi_n_343);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5536(csa_tree_add_101_22_pad_groupi_n_343 ,csa_tree_add_101_22_pad_groupi_n_356);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5538(csa_tree_add_101_22_pad_groupi_n_342 ,csa_tree_add_101_22_pad_groupi_n_340);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5539(csa_tree_add_101_22_pad_groupi_n_341 ,csa_tree_add_101_22_pad_groupi_n_340);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5540(csa_tree_add_101_22_pad_groupi_n_340 ,csa_tree_add_101_22_pad_groupi_n_422);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5542(csa_tree_add_101_22_pad_groupi_n_339 ,csa_tree_add_101_22_pad_groupi_n_337);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5543(csa_tree_add_101_22_pad_groupi_n_338 ,csa_tree_add_101_22_pad_groupi_n_337);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5544(csa_tree_add_101_22_pad_groupi_n_337 ,csa_tree_add_101_22_pad_groupi_n_413);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5546(csa_tree_add_101_22_pad_groupi_n_336 ,csa_tree_add_101_22_pad_groupi_n_334);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5547(csa_tree_add_101_22_pad_groupi_n_335 ,csa_tree_add_101_22_pad_groupi_n_334);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5548(csa_tree_add_101_22_pad_groupi_n_334 ,csa_tree_add_101_22_pad_groupi_n_348);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5550(csa_tree_add_101_22_pad_groupi_n_333 ,csa_tree_add_101_22_pad_groupi_n_331);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5551(csa_tree_add_101_22_pad_groupi_n_332 ,csa_tree_add_101_22_pad_groupi_n_331);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5552(csa_tree_add_101_22_pad_groupi_n_331 ,csa_tree_add_101_22_pad_groupi_n_411);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5554(csa_tree_add_101_22_pad_groupi_n_330 ,csa_tree_add_101_22_pad_groupi_n_328);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5555(csa_tree_add_101_22_pad_groupi_n_329 ,csa_tree_add_101_22_pad_groupi_n_328);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5556(csa_tree_add_101_22_pad_groupi_n_328 ,csa_tree_add_101_22_pad_groupi_n_410);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5558(csa_tree_add_101_22_pad_groupi_n_327 ,csa_tree_add_101_22_pad_groupi_n_325);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5559(csa_tree_add_101_22_pad_groupi_n_326 ,csa_tree_add_101_22_pad_groupi_n_325);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5560(csa_tree_add_101_22_pad_groupi_n_325 ,csa_tree_add_101_22_pad_groupi_n_350);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5562(csa_tree_add_101_22_pad_groupi_n_324 ,csa_tree_add_101_22_pad_groupi_n_322);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5563(csa_tree_add_101_22_pad_groupi_n_323 ,csa_tree_add_101_22_pad_groupi_n_322);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5564(csa_tree_add_101_22_pad_groupi_n_322 ,csa_tree_add_101_22_pad_groupi_n_419);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5566(csa_tree_add_101_22_pad_groupi_n_321 ,csa_tree_add_101_22_pad_groupi_n_319);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5567(csa_tree_add_101_22_pad_groupi_n_320 ,csa_tree_add_101_22_pad_groupi_n_319);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5568(csa_tree_add_101_22_pad_groupi_n_319 ,csa_tree_add_101_22_pad_groupi_n_416);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5570(csa_tree_add_101_22_pad_groupi_n_318 ,csa_tree_add_101_22_pad_groupi_n_316);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5571(csa_tree_add_101_22_pad_groupi_n_317 ,csa_tree_add_101_22_pad_groupi_n_316);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5572(csa_tree_add_101_22_pad_groupi_n_316 ,csa_tree_add_101_22_pad_groupi_n_351);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5574(csa_tree_add_101_22_pad_groupi_n_315 ,csa_tree_add_101_22_pad_groupi_n_313);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5575(csa_tree_add_101_22_pad_groupi_n_314 ,csa_tree_add_101_22_pad_groupi_n_313);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5576(csa_tree_add_101_22_pad_groupi_n_313 ,csa_tree_add_101_22_pad_groupi_n_415);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5578(csa_tree_add_101_22_pad_groupi_n_312 ,csa_tree_add_101_22_pad_groupi_n_310);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5579(csa_tree_add_101_22_pad_groupi_n_311 ,csa_tree_add_101_22_pad_groupi_n_310);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5580(csa_tree_add_101_22_pad_groupi_n_310 ,csa_tree_add_101_22_pad_groupi_n_423);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5582(csa_tree_add_101_22_pad_groupi_n_309 ,csa_tree_add_101_22_pad_groupi_n_307);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5583(csa_tree_add_101_22_pad_groupi_n_308 ,csa_tree_add_101_22_pad_groupi_n_307);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5584(csa_tree_add_101_22_pad_groupi_n_307 ,csa_tree_add_101_22_pad_groupi_n_414);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5586(csa_tree_add_101_22_pad_groupi_n_306 ,csa_tree_add_101_22_pad_groupi_n_304);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5587(csa_tree_add_101_22_pad_groupi_n_305 ,csa_tree_add_101_22_pad_groupi_n_304);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5588(csa_tree_add_101_22_pad_groupi_n_304 ,csa_tree_add_101_22_pad_groupi_n_353);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5590(csa_tree_add_101_22_pad_groupi_n_303 ,csa_tree_add_101_22_pad_groupi_n_301);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5591(csa_tree_add_101_22_pad_groupi_n_302 ,csa_tree_add_101_22_pad_groupi_n_301);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5592(csa_tree_add_101_22_pad_groupi_n_301 ,csa_tree_add_101_22_pad_groupi_n_418);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5594(csa_tree_add_101_22_pad_groupi_n_300 ,csa_tree_add_101_22_pad_groupi_n_298);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5595(csa_tree_add_101_22_pad_groupi_n_299 ,csa_tree_add_101_22_pad_groupi_n_298);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5596(csa_tree_add_101_22_pad_groupi_n_298 ,csa_tree_add_101_22_pad_groupi_n_397);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5598(csa_tree_add_101_22_pad_groupi_n_297 ,csa_tree_add_101_22_pad_groupi_n_295);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5599(csa_tree_add_101_22_pad_groupi_n_296 ,csa_tree_add_101_22_pad_groupi_n_295);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5600(csa_tree_add_101_22_pad_groupi_n_295 ,csa_tree_add_101_22_pad_groupi_n_346);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5602(csa_tree_add_101_22_pad_groupi_n_294 ,csa_tree_add_101_22_pad_groupi_n_292);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5603(csa_tree_add_101_22_pad_groupi_n_293 ,csa_tree_add_101_22_pad_groupi_n_292);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5604(csa_tree_add_101_22_pad_groupi_n_292 ,csa_tree_add_101_22_pad_groupi_n_398);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5606(csa_tree_add_101_22_pad_groupi_n_291 ,csa_tree_add_101_22_pad_groupi_n_289);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5607(csa_tree_add_101_22_pad_groupi_n_290 ,csa_tree_add_101_22_pad_groupi_n_289);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5608(csa_tree_add_101_22_pad_groupi_n_289 ,csa_tree_add_101_22_pad_groupi_n_397);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5610(csa_tree_add_101_22_pad_groupi_n_288 ,csa_tree_add_101_22_pad_groupi_n_286);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5611(csa_tree_add_101_22_pad_groupi_n_287 ,csa_tree_add_101_22_pad_groupi_n_286);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5612(csa_tree_add_101_22_pad_groupi_n_286 ,csa_tree_add_101_22_pad_groupi_n_509);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5614(csa_tree_add_101_22_pad_groupi_n_285 ,csa_tree_add_101_22_pad_groupi_n_283);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5615(csa_tree_add_101_22_pad_groupi_n_284 ,csa_tree_add_101_22_pad_groupi_n_283);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5616(csa_tree_add_101_22_pad_groupi_n_283 ,csa_tree_add_101_22_pad_groupi_n_503);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5620(csa_tree_add_101_22_pad_groupi_n_358 ,csa_tree_add_101_22_pad_groupi_n_581);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5623(csa_tree_add_101_22_pad_groupi_n_282 ,csa_tree_add_101_22_pad_groupi_n_281);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5624(csa_tree_add_101_22_pad_groupi_n_281 ,csa_tree_add_101_22_pad_groupi_n_579);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5627(csa_tree_add_101_22_pad_groupi_n_280 ,csa_tree_add_101_22_pad_groupi_n_279);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5628(csa_tree_add_101_22_pad_groupi_n_279 ,csa_tree_add_101_22_pad_groupi_n_582);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5632(csa_tree_add_101_22_pad_groupi_n_357 ,csa_tree_add_101_22_pad_groupi_n_580);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5635(csa_tree_add_101_22_pad_groupi_n_278 ,csa_tree_add_101_22_pad_groupi_n_277);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5636(csa_tree_add_101_22_pad_groupi_n_277 ,csa_tree_add_101_22_pad_groupi_n_497);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5639(csa_tree_add_101_22_pad_groupi_n_276 ,csa_tree_add_101_22_pad_groupi_n_359);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5640(csa_tree_add_101_22_pad_groupi_n_359 ,csa_tree_add_101_22_pad_groupi_n_934);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5642(csa_tree_add_101_22_pad_groupi_n_275 ,csa_tree_add_101_22_pad_groupi_n_273);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5643(csa_tree_add_101_22_pad_groupi_n_274 ,csa_tree_add_101_22_pad_groupi_n_273);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5644(csa_tree_add_101_22_pad_groupi_n_273 ,csa_tree_add_101_22_pad_groupi_n_355);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5646(csa_tree_add_101_22_pad_groupi_n_272 ,csa_tree_add_101_22_pad_groupi_n_270);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5647(csa_tree_add_101_22_pad_groupi_n_271 ,csa_tree_add_101_22_pad_groupi_n_270);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5648(csa_tree_add_101_22_pad_groupi_n_270 ,csa_tree_add_101_22_pad_groupi_n_349);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5650(csa_tree_add_101_22_pad_groupi_n_269 ,csa_tree_add_101_22_pad_groupi_n_267);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5651(csa_tree_add_101_22_pad_groupi_n_268 ,csa_tree_add_101_22_pad_groupi_n_267);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5652(csa_tree_add_101_22_pad_groupi_n_267 ,csa_tree_add_101_22_pad_groupi_n_347);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5654(csa_tree_add_101_22_pad_groupi_n_266 ,csa_tree_add_101_22_pad_groupi_n_264);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5655(csa_tree_add_101_22_pad_groupi_n_265 ,csa_tree_add_101_22_pad_groupi_n_264);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5656(csa_tree_add_101_22_pad_groupi_n_264 ,csa_tree_add_101_22_pad_groupi_n_354);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5658(csa_tree_add_101_22_pad_groupi_n_263 ,csa_tree_add_101_22_pad_groupi_n_261);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5659(csa_tree_add_101_22_pad_groupi_n_262 ,csa_tree_add_101_22_pad_groupi_n_261);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5660(csa_tree_add_101_22_pad_groupi_n_261 ,csa_tree_add_101_22_pad_groupi_n_352);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5662(csa_tree_add_101_22_pad_groupi_n_260 ,csa_tree_add_101_22_pad_groupi_n_259);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5664(csa_tree_add_101_22_pad_groupi_n_259 ,csa_tree_add_101_22_pad_groupi_n_399);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5686(csa_tree_add_101_22_pad_groupi_n_258 ,csa_tree_add_101_22_pad_groupi_n_346);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5688(csa_tree_add_101_22_pad_groupi_n_346 ,csa_tree_add_101_22_pad_groupi_n_398);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5690(csa_tree_add_101_22_pad_groupi_n_257 ,csa_tree_add_101_22_pad_groupi_n_256);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5692(csa_tree_add_101_22_pad_groupi_n_256 ,csa_tree_add_101_22_pad_groupi_n_507);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5694(csa_tree_add_101_22_pad_groupi_n_255 ,csa_tree_add_101_22_pad_groupi_n_254);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5696(csa_tree_add_101_22_pad_groupi_n_254 ,csa_tree_add_101_22_pad_groupi_n_501);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5709(csa_tree_add_101_22_pad_groupi_n_253 ,csa_tree_add_101_22_pad_groupi_n_251);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5710(csa_tree_add_101_22_pad_groupi_n_252 ,csa_tree_add_101_22_pad_groupi_n_251);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5711(csa_tree_add_101_22_pad_groupi_n_251 ,csa_tree_add_101_22_pad_groupi_n_511);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5713(csa_tree_add_101_22_pad_groupi_n_250 ,csa_tree_add_101_22_pad_groupi_n_248);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5714(csa_tree_add_101_22_pad_groupi_n_249 ,csa_tree_add_101_22_pad_groupi_n_248);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5715(csa_tree_add_101_22_pad_groupi_n_248 ,csa_tree_add_101_22_pad_groupi_n_401);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5721(csa_tree_add_101_22_pad_groupi_n_247 ,csa_tree_add_101_22_pad_groupi_n_245);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5722(csa_tree_add_101_22_pad_groupi_n_246 ,csa_tree_add_101_22_pad_groupi_n_245);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5723(csa_tree_add_101_22_pad_groupi_n_245 ,csa_tree_add_101_22_pad_groupi_n_385);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5733(csa_tree_add_101_22_pad_groupi_n_244 ,csa_tree_add_101_22_pad_groupi_n_242);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5734(csa_tree_add_101_22_pad_groupi_n_243 ,csa_tree_add_101_22_pad_groupi_n_242);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5735(csa_tree_add_101_22_pad_groupi_n_242 ,csa_tree_add_101_22_pad_groupi_n_368);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5737(csa_tree_add_101_22_pad_groupi_n_241 ,csa_tree_add_101_22_pad_groupi_n_239);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5738(csa_tree_add_101_22_pad_groupi_n_240 ,csa_tree_add_101_22_pad_groupi_n_239);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5739(csa_tree_add_101_22_pad_groupi_n_239 ,csa_tree_add_101_22_pad_groupi_n_396);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5741(csa_tree_add_101_22_pad_groupi_n_238 ,csa_tree_add_101_22_pad_groupi_n_236);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5742(csa_tree_add_101_22_pad_groupi_n_237 ,csa_tree_add_101_22_pad_groupi_n_236);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5743(csa_tree_add_101_22_pad_groupi_n_236 ,csa_tree_add_101_22_pad_groupi_n_396);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5746(csa_tree_add_101_22_pad_groupi_n_235 ,csa_tree_add_101_22_pad_groupi_n_234);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5747(csa_tree_add_101_22_pad_groupi_n_234 ,csa_tree_add_101_22_pad_groupi_n_381);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5750(csa_tree_add_101_22_pad_groupi_n_233 ,csa_tree_add_101_22_pad_groupi_n_232);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5751(csa_tree_add_101_22_pad_groupi_n_232 ,csa_tree_add_101_22_pad_groupi_n_366);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5754(csa_tree_add_101_22_pad_groupi_n_231 ,csa_tree_add_101_22_pad_groupi_n_230);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5755(csa_tree_add_101_22_pad_groupi_n_230 ,csa_tree_add_101_22_pad_groupi_n_382);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5758(csa_tree_add_101_22_pad_groupi_n_229 ,csa_tree_add_101_22_pad_groupi_n_228);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5759(csa_tree_add_101_22_pad_groupi_n_228 ,csa_tree_add_101_22_pad_groupi_n_383);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5762(csa_tree_add_101_22_pad_groupi_n_227 ,csa_tree_add_101_22_pad_groupi_n_226);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5763(csa_tree_add_101_22_pad_groupi_n_226 ,csa_tree_add_101_22_pad_groupi_n_365);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5766(csa_tree_add_101_22_pad_groupi_n_225 ,csa_tree_add_101_22_pad_groupi_n_224);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5767(csa_tree_add_101_22_pad_groupi_n_224 ,csa_tree_add_101_22_pad_groupi_n_363);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5769(csa_tree_add_101_22_pad_groupi_n_223 ,csa_tree_add_101_22_pad_groupi_n_221);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5770(csa_tree_add_101_22_pad_groupi_n_222 ,csa_tree_add_101_22_pad_groupi_n_221);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5771(csa_tree_add_101_22_pad_groupi_n_221 ,csa_tree_add_101_22_pad_groupi_n_366);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5774(csa_tree_add_101_22_pad_groupi_n_220 ,csa_tree_add_101_22_pad_groupi_n_219);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5775(csa_tree_add_101_22_pad_groupi_n_219 ,csa_tree_add_101_22_pad_groupi_n_362);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5777(csa_tree_add_101_22_pad_groupi_n_218 ,csa_tree_add_101_22_pad_groupi_n_216);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5778(csa_tree_add_101_22_pad_groupi_n_217 ,csa_tree_add_101_22_pad_groupi_n_216);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5779(csa_tree_add_101_22_pad_groupi_n_216 ,csa_tree_add_101_22_pad_groupi_n_380);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5781(csa_tree_add_101_22_pad_groupi_n_215 ,csa_tree_add_101_22_pad_groupi_n_213);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5782(csa_tree_add_101_22_pad_groupi_n_214 ,csa_tree_add_101_22_pad_groupi_n_213);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5783(csa_tree_add_101_22_pad_groupi_n_213 ,csa_tree_add_101_22_pad_groupi_n_381);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5785(csa_tree_add_101_22_pad_groupi_n_212 ,csa_tree_add_101_22_pad_groupi_n_210);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5786(csa_tree_add_101_22_pad_groupi_n_211 ,csa_tree_add_101_22_pad_groupi_n_210);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5787(csa_tree_add_101_22_pad_groupi_n_210 ,csa_tree_add_101_22_pad_groupi_n_362);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5790(csa_tree_add_101_22_pad_groupi_n_209 ,csa_tree_add_101_22_pad_groupi_n_208);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5791(csa_tree_add_101_22_pad_groupi_n_208 ,csa_tree_add_101_22_pad_groupi_n_379);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5793(csa_tree_add_101_22_pad_groupi_n_207 ,csa_tree_add_101_22_pad_groupi_n_205);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5794(csa_tree_add_101_22_pad_groupi_n_206 ,csa_tree_add_101_22_pad_groupi_n_205);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5795(csa_tree_add_101_22_pad_groupi_n_205 ,csa_tree_add_101_22_pad_groupi_n_379);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5798(csa_tree_add_101_22_pad_groupi_n_204 ,csa_tree_add_101_22_pad_groupi_n_203);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5799(csa_tree_add_101_22_pad_groupi_n_203 ,csa_tree_add_101_22_pad_groupi_n_384);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5801(csa_tree_add_101_22_pad_groupi_n_202 ,csa_tree_add_101_22_pad_groupi_n_200);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5802(csa_tree_add_101_22_pad_groupi_n_201 ,csa_tree_add_101_22_pad_groupi_n_200);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5803(csa_tree_add_101_22_pad_groupi_n_200 ,csa_tree_add_101_22_pad_groupi_n_382);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5807(csa_tree_add_101_22_pad_groupi_n_198 ,csa_tree_add_101_22_pad_groupi_n_361);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5809(csa_tree_add_101_22_pad_groupi_n_197 ,csa_tree_add_101_22_pad_groupi_n_195);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5810(csa_tree_add_101_22_pad_groupi_n_196 ,csa_tree_add_101_22_pad_groupi_n_195);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5811(csa_tree_add_101_22_pad_groupi_n_195 ,csa_tree_add_101_22_pad_groupi_n_384);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5813(csa_tree_add_101_22_pad_groupi_n_194 ,csa_tree_add_101_22_pad_groupi_n_192);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5814(csa_tree_add_101_22_pad_groupi_n_193 ,csa_tree_add_101_22_pad_groupi_n_192);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5815(csa_tree_add_101_22_pad_groupi_n_192 ,csa_tree_add_101_22_pad_groupi_n_361);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5817(csa_tree_add_101_22_pad_groupi_n_191 ,csa_tree_add_101_22_pad_groupi_n_190);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5819(csa_tree_add_101_22_pad_groupi_n_190 ,csa_tree_add_101_22_pad_groupi_n_364);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5822(csa_tree_add_101_22_pad_groupi_n_189 ,csa_tree_add_101_22_pad_groupi_n_188);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5823(csa_tree_add_101_22_pad_groupi_n_188 ,csa_tree_add_101_22_pad_groupi_n_367);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5825(csa_tree_add_101_22_pad_groupi_n_187 ,csa_tree_add_101_22_pad_groupi_n_185);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5826(csa_tree_add_101_22_pad_groupi_n_186 ,csa_tree_add_101_22_pad_groupi_n_185);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5827(csa_tree_add_101_22_pad_groupi_n_185 ,csa_tree_add_101_22_pad_groupi_n_383);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5829(csa_tree_add_101_22_pad_groupi_n_184 ,csa_tree_add_101_22_pad_groupi_n_182);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5830(csa_tree_add_101_22_pad_groupi_n_183 ,csa_tree_add_101_22_pad_groupi_n_182);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5831(csa_tree_add_101_22_pad_groupi_n_182 ,csa_tree_add_101_22_pad_groupi_n_364);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5833(csa_tree_add_101_22_pad_groupi_n_181 ,csa_tree_add_101_22_pad_groupi_n_179);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5834(csa_tree_add_101_22_pad_groupi_n_180 ,csa_tree_add_101_22_pad_groupi_n_179);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5835(csa_tree_add_101_22_pad_groupi_n_179 ,csa_tree_add_101_22_pad_groupi_n_365);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5837(csa_tree_add_101_22_pad_groupi_n_178 ,csa_tree_add_101_22_pad_groupi_n_176);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5838(csa_tree_add_101_22_pad_groupi_n_177 ,csa_tree_add_101_22_pad_groupi_n_176);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5839(csa_tree_add_101_22_pad_groupi_n_176 ,csa_tree_add_101_22_pad_groupi_n_363);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5841(csa_tree_add_101_22_pad_groupi_n_175 ,csa_tree_add_101_22_pad_groupi_n_173);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5842(csa_tree_add_101_22_pad_groupi_n_174 ,csa_tree_add_101_22_pad_groupi_n_173);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5843(csa_tree_add_101_22_pad_groupi_n_173 ,csa_tree_add_101_22_pad_groupi_n_367);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5845(csa_tree_add_101_22_pad_groupi_n_172 ,csa_tree_add_101_22_pad_groupi_n_170);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5846(csa_tree_add_101_22_pad_groupi_n_171 ,csa_tree_add_101_22_pad_groupi_n_170);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5847(csa_tree_add_101_22_pad_groupi_n_170 ,csa_tree_add_101_22_pad_groupi_n_495);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5849(csa_tree_add_101_22_pad_groupi_n_169 ,csa_tree_add_101_22_pad_groupi_n_167);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5850(csa_tree_add_101_22_pad_groupi_n_168 ,csa_tree_add_101_22_pad_groupi_n_167);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5851(csa_tree_add_101_22_pad_groupi_n_167 ,csa_tree_add_101_22_pad_groupi_n_495);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5853(csa_tree_add_101_22_pad_groupi_n_166 ,csa_tree_add_101_22_pad_groupi_n_164);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5854(csa_tree_add_101_22_pad_groupi_n_165 ,csa_tree_add_101_22_pad_groupi_n_164);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5855(csa_tree_add_101_22_pad_groupi_n_164 ,csa_tree_add_101_22_pad_groupi_n_498);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5857(csa_tree_add_101_22_pad_groupi_n_163 ,csa_tree_add_101_22_pad_groupi_n_161);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5858(csa_tree_add_101_22_pad_groupi_n_162 ,csa_tree_add_101_22_pad_groupi_n_161);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5859(csa_tree_add_101_22_pad_groupi_n_161 ,csa_tree_add_101_22_pad_groupi_n_386);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5861(csa_tree_add_101_22_pad_groupi_n_160 ,csa_tree_add_101_22_pad_groupi_n_350);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5863(csa_tree_add_101_22_pad_groupi_n_350 ,csa_tree_add_101_22_pad_groupi_n_412);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5865(csa_tree_add_101_22_pad_groupi_n_159 ,csa_tree_add_101_22_pad_groupi_n_348);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5867(csa_tree_add_101_22_pad_groupi_n_348 ,csa_tree_add_101_22_pad_groupi_n_409);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5869(csa_tree_add_101_22_pad_groupi_n_158 ,csa_tree_add_101_22_pad_groupi_n_356);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5871(csa_tree_add_101_22_pad_groupi_n_356 ,csa_tree_add_101_22_pad_groupi_n_421);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5877(csa_tree_add_101_22_pad_groupi_n_155 ,csa_tree_add_101_22_pad_groupi_n_355);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5879(csa_tree_add_101_22_pad_groupi_n_355 ,csa_tree_add_101_22_pad_groupi_n_421);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5881(csa_tree_add_101_22_pad_groupi_n_154 ,csa_tree_add_101_22_pad_groupi_n_353);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5883(csa_tree_add_101_22_pad_groupi_n_353 ,csa_tree_add_101_22_pad_groupi_n_420);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5885(csa_tree_add_101_22_pad_groupi_n_153 ,csa_tree_add_101_22_pad_groupi_n_349);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5887(csa_tree_add_101_22_pad_groupi_n_349 ,csa_tree_add_101_22_pad_groupi_n_412);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5889(csa_tree_add_101_22_pad_groupi_n_152 ,csa_tree_add_101_22_pad_groupi_n_351);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5891(csa_tree_add_101_22_pad_groupi_n_351 ,csa_tree_add_101_22_pad_groupi_n_417);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5893(csa_tree_add_101_22_pad_groupi_n_151 ,csa_tree_add_101_22_pad_groupi_n_352);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5895(csa_tree_add_101_22_pad_groupi_n_352 ,csa_tree_add_101_22_pad_groupi_n_417);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5897(csa_tree_add_101_22_pad_groupi_n_150 ,csa_tree_add_101_22_pad_groupi_n_347);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5899(csa_tree_add_101_22_pad_groupi_n_347 ,csa_tree_add_101_22_pad_groupi_n_409);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5901(csa_tree_add_101_22_pad_groupi_n_149 ,csa_tree_add_101_22_pad_groupi_n_354);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5903(csa_tree_add_101_22_pad_groupi_n_354 ,csa_tree_add_101_22_pad_groupi_n_420);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5905(csa_tree_add_101_22_pad_groupi_n_148 ,csa_tree_add_101_22_pad_groupi_n_146);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5906(csa_tree_add_101_22_pad_groupi_n_147 ,csa_tree_add_101_22_pad_groupi_n_146);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5907(csa_tree_add_101_22_pad_groupi_n_146 ,csa_tree_add_101_22_pad_groupi_n_504);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5909(csa_tree_add_101_22_pad_groupi_n_145 ,csa_tree_add_101_22_pad_groupi_n_143);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5910(csa_tree_add_101_22_pad_groupi_n_144 ,csa_tree_add_101_22_pad_groupi_n_143);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5911(csa_tree_add_101_22_pad_groupi_n_143 ,csa_tree_add_101_22_pad_groupi_n_510);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5913(csa_tree_add_101_22_pad_groupi_n_142 ,csa_tree_add_101_22_pad_groupi_n_140);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5914(csa_tree_add_101_22_pad_groupi_n_141 ,csa_tree_add_101_22_pad_groupi_n_140);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5915(csa_tree_add_101_22_pad_groupi_n_140 ,csa_tree_add_101_22_pad_groupi_n_510);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5917(csa_tree_add_101_22_pad_groupi_n_139 ,csa_tree_add_101_22_pad_groupi_n_137);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5918(csa_tree_add_101_22_pad_groupi_n_138 ,csa_tree_add_101_22_pad_groupi_n_137);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5919(csa_tree_add_101_22_pad_groupi_n_137 ,csa_tree_add_101_22_pad_groupi_n_494);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5921(csa_tree_add_101_22_pad_groupi_n_136 ,csa_tree_add_101_22_pad_groupi_n_134);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5922(csa_tree_add_101_22_pad_groupi_n_135 ,csa_tree_add_101_22_pad_groupi_n_134);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5923(csa_tree_add_101_22_pad_groupi_n_134 ,csa_tree_add_101_22_pad_groupi_n_494);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5925(csa_tree_add_101_22_pad_groupi_n_133 ,csa_tree_add_101_22_pad_groupi_n_131);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5926(csa_tree_add_101_22_pad_groupi_n_132 ,csa_tree_add_101_22_pad_groupi_n_131);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5927(csa_tree_add_101_22_pad_groupi_n_131 ,csa_tree_add_101_22_pad_groupi_n_504);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5929(csa_tree_add_101_22_pad_groupi_n_130 ,csa_tree_add_101_22_pad_groupi_n_128);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5930(csa_tree_add_101_22_pad_groupi_n_129 ,csa_tree_add_101_22_pad_groupi_n_128);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5931(csa_tree_add_101_22_pad_groupi_n_128 ,csa_tree_add_101_22_pad_groupi_n_498);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5933(csa_tree_add_101_22_pad_groupi_n_127 ,csa_tree_add_101_22_pad_groupi_n_125);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5934(csa_tree_add_101_22_pad_groupi_n_126 ,csa_tree_add_101_22_pad_groupi_n_125);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5935(csa_tree_add_101_22_pad_groupi_n_125 ,csa_tree_add_101_22_pad_groupi_n_496);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5937(csa_tree_add_101_22_pad_groupi_n_124 ,csa_tree_add_101_22_pad_groupi_n_122);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5938(csa_tree_add_101_22_pad_groupi_n_123 ,csa_tree_add_101_22_pad_groupi_n_122);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5939(csa_tree_add_101_22_pad_groupi_n_122 ,csa_tree_add_101_22_pad_groupi_n_496);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5941(csa_tree_add_101_22_pad_groupi_n_121 ,csa_tree_add_101_22_pad_groupi_n_120);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5943(csa_tree_add_101_22_pad_groupi_n_120 ,csa_tree_add_101_22_pad_groupi_n_386);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5945(csa_tree_add_101_22_pad_groupi_n_119 ,csa_tree_add_101_22_pad_groupi_n_117);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5946(csa_tree_add_101_22_pad_groupi_n_118 ,csa_tree_add_101_22_pad_groupi_n_117);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5947(csa_tree_add_101_22_pad_groupi_n_117 ,csa_tree_add_101_22_pad_groupi_n_511);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5949(csa_tree_add_101_22_pad_groupi_n_116 ,csa_tree_add_101_22_pad_groupi_n_114);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5950(csa_tree_add_101_22_pad_groupi_n_115 ,csa_tree_add_101_22_pad_groupi_n_114);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5951(csa_tree_add_101_22_pad_groupi_n_114 ,csa_tree_add_101_22_pad_groupi_n_511);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5953(csa_tree_add_101_22_pad_groupi_n_113 ,csa_tree_add_101_22_pad_groupi_n_111);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5954(csa_tree_add_101_22_pad_groupi_n_112 ,csa_tree_add_101_22_pad_groupi_n_111);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5955(csa_tree_add_101_22_pad_groupi_n_111 ,csa_tree_add_101_22_pad_groupi_n_253);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5957(csa_tree_add_101_22_pad_groupi_n_110 ,csa_tree_add_101_22_pad_groupi_n_108);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5958(csa_tree_add_101_22_pad_groupi_n_109 ,csa_tree_add_101_22_pad_groupi_n_108);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5959(csa_tree_add_101_22_pad_groupi_n_108 ,csa_tree_add_101_22_pad_groupi_n_401);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5961(csa_tree_add_101_22_pad_groupi_n_107 ,csa_tree_add_101_22_pad_groupi_n_105);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5962(csa_tree_add_101_22_pad_groupi_n_106 ,csa_tree_add_101_22_pad_groupi_n_105);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5963(csa_tree_add_101_22_pad_groupi_n_105 ,csa_tree_add_101_22_pad_groupi_n_401);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5965(csa_tree_add_101_22_pad_groupi_n_104 ,csa_tree_add_101_22_pad_groupi_n_102);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5966(csa_tree_add_101_22_pad_groupi_n_103 ,csa_tree_add_101_22_pad_groupi_n_102);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5967(csa_tree_add_101_22_pad_groupi_n_102 ,csa_tree_add_101_22_pad_groupi_n_250);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5969(csa_tree_add_101_22_pad_groupi_n_101 ,csa_tree_add_101_22_pad_groupi_n_99);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5970(csa_tree_add_101_22_pad_groupi_n_100 ,csa_tree_add_101_22_pad_groupi_n_99);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5971(csa_tree_add_101_22_pad_groupi_n_99 ,csa_tree_add_101_22_pad_groupi_n_385);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5973(csa_tree_add_101_22_pad_groupi_n_98 ,csa_tree_add_101_22_pad_groupi_n_97);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5975(csa_tree_add_101_22_pad_groupi_n_97 ,csa_tree_add_101_22_pad_groupi_n_247);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5977(csa_tree_add_101_22_pad_groupi_n_96 ,csa_tree_add_101_22_pad_groupi_n_94);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5978(csa_tree_add_101_22_pad_groupi_n_95 ,csa_tree_add_101_22_pad_groupi_n_94);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5979(csa_tree_add_101_22_pad_groupi_n_94 ,csa_tree_add_101_22_pad_groupi_n_381);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5981(csa_tree_add_101_22_pad_groupi_n_93 ,csa_tree_add_101_22_pad_groupi_n_92);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5983(csa_tree_add_101_22_pad_groupi_n_92 ,csa_tree_add_101_22_pad_groupi_n_252);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5985(csa_tree_add_101_22_pad_groupi_n_91 ,csa_tree_add_101_22_pad_groupi_n_89);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5986(csa_tree_add_101_22_pad_groupi_n_90 ,csa_tree_add_101_22_pad_groupi_n_89);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5987(csa_tree_add_101_22_pad_groupi_n_89 ,csa_tree_add_101_22_pad_groupi_n_366);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5989(csa_tree_add_101_22_pad_groupi_n_88 ,csa_tree_add_101_22_pad_groupi_n_86);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5990(csa_tree_add_101_22_pad_groupi_n_87 ,csa_tree_add_101_22_pad_groupi_n_86);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5991(csa_tree_add_101_22_pad_groupi_n_86 ,csa_tree_add_101_22_pad_groupi_n_382);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5993(csa_tree_add_101_22_pad_groupi_n_85 ,csa_tree_add_101_22_pad_groupi_n_83);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5994(csa_tree_add_101_22_pad_groupi_n_84 ,csa_tree_add_101_22_pad_groupi_n_83);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5995(csa_tree_add_101_22_pad_groupi_n_83 ,csa_tree_add_101_22_pad_groupi_n_383);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5997(csa_tree_add_101_22_pad_groupi_n_82 ,csa_tree_add_101_22_pad_groupi_n_80);
  not csa_tree_add_101_22_pad_groupi_drc_bufs5999(csa_tree_add_101_22_pad_groupi_n_80 ,csa_tree_add_101_22_pad_groupi_n_365);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6001(csa_tree_add_101_22_pad_groupi_n_79 ,csa_tree_add_101_22_pad_groupi_n_77);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6002(csa_tree_add_101_22_pad_groupi_n_78 ,csa_tree_add_101_22_pad_groupi_n_77);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6003(csa_tree_add_101_22_pad_groupi_n_77 ,csa_tree_add_101_22_pad_groupi_n_363);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6005(csa_tree_add_101_22_pad_groupi_n_76 ,csa_tree_add_101_22_pad_groupi_n_75);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6007(csa_tree_add_101_22_pad_groupi_n_75 ,csa_tree_add_101_22_pad_groupi_n_215);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6009(csa_tree_add_101_22_pad_groupi_n_74 ,csa_tree_add_101_22_pad_groupi_n_72);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6010(csa_tree_add_101_22_pad_groupi_n_73 ,csa_tree_add_101_22_pad_groupi_n_72);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6011(csa_tree_add_101_22_pad_groupi_n_72 ,csa_tree_add_101_22_pad_groupi_n_385);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6013(csa_tree_add_101_22_pad_groupi_n_71 ,csa_tree_add_101_22_pad_groupi_n_70);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6015(csa_tree_add_101_22_pad_groupi_n_70 ,csa_tree_add_101_22_pad_groupi_n_218);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6017(csa_tree_add_101_22_pad_groupi_n_69 ,csa_tree_add_101_22_pad_groupi_n_68);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6019(csa_tree_add_101_22_pad_groupi_n_68 ,csa_tree_add_101_22_pad_groupi_n_223);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6021(csa_tree_add_101_22_pad_groupi_n_67 ,csa_tree_add_101_22_pad_groupi_n_65);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6022(csa_tree_add_101_22_pad_groupi_n_66 ,csa_tree_add_101_22_pad_groupi_n_65);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6023(csa_tree_add_101_22_pad_groupi_n_65 ,csa_tree_add_101_22_pad_groupi_n_362);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6025(csa_tree_add_101_22_pad_groupi_n_64 ,csa_tree_add_101_22_pad_groupi_n_62);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6027(csa_tree_add_101_22_pad_groupi_n_62 ,csa_tree_add_101_22_pad_groupi_n_380);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6029(csa_tree_add_101_22_pad_groupi_n_61 ,csa_tree_add_101_22_pad_groupi_n_60);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6031(csa_tree_add_101_22_pad_groupi_n_60 ,csa_tree_add_101_22_pad_groupi_n_249);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6033(csa_tree_add_101_22_pad_groupi_n_59 ,csa_tree_add_101_22_pad_groupi_n_58);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6035(csa_tree_add_101_22_pad_groupi_n_58 ,csa_tree_add_101_22_pad_groupi_n_212);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6037(csa_tree_add_101_22_pad_groupi_n_57 ,csa_tree_add_101_22_pad_groupi_n_56);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6039(csa_tree_add_101_22_pad_groupi_n_56 ,csa_tree_add_101_22_pad_groupi_n_244);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6041(csa_tree_add_101_22_pad_groupi_n_55 ,csa_tree_add_101_22_pad_groupi_n_54);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6043(csa_tree_add_101_22_pad_groupi_n_54 ,csa_tree_add_101_22_pad_groupi_n_207);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6045(csa_tree_add_101_22_pad_groupi_n_53 ,csa_tree_add_101_22_pad_groupi_n_51);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6046(csa_tree_add_101_22_pad_groupi_n_52 ,csa_tree_add_101_22_pad_groupi_n_51);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6047(csa_tree_add_101_22_pad_groupi_n_51 ,csa_tree_add_101_22_pad_groupi_n_384);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6049(csa_tree_add_101_22_pad_groupi_n_50 ,csa_tree_add_101_22_pad_groupi_n_48);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6051(csa_tree_add_101_22_pad_groupi_n_48 ,csa_tree_add_101_22_pad_groupi_n_379);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6053(csa_tree_add_101_22_pad_groupi_n_47 ,csa_tree_add_101_22_pad_groupi_n_46);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6055(csa_tree_add_101_22_pad_groupi_n_46 ,csa_tree_add_101_22_pad_groupi_n_246);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6057(csa_tree_add_101_22_pad_groupi_n_45 ,csa_tree_add_101_22_pad_groupi_n_43);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6059(csa_tree_add_101_22_pad_groupi_n_43 ,csa_tree_add_101_22_pad_groupi_n_380);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6061(csa_tree_add_101_22_pad_groupi_n_42 ,csa_tree_add_101_22_pad_groupi_n_40);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6062(csa_tree_add_101_22_pad_groupi_n_41 ,csa_tree_add_101_22_pad_groupi_n_40);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6063(csa_tree_add_101_22_pad_groupi_n_40 ,csa_tree_add_101_22_pad_groupi_n_368);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6065(csa_tree_add_101_22_pad_groupi_n_39 ,csa_tree_add_101_22_pad_groupi_n_37);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6066(csa_tree_add_101_22_pad_groupi_n_38 ,csa_tree_add_101_22_pad_groupi_n_37);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6067(csa_tree_add_101_22_pad_groupi_n_37 ,csa_tree_add_101_22_pad_groupi_n_361);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6069(csa_tree_add_101_22_pad_groupi_n_36 ,csa_tree_add_101_22_pad_groupi_n_35);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6071(csa_tree_add_101_22_pad_groupi_n_35 ,csa_tree_add_101_22_pad_groupi_n_202);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6073(csa_tree_add_101_22_pad_groupi_n_34 ,csa_tree_add_101_22_pad_groupi_n_33);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6075(csa_tree_add_101_22_pad_groupi_n_33 ,csa_tree_add_101_22_pad_groupi_n_238);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6077(csa_tree_add_101_22_pad_groupi_n_32 ,csa_tree_add_101_22_pad_groupi_n_31);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6079(csa_tree_add_101_22_pad_groupi_n_31 ,csa_tree_add_101_22_pad_groupi_n_241);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6082(csa_tree_add_101_22_pad_groupi_n_30 ,csa_tree_add_101_22_pad_groupi_n_29);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6083(csa_tree_add_101_22_pad_groupi_n_29 ,csa_tree_add_101_22_pad_groupi_n_193);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6085(csa_tree_add_101_22_pad_groupi_n_28 ,csa_tree_add_101_22_pad_groupi_n_26);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6086(csa_tree_add_101_22_pad_groupi_n_27 ,csa_tree_add_101_22_pad_groupi_n_26);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6087(csa_tree_add_101_22_pad_groupi_n_26 ,csa_tree_add_101_22_pad_groupi_n_367);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6089(csa_tree_add_101_22_pad_groupi_n_25 ,csa_tree_add_101_22_pad_groupi_n_23);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6090(csa_tree_add_101_22_pad_groupi_n_24 ,csa_tree_add_101_22_pad_groupi_n_23);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6091(csa_tree_add_101_22_pad_groupi_n_23 ,csa_tree_add_101_22_pad_groupi_n_368);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6093(csa_tree_add_101_22_pad_groupi_n_22 ,csa_tree_add_101_22_pad_groupi_n_20);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6094(csa_tree_add_101_22_pad_groupi_n_21 ,csa_tree_add_101_22_pad_groupi_n_20);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6095(csa_tree_add_101_22_pad_groupi_n_20 ,csa_tree_add_101_22_pad_groupi_n_364);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6098(csa_tree_add_101_22_pad_groupi_n_19 ,csa_tree_add_101_22_pad_groupi_n_18);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6099(csa_tree_add_101_22_pad_groupi_n_18 ,csa_tree_add_101_22_pad_groupi_n_243);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6102(csa_tree_add_101_22_pad_groupi_n_17 ,csa_tree_add_101_22_pad_groupi_n_16);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6103(csa_tree_add_101_22_pad_groupi_n_16 ,csa_tree_add_101_22_pad_groupi_n_196);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6106(csa_tree_add_101_22_pad_groupi_n_15 ,csa_tree_add_101_22_pad_groupi_n_14);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6107(csa_tree_add_101_22_pad_groupi_n_14 ,csa_tree_add_101_22_pad_groupi_n_237);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6110(csa_tree_add_101_22_pad_groupi_n_13 ,csa_tree_add_101_22_pad_groupi_n_12);
  not csa_tree_add_101_22_pad_groupi_drc_bufs6111(csa_tree_add_101_22_pad_groupi_n_12 ,csa_tree_add_101_22_pad_groupi_n_240);
  xor csa_tree_add_101_22_pad_groupi_g2(n_231 ,csa_tree_add_101_22_pad_groupi_n_1537 ,csa_tree_add_101_22_pad_groupi_n_1520);
  xor csa_tree_add_101_22_pad_groupi_g6113(n_229 ,csa_tree_add_101_22_pad_groupi_n_1532 ,csa_tree_add_101_22_pad_groupi_n_1518);
  xor csa_tree_add_101_22_pad_groupi_g6114(n_226 ,csa_tree_add_101_22_pad_groupi_n_1524 ,csa_tree_add_101_22_pad_groupi_n_1482);
  xor csa_tree_add_101_22_pad_groupi_g6115(n_225 ,csa_tree_add_101_22_pad_groupi_n_1522 ,csa_tree_add_101_22_pad_groupi_n_1502);
  xor csa_tree_add_101_22_pad_groupi_g6116(n_224 ,csa_tree_add_101_22_pad_groupi_n_1515 ,csa_tree_add_101_22_pad_groupi_n_1461);
  xor csa_tree_add_101_22_pad_groupi_g6117(csa_tree_add_101_22_pad_groupi_n_6 ,csa_tree_add_101_22_pad_groupi_n_1368 ,csa_tree_add_101_22_pad_groupi_n_1406);
  xor csa_tree_add_101_22_pad_groupi_g6118(csa_tree_add_101_22_pad_groupi_n_5 ,csa_tree_add_101_22_pad_groupi_n_1332 ,csa_tree_add_101_22_pad_groupi_n_1350);
  xor csa_tree_add_101_22_pad_groupi_g6119(csa_tree_add_101_22_pad_groupi_n_4 ,csa_tree_add_101_22_pad_groupi_n_836 ,csa_tree_add_101_22_pad_groupi_n_0);
  xor csa_tree_add_101_22_pad_groupi_g6120(csa_tree_add_101_22_pad_groupi_n_3 ,csa_tree_add_101_22_pad_groupi_n_835 ,csa_tree_add_101_22_pad_groupi_n_948);
  xor csa_tree_add_101_22_pad_groupi_g6122(csa_tree_add_101_22_pad_groupi_n_1 ,csa_tree_add_101_22_pad_groupi_n_358 ,in21[9]);
  xor csa_tree_add_101_22_pad_groupi_g6123(csa_tree_add_101_22_pad_groupi_n_0 ,csa_tree_add_101_22_pad_groupi_n_357 ,in21[11]);
  xnor csa_tree_add_107_22_pad_groupi_g4151(n_270 ,csa_tree_add_107_22_pad_groupi_n_1336 ,csa_tree_add_107_22_pad_groupi_n_1558);
  or csa_tree_add_107_22_pad_groupi_g4152(csa_tree_add_107_22_pad_groupi_n_1558 ,csa_tree_add_107_22_pad_groupi_n_1393 ,csa_tree_add_107_22_pad_groupi_n_1556);
  xnor csa_tree_add_107_22_pad_groupi_g4153(n_269 ,csa_tree_add_107_22_pad_groupi_n_1555 ,csa_tree_add_107_22_pad_groupi_n_1404);
  and csa_tree_add_107_22_pad_groupi_g4154(csa_tree_add_107_22_pad_groupi_n_1556 ,csa_tree_add_107_22_pad_groupi_n_1389 ,csa_tree_add_107_22_pad_groupi_n_1555);
  or csa_tree_add_107_22_pad_groupi_g4155(csa_tree_add_107_22_pad_groupi_n_1555 ,csa_tree_add_107_22_pad_groupi_n_1407 ,csa_tree_add_107_22_pad_groupi_n_1553);
  xnor csa_tree_add_107_22_pad_groupi_g4156(n_268 ,csa_tree_add_107_22_pad_groupi_n_1552 ,csa_tree_add_107_22_pad_groupi_n_1434);
  and csa_tree_add_107_22_pad_groupi_g4157(csa_tree_add_107_22_pad_groupi_n_1553 ,csa_tree_add_107_22_pad_groupi_n_1410 ,csa_tree_add_107_22_pad_groupi_n_1552);
  or csa_tree_add_107_22_pad_groupi_g4158(csa_tree_add_107_22_pad_groupi_n_1552 ,csa_tree_add_107_22_pad_groupi_n_1453 ,csa_tree_add_107_22_pad_groupi_n_1550);
  xnor csa_tree_add_107_22_pad_groupi_g4159(n_267 ,csa_tree_add_107_22_pad_groupi_n_1549 ,csa_tree_add_107_22_pad_groupi_n_1462);
  and csa_tree_add_107_22_pad_groupi_g4160(csa_tree_add_107_22_pad_groupi_n_1550 ,csa_tree_add_107_22_pad_groupi_n_1459 ,csa_tree_add_107_22_pad_groupi_n_1549);
  or csa_tree_add_107_22_pad_groupi_g4161(csa_tree_add_107_22_pad_groupi_n_1549 ,csa_tree_add_107_22_pad_groupi_n_1463 ,csa_tree_add_107_22_pad_groupi_n_1547);
  xnor csa_tree_add_107_22_pad_groupi_g4162(n_266 ,csa_tree_add_107_22_pad_groupi_n_1546 ,csa_tree_add_107_22_pad_groupi_n_1483);
  nor csa_tree_add_107_22_pad_groupi_g4163(csa_tree_add_107_22_pad_groupi_n_1547 ,csa_tree_add_107_22_pad_groupi_n_1546 ,csa_tree_add_107_22_pad_groupi_n_1464);
  and csa_tree_add_107_22_pad_groupi_g4164(csa_tree_add_107_22_pad_groupi_n_1546 ,csa_tree_add_107_22_pad_groupi_n_1500 ,csa_tree_add_107_22_pad_groupi_n_1544);
  xnor csa_tree_add_107_22_pad_groupi_g4165(n_265 ,csa_tree_add_107_22_pad_groupi_n_1542 ,csa_tree_add_107_22_pad_groupi_n_1501);
  or csa_tree_add_107_22_pad_groupi_g4166(csa_tree_add_107_22_pad_groupi_n_1544 ,csa_tree_add_107_22_pad_groupi_n_1494 ,csa_tree_add_107_22_pad_groupi_n_1543);
  not csa_tree_add_107_22_pad_groupi_g4167(csa_tree_add_107_22_pad_groupi_n_1543 ,csa_tree_add_107_22_pad_groupi_n_1542);
  or csa_tree_add_107_22_pad_groupi_g4168(csa_tree_add_107_22_pad_groupi_n_1542 ,csa_tree_add_107_22_pad_groupi_n_1499 ,csa_tree_add_107_22_pad_groupi_n_1540);
  xnor csa_tree_add_107_22_pad_groupi_g4169(n_264 ,csa_tree_add_107_22_pad_groupi_n_1539 ,csa_tree_add_107_22_pad_groupi_n_1503);
  nor csa_tree_add_107_22_pad_groupi_g4170(csa_tree_add_107_22_pad_groupi_n_1540 ,csa_tree_add_107_22_pad_groupi_n_1496 ,csa_tree_add_107_22_pad_groupi_n_1539);
  and csa_tree_add_107_22_pad_groupi_g4171(csa_tree_add_107_22_pad_groupi_n_1539 ,csa_tree_add_107_22_pad_groupi_n_1538 ,csa_tree_add_107_22_pad_groupi_n_1510);
  or csa_tree_add_107_22_pad_groupi_g4173(csa_tree_add_107_22_pad_groupi_n_1538 ,csa_tree_add_107_22_pad_groupi_n_1513 ,csa_tree_add_107_22_pad_groupi_n_1537);
  and csa_tree_add_107_22_pad_groupi_g4175(csa_tree_add_107_22_pad_groupi_n_1537 ,csa_tree_add_107_22_pad_groupi_n_1512 ,csa_tree_add_107_22_pad_groupi_n_1535);
  xnor csa_tree_add_107_22_pad_groupi_g4176(n_262 ,csa_tree_add_107_22_pad_groupi_n_1534 ,csa_tree_add_107_22_pad_groupi_n_1519);
  or csa_tree_add_107_22_pad_groupi_g4177(csa_tree_add_107_22_pad_groupi_n_1535 ,csa_tree_add_107_22_pad_groupi_n_1514 ,csa_tree_add_107_22_pad_groupi_n_1534);
  and csa_tree_add_107_22_pad_groupi_g4178(csa_tree_add_107_22_pad_groupi_n_1534 ,csa_tree_add_107_22_pad_groupi_n_1533 ,csa_tree_add_107_22_pad_groupi_n_1511);
  or csa_tree_add_107_22_pad_groupi_g4180(csa_tree_add_107_22_pad_groupi_n_1533 ,csa_tree_add_107_22_pad_groupi_n_1505 ,csa_tree_add_107_22_pad_groupi_n_1532);
  and csa_tree_add_107_22_pad_groupi_g4182(csa_tree_add_107_22_pad_groupi_n_1532 ,csa_tree_add_107_22_pad_groupi_n_1506 ,csa_tree_add_107_22_pad_groupi_n_1530);
  xnor csa_tree_add_107_22_pad_groupi_g4183(n_260 ,csa_tree_add_107_22_pad_groupi_n_1529 ,csa_tree_add_107_22_pad_groupi_n_1517);
  or csa_tree_add_107_22_pad_groupi_g4184(csa_tree_add_107_22_pad_groupi_n_1530 ,csa_tree_add_107_22_pad_groupi_n_1507 ,csa_tree_add_107_22_pad_groupi_n_1529);
  and csa_tree_add_107_22_pad_groupi_g4185(csa_tree_add_107_22_pad_groupi_n_1529 ,csa_tree_add_107_22_pad_groupi_n_1508 ,csa_tree_add_107_22_pad_groupi_n_1527);
  xnor csa_tree_add_107_22_pad_groupi_g4186(n_259 ,csa_tree_add_107_22_pad_groupi_n_1526 ,csa_tree_add_107_22_pad_groupi_n_1516);
  or csa_tree_add_107_22_pad_groupi_g4187(csa_tree_add_107_22_pad_groupi_n_1527 ,csa_tree_add_107_22_pad_groupi_n_1526 ,csa_tree_add_107_22_pad_groupi_n_1509);
  and csa_tree_add_107_22_pad_groupi_g4188(csa_tree_add_107_22_pad_groupi_n_1526 ,csa_tree_add_107_22_pad_groupi_n_1471 ,csa_tree_add_107_22_pad_groupi_n_1525);
  or csa_tree_add_107_22_pad_groupi_g4190(csa_tree_add_107_22_pad_groupi_n_1525 ,csa_tree_add_107_22_pad_groupi_n_1470 ,csa_tree_add_107_22_pad_groupi_n_1524);
  and csa_tree_add_107_22_pad_groupi_g4192(csa_tree_add_107_22_pad_groupi_n_1524 ,csa_tree_add_107_22_pad_groupi_n_1498 ,csa_tree_add_107_22_pad_groupi_n_1523);
  or csa_tree_add_107_22_pad_groupi_g4194(csa_tree_add_107_22_pad_groupi_n_1523 ,csa_tree_add_107_22_pad_groupi_n_1497 ,csa_tree_add_107_22_pad_groupi_n_1522);
  and csa_tree_add_107_22_pad_groupi_g4196(csa_tree_add_107_22_pad_groupi_n_1522 ,csa_tree_add_107_22_pad_groupi_n_1452 ,csa_tree_add_107_22_pad_groupi_n_1521);
  or csa_tree_add_107_22_pad_groupi_g4198(csa_tree_add_107_22_pad_groupi_n_1521 ,csa_tree_add_107_22_pad_groupi_n_1451 ,csa_tree_add_107_22_pad_groupi_n_1515);
  xnor csa_tree_add_107_22_pad_groupi_g4199(csa_tree_add_107_22_pad_groupi_n_1520 ,csa_tree_add_107_22_pad_groupi_n_1475 ,csa_tree_add_107_22_pad_groupi_n_1491);
  xnor csa_tree_add_107_22_pad_groupi_g4200(csa_tree_add_107_22_pad_groupi_n_1519 ,csa_tree_add_107_22_pad_groupi_n_1473 ,csa_tree_add_107_22_pad_groupi_n_1489);
  xnor csa_tree_add_107_22_pad_groupi_g4201(csa_tree_add_107_22_pad_groupi_n_1518 ,csa_tree_add_107_22_pad_groupi_n_1480 ,csa_tree_add_107_22_pad_groupi_n_1487);
  xnor csa_tree_add_107_22_pad_groupi_g4202(csa_tree_add_107_22_pad_groupi_n_1517 ,csa_tree_add_107_22_pad_groupi_n_1477 ,csa_tree_add_107_22_pad_groupi_n_1493);
  xnor csa_tree_add_107_22_pad_groupi_g4203(csa_tree_add_107_22_pad_groupi_n_1516 ,csa_tree_add_107_22_pad_groupi_n_1448 ,csa_tree_add_107_22_pad_groupi_n_1485);
  nor csa_tree_add_107_22_pad_groupi_g4205(csa_tree_add_107_22_pad_groupi_n_1514 ,csa_tree_add_107_22_pad_groupi_n_1472 ,csa_tree_add_107_22_pad_groupi_n_1489);
  nor csa_tree_add_107_22_pad_groupi_g4206(csa_tree_add_107_22_pad_groupi_n_1513 ,csa_tree_add_107_22_pad_groupi_n_1475 ,csa_tree_add_107_22_pad_groupi_n_1491);
  or csa_tree_add_107_22_pad_groupi_g4207(csa_tree_add_107_22_pad_groupi_n_1512 ,csa_tree_add_107_22_pad_groupi_n_1473 ,csa_tree_add_107_22_pad_groupi_n_1488);
  or csa_tree_add_107_22_pad_groupi_g4208(csa_tree_add_107_22_pad_groupi_n_1511 ,csa_tree_add_107_22_pad_groupi_n_1479 ,csa_tree_add_107_22_pad_groupi_n_1486);
  or csa_tree_add_107_22_pad_groupi_g4209(csa_tree_add_107_22_pad_groupi_n_1510 ,csa_tree_add_107_22_pad_groupi_n_1474 ,csa_tree_add_107_22_pad_groupi_n_1490);
  nor csa_tree_add_107_22_pad_groupi_g4210(csa_tree_add_107_22_pad_groupi_n_1509 ,csa_tree_add_107_22_pad_groupi_n_1447 ,csa_tree_add_107_22_pad_groupi_n_1485);
  and csa_tree_add_107_22_pad_groupi_g4211(csa_tree_add_107_22_pad_groupi_n_1515 ,csa_tree_add_107_22_pad_groupi_n_1450 ,csa_tree_add_107_22_pad_groupi_n_1495);
  or csa_tree_add_107_22_pad_groupi_g4212(csa_tree_add_107_22_pad_groupi_n_1508 ,csa_tree_add_107_22_pad_groupi_n_1448 ,csa_tree_add_107_22_pad_groupi_n_1484);
  nor csa_tree_add_107_22_pad_groupi_g4213(csa_tree_add_107_22_pad_groupi_n_1507 ,csa_tree_add_107_22_pad_groupi_n_1476 ,csa_tree_add_107_22_pad_groupi_n_1493);
  or csa_tree_add_107_22_pad_groupi_g4214(csa_tree_add_107_22_pad_groupi_n_1506 ,csa_tree_add_107_22_pad_groupi_n_1477 ,csa_tree_add_107_22_pad_groupi_n_1492);
  nor csa_tree_add_107_22_pad_groupi_g4215(csa_tree_add_107_22_pad_groupi_n_1505 ,csa_tree_add_107_22_pad_groupi_n_1480 ,csa_tree_add_107_22_pad_groupi_n_1487);
  xnor csa_tree_add_107_22_pad_groupi_g4216(n_255 ,csa_tree_add_107_22_pad_groupi_n_1481 ,csa_tree_add_107_22_pad_groupi_n_1460);
  xnor csa_tree_add_107_22_pad_groupi_g4217(csa_tree_add_107_22_pad_groupi_n_1503 ,csa_tree_add_107_22_pad_groupi_n_1478 ,csa_tree_add_107_22_pad_groupi_n_1467);
  xnor csa_tree_add_107_22_pad_groupi_g4218(csa_tree_add_107_22_pad_groupi_n_1502 ,csa_tree_add_107_22_pad_groupi_n_1412 ,csa_tree_add_107_22_pad_groupi_n_1466);
  xnor csa_tree_add_107_22_pad_groupi_g4219(csa_tree_add_107_22_pad_groupi_n_1501 ,csa_tree_add_107_22_pad_groupi_n_1442 ,csa_tree_add_107_22_pad_groupi_n_1469);
  or csa_tree_add_107_22_pad_groupi_g4220(csa_tree_add_107_22_pad_groupi_n_1500 ,csa_tree_add_107_22_pad_groupi_n_1441 ,csa_tree_add_107_22_pad_groupi_n_6);
  nor csa_tree_add_107_22_pad_groupi_g4221(csa_tree_add_107_22_pad_groupi_n_1499 ,csa_tree_add_107_22_pad_groupi_n_1478 ,csa_tree_add_107_22_pad_groupi_n_1468);
  or csa_tree_add_107_22_pad_groupi_g4222(csa_tree_add_107_22_pad_groupi_n_1498 ,csa_tree_add_107_22_pad_groupi_n_1411 ,csa_tree_add_107_22_pad_groupi_n_1465);
  nor csa_tree_add_107_22_pad_groupi_g4223(csa_tree_add_107_22_pad_groupi_n_1497 ,csa_tree_add_107_22_pad_groupi_n_1412 ,csa_tree_add_107_22_pad_groupi_n_1466);
  and csa_tree_add_107_22_pad_groupi_g4224(csa_tree_add_107_22_pad_groupi_n_1496 ,csa_tree_add_107_22_pad_groupi_n_1478 ,csa_tree_add_107_22_pad_groupi_n_1468);
  or csa_tree_add_107_22_pad_groupi_g4225(csa_tree_add_107_22_pad_groupi_n_1495 ,csa_tree_add_107_22_pad_groupi_n_1449 ,csa_tree_add_107_22_pad_groupi_n_1481);
  nor csa_tree_add_107_22_pad_groupi_g4226(csa_tree_add_107_22_pad_groupi_n_1494 ,csa_tree_add_107_22_pad_groupi_n_1442 ,csa_tree_add_107_22_pad_groupi_n_1469);
  not csa_tree_add_107_22_pad_groupi_g4227(csa_tree_add_107_22_pad_groupi_n_1493 ,csa_tree_add_107_22_pad_groupi_n_1492);
  not csa_tree_add_107_22_pad_groupi_g4228(csa_tree_add_107_22_pad_groupi_n_1491 ,csa_tree_add_107_22_pad_groupi_n_1490);
  not csa_tree_add_107_22_pad_groupi_g4229(csa_tree_add_107_22_pad_groupi_n_1489 ,csa_tree_add_107_22_pad_groupi_n_1488);
  not csa_tree_add_107_22_pad_groupi_g4230(csa_tree_add_107_22_pad_groupi_n_1487 ,csa_tree_add_107_22_pad_groupi_n_1486);
  not csa_tree_add_107_22_pad_groupi_g4231(csa_tree_add_107_22_pad_groupi_n_1485 ,csa_tree_add_107_22_pad_groupi_n_1484);
  xnor csa_tree_add_107_22_pad_groupi_g4232(csa_tree_add_107_22_pad_groupi_n_1483 ,csa_tree_add_107_22_pad_groupi_n_1440 ,csa_tree_add_107_22_pad_groupi_n_1445);
  xnor csa_tree_add_107_22_pad_groupi_g4233(csa_tree_add_107_22_pad_groupi_n_1482 ,csa_tree_add_107_22_pad_groupi_n_1419 ,csa_tree_add_107_22_pad_groupi_n_1444);
  xnor csa_tree_add_107_22_pad_groupi_g4234(csa_tree_add_107_22_pad_groupi_n_1492 ,csa_tree_add_107_22_pad_groupi_n_1387 ,csa_tree_add_107_22_pad_groupi_n_1438);
  xnor csa_tree_add_107_22_pad_groupi_g4235(csa_tree_add_107_22_pad_groupi_n_1490 ,csa_tree_add_107_22_pad_groupi_n_1400 ,csa_tree_add_107_22_pad_groupi_n_1433);
  xnor csa_tree_add_107_22_pad_groupi_g4236(csa_tree_add_107_22_pad_groupi_n_1488 ,csa_tree_add_107_22_pad_groupi_n_1401 ,csa_tree_add_107_22_pad_groupi_n_1436);
  xnor csa_tree_add_107_22_pad_groupi_g4237(csa_tree_add_107_22_pad_groupi_n_1486 ,csa_tree_add_107_22_pad_groupi_n_1402 ,csa_tree_add_107_22_pad_groupi_n_1437);
  xnor csa_tree_add_107_22_pad_groupi_g4238(csa_tree_add_107_22_pad_groupi_n_1484 ,csa_tree_add_107_22_pad_groupi_n_1403 ,csa_tree_add_107_22_pad_groupi_n_1435);
  not csa_tree_add_107_22_pad_groupi_g4239(csa_tree_add_107_22_pad_groupi_n_1479 ,csa_tree_add_107_22_pad_groupi_n_1480);
  not csa_tree_add_107_22_pad_groupi_g4240(csa_tree_add_107_22_pad_groupi_n_1477 ,csa_tree_add_107_22_pad_groupi_n_1476);
  not csa_tree_add_107_22_pad_groupi_g4241(csa_tree_add_107_22_pad_groupi_n_1474 ,csa_tree_add_107_22_pad_groupi_n_1475);
  not csa_tree_add_107_22_pad_groupi_g4242(csa_tree_add_107_22_pad_groupi_n_1473 ,csa_tree_add_107_22_pad_groupi_n_1472);
  or csa_tree_add_107_22_pad_groupi_g4243(csa_tree_add_107_22_pad_groupi_n_1471 ,csa_tree_add_107_22_pad_groupi_n_1418 ,csa_tree_add_107_22_pad_groupi_n_1443);
  nor csa_tree_add_107_22_pad_groupi_g4244(csa_tree_add_107_22_pad_groupi_n_1470 ,csa_tree_add_107_22_pad_groupi_n_1419 ,csa_tree_add_107_22_pad_groupi_n_1444);
  and csa_tree_add_107_22_pad_groupi_g4245(csa_tree_add_107_22_pad_groupi_n_1481 ,csa_tree_add_107_22_pad_groupi_n_1371 ,csa_tree_add_107_22_pad_groupi_n_1439);
  or csa_tree_add_107_22_pad_groupi_g4246(csa_tree_add_107_22_pad_groupi_n_1480 ,csa_tree_add_107_22_pad_groupi_n_1424 ,csa_tree_add_107_22_pad_groupi_n_1456);
  and csa_tree_add_107_22_pad_groupi_g4247(csa_tree_add_107_22_pad_groupi_n_1478 ,csa_tree_add_107_22_pad_groupi_n_1431 ,csa_tree_add_107_22_pad_groupi_n_1454);
  or csa_tree_add_107_22_pad_groupi_g4248(csa_tree_add_107_22_pad_groupi_n_1476 ,csa_tree_add_107_22_pad_groupi_n_1422 ,csa_tree_add_107_22_pad_groupi_n_1455);
  or csa_tree_add_107_22_pad_groupi_g4249(csa_tree_add_107_22_pad_groupi_n_1475 ,csa_tree_add_107_22_pad_groupi_n_1429 ,csa_tree_add_107_22_pad_groupi_n_1458);
  or csa_tree_add_107_22_pad_groupi_g4250(csa_tree_add_107_22_pad_groupi_n_1472 ,csa_tree_add_107_22_pad_groupi_n_1426 ,csa_tree_add_107_22_pad_groupi_n_1457);
  not csa_tree_add_107_22_pad_groupi_g4251(csa_tree_add_107_22_pad_groupi_n_1469 ,csa_tree_add_107_22_pad_groupi_n_6);
  not csa_tree_add_107_22_pad_groupi_g4252(csa_tree_add_107_22_pad_groupi_n_1468 ,csa_tree_add_107_22_pad_groupi_n_1467);
  not csa_tree_add_107_22_pad_groupi_g4253(csa_tree_add_107_22_pad_groupi_n_1466 ,csa_tree_add_107_22_pad_groupi_n_1465);
  and csa_tree_add_107_22_pad_groupi_g4254(csa_tree_add_107_22_pad_groupi_n_1464 ,csa_tree_add_107_22_pad_groupi_n_1440 ,csa_tree_add_107_22_pad_groupi_n_1446);
  nor csa_tree_add_107_22_pad_groupi_g4255(csa_tree_add_107_22_pad_groupi_n_1463 ,csa_tree_add_107_22_pad_groupi_n_1440 ,csa_tree_add_107_22_pad_groupi_n_1446);
  xnor csa_tree_add_107_22_pad_groupi_g4256(csa_tree_add_107_22_pad_groupi_n_1462 ,csa_tree_add_107_22_pad_groupi_n_1432 ,csa_tree_add_107_22_pad_groupi_n_1413);
  xnor csa_tree_add_107_22_pad_groupi_g4257(csa_tree_add_107_22_pad_groupi_n_1461 ,csa_tree_add_107_22_pad_groupi_n_1397 ,csa_tree_add_107_22_pad_groupi_n_1417);
  xnor csa_tree_add_107_22_pad_groupi_g4258(csa_tree_add_107_22_pad_groupi_n_1460 ,csa_tree_add_107_22_pad_groupi_n_1367 ,csa_tree_add_107_22_pad_groupi_n_1415);
  xnor csa_tree_add_107_22_pad_groupi_g4260(csa_tree_add_107_22_pad_groupi_n_1467 ,csa_tree_add_107_22_pad_groupi_n_1384 ,csa_tree_add_107_22_pad_groupi_n_1405);
  xnor csa_tree_add_107_22_pad_groupi_g4261(csa_tree_add_107_22_pad_groupi_n_1465 ,csa_tree_add_107_22_pad_groupi_n_1295 ,csa_tree_add_107_22_pad_groupi_n_5);
  or csa_tree_add_107_22_pad_groupi_g4262(csa_tree_add_107_22_pad_groupi_n_1459 ,csa_tree_add_107_22_pad_groupi_n_1432 ,csa_tree_add_107_22_pad_groupi_n_1413);
  and csa_tree_add_107_22_pad_groupi_g4263(csa_tree_add_107_22_pad_groupi_n_1458 ,csa_tree_add_107_22_pad_groupi_n_1401 ,csa_tree_add_107_22_pad_groupi_n_1427);
  and csa_tree_add_107_22_pad_groupi_g4264(csa_tree_add_107_22_pad_groupi_n_1457 ,csa_tree_add_107_22_pad_groupi_n_1402 ,csa_tree_add_107_22_pad_groupi_n_1425);
  and csa_tree_add_107_22_pad_groupi_g4265(csa_tree_add_107_22_pad_groupi_n_1456 ,csa_tree_add_107_22_pad_groupi_n_1387 ,csa_tree_add_107_22_pad_groupi_n_1423);
  and csa_tree_add_107_22_pad_groupi_g4266(csa_tree_add_107_22_pad_groupi_n_1455 ,csa_tree_add_107_22_pad_groupi_n_1403 ,csa_tree_add_107_22_pad_groupi_n_1421);
  or csa_tree_add_107_22_pad_groupi_g4267(csa_tree_add_107_22_pad_groupi_n_1454 ,csa_tree_add_107_22_pad_groupi_n_1430 ,csa_tree_add_107_22_pad_groupi_n_1386);
  and csa_tree_add_107_22_pad_groupi_g4268(csa_tree_add_107_22_pad_groupi_n_1453 ,csa_tree_add_107_22_pad_groupi_n_1432 ,csa_tree_add_107_22_pad_groupi_n_1413);
  or csa_tree_add_107_22_pad_groupi_g4269(csa_tree_add_107_22_pad_groupi_n_1452 ,csa_tree_add_107_22_pad_groupi_n_1396 ,csa_tree_add_107_22_pad_groupi_n_1416);
  nor csa_tree_add_107_22_pad_groupi_g4270(csa_tree_add_107_22_pad_groupi_n_1451 ,csa_tree_add_107_22_pad_groupi_n_1397 ,csa_tree_add_107_22_pad_groupi_n_1417);
  or csa_tree_add_107_22_pad_groupi_g4271(csa_tree_add_107_22_pad_groupi_n_1450 ,csa_tree_add_107_22_pad_groupi_n_1367 ,csa_tree_add_107_22_pad_groupi_n_1414);
  nor csa_tree_add_107_22_pad_groupi_g4272(csa_tree_add_107_22_pad_groupi_n_1449 ,csa_tree_add_107_22_pad_groupi_n_1366 ,csa_tree_add_107_22_pad_groupi_n_1415);
  not csa_tree_add_107_22_pad_groupi_g4273(csa_tree_add_107_22_pad_groupi_n_1448 ,csa_tree_add_107_22_pad_groupi_n_1447);
  not csa_tree_add_107_22_pad_groupi_g4274(csa_tree_add_107_22_pad_groupi_n_1446 ,csa_tree_add_107_22_pad_groupi_n_1445);
  not csa_tree_add_107_22_pad_groupi_g4275(csa_tree_add_107_22_pad_groupi_n_1444 ,csa_tree_add_107_22_pad_groupi_n_1443);
  not csa_tree_add_107_22_pad_groupi_g4276(csa_tree_add_107_22_pad_groupi_n_1441 ,csa_tree_add_107_22_pad_groupi_n_1442);
  or csa_tree_add_107_22_pad_groupi_g4277(csa_tree_add_107_22_pad_groupi_n_1439 ,csa_tree_add_107_22_pad_groupi_n_1372 ,csa_tree_add_107_22_pad_groupi_n_1428);
  xnor csa_tree_add_107_22_pad_groupi_g4278(csa_tree_add_107_22_pad_groupi_n_1438 ,csa_tree_add_107_22_pad_groupi_n_1291 ,csa_tree_add_107_22_pad_groupi_n_1379);
  xnor csa_tree_add_107_22_pad_groupi_g4279(csa_tree_add_107_22_pad_groupi_n_1437 ,csa_tree_add_107_22_pad_groupi_n_1293 ,csa_tree_add_107_22_pad_groupi_n_1381);
  xnor csa_tree_add_107_22_pad_groupi_g4280(csa_tree_add_107_22_pad_groupi_n_1436 ,csa_tree_add_107_22_pad_groupi_n_1301 ,csa_tree_add_107_22_pad_groupi_n_1376);
  xnor csa_tree_add_107_22_pad_groupi_g4281(csa_tree_add_107_22_pad_groupi_n_1435 ,csa_tree_add_107_22_pad_groupi_n_1303 ,csa_tree_add_107_22_pad_groupi_n_1383);
  xnor csa_tree_add_107_22_pad_groupi_g4282(csa_tree_add_107_22_pad_groupi_n_1434 ,csa_tree_add_107_22_pad_groupi_n_1377 ,csa_tree_add_107_22_pad_groupi_n_1398);
  xnor csa_tree_add_107_22_pad_groupi_g4283(csa_tree_add_107_22_pad_groupi_n_1433 ,csa_tree_add_107_22_pad_groupi_n_1298 ,csa_tree_add_107_22_pad_groupi_n_1386);
  or csa_tree_add_107_22_pad_groupi_g4284(csa_tree_add_107_22_pad_groupi_n_1447 ,csa_tree_add_107_22_pad_groupi_n_1340 ,csa_tree_add_107_22_pad_groupi_n_1420);
  xnor csa_tree_add_107_22_pad_groupi_g4285(csa_tree_add_107_22_pad_groupi_n_1445 ,csa_tree_add_107_22_pad_groupi_n_1334 ,csa_tree_add_107_22_pad_groupi_n_1370);
  xnor csa_tree_add_107_22_pad_groupi_g4286(csa_tree_add_107_22_pad_groupi_n_1443 ,csa_tree_add_107_22_pad_groupi_n_1385 ,csa_tree_add_107_22_pad_groupi_n_1369);
  or csa_tree_add_107_22_pad_groupi_g4287(csa_tree_add_107_22_pad_groupi_n_1442 ,csa_tree_add_107_22_pad_groupi_n_1374 ,csa_tree_add_107_22_pad_groupi_n_1409);
  and csa_tree_add_107_22_pad_groupi_g4288(csa_tree_add_107_22_pad_groupi_n_1440 ,csa_tree_add_107_22_pad_groupi_n_1395 ,csa_tree_add_107_22_pad_groupi_n_1408);
  or csa_tree_add_107_22_pad_groupi_g4289(csa_tree_add_107_22_pad_groupi_n_1431 ,csa_tree_add_107_22_pad_groupi_n_1297 ,csa_tree_add_107_22_pad_groupi_n_1399);
  nor csa_tree_add_107_22_pad_groupi_g4290(csa_tree_add_107_22_pad_groupi_n_1430 ,csa_tree_add_107_22_pad_groupi_n_1298 ,csa_tree_add_107_22_pad_groupi_n_1400);
  nor csa_tree_add_107_22_pad_groupi_g4291(csa_tree_add_107_22_pad_groupi_n_1429 ,csa_tree_add_107_22_pad_groupi_n_1300 ,csa_tree_add_107_22_pad_groupi_n_1376);
  nor csa_tree_add_107_22_pad_groupi_g4292(csa_tree_add_107_22_pad_groupi_n_1428 ,csa_tree_add_107_22_pad_groupi_n_1363 ,csa_tree_add_107_22_pad_groupi_n_1394);
  or csa_tree_add_107_22_pad_groupi_g4293(csa_tree_add_107_22_pad_groupi_n_1427 ,csa_tree_add_107_22_pad_groupi_n_1301 ,csa_tree_add_107_22_pad_groupi_n_1375);
  nor csa_tree_add_107_22_pad_groupi_g4294(csa_tree_add_107_22_pad_groupi_n_1426 ,csa_tree_add_107_22_pad_groupi_n_1292 ,csa_tree_add_107_22_pad_groupi_n_1381);
  or csa_tree_add_107_22_pad_groupi_g4295(csa_tree_add_107_22_pad_groupi_n_1425 ,csa_tree_add_107_22_pad_groupi_n_1293 ,csa_tree_add_107_22_pad_groupi_n_1380);
  nor csa_tree_add_107_22_pad_groupi_g4296(csa_tree_add_107_22_pad_groupi_n_1424 ,csa_tree_add_107_22_pad_groupi_n_1290 ,csa_tree_add_107_22_pad_groupi_n_1379);
  or csa_tree_add_107_22_pad_groupi_g4297(csa_tree_add_107_22_pad_groupi_n_1423 ,csa_tree_add_107_22_pad_groupi_n_1291 ,csa_tree_add_107_22_pad_groupi_n_1378);
  nor csa_tree_add_107_22_pad_groupi_g4298(csa_tree_add_107_22_pad_groupi_n_1422 ,csa_tree_add_107_22_pad_groupi_n_1302 ,csa_tree_add_107_22_pad_groupi_n_1383);
  or csa_tree_add_107_22_pad_groupi_g4299(csa_tree_add_107_22_pad_groupi_n_1421 ,csa_tree_add_107_22_pad_groupi_n_1303 ,csa_tree_add_107_22_pad_groupi_n_1382);
  nor csa_tree_add_107_22_pad_groupi_g4300(csa_tree_add_107_22_pad_groupi_n_1420 ,csa_tree_add_107_22_pad_groupi_n_1355 ,csa_tree_add_107_22_pad_groupi_n_1385);
  or csa_tree_add_107_22_pad_groupi_g4301(csa_tree_add_107_22_pad_groupi_n_1432 ,csa_tree_add_107_22_pad_groupi_n_1365 ,csa_tree_add_107_22_pad_groupi_n_1391);
  not csa_tree_add_107_22_pad_groupi_g4302(csa_tree_add_107_22_pad_groupi_n_1419 ,csa_tree_add_107_22_pad_groupi_n_1418);
  not csa_tree_add_107_22_pad_groupi_g4303(csa_tree_add_107_22_pad_groupi_n_1417 ,csa_tree_add_107_22_pad_groupi_n_1416);
  not csa_tree_add_107_22_pad_groupi_g4304(csa_tree_add_107_22_pad_groupi_n_1415 ,csa_tree_add_107_22_pad_groupi_n_1414);
  not csa_tree_add_107_22_pad_groupi_g4305(csa_tree_add_107_22_pad_groupi_n_1412 ,csa_tree_add_107_22_pad_groupi_n_1411);
  or csa_tree_add_107_22_pad_groupi_g4306(csa_tree_add_107_22_pad_groupi_n_1410 ,csa_tree_add_107_22_pad_groupi_n_1377 ,csa_tree_add_107_22_pad_groupi_n_1398);
  nor csa_tree_add_107_22_pad_groupi_g4307(csa_tree_add_107_22_pad_groupi_n_1409 ,csa_tree_add_107_22_pad_groupi_n_1384 ,csa_tree_add_107_22_pad_groupi_n_1392);
  or csa_tree_add_107_22_pad_groupi_g4308(csa_tree_add_107_22_pad_groupi_n_1408 ,csa_tree_add_107_22_pad_groupi_n_1368 ,csa_tree_add_107_22_pad_groupi_n_1373);
  and csa_tree_add_107_22_pad_groupi_g4309(csa_tree_add_107_22_pad_groupi_n_1407 ,csa_tree_add_107_22_pad_groupi_n_1377 ,csa_tree_add_107_22_pad_groupi_n_1398);
  xnor csa_tree_add_107_22_pad_groupi_g4310(csa_tree_add_107_22_pad_groupi_n_1406 ,csa_tree_add_107_22_pad_groupi_n_1280 ,csa_tree_add_107_22_pad_groupi_n_1346);
  xnor csa_tree_add_107_22_pad_groupi_g4312(csa_tree_add_107_22_pad_groupi_n_1405 ,csa_tree_add_107_22_pad_groupi_n_1304 ,csa_tree_add_107_22_pad_groupi_n_1348);
  xnor csa_tree_add_107_22_pad_groupi_g4313(csa_tree_add_107_22_pad_groupi_n_1404 ,csa_tree_add_107_22_pad_groupi_n_1309 ,csa_tree_add_107_22_pad_groupi_n_1345);
  and csa_tree_add_107_22_pad_groupi_g4314(csa_tree_add_107_22_pad_groupi_n_1418 ,csa_tree_add_107_22_pad_groupi_n_1354 ,csa_tree_add_107_22_pad_groupi_n_1390);
  xnor csa_tree_add_107_22_pad_groupi_g4315(csa_tree_add_107_22_pad_groupi_n_1416 ,csa_tree_add_107_22_pad_groupi_n_1311 ,csa_tree_add_107_22_pad_groupi_n_1337);
  xnor csa_tree_add_107_22_pad_groupi_g4316(csa_tree_add_107_22_pad_groupi_n_1414 ,csa_tree_add_107_22_pad_groupi_n_1320 ,csa_tree_add_107_22_pad_groupi_n_1335);
  xnor csa_tree_add_107_22_pad_groupi_g4317(csa_tree_add_107_22_pad_groupi_n_1413 ,csa_tree_add_107_22_pad_groupi_n_1333 ,csa_tree_add_107_22_pad_groupi_n_1338);
  and csa_tree_add_107_22_pad_groupi_g4318(csa_tree_add_107_22_pad_groupi_n_1411 ,csa_tree_add_107_22_pad_groupi_n_1356 ,csa_tree_add_107_22_pad_groupi_n_1388);
  not csa_tree_add_107_22_pad_groupi_g4319(csa_tree_add_107_22_pad_groupi_n_1400 ,csa_tree_add_107_22_pad_groupi_n_1399);
  not csa_tree_add_107_22_pad_groupi_g4320(csa_tree_add_107_22_pad_groupi_n_1396 ,csa_tree_add_107_22_pad_groupi_n_1397);
  or csa_tree_add_107_22_pad_groupi_g4321(csa_tree_add_107_22_pad_groupi_n_1395 ,csa_tree_add_107_22_pad_groupi_n_1280 ,csa_tree_add_107_22_pad_groupi_n_1347);
  nor csa_tree_add_107_22_pad_groupi_g4322(csa_tree_add_107_22_pad_groupi_n_1394 ,csa_tree_add_107_22_pad_groupi_n_1362 ,csa_tree_add_107_22_pad_groupi_n_1361);
  and csa_tree_add_107_22_pad_groupi_g4323(csa_tree_add_107_22_pad_groupi_n_1393 ,csa_tree_add_107_22_pad_groupi_n_1309 ,csa_tree_add_107_22_pad_groupi_n_1345);
  and csa_tree_add_107_22_pad_groupi_g4324(csa_tree_add_107_22_pad_groupi_n_1392 ,csa_tree_add_107_22_pad_groupi_n_1304 ,csa_tree_add_107_22_pad_groupi_n_1349);
  and csa_tree_add_107_22_pad_groupi_g4325(csa_tree_add_107_22_pad_groupi_n_1391 ,csa_tree_add_107_22_pad_groupi_n_1334 ,csa_tree_add_107_22_pad_groupi_n_1360);
  or csa_tree_add_107_22_pad_groupi_g4326(csa_tree_add_107_22_pad_groupi_n_1390 ,csa_tree_add_107_22_pad_groupi_n_1353 ,csa_tree_add_107_22_pad_groupi_n_1350);
  or csa_tree_add_107_22_pad_groupi_g4327(csa_tree_add_107_22_pad_groupi_n_1389 ,csa_tree_add_107_22_pad_groupi_n_1309 ,csa_tree_add_107_22_pad_groupi_n_1345);
  or csa_tree_add_107_22_pad_groupi_g4328(csa_tree_add_107_22_pad_groupi_n_1388 ,csa_tree_add_107_22_pad_groupi_n_1305 ,csa_tree_add_107_22_pad_groupi_n_1342);
  or csa_tree_add_107_22_pad_groupi_g4329(csa_tree_add_107_22_pad_groupi_n_1403 ,csa_tree_add_107_22_pad_groupi_n_1246 ,csa_tree_add_107_22_pad_groupi_n_1359);
  or csa_tree_add_107_22_pad_groupi_g4330(csa_tree_add_107_22_pad_groupi_n_1402 ,csa_tree_add_107_22_pad_groupi_n_1230 ,csa_tree_add_107_22_pad_groupi_n_1343);
  or csa_tree_add_107_22_pad_groupi_g4331(csa_tree_add_107_22_pad_groupi_n_1401 ,csa_tree_add_107_22_pad_groupi_n_1232 ,csa_tree_add_107_22_pad_groupi_n_1339);
  and csa_tree_add_107_22_pad_groupi_g4332(csa_tree_add_107_22_pad_groupi_n_1399 ,csa_tree_add_107_22_pad_groupi_n_1254 ,csa_tree_add_107_22_pad_groupi_n_1364);
  or csa_tree_add_107_22_pad_groupi_g4333(csa_tree_add_107_22_pad_groupi_n_1398 ,csa_tree_add_107_22_pad_groupi_n_1329 ,csa_tree_add_107_22_pad_groupi_n_1357);
  or csa_tree_add_107_22_pad_groupi_g4334(csa_tree_add_107_22_pad_groupi_n_1397 ,csa_tree_add_107_22_pad_groupi_n_1323 ,csa_tree_add_107_22_pad_groupi_n_1358);
  not csa_tree_add_107_22_pad_groupi_g4335(csa_tree_add_107_22_pad_groupi_n_1383 ,csa_tree_add_107_22_pad_groupi_n_1382);
  not csa_tree_add_107_22_pad_groupi_g4336(csa_tree_add_107_22_pad_groupi_n_1381 ,csa_tree_add_107_22_pad_groupi_n_1380);
  not csa_tree_add_107_22_pad_groupi_g4337(csa_tree_add_107_22_pad_groupi_n_1379 ,csa_tree_add_107_22_pad_groupi_n_1378);
  not csa_tree_add_107_22_pad_groupi_g4338(csa_tree_add_107_22_pad_groupi_n_1376 ,csa_tree_add_107_22_pad_groupi_n_1375);
  nor csa_tree_add_107_22_pad_groupi_g4339(csa_tree_add_107_22_pad_groupi_n_1374 ,csa_tree_add_107_22_pad_groupi_n_1304 ,csa_tree_add_107_22_pad_groupi_n_1349);
  and csa_tree_add_107_22_pad_groupi_g4340(csa_tree_add_107_22_pad_groupi_n_1373 ,csa_tree_add_107_22_pad_groupi_n_1280 ,csa_tree_add_107_22_pad_groupi_n_1347);
  nor csa_tree_add_107_22_pad_groupi_g4341(csa_tree_add_107_22_pad_groupi_n_1372 ,csa_tree_add_107_22_pad_groupi_n_1306 ,csa_tree_add_107_22_pad_groupi_n_1352);
  or csa_tree_add_107_22_pad_groupi_g4342(csa_tree_add_107_22_pad_groupi_n_1371 ,csa_tree_add_107_22_pad_groupi_n_1307 ,csa_tree_add_107_22_pad_groupi_n_1351);
  xnor csa_tree_add_107_22_pad_groupi_g4343(csa_tree_add_107_22_pad_groupi_n_1370 ,csa_tree_add_107_22_pad_groupi_n_1261 ,csa_tree_add_107_22_pad_groupi_n_1310);
  xnor csa_tree_add_107_22_pad_groupi_g4344(csa_tree_add_107_22_pad_groupi_n_1369 ,csa_tree_add_107_22_pad_groupi_n_1299 ,csa_tree_add_107_22_pad_groupi_n_1330);
  or csa_tree_add_107_22_pad_groupi_g4345(csa_tree_add_107_22_pad_groupi_n_1387 ,csa_tree_add_107_22_pad_groupi_n_1227 ,csa_tree_add_107_22_pad_groupi_n_1341);
  xnor csa_tree_add_107_22_pad_groupi_g4346(csa_tree_add_107_22_pad_groupi_n_1386 ,csa_tree_add_107_22_pad_groupi_n_1317 ,csa_tree_add_107_22_pad_groupi_n_1273);
  xnor csa_tree_add_107_22_pad_groupi_g4347(csa_tree_add_107_22_pad_groupi_n_1385 ,csa_tree_add_107_22_pad_groupi_n_1316 ,csa_tree_add_107_22_pad_groupi_n_1268);
  and csa_tree_add_107_22_pad_groupi_g4348(csa_tree_add_107_22_pad_groupi_n_1384 ,csa_tree_add_107_22_pad_groupi_n_1225 ,csa_tree_add_107_22_pad_groupi_n_1344);
  xnor csa_tree_add_107_22_pad_groupi_g4349(csa_tree_add_107_22_pad_groupi_n_1382 ,csa_tree_add_107_22_pad_groupi_n_1313 ,csa_tree_add_107_22_pad_groupi_n_1266);
  xnor csa_tree_add_107_22_pad_groupi_g4350(csa_tree_add_107_22_pad_groupi_n_1380 ,csa_tree_add_107_22_pad_groupi_n_1315 ,csa_tree_add_107_22_pad_groupi_n_1270);
  xnor csa_tree_add_107_22_pad_groupi_g4351(csa_tree_add_107_22_pad_groupi_n_1378 ,csa_tree_add_107_22_pad_groupi_n_1314 ,csa_tree_add_107_22_pad_groupi_n_1267);
  xnor csa_tree_add_107_22_pad_groupi_g4352(csa_tree_add_107_22_pad_groupi_n_1377 ,csa_tree_add_107_22_pad_groupi_n_1262 ,csa_tree_add_107_22_pad_groupi_n_1308);
  xnor csa_tree_add_107_22_pad_groupi_g4353(csa_tree_add_107_22_pad_groupi_n_1375 ,csa_tree_add_107_22_pad_groupi_n_1318 ,csa_tree_add_107_22_pad_groupi_n_1271);
  not csa_tree_add_107_22_pad_groupi_g4355(csa_tree_add_107_22_pad_groupi_n_1367 ,csa_tree_add_107_22_pad_groupi_n_1366);
  and csa_tree_add_107_22_pad_groupi_g4356(csa_tree_add_107_22_pad_groupi_n_1365 ,csa_tree_add_107_22_pad_groupi_n_1261 ,csa_tree_add_107_22_pad_groupi_n_1310);
  or csa_tree_add_107_22_pad_groupi_g4357(csa_tree_add_107_22_pad_groupi_n_1364 ,csa_tree_add_107_22_pad_groupi_n_1224 ,csa_tree_add_107_22_pad_groupi_n_1319);
  and csa_tree_add_107_22_pad_groupi_g4358(csa_tree_add_107_22_pad_groupi_n_1363 ,csa_tree_add_107_22_pad_groupi_n_1265 ,csa_tree_add_107_22_pad_groupi_n_1321);
  nor csa_tree_add_107_22_pad_groupi_g4359(csa_tree_add_107_22_pad_groupi_n_1362 ,csa_tree_add_107_22_pad_groupi_n_1265 ,csa_tree_add_107_22_pad_groupi_n_1321);
  nor csa_tree_add_107_22_pad_groupi_g4360(csa_tree_add_107_22_pad_groupi_n_1361 ,csa_tree_add_107_22_pad_groupi_n_1285 ,csa_tree_add_107_22_pad_groupi_n_1326);
  or csa_tree_add_107_22_pad_groupi_g4361(csa_tree_add_107_22_pad_groupi_n_1360 ,csa_tree_add_107_22_pad_groupi_n_1261 ,csa_tree_add_107_22_pad_groupi_n_1310);
  nor csa_tree_add_107_22_pad_groupi_g4362(csa_tree_add_107_22_pad_groupi_n_1359 ,csa_tree_add_107_22_pad_groupi_n_1245 ,csa_tree_add_107_22_pad_groupi_n_1316);
  nor csa_tree_add_107_22_pad_groupi_g4363(csa_tree_add_107_22_pad_groupi_n_1358 ,csa_tree_add_107_22_pad_groupi_n_1328 ,csa_tree_add_107_22_pad_groupi_n_1320);
  nor csa_tree_add_107_22_pad_groupi_g4364(csa_tree_add_107_22_pad_groupi_n_1357 ,csa_tree_add_107_22_pad_groupi_n_1333 ,csa_tree_add_107_22_pad_groupi_n_1322);
  or csa_tree_add_107_22_pad_groupi_g4365(csa_tree_add_107_22_pad_groupi_n_1356 ,csa_tree_add_107_22_pad_groupi_n_1278 ,csa_tree_add_107_22_pad_groupi_n_1312);
  nor csa_tree_add_107_22_pad_groupi_g4366(csa_tree_add_107_22_pad_groupi_n_1355 ,csa_tree_add_107_22_pad_groupi_n_1299 ,csa_tree_add_107_22_pad_groupi_n_1330);
  or csa_tree_add_107_22_pad_groupi_g4367(csa_tree_add_107_22_pad_groupi_n_1354 ,csa_tree_add_107_22_pad_groupi_n_1294 ,csa_tree_add_107_22_pad_groupi_n_1332);
  nor csa_tree_add_107_22_pad_groupi_g4368(csa_tree_add_107_22_pad_groupi_n_1353 ,csa_tree_add_107_22_pad_groupi_n_1295 ,csa_tree_add_107_22_pad_groupi_n_1331);
  and csa_tree_add_107_22_pad_groupi_g4369(csa_tree_add_107_22_pad_groupi_n_1368 ,csa_tree_add_107_22_pad_groupi_n_1243 ,csa_tree_add_107_22_pad_groupi_n_1324);
  or csa_tree_add_107_22_pad_groupi_g4370(csa_tree_add_107_22_pad_groupi_n_1366 ,csa_tree_add_107_22_pad_groupi_n_1185 ,csa_tree_add_107_22_pad_groupi_n_1327);
  not csa_tree_add_107_22_pad_groupi_g4371(csa_tree_add_107_22_pad_groupi_n_1352 ,csa_tree_add_107_22_pad_groupi_n_1351);
  not csa_tree_add_107_22_pad_groupi_g4373(csa_tree_add_107_22_pad_groupi_n_1349 ,csa_tree_add_107_22_pad_groupi_n_1348);
  not csa_tree_add_107_22_pad_groupi_g4374(csa_tree_add_107_22_pad_groupi_n_1347 ,csa_tree_add_107_22_pad_groupi_n_1346);
  or csa_tree_add_107_22_pad_groupi_g4375(csa_tree_add_107_22_pad_groupi_n_1344 ,csa_tree_add_107_22_pad_groupi_n_1223 ,csa_tree_add_107_22_pad_groupi_n_1317);
  and csa_tree_add_107_22_pad_groupi_g4376(csa_tree_add_107_22_pad_groupi_n_1343 ,csa_tree_add_107_22_pad_groupi_n_1228 ,csa_tree_add_107_22_pad_groupi_n_1314);
  and csa_tree_add_107_22_pad_groupi_g4377(csa_tree_add_107_22_pad_groupi_n_1342 ,csa_tree_add_107_22_pad_groupi_n_1278 ,csa_tree_add_107_22_pad_groupi_n_1312);
  and csa_tree_add_107_22_pad_groupi_g4378(csa_tree_add_107_22_pad_groupi_n_1341 ,csa_tree_add_107_22_pad_groupi_n_1226 ,csa_tree_add_107_22_pad_groupi_n_1313);
  and csa_tree_add_107_22_pad_groupi_g4379(csa_tree_add_107_22_pad_groupi_n_1340 ,csa_tree_add_107_22_pad_groupi_n_1299 ,csa_tree_add_107_22_pad_groupi_n_1330);
  and csa_tree_add_107_22_pad_groupi_g4380(csa_tree_add_107_22_pad_groupi_n_1339 ,csa_tree_add_107_22_pad_groupi_n_1231 ,csa_tree_add_107_22_pad_groupi_n_1315);
  xnor csa_tree_add_107_22_pad_groupi_g4381(csa_tree_add_107_22_pad_groupi_n_1338 ,csa_tree_add_107_22_pad_groupi_n_1201 ,csa_tree_add_107_22_pad_groupi_n_1279);
  xnor csa_tree_add_107_22_pad_groupi_g4382(csa_tree_add_107_22_pad_groupi_n_1351 ,csa_tree_add_107_22_pad_groupi_n_1281 ,csa_tree_add_107_22_pad_groupi_n_1211);
  xor csa_tree_add_107_22_pad_groupi_g4383(csa_tree_add_107_22_pad_groupi_n_1337 ,csa_tree_add_107_22_pad_groupi_n_1278 ,csa_tree_add_107_22_pad_groupi_n_1305);
  xnor csa_tree_add_107_22_pad_groupi_g4384(csa_tree_add_107_22_pad_groupi_n_1336 ,csa_tree_add_107_22_pad_groupi_n_1075 ,csa_tree_add_107_22_pad_groupi_n_1274);
  xnor csa_tree_add_107_22_pad_groupi_g4385(csa_tree_add_107_22_pad_groupi_n_1335 ,csa_tree_add_107_22_pad_groupi_n_1235 ,csa_tree_add_107_22_pad_groupi_n_1296);
  xnor csa_tree_add_107_22_pad_groupi_g4386(csa_tree_add_107_22_pad_groupi_n_1350 ,csa_tree_add_107_22_pad_groupi_n_1264 ,csa_tree_add_107_22_pad_groupi_n_1272);
  xnor csa_tree_add_107_22_pad_groupi_g4387(csa_tree_add_107_22_pad_groupi_n_1348 ,csa_tree_add_107_22_pad_groupi_n_1282 ,csa_tree_add_107_22_pad_groupi_n_1269);
  xnor csa_tree_add_107_22_pad_groupi_g4388(csa_tree_add_107_22_pad_groupi_n_1346 ,csa_tree_add_107_22_pad_groupi_n_1263 ,csa_tree_add_107_22_pad_groupi_n_1275);
  or csa_tree_add_107_22_pad_groupi_g4389(csa_tree_add_107_22_pad_groupi_n_1345 ,csa_tree_add_107_22_pad_groupi_n_1277 ,csa_tree_add_107_22_pad_groupi_n_1325);
  not csa_tree_add_107_22_pad_groupi_g4390(csa_tree_add_107_22_pad_groupi_n_1332 ,csa_tree_add_107_22_pad_groupi_n_1331);
  nor csa_tree_add_107_22_pad_groupi_g4391(csa_tree_add_107_22_pad_groupi_n_1329 ,csa_tree_add_107_22_pad_groupi_n_1202 ,csa_tree_add_107_22_pad_groupi_n_1279);
  nor csa_tree_add_107_22_pad_groupi_g4392(csa_tree_add_107_22_pad_groupi_n_1328 ,csa_tree_add_107_22_pad_groupi_n_1235 ,csa_tree_add_107_22_pad_groupi_n_1296);
  nor csa_tree_add_107_22_pad_groupi_g4393(csa_tree_add_107_22_pad_groupi_n_1327 ,csa_tree_add_107_22_pad_groupi_n_1184 ,csa_tree_add_107_22_pad_groupi_n_1281);
  nor csa_tree_add_107_22_pad_groupi_g4394(csa_tree_add_107_22_pad_groupi_n_1326 ,csa_tree_add_107_22_pad_groupi_n_1287 ,csa_tree_add_107_22_pad_groupi_n_1288);
  nor csa_tree_add_107_22_pad_groupi_g4395(csa_tree_add_107_22_pad_groupi_n_1325 ,csa_tree_add_107_22_pad_groupi_n_1276 ,csa_tree_add_107_22_pad_groupi_n_1262);
  or csa_tree_add_107_22_pad_groupi_g4396(csa_tree_add_107_22_pad_groupi_n_1324 ,csa_tree_add_107_22_pad_groupi_n_1252 ,csa_tree_add_107_22_pad_groupi_n_1283);
  and csa_tree_add_107_22_pad_groupi_g4397(csa_tree_add_107_22_pad_groupi_n_1323 ,csa_tree_add_107_22_pad_groupi_n_1235 ,csa_tree_add_107_22_pad_groupi_n_1296);
  and csa_tree_add_107_22_pad_groupi_g4398(csa_tree_add_107_22_pad_groupi_n_1322 ,csa_tree_add_107_22_pad_groupi_n_1202 ,csa_tree_add_107_22_pad_groupi_n_1279);
  or csa_tree_add_107_22_pad_groupi_g4399(csa_tree_add_107_22_pad_groupi_n_1334 ,csa_tree_add_107_22_pad_groupi_n_1240 ,csa_tree_add_107_22_pad_groupi_n_1284);
  and csa_tree_add_107_22_pad_groupi_g4400(csa_tree_add_107_22_pad_groupi_n_1333 ,csa_tree_add_107_22_pad_groupi_n_1156 ,csa_tree_add_107_22_pad_groupi_n_1286);
  xnor csa_tree_add_107_22_pad_groupi_g4401(csa_tree_add_107_22_pad_groupi_n_1331 ,csa_tree_add_107_22_pad_groupi_n_1039 ,csa_tree_add_107_22_pad_groupi_n_1216);
  or csa_tree_add_107_22_pad_groupi_g4402(csa_tree_add_107_22_pad_groupi_n_1330 ,csa_tree_add_107_22_pad_groupi_n_1242 ,csa_tree_add_107_22_pad_groupi_n_1289);
  not csa_tree_add_107_22_pad_groupi_g4403(csa_tree_add_107_22_pad_groupi_n_1319 ,csa_tree_add_107_22_pad_groupi_n_1318);
  not csa_tree_add_107_22_pad_groupi_g4404(csa_tree_add_107_22_pad_groupi_n_1312 ,csa_tree_add_107_22_pad_groupi_n_1311);
  xnor csa_tree_add_107_22_pad_groupi_g4405(csa_tree_add_107_22_pad_groupi_n_1321 ,csa_tree_add_107_22_pad_groupi_n_1176 ,csa_tree_add_107_22_pad_groupi_n_1210);
  xnor csa_tree_add_107_22_pad_groupi_g4406(csa_tree_add_107_22_pad_groupi_n_1308 ,csa_tree_add_107_22_pad_groupi_n_1132 ,csa_tree_add_107_22_pad_groupi_n_1233);
  xnor csa_tree_add_107_22_pad_groupi_g4407(csa_tree_add_107_22_pad_groupi_n_1320 ,csa_tree_add_107_22_pad_groupi_n_1084 ,csa_tree_add_107_22_pad_groupi_n_1220);
  xnor csa_tree_add_107_22_pad_groupi_g4408(csa_tree_add_107_22_pad_groupi_n_1318 ,csa_tree_add_107_22_pad_groupi_n_1138 ,csa_tree_add_107_22_pad_groupi_n_1221);
  xnor csa_tree_add_107_22_pad_groupi_g4409(csa_tree_add_107_22_pad_groupi_n_1317 ,csa_tree_add_107_22_pad_groupi_n_1092 ,csa_tree_add_107_22_pad_groupi_n_1213);
  xnor csa_tree_add_107_22_pad_groupi_g4410(csa_tree_add_107_22_pad_groupi_n_1316 ,csa_tree_add_107_22_pad_groupi_n_1088 ,csa_tree_add_107_22_pad_groupi_n_1214);
  xnor csa_tree_add_107_22_pad_groupi_g4411(csa_tree_add_107_22_pad_groupi_n_1315 ,csa_tree_add_107_22_pad_groupi_n_1141 ,csa_tree_add_107_22_pad_groupi_n_1218);
  xnor csa_tree_add_107_22_pad_groupi_g4412(csa_tree_add_107_22_pad_groupi_n_1314 ,csa_tree_add_107_22_pad_groupi_n_1102 ,csa_tree_add_107_22_pad_groupi_n_1217);
  xnor csa_tree_add_107_22_pad_groupi_g4413(csa_tree_add_107_22_pad_groupi_n_1313 ,csa_tree_add_107_22_pad_groupi_n_1107 ,csa_tree_add_107_22_pad_groupi_n_1222);
  xnor csa_tree_add_107_22_pad_groupi_g4414(csa_tree_add_107_22_pad_groupi_n_1311 ,csa_tree_add_107_22_pad_groupi_n_1209 ,csa_tree_add_107_22_pad_groupi_n_1215);
  xnor csa_tree_add_107_22_pad_groupi_g4415(csa_tree_add_107_22_pad_groupi_n_1310 ,csa_tree_add_107_22_pad_groupi_n_1236 ,csa_tree_add_107_22_pad_groupi_n_1212);
  xnor csa_tree_add_107_22_pad_groupi_g4416(csa_tree_add_107_22_pad_groupi_n_1309 ,csa_tree_add_107_22_pad_groupi_n_1175 ,csa_tree_add_107_22_pad_groupi_n_1219);
  not csa_tree_add_107_22_pad_groupi_g4417(csa_tree_add_107_22_pad_groupi_n_1307 ,csa_tree_add_107_22_pad_groupi_n_1306);
  not csa_tree_add_107_22_pad_groupi_g4418(csa_tree_add_107_22_pad_groupi_n_1302 ,csa_tree_add_107_22_pad_groupi_n_1303);
  not csa_tree_add_107_22_pad_groupi_g4419(csa_tree_add_107_22_pad_groupi_n_1300 ,csa_tree_add_107_22_pad_groupi_n_1301);
  not csa_tree_add_107_22_pad_groupi_g4420(csa_tree_add_107_22_pad_groupi_n_1297 ,csa_tree_add_107_22_pad_groupi_n_1298);
  not csa_tree_add_107_22_pad_groupi_g4421(csa_tree_add_107_22_pad_groupi_n_1295 ,csa_tree_add_107_22_pad_groupi_n_1294);
  not csa_tree_add_107_22_pad_groupi_g4422(csa_tree_add_107_22_pad_groupi_n_1292 ,csa_tree_add_107_22_pad_groupi_n_1293);
  not csa_tree_add_107_22_pad_groupi_g4423(csa_tree_add_107_22_pad_groupi_n_1290 ,csa_tree_add_107_22_pad_groupi_n_1291);
  nor csa_tree_add_107_22_pad_groupi_g4424(csa_tree_add_107_22_pad_groupi_n_1289 ,csa_tree_add_107_22_pad_groupi_n_1247 ,csa_tree_add_107_22_pad_groupi_n_1264);
  nor csa_tree_add_107_22_pad_groupi_g4425(csa_tree_add_107_22_pad_groupi_n_1288 ,csa_tree_add_107_22_pad_groupi_n_1048 ,csa_tree_add_107_22_pad_groupi_n_1238);
  nor csa_tree_add_107_22_pad_groupi_g4426(csa_tree_add_107_22_pad_groupi_n_1287 ,csa_tree_add_107_22_pad_groupi_n_1178 ,csa_tree_add_107_22_pad_groupi_n_1251);
  or csa_tree_add_107_22_pad_groupi_g4427(csa_tree_add_107_22_pad_groupi_n_1286 ,csa_tree_add_107_22_pad_groupi_n_1150 ,csa_tree_add_107_22_pad_groupi_n_1237);
  nor csa_tree_add_107_22_pad_groupi_g4428(csa_tree_add_107_22_pad_groupi_n_1285 ,csa_tree_add_107_22_pad_groupi_n_1047 ,csa_tree_add_107_22_pad_groupi_n_1239);
  and csa_tree_add_107_22_pad_groupi_g4429(csa_tree_add_107_22_pad_groupi_n_1284 ,csa_tree_add_107_22_pad_groupi_n_1241 ,csa_tree_add_107_22_pad_groupi_n_1263);
  or csa_tree_add_107_22_pad_groupi_g4430(csa_tree_add_107_22_pad_groupi_n_1306 ,csa_tree_add_107_22_pad_groupi_n_1183 ,csa_tree_add_107_22_pad_groupi_n_1253);
  and csa_tree_add_107_22_pad_groupi_g4431(csa_tree_add_107_22_pad_groupi_n_1305 ,csa_tree_add_107_22_pad_groupi_n_1192 ,csa_tree_add_107_22_pad_groupi_n_1257);
  and csa_tree_add_107_22_pad_groupi_g4432(csa_tree_add_107_22_pad_groupi_n_1304 ,csa_tree_add_107_22_pad_groupi_n_1155 ,csa_tree_add_107_22_pad_groupi_n_1260);
  or csa_tree_add_107_22_pad_groupi_g4433(csa_tree_add_107_22_pad_groupi_n_1303 ,csa_tree_add_107_22_pad_groupi_n_1154 ,csa_tree_add_107_22_pad_groupi_n_1248);
  or csa_tree_add_107_22_pad_groupi_g4434(csa_tree_add_107_22_pad_groupi_n_1301 ,csa_tree_add_107_22_pad_groupi_n_1187 ,csa_tree_add_107_22_pad_groupi_n_1255);
  or csa_tree_add_107_22_pad_groupi_g4435(csa_tree_add_107_22_pad_groupi_n_1299 ,csa_tree_add_107_22_pad_groupi_n_1147 ,csa_tree_add_107_22_pad_groupi_n_1244);
  or csa_tree_add_107_22_pad_groupi_g4436(csa_tree_add_107_22_pad_groupi_n_1298 ,csa_tree_add_107_22_pad_groupi_n_1198 ,csa_tree_add_107_22_pad_groupi_n_1258);
  or csa_tree_add_107_22_pad_groupi_g4437(csa_tree_add_107_22_pad_groupi_n_1296 ,csa_tree_add_107_22_pad_groupi_n_1188 ,csa_tree_add_107_22_pad_groupi_n_1256);
  and csa_tree_add_107_22_pad_groupi_g4438(csa_tree_add_107_22_pad_groupi_n_1294 ,csa_tree_add_107_22_pad_groupi_n_1197 ,csa_tree_add_107_22_pad_groupi_n_1259);
  or csa_tree_add_107_22_pad_groupi_g4439(csa_tree_add_107_22_pad_groupi_n_1293 ,csa_tree_add_107_22_pad_groupi_n_1179 ,csa_tree_add_107_22_pad_groupi_n_1250);
  or csa_tree_add_107_22_pad_groupi_g4440(csa_tree_add_107_22_pad_groupi_n_1291 ,csa_tree_add_107_22_pad_groupi_n_1200 ,csa_tree_add_107_22_pad_groupi_n_1249);
  not csa_tree_add_107_22_pad_groupi_g4441(csa_tree_add_107_22_pad_groupi_n_1283 ,csa_tree_add_107_22_pad_groupi_n_1282);
  nor csa_tree_add_107_22_pad_groupi_g4442(csa_tree_add_107_22_pad_groupi_n_1277 ,csa_tree_add_107_22_pad_groupi_n_1132 ,csa_tree_add_107_22_pad_groupi_n_1234);
  and csa_tree_add_107_22_pad_groupi_g4443(csa_tree_add_107_22_pad_groupi_n_1276 ,csa_tree_add_107_22_pad_groupi_n_1132 ,csa_tree_add_107_22_pad_groupi_n_1234);
  xnor csa_tree_add_107_22_pad_groupi_g4444(csa_tree_add_107_22_pad_groupi_n_1275 ,csa_tree_add_107_22_pad_groupi_n_1207 ,csa_tree_add_107_22_pad_groupi_n_1098);
  nor csa_tree_add_107_22_pad_groupi_g4445(csa_tree_add_107_22_pad_groupi_n_1274 ,csa_tree_add_107_22_pad_groupi_n_1157 ,csa_tree_add_107_22_pad_groupi_n_1229);
  xnor csa_tree_add_107_22_pad_groupi_g4446(csa_tree_add_107_22_pad_groupi_n_1273 ,csa_tree_add_107_22_pad_groupi_n_1163 ,csa_tree_add_107_22_pad_groupi_n_1166);
  xnor csa_tree_add_107_22_pad_groupi_g4447(csa_tree_add_107_22_pad_groupi_n_1272 ,csa_tree_add_107_22_pad_groupi_n_1099 ,csa_tree_add_107_22_pad_groupi_n_1169);
  xnor csa_tree_add_107_22_pad_groupi_g4448(csa_tree_add_107_22_pad_groupi_n_1271 ,csa_tree_add_107_22_pad_groupi_n_1204 ,csa_tree_add_107_22_pad_groupi_n_1160);
  xnor csa_tree_add_107_22_pad_groupi_g4449(csa_tree_add_107_22_pad_groupi_n_1270 ,csa_tree_add_107_22_pad_groupi_n_1208 ,csa_tree_add_107_22_pad_groupi_n_1174);
  xnor csa_tree_add_107_22_pad_groupi_g4450(csa_tree_add_107_22_pad_groupi_n_1269 ,csa_tree_add_107_22_pad_groupi_n_1206 ,csa_tree_add_107_22_pad_groupi_n_1171);
  xnor csa_tree_add_107_22_pad_groupi_g4451(csa_tree_add_107_22_pad_groupi_n_1268 ,csa_tree_add_107_22_pad_groupi_n_1164 ,csa_tree_add_107_22_pad_groupi_n_1167);
  xnor csa_tree_add_107_22_pad_groupi_g4452(csa_tree_add_107_22_pad_groupi_n_1267 ,csa_tree_add_107_22_pad_groupi_n_1173 ,csa_tree_add_107_22_pad_groupi_n_1172);
  xnor csa_tree_add_107_22_pad_groupi_g4453(csa_tree_add_107_22_pad_groupi_n_1266 ,csa_tree_add_107_22_pad_groupi_n_1161 ,csa_tree_add_107_22_pad_groupi_n_1168);
  xnor csa_tree_add_107_22_pad_groupi_g4454(csa_tree_add_107_22_pad_groupi_n_1282 ,csa_tree_add_107_22_pad_groupi_n_1106 ,csa_tree_add_107_22_pad_groupi_n_1143);
  xnor csa_tree_add_107_22_pad_groupi_g4455(csa_tree_add_107_22_pad_groupi_n_1281 ,csa_tree_add_107_22_pad_groupi_n_1080 ,csa_tree_add_107_22_pad_groupi_n_1145);
  xnor csa_tree_add_107_22_pad_groupi_g4456(csa_tree_add_107_22_pad_groupi_n_1280 ,csa_tree_add_107_22_pad_groupi_n_1103 ,csa_tree_add_107_22_pad_groupi_n_1146);
  xnor csa_tree_add_107_22_pad_groupi_g4457(csa_tree_add_107_22_pad_groupi_n_1279 ,csa_tree_add_107_22_pad_groupi_n_1101 ,csa_tree_add_107_22_pad_groupi_n_1142);
  xnor csa_tree_add_107_22_pad_groupi_g4458(csa_tree_add_107_22_pad_groupi_n_1278 ,csa_tree_add_107_22_pad_groupi_n_1105 ,csa_tree_add_107_22_pad_groupi_n_1144);
  or csa_tree_add_107_22_pad_groupi_g4459(csa_tree_add_107_22_pad_groupi_n_1260 ,csa_tree_add_107_22_pad_groupi_n_1104 ,csa_tree_add_107_22_pad_groupi_n_1151);
  or csa_tree_add_107_22_pad_groupi_g4460(csa_tree_add_107_22_pad_groupi_n_1259 ,csa_tree_add_107_22_pad_groupi_n_1209 ,csa_tree_add_107_22_pad_groupi_n_1193);
  nor csa_tree_add_107_22_pad_groupi_g4461(csa_tree_add_107_22_pad_groupi_n_1258 ,csa_tree_add_107_22_pad_groupi_n_1074 ,csa_tree_add_107_22_pad_groupi_n_1195);
  or csa_tree_add_107_22_pad_groupi_g4462(csa_tree_add_107_22_pad_groupi_n_1257 ,csa_tree_add_107_22_pad_groupi_n_1072 ,csa_tree_add_107_22_pad_groupi_n_1190);
  nor csa_tree_add_107_22_pad_groupi_g4463(csa_tree_add_107_22_pad_groupi_n_1256 ,csa_tree_add_107_22_pad_groupi_n_1067 ,csa_tree_add_107_22_pad_groupi_n_1186);
  and csa_tree_add_107_22_pad_groupi_g4464(csa_tree_add_107_22_pad_groupi_n_1255 ,csa_tree_add_107_22_pad_groupi_n_1141 ,csa_tree_add_107_22_pad_groupi_n_1189);
  or csa_tree_add_107_22_pad_groupi_g4465(csa_tree_add_107_22_pad_groupi_n_1254 ,csa_tree_add_107_22_pad_groupi_n_1203 ,csa_tree_add_107_22_pad_groupi_n_1159);
  and csa_tree_add_107_22_pad_groupi_g4466(csa_tree_add_107_22_pad_groupi_n_1253 ,csa_tree_add_107_22_pad_groupi_n_1181 ,csa_tree_add_107_22_pad_groupi_n_1176);
  nor csa_tree_add_107_22_pad_groupi_g4467(csa_tree_add_107_22_pad_groupi_n_1252 ,csa_tree_add_107_22_pad_groupi_n_1206 ,csa_tree_add_107_22_pad_groupi_n_1171);
  nor csa_tree_add_107_22_pad_groupi_g4468(csa_tree_add_107_22_pad_groupi_n_1251 ,csa_tree_add_107_22_pad_groupi_n_1177 ,csa_tree_add_107_22_pad_groupi_n_1191);
  and csa_tree_add_107_22_pad_groupi_g4469(csa_tree_add_107_22_pad_groupi_n_1250 ,csa_tree_add_107_22_pad_groupi_n_1102 ,csa_tree_add_107_22_pad_groupi_n_1194);
  and csa_tree_add_107_22_pad_groupi_g4470(csa_tree_add_107_22_pad_groupi_n_1249 ,csa_tree_add_107_22_pad_groupi_n_1107 ,csa_tree_add_107_22_pad_groupi_n_1158);
  nor csa_tree_add_107_22_pad_groupi_g4471(csa_tree_add_107_22_pad_groupi_n_1248 ,csa_tree_add_107_22_pad_groupi_n_1042 ,csa_tree_add_107_22_pad_groupi_n_1153);
  nor csa_tree_add_107_22_pad_groupi_g4472(csa_tree_add_107_22_pad_groupi_n_1247 ,csa_tree_add_107_22_pad_groupi_n_1099 ,csa_tree_add_107_22_pad_groupi_n_1169);
  and csa_tree_add_107_22_pad_groupi_g4473(csa_tree_add_107_22_pad_groupi_n_1246 ,csa_tree_add_107_22_pad_groupi_n_1164 ,csa_tree_add_107_22_pad_groupi_n_1167);
  nor csa_tree_add_107_22_pad_groupi_g4474(csa_tree_add_107_22_pad_groupi_n_1245 ,csa_tree_add_107_22_pad_groupi_n_1164 ,csa_tree_add_107_22_pad_groupi_n_1167);
  nor csa_tree_add_107_22_pad_groupi_g4475(csa_tree_add_107_22_pad_groupi_n_1244 ,csa_tree_add_107_22_pad_groupi_n_1039 ,csa_tree_add_107_22_pad_groupi_n_1148);
  or csa_tree_add_107_22_pad_groupi_g4476(csa_tree_add_107_22_pad_groupi_n_1243 ,csa_tree_add_107_22_pad_groupi_n_1205 ,csa_tree_add_107_22_pad_groupi_n_1170);
  and csa_tree_add_107_22_pad_groupi_g4477(csa_tree_add_107_22_pad_groupi_n_1242 ,csa_tree_add_107_22_pad_groupi_n_1099 ,csa_tree_add_107_22_pad_groupi_n_1169);
  or csa_tree_add_107_22_pad_groupi_g4478(csa_tree_add_107_22_pad_groupi_n_1241 ,csa_tree_add_107_22_pad_groupi_n_1207 ,csa_tree_add_107_22_pad_groupi_n_1098);
  and csa_tree_add_107_22_pad_groupi_g4479(csa_tree_add_107_22_pad_groupi_n_1240 ,csa_tree_add_107_22_pad_groupi_n_1207 ,csa_tree_add_107_22_pad_groupi_n_1098);
  or csa_tree_add_107_22_pad_groupi_g4480(csa_tree_add_107_22_pad_groupi_n_1265 ,csa_tree_add_107_22_pad_groupi_n_1051 ,csa_tree_add_107_22_pad_groupi_n_1180);
  and csa_tree_add_107_22_pad_groupi_g4481(csa_tree_add_107_22_pad_groupi_n_1264 ,csa_tree_add_107_22_pad_groupi_n_1115 ,csa_tree_add_107_22_pad_groupi_n_1199);
  or csa_tree_add_107_22_pad_groupi_g4482(csa_tree_add_107_22_pad_groupi_n_1263 ,csa_tree_add_107_22_pad_groupi_n_1123 ,csa_tree_add_107_22_pad_groupi_n_1182);
  and csa_tree_add_107_22_pad_groupi_g4483(csa_tree_add_107_22_pad_groupi_n_1262 ,csa_tree_add_107_22_pad_groupi_n_1114 ,csa_tree_add_107_22_pad_groupi_n_1149);
  or csa_tree_add_107_22_pad_groupi_g4484(csa_tree_add_107_22_pad_groupi_n_1261 ,csa_tree_add_107_22_pad_groupi_n_1124 ,csa_tree_add_107_22_pad_groupi_n_1196);
  not csa_tree_add_107_22_pad_groupi_g4485(csa_tree_add_107_22_pad_groupi_n_1239 ,csa_tree_add_107_22_pad_groupi_n_1238);
  not csa_tree_add_107_22_pad_groupi_g4486(csa_tree_add_107_22_pad_groupi_n_1237 ,csa_tree_add_107_22_pad_groupi_n_1236);
  not csa_tree_add_107_22_pad_groupi_g4487(csa_tree_add_107_22_pad_groupi_n_1234 ,csa_tree_add_107_22_pad_groupi_n_1233);
  and csa_tree_add_107_22_pad_groupi_g4488(csa_tree_add_107_22_pad_groupi_n_1232 ,csa_tree_add_107_22_pad_groupi_n_1208 ,csa_tree_add_107_22_pad_groupi_n_1174);
  or csa_tree_add_107_22_pad_groupi_g4489(csa_tree_add_107_22_pad_groupi_n_1231 ,csa_tree_add_107_22_pad_groupi_n_1208 ,csa_tree_add_107_22_pad_groupi_n_1174);
  and csa_tree_add_107_22_pad_groupi_g4490(csa_tree_add_107_22_pad_groupi_n_1230 ,csa_tree_add_107_22_pad_groupi_n_1173 ,csa_tree_add_107_22_pad_groupi_n_1172);
  nor csa_tree_add_107_22_pad_groupi_g4491(csa_tree_add_107_22_pad_groupi_n_1229 ,csa_tree_add_107_22_pad_groupi_n_1152 ,csa_tree_add_107_22_pad_groupi_n_1175);
  or csa_tree_add_107_22_pad_groupi_g4492(csa_tree_add_107_22_pad_groupi_n_1228 ,csa_tree_add_107_22_pad_groupi_n_1173 ,csa_tree_add_107_22_pad_groupi_n_1172);
  and csa_tree_add_107_22_pad_groupi_g4493(csa_tree_add_107_22_pad_groupi_n_1227 ,csa_tree_add_107_22_pad_groupi_n_1161 ,csa_tree_add_107_22_pad_groupi_n_1168);
  or csa_tree_add_107_22_pad_groupi_g4494(csa_tree_add_107_22_pad_groupi_n_1226 ,csa_tree_add_107_22_pad_groupi_n_1161 ,csa_tree_add_107_22_pad_groupi_n_1168);
  or csa_tree_add_107_22_pad_groupi_g4495(csa_tree_add_107_22_pad_groupi_n_1225 ,csa_tree_add_107_22_pad_groupi_n_1162 ,csa_tree_add_107_22_pad_groupi_n_1165);
  nor csa_tree_add_107_22_pad_groupi_g4496(csa_tree_add_107_22_pad_groupi_n_1224 ,csa_tree_add_107_22_pad_groupi_n_1204 ,csa_tree_add_107_22_pad_groupi_n_1160);
  nor csa_tree_add_107_22_pad_groupi_g4497(csa_tree_add_107_22_pad_groupi_n_1223 ,csa_tree_add_107_22_pad_groupi_n_1163 ,csa_tree_add_107_22_pad_groupi_n_1166);
  xnor csa_tree_add_107_22_pad_groupi_g4498(csa_tree_add_107_22_pad_groupi_n_1222 ,csa_tree_add_107_22_pad_groupi_n_1035 ,csa_tree_add_107_22_pad_groupi_n_1094);
  xnor csa_tree_add_107_22_pad_groupi_g4499(csa_tree_add_107_22_pad_groupi_n_1221 ,csa_tree_add_107_22_pad_groupi_n_1100 ,csa_tree_add_107_22_pad_groupi_n_1074);
  xnor csa_tree_add_107_22_pad_groupi_g4500(csa_tree_add_107_22_pad_groupi_n_1220 ,csa_tree_add_107_22_pad_groupi_n_1072 ,csa_tree_add_107_22_pad_groupi_n_1090);
  xnor csa_tree_add_107_22_pad_groupi_g4501(csa_tree_add_107_22_pad_groupi_n_1219 ,csa_tree_add_107_22_pad_groupi_n_1016 ,csa_tree_add_107_22_pad_groupi_n_1097);
  xnor csa_tree_add_107_22_pad_groupi_g4502(csa_tree_add_107_22_pad_groupi_n_1218 ,csa_tree_add_107_22_pad_groupi_n_1056 ,csa_tree_add_107_22_pad_groupi_n_3);
  xnor csa_tree_add_107_22_pad_groupi_g4503(csa_tree_add_107_22_pad_groupi_n_1238 ,csa_tree_add_107_22_pad_groupi_n_1140 ,csa_tree_add_107_22_pad_groupi_n_1076);
  xnor csa_tree_add_107_22_pad_groupi_g4504(csa_tree_add_107_22_pad_groupi_n_1217 ,csa_tree_add_107_22_pad_groupi_n_1055 ,csa_tree_add_107_22_pad_groupi_n_1095);
  xnor csa_tree_add_107_22_pad_groupi_g4505(csa_tree_add_107_22_pad_groupi_n_1216 ,csa_tree_add_107_22_pad_groupi_n_1036 ,csa_tree_add_107_22_pad_groupi_n_1087);
  xnor csa_tree_add_107_22_pad_groupi_g4506(csa_tree_add_107_22_pad_groupi_n_1215 ,csa_tree_add_107_22_pad_groupi_n_1137 ,csa_tree_add_107_22_pad_groupi_n_1086);
  xnor csa_tree_add_107_22_pad_groupi_g4507(csa_tree_add_107_22_pad_groupi_n_1214 ,csa_tree_add_107_22_pad_groupi_n_1042 ,csa_tree_add_107_22_pad_groupi_n_1093);
  xnor csa_tree_add_107_22_pad_groupi_g4508(csa_tree_add_107_22_pad_groupi_n_1213 ,csa_tree_add_107_22_pad_groupi_n_1034 ,csa_tree_add_107_22_pad_groupi_n_1104);
  xnor csa_tree_add_107_22_pad_groupi_g4509(csa_tree_add_107_22_pad_groupi_n_1212 ,csa_tree_add_107_22_pad_groupi_n_1131 ,csa_tree_add_107_22_pad_groupi_n_1082);
  xnor csa_tree_add_107_22_pad_groupi_g4510(csa_tree_add_107_22_pad_groupi_n_1211 ,csa_tree_add_107_22_pad_groupi_n_1134 ,csa_tree_add_107_22_pad_groupi_n_1135);
  xnor csa_tree_add_107_22_pad_groupi_g4511(csa_tree_add_107_22_pad_groupi_n_1210 ,csa_tree_add_107_22_pad_groupi_n_1062 ,csa_tree_add_107_22_pad_groupi_n_1133);
  xnor csa_tree_add_107_22_pad_groupi_g4512(csa_tree_add_107_22_pad_groupi_n_1236 ,csa_tree_add_107_22_pad_groupi_n_1043 ,csa_tree_add_107_22_pad_groupi_n_1078);
  xnor csa_tree_add_107_22_pad_groupi_g4513(csa_tree_add_107_22_pad_groupi_n_1235 ,csa_tree_add_107_22_pad_groupi_n_1070 ,csa_tree_add_107_22_pad_groupi_n_1079);
  xnor csa_tree_add_107_22_pad_groupi_g4514(csa_tree_add_107_22_pad_groupi_n_1233 ,csa_tree_add_107_22_pad_groupi_n_976 ,csa_tree_add_107_22_pad_groupi_n_1077);
  not csa_tree_add_107_22_pad_groupi_g4515(csa_tree_add_107_22_pad_groupi_n_1206 ,csa_tree_add_107_22_pad_groupi_n_1205);
  not csa_tree_add_107_22_pad_groupi_g4516(csa_tree_add_107_22_pad_groupi_n_1204 ,csa_tree_add_107_22_pad_groupi_n_1203);
  not csa_tree_add_107_22_pad_groupi_g4517(csa_tree_add_107_22_pad_groupi_n_1202 ,csa_tree_add_107_22_pad_groupi_n_1201);
  and csa_tree_add_107_22_pad_groupi_g4518(csa_tree_add_107_22_pad_groupi_n_1200 ,csa_tree_add_107_22_pad_groupi_n_1035 ,csa_tree_add_107_22_pad_groupi_n_1094);
  or csa_tree_add_107_22_pad_groupi_g4519(csa_tree_add_107_22_pad_groupi_n_1199 ,csa_tree_add_107_22_pad_groupi_n_1105 ,csa_tree_add_107_22_pad_groupi_n_1128);
  nor csa_tree_add_107_22_pad_groupi_g4520(csa_tree_add_107_22_pad_groupi_n_1198 ,csa_tree_add_107_22_pad_groupi_n_1100 ,csa_tree_add_107_22_pad_groupi_n_1139);
  or csa_tree_add_107_22_pad_groupi_g4521(csa_tree_add_107_22_pad_groupi_n_1197 ,csa_tree_add_107_22_pad_groupi_n_1136 ,csa_tree_add_107_22_pad_groupi_n_1086);
  and csa_tree_add_107_22_pad_groupi_g4522(csa_tree_add_107_22_pad_groupi_n_1196 ,csa_tree_add_107_22_pad_groupi_n_1118 ,csa_tree_add_107_22_pad_groupi_n_1103);
  and csa_tree_add_107_22_pad_groupi_g4523(csa_tree_add_107_22_pad_groupi_n_1195 ,csa_tree_add_107_22_pad_groupi_n_1100 ,csa_tree_add_107_22_pad_groupi_n_1139);
  or csa_tree_add_107_22_pad_groupi_g4524(csa_tree_add_107_22_pad_groupi_n_1194 ,csa_tree_add_107_22_pad_groupi_n_1055 ,csa_tree_add_107_22_pad_groupi_n_1095);
  nor csa_tree_add_107_22_pad_groupi_g4525(csa_tree_add_107_22_pad_groupi_n_1193 ,csa_tree_add_107_22_pad_groupi_n_1137 ,csa_tree_add_107_22_pad_groupi_n_1085);
  or csa_tree_add_107_22_pad_groupi_g4526(csa_tree_add_107_22_pad_groupi_n_1192 ,csa_tree_add_107_22_pad_groupi_n_1083 ,csa_tree_add_107_22_pad_groupi_n_1089);
  nor csa_tree_add_107_22_pad_groupi_g4527(csa_tree_add_107_22_pad_groupi_n_1191 ,csa_tree_add_107_22_pad_groupi_n_1022 ,csa_tree_add_107_22_pad_groupi_n_1109);
  nor csa_tree_add_107_22_pad_groupi_g4528(csa_tree_add_107_22_pad_groupi_n_1190 ,csa_tree_add_107_22_pad_groupi_n_1084 ,csa_tree_add_107_22_pad_groupi_n_1090);
  or csa_tree_add_107_22_pad_groupi_g4529(csa_tree_add_107_22_pad_groupi_n_1189 ,csa_tree_add_107_22_pad_groupi_n_1056 ,csa_tree_add_107_22_pad_groupi_n_3);
  nor csa_tree_add_107_22_pad_groupi_g4530(csa_tree_add_107_22_pad_groupi_n_1188 ,csa_tree_add_107_22_pad_groupi_n_1019 ,csa_tree_add_107_22_pad_groupi_n_1080);
  and csa_tree_add_107_22_pad_groupi_g4531(csa_tree_add_107_22_pad_groupi_n_1187 ,csa_tree_add_107_22_pad_groupi_n_1056 ,csa_tree_add_107_22_pad_groupi_n_3);
  and csa_tree_add_107_22_pad_groupi_g4532(csa_tree_add_107_22_pad_groupi_n_1186 ,csa_tree_add_107_22_pad_groupi_n_1019 ,csa_tree_add_107_22_pad_groupi_n_1080);
  and csa_tree_add_107_22_pad_groupi_g4533(csa_tree_add_107_22_pad_groupi_n_1185 ,csa_tree_add_107_22_pad_groupi_n_1134 ,csa_tree_add_107_22_pad_groupi_n_1135);
  nor csa_tree_add_107_22_pad_groupi_g4534(csa_tree_add_107_22_pad_groupi_n_1184 ,csa_tree_add_107_22_pad_groupi_n_1134 ,csa_tree_add_107_22_pad_groupi_n_1135);
  and csa_tree_add_107_22_pad_groupi_g4535(csa_tree_add_107_22_pad_groupi_n_1183 ,csa_tree_add_107_22_pad_groupi_n_1062 ,csa_tree_add_107_22_pad_groupi_n_1133);
  and csa_tree_add_107_22_pad_groupi_g4536(csa_tree_add_107_22_pad_groupi_n_1182 ,csa_tree_add_107_22_pad_groupi_n_1120 ,csa_tree_add_107_22_pad_groupi_n_1106);
  or csa_tree_add_107_22_pad_groupi_g4537(csa_tree_add_107_22_pad_groupi_n_1181 ,csa_tree_add_107_22_pad_groupi_n_1062 ,csa_tree_add_107_22_pad_groupi_n_1133);
  and csa_tree_add_107_22_pad_groupi_g4538(csa_tree_add_107_22_pad_groupi_n_1180 ,csa_tree_add_107_22_pad_groupi_n_1050 ,csa_tree_add_107_22_pad_groupi_n_1140);
  and csa_tree_add_107_22_pad_groupi_g4539(csa_tree_add_107_22_pad_groupi_n_1179 ,csa_tree_add_107_22_pad_groupi_n_1055 ,csa_tree_add_107_22_pad_groupi_n_1095);
  nor csa_tree_add_107_22_pad_groupi_g4540(csa_tree_add_107_22_pad_groupi_n_1178 ,csa_tree_add_107_22_pad_groupi_n_1023 ,csa_tree_add_107_22_pad_groupi_n_1108);
  nor csa_tree_add_107_22_pad_groupi_g4541(csa_tree_add_107_22_pad_groupi_n_1177 ,csa_tree_add_107_22_pad_groupi_n_1031 ,csa_tree_add_107_22_pad_groupi_n_1119);
  and csa_tree_add_107_22_pad_groupi_g4542(csa_tree_add_107_22_pad_groupi_n_1209 ,csa_tree_add_107_22_pad_groupi_n_1054 ,csa_tree_add_107_22_pad_groupi_n_1127);
  or csa_tree_add_107_22_pad_groupi_g4543(csa_tree_add_107_22_pad_groupi_n_1208 ,csa_tree_add_107_22_pad_groupi_n_901 ,csa_tree_add_107_22_pad_groupi_n_1122);
  or csa_tree_add_107_22_pad_groupi_g4544(csa_tree_add_107_22_pad_groupi_n_1207 ,csa_tree_add_107_22_pad_groupi_n_914 ,csa_tree_add_107_22_pad_groupi_n_1125);
  and csa_tree_add_107_22_pad_groupi_g4545(csa_tree_add_107_22_pad_groupi_n_1205 ,csa_tree_add_107_22_pad_groupi_n_884 ,csa_tree_add_107_22_pad_groupi_n_1116);
  and csa_tree_add_107_22_pad_groupi_g4546(csa_tree_add_107_22_pad_groupi_n_1203 ,csa_tree_add_107_22_pad_groupi_n_921 ,csa_tree_add_107_22_pad_groupi_n_1126);
  or csa_tree_add_107_22_pad_groupi_g4547(csa_tree_add_107_22_pad_groupi_n_1201 ,csa_tree_add_107_22_pad_groupi_n_1049 ,csa_tree_add_107_22_pad_groupi_n_1117);
  not csa_tree_add_107_22_pad_groupi_g4548(csa_tree_add_107_22_pad_groupi_n_1170 ,csa_tree_add_107_22_pad_groupi_n_1171);
  not csa_tree_add_107_22_pad_groupi_g4549(csa_tree_add_107_22_pad_groupi_n_1166 ,csa_tree_add_107_22_pad_groupi_n_1165);
  not csa_tree_add_107_22_pad_groupi_g4550(csa_tree_add_107_22_pad_groupi_n_1163 ,csa_tree_add_107_22_pad_groupi_n_1162);
  not csa_tree_add_107_22_pad_groupi_g4551(csa_tree_add_107_22_pad_groupi_n_1160 ,csa_tree_add_107_22_pad_groupi_n_1159);
  or csa_tree_add_107_22_pad_groupi_g4552(csa_tree_add_107_22_pad_groupi_n_1158 ,csa_tree_add_107_22_pad_groupi_n_1035 ,csa_tree_add_107_22_pad_groupi_n_1094);
  and csa_tree_add_107_22_pad_groupi_g4553(csa_tree_add_107_22_pad_groupi_n_1157 ,csa_tree_add_107_22_pad_groupi_n_1015 ,csa_tree_add_107_22_pad_groupi_n_1097);
  or csa_tree_add_107_22_pad_groupi_g4554(csa_tree_add_107_22_pad_groupi_n_1156 ,csa_tree_add_107_22_pad_groupi_n_1130 ,csa_tree_add_107_22_pad_groupi_n_1081);
  or csa_tree_add_107_22_pad_groupi_g4555(csa_tree_add_107_22_pad_groupi_n_1155 ,csa_tree_add_107_22_pad_groupi_n_1033 ,csa_tree_add_107_22_pad_groupi_n_1091);
  and csa_tree_add_107_22_pad_groupi_g4556(csa_tree_add_107_22_pad_groupi_n_1154 ,csa_tree_add_107_22_pad_groupi_n_1093 ,csa_tree_add_107_22_pad_groupi_n_1088);
  nor csa_tree_add_107_22_pad_groupi_g4557(csa_tree_add_107_22_pad_groupi_n_1153 ,csa_tree_add_107_22_pad_groupi_n_1093 ,csa_tree_add_107_22_pad_groupi_n_1088);
  and csa_tree_add_107_22_pad_groupi_g4558(csa_tree_add_107_22_pad_groupi_n_1152 ,csa_tree_add_107_22_pad_groupi_n_1016 ,csa_tree_add_107_22_pad_groupi_n_1096);
  nor csa_tree_add_107_22_pad_groupi_g4559(csa_tree_add_107_22_pad_groupi_n_1151 ,csa_tree_add_107_22_pad_groupi_n_1034 ,csa_tree_add_107_22_pad_groupi_n_1092);
  nor csa_tree_add_107_22_pad_groupi_g4560(csa_tree_add_107_22_pad_groupi_n_1150 ,csa_tree_add_107_22_pad_groupi_n_1131 ,csa_tree_add_107_22_pad_groupi_n_1082);
  or csa_tree_add_107_22_pad_groupi_g4561(csa_tree_add_107_22_pad_groupi_n_1149 ,csa_tree_add_107_22_pad_groupi_n_1110 ,csa_tree_add_107_22_pad_groupi_n_1101);
  and csa_tree_add_107_22_pad_groupi_g4562(csa_tree_add_107_22_pad_groupi_n_1148 ,csa_tree_add_107_22_pad_groupi_n_1037 ,csa_tree_add_107_22_pad_groupi_n_1087);
  nor csa_tree_add_107_22_pad_groupi_g4563(csa_tree_add_107_22_pad_groupi_n_1147 ,csa_tree_add_107_22_pad_groupi_n_1037 ,csa_tree_add_107_22_pad_groupi_n_1087);
  xnor csa_tree_add_107_22_pad_groupi_g4564(csa_tree_add_107_22_pad_groupi_n_1146 ,csa_tree_add_107_22_pad_groupi_n_1010 ,csa_tree_add_107_22_pad_groupi_n_1064);
  xnor csa_tree_add_107_22_pad_groupi_g4565(csa_tree_add_107_22_pad_groupi_n_1145 ,csa_tree_add_107_22_pad_groupi_n_1067 ,csa_tree_add_107_22_pad_groupi_n_1019);
  xnor csa_tree_add_107_22_pad_groupi_g4566(csa_tree_add_107_22_pad_groupi_n_1144 ,csa_tree_add_107_22_pad_groupi_n_1058 ,csa_tree_add_107_22_pad_groupi_n_1061);
  xnor csa_tree_add_107_22_pad_groupi_g4567(csa_tree_add_107_22_pad_groupi_n_1143 ,csa_tree_add_107_22_pad_groupi_n_1011 ,csa_tree_add_107_22_pad_groupi_n_1059);
  xnor csa_tree_add_107_22_pad_groupi_g4568(csa_tree_add_107_22_pad_groupi_n_1142 ,csa_tree_add_107_22_pad_groupi_n_1018 ,csa_tree_add_107_22_pad_groupi_n_1066);
  xnor csa_tree_add_107_22_pad_groupi_g4569(csa_tree_add_107_22_pad_groupi_n_1176 ,csa_tree_add_107_22_pad_groupi_n_1020 ,csa_tree_add_107_22_pad_groupi_n_1025);
  and csa_tree_add_107_22_pad_groupi_g4570(csa_tree_add_107_22_pad_groupi_n_1175 ,csa_tree_add_107_22_pad_groupi_n_1030 ,csa_tree_add_107_22_pad_groupi_n_1111);
  xnor csa_tree_add_107_22_pad_groupi_g4571(csa_tree_add_107_22_pad_groupi_n_1174 ,csa_tree_add_107_22_pad_groupi_n_1068 ,csa_tree_add_107_22_pad_groupi_n_950);
  or csa_tree_add_107_22_pad_groupi_g4572(csa_tree_add_107_22_pad_groupi_n_1173 ,csa_tree_add_107_22_pad_groupi_n_908 ,csa_tree_add_107_22_pad_groupi_n_1121);
  xnor csa_tree_add_107_22_pad_groupi_g4573(csa_tree_add_107_22_pad_groupi_n_1172 ,csa_tree_add_107_22_pad_groupi_n_1045 ,csa_tree_add_107_22_pad_groupi_n_944);
  xnor csa_tree_add_107_22_pad_groupi_g4574(csa_tree_add_107_22_pad_groupi_n_1171 ,csa_tree_add_107_22_pad_groupi_n_1073 ,csa_tree_add_107_22_pad_groupi_n_941);
  xnor csa_tree_add_107_22_pad_groupi_g4575(csa_tree_add_107_22_pad_groupi_n_1169 ,csa_tree_add_107_22_pad_groupi_n_1041 ,csa_tree_add_107_22_pad_groupi_n_974);
  xnor csa_tree_add_107_22_pad_groupi_g4576(csa_tree_add_107_22_pad_groupi_n_1168 ,csa_tree_add_107_22_pad_groupi_n_1044 ,csa_tree_add_107_22_pad_groupi_n_939);
  xnor csa_tree_add_107_22_pad_groupi_g4577(csa_tree_add_107_22_pad_groupi_n_1167 ,csa_tree_add_107_22_pad_groupi_n_1040 ,csa_tree_add_107_22_pad_groupi_n_969);
  xnor csa_tree_add_107_22_pad_groupi_g4578(csa_tree_add_107_22_pad_groupi_n_1165 ,csa_tree_add_107_22_pad_groupi_n_1038 ,csa_tree_add_107_22_pad_groupi_n_970);
  or csa_tree_add_107_22_pad_groupi_g4579(csa_tree_add_107_22_pad_groupi_n_1164 ,csa_tree_add_107_22_pad_groupi_n_858 ,csa_tree_add_107_22_pad_groupi_n_1113);
  and csa_tree_add_107_22_pad_groupi_g4580(csa_tree_add_107_22_pad_groupi_n_1162 ,csa_tree_add_107_22_pad_groupi_n_857 ,csa_tree_add_107_22_pad_groupi_n_1112);
  or csa_tree_add_107_22_pad_groupi_g4581(csa_tree_add_107_22_pad_groupi_n_1161 ,csa_tree_add_107_22_pad_groupi_n_873 ,csa_tree_add_107_22_pad_groupi_n_1129);
  xnor csa_tree_add_107_22_pad_groupi_g4582(csa_tree_add_107_22_pad_groupi_n_1159 ,csa_tree_add_107_22_pad_groupi_n_1046 ,csa_tree_add_107_22_pad_groupi_n_955);
  not csa_tree_add_107_22_pad_groupi_g4583(csa_tree_add_107_22_pad_groupi_n_1139 ,csa_tree_add_107_22_pad_groupi_n_1138);
  not csa_tree_add_107_22_pad_groupi_g4584(csa_tree_add_107_22_pad_groupi_n_1136 ,csa_tree_add_107_22_pad_groupi_n_1137);
  not csa_tree_add_107_22_pad_groupi_g4585(csa_tree_add_107_22_pad_groupi_n_1130 ,csa_tree_add_107_22_pad_groupi_n_1131);
  and csa_tree_add_107_22_pad_groupi_g4586(csa_tree_add_107_22_pad_groupi_n_1129 ,csa_tree_add_107_22_pad_groupi_n_871 ,csa_tree_add_107_22_pad_groupi_n_1040);
  nor csa_tree_add_107_22_pad_groupi_g4587(csa_tree_add_107_22_pad_groupi_n_1128 ,csa_tree_add_107_22_pad_groupi_n_1058 ,csa_tree_add_107_22_pad_groupi_n_1061);
  or csa_tree_add_107_22_pad_groupi_g4588(csa_tree_add_107_22_pad_groupi_n_1127 ,csa_tree_add_107_22_pad_groupi_n_1053 ,csa_tree_add_107_22_pad_groupi_n_1071);
  or csa_tree_add_107_22_pad_groupi_g4589(csa_tree_add_107_22_pad_groupi_n_1126 ,csa_tree_add_107_22_pad_groupi_n_918 ,csa_tree_add_107_22_pad_groupi_n_1069);
  and csa_tree_add_107_22_pad_groupi_g4590(csa_tree_add_107_22_pad_groupi_n_1125 ,csa_tree_add_107_22_pad_groupi_n_932 ,csa_tree_add_107_22_pad_groupi_n_1073);
  nor csa_tree_add_107_22_pad_groupi_g4591(csa_tree_add_107_22_pad_groupi_n_1124 ,csa_tree_add_107_22_pad_groupi_n_1010 ,csa_tree_add_107_22_pad_groupi_n_1063);
  and csa_tree_add_107_22_pad_groupi_g4592(csa_tree_add_107_22_pad_groupi_n_1123 ,csa_tree_add_107_22_pad_groupi_n_1011 ,csa_tree_add_107_22_pad_groupi_n_1059);
  and csa_tree_add_107_22_pad_groupi_g4593(csa_tree_add_107_22_pad_groupi_n_1122 ,csa_tree_add_107_22_pad_groupi_n_880 ,csa_tree_add_107_22_pad_groupi_n_1045);
  and csa_tree_add_107_22_pad_groupi_g4594(csa_tree_add_107_22_pad_groupi_n_1121 ,csa_tree_add_107_22_pad_groupi_n_867 ,csa_tree_add_107_22_pad_groupi_n_1044);
  or csa_tree_add_107_22_pad_groupi_g4595(csa_tree_add_107_22_pad_groupi_n_1120 ,csa_tree_add_107_22_pad_groupi_n_1011 ,csa_tree_add_107_22_pad_groupi_n_1059);
  nor csa_tree_add_107_22_pad_groupi_g4596(csa_tree_add_107_22_pad_groupi_n_1119 ,csa_tree_add_107_22_pad_groupi_n_1026 ,csa_tree_add_107_22_pad_groupi_n_980);
  or csa_tree_add_107_22_pad_groupi_g4597(csa_tree_add_107_22_pad_groupi_n_1118 ,csa_tree_add_107_22_pad_groupi_n_1009 ,csa_tree_add_107_22_pad_groupi_n_1064);
  and csa_tree_add_107_22_pad_groupi_g4598(csa_tree_add_107_22_pad_groupi_n_1117 ,csa_tree_add_107_22_pad_groupi_n_1029 ,csa_tree_add_107_22_pad_groupi_n_1043);
  or csa_tree_add_107_22_pad_groupi_g4599(csa_tree_add_107_22_pad_groupi_n_1116 ,csa_tree_add_107_22_pad_groupi_n_882 ,csa_tree_add_107_22_pad_groupi_n_1038);
  or csa_tree_add_107_22_pad_groupi_g4600(csa_tree_add_107_22_pad_groupi_n_1115 ,csa_tree_add_107_22_pad_groupi_n_1057 ,csa_tree_add_107_22_pad_groupi_n_1060);
  or csa_tree_add_107_22_pad_groupi_g4601(csa_tree_add_107_22_pad_groupi_n_1114 ,csa_tree_add_107_22_pad_groupi_n_1017 ,csa_tree_add_107_22_pad_groupi_n_1065);
  and csa_tree_add_107_22_pad_groupi_g4602(csa_tree_add_107_22_pad_groupi_n_1113 ,csa_tree_add_107_22_pad_groupi_n_860 ,csa_tree_add_107_22_pad_groupi_n_1041);
  or csa_tree_add_107_22_pad_groupi_g4603(csa_tree_add_107_22_pad_groupi_n_1112 ,csa_tree_add_107_22_pad_groupi_n_854 ,csa_tree_add_107_22_pad_groupi_n_1046);
  or csa_tree_add_107_22_pad_groupi_g4604(csa_tree_add_107_22_pad_groupi_n_1111 ,csa_tree_add_107_22_pad_groupi_n_1028 ,csa_tree_add_107_22_pad_groupi_n_976);
  nor csa_tree_add_107_22_pad_groupi_g4605(csa_tree_add_107_22_pad_groupi_n_1110 ,csa_tree_add_107_22_pad_groupi_n_1018 ,csa_tree_add_107_22_pad_groupi_n_1066);
  xnor csa_tree_add_107_22_pad_groupi_g4606(csa_tree_add_107_22_pad_groupi_n_1141 ,csa_tree_add_107_22_pad_groupi_n_842 ,csa_tree_add_107_22_pad_groupi_n_951);
  xnor csa_tree_add_107_22_pad_groupi_g4607(csa_tree_add_107_22_pad_groupi_n_1140 ,csa_tree_add_107_22_pad_groupi_n_803 ,csa_tree_add_107_22_pad_groupi_n_964);
  xnor csa_tree_add_107_22_pad_groupi_g4608(csa_tree_add_107_22_pad_groupi_n_1138 ,csa_tree_add_107_22_pad_groupi_n_773 ,csa_tree_add_107_22_pad_groupi_n_962);
  xnor csa_tree_add_107_22_pad_groupi_g4609(csa_tree_add_107_22_pad_groupi_n_1137 ,csa_tree_add_107_22_pad_groupi_n_783 ,csa_tree_add_107_22_pad_groupi_n_960);
  xnor csa_tree_add_107_22_pad_groupi_g4610(csa_tree_add_107_22_pad_groupi_n_1135 ,csa_tree_add_107_22_pad_groupi_n_840 ,csa_tree_add_107_22_pad_groupi_n_965);
  or csa_tree_add_107_22_pad_groupi_g4611(csa_tree_add_107_22_pad_groupi_n_1134 ,csa_tree_add_107_22_pad_groupi_n_1000 ,csa_tree_add_107_22_pad_groupi_n_1052);
  xnor csa_tree_add_107_22_pad_groupi_g4612(csa_tree_add_107_22_pad_groupi_n_1133 ,csa_tree_add_107_22_pad_groupi_n_778 ,csa_tree_add_107_22_pad_groupi_n_949);
  and csa_tree_add_107_22_pad_groupi_g4613(csa_tree_add_107_22_pad_groupi_n_1132 ,csa_tree_add_107_22_pad_groupi_n_888 ,csa_tree_add_107_22_pad_groupi_n_1032);
  or csa_tree_add_107_22_pad_groupi_g4614(csa_tree_add_107_22_pad_groupi_n_1131 ,csa_tree_add_107_22_pad_groupi_n_868 ,csa_tree_add_107_22_pad_groupi_n_1027);
  not csa_tree_add_107_22_pad_groupi_g4615(csa_tree_add_107_22_pad_groupi_n_1109 ,csa_tree_add_107_22_pad_groupi_n_1108);
  not csa_tree_add_107_22_pad_groupi_g4616(csa_tree_add_107_22_pad_groupi_n_1097 ,csa_tree_add_107_22_pad_groupi_n_1096);
  not csa_tree_add_107_22_pad_groupi_g4617(csa_tree_add_107_22_pad_groupi_n_1091 ,csa_tree_add_107_22_pad_groupi_n_1092);
  not csa_tree_add_107_22_pad_groupi_g4618(csa_tree_add_107_22_pad_groupi_n_1090 ,csa_tree_add_107_22_pad_groupi_n_1089);
  not csa_tree_add_107_22_pad_groupi_g4619(csa_tree_add_107_22_pad_groupi_n_1085 ,csa_tree_add_107_22_pad_groupi_n_1086);
  not csa_tree_add_107_22_pad_groupi_g4620(csa_tree_add_107_22_pad_groupi_n_1083 ,csa_tree_add_107_22_pad_groupi_n_1084);
  not csa_tree_add_107_22_pad_groupi_g4621(csa_tree_add_107_22_pad_groupi_n_1081 ,csa_tree_add_107_22_pad_groupi_n_1082);
  xnor csa_tree_add_107_22_pad_groupi_g4622(csa_tree_add_107_22_pad_groupi_n_1079 ,csa_tree_add_107_22_pad_groupi_n_975 ,csa_tree_add_107_22_pad_groupi_n_934);
  xnor csa_tree_add_107_22_pad_groupi_g4623(csa_tree_add_107_22_pad_groupi_n_1108 ,csa_tree_add_107_22_pad_groupi_n_892 ,csa_tree_add_107_22_pad_groupi_n_961);
  xnor csa_tree_add_107_22_pad_groupi_g4624(csa_tree_add_107_22_pad_groupi_n_1078 ,csa_tree_add_107_22_pad_groupi_n_797 ,csa_tree_add_107_22_pad_groupi_n_4);
  xnor csa_tree_add_107_22_pad_groupi_g4625(csa_tree_add_107_22_pad_groupi_n_1077 ,csa_tree_add_107_22_pad_groupi_n_746 ,csa_tree_add_107_22_pad_groupi_n_1014);
  xnor csa_tree_add_107_22_pad_groupi_g4626(csa_tree_add_107_22_pad_groupi_n_1076 ,csa_tree_add_107_22_pad_groupi_n_1012 ,csa_tree_add_107_22_pad_groupi_n_933);
  xnor csa_tree_add_107_22_pad_groupi_g4628(csa_tree_add_107_22_pad_groupi_n_1107 ,csa_tree_add_107_22_pad_groupi_n_768 ,csa_tree_add_107_22_pad_groupi_n_942);
  xnor csa_tree_add_107_22_pad_groupi_g4629(csa_tree_add_107_22_pad_groupi_n_1106 ,csa_tree_add_107_22_pad_groupi_n_764 ,csa_tree_add_107_22_pad_groupi_n_968);
  xnor csa_tree_add_107_22_pad_groupi_g4630(csa_tree_add_107_22_pad_groupi_n_1105 ,csa_tree_add_107_22_pad_groupi_n_740 ,csa_tree_add_107_22_pad_groupi_n_963);
  xnor csa_tree_add_107_22_pad_groupi_g4631(csa_tree_add_107_22_pad_groupi_n_1104 ,csa_tree_add_107_22_pad_groupi_n_782 ,csa_tree_add_107_22_pad_groupi_n_967);
  xnor csa_tree_add_107_22_pad_groupi_g4632(csa_tree_add_107_22_pad_groupi_n_1103 ,csa_tree_add_107_22_pad_groupi_n_1021 ,csa_tree_add_107_22_pad_groupi_n_957);
  xnor csa_tree_add_107_22_pad_groupi_g4633(csa_tree_add_107_22_pad_groupi_n_1102 ,csa_tree_add_107_22_pad_groupi_n_769 ,csa_tree_add_107_22_pad_groupi_n_945);
  xnor csa_tree_add_107_22_pad_groupi_g4634(csa_tree_add_107_22_pad_groupi_n_1101 ,csa_tree_add_107_22_pad_groupi_n_977 ,csa_tree_add_107_22_pad_groupi_n_966);
  xnor csa_tree_add_107_22_pad_groupi_g4635(csa_tree_add_107_22_pad_groupi_n_1100 ,csa_tree_add_107_22_pad_groupi_n_838 ,csa_tree_add_107_22_pad_groupi_n_946);
  xnor csa_tree_add_107_22_pad_groupi_g4637(csa_tree_add_107_22_pad_groupi_n_1099 ,csa_tree_add_107_22_pad_groupi_n_750 ,csa_tree_add_107_22_pad_groupi_n_952);
  xnor csa_tree_add_107_22_pad_groupi_g4638(csa_tree_add_107_22_pad_groupi_n_1098 ,csa_tree_add_107_22_pad_groupi_n_743 ,csa_tree_add_107_22_pad_groupi_n_972);
  xnor csa_tree_add_107_22_pad_groupi_g4639(csa_tree_add_107_22_pad_groupi_n_1096 ,csa_tree_add_107_22_pad_groupi_n_971 ,csa_tree_add_107_22_pad_groupi_n_578);
  xnor csa_tree_add_107_22_pad_groupi_g4640(csa_tree_add_107_22_pad_groupi_n_1095 ,csa_tree_add_107_22_pad_groupi_n_770 ,csa_tree_add_107_22_pad_groupi_n_947);
  xnor csa_tree_add_107_22_pad_groupi_g4641(csa_tree_add_107_22_pad_groupi_n_1094 ,csa_tree_add_107_22_pad_groupi_n_830 ,csa_tree_add_107_22_pad_groupi_n_943);
  xnor csa_tree_add_107_22_pad_groupi_g4642(csa_tree_add_107_22_pad_groupi_n_1093 ,csa_tree_add_107_22_pad_groupi_n_780 ,csa_tree_add_107_22_pad_groupi_n_938);
  xnor csa_tree_add_107_22_pad_groupi_g4643(csa_tree_add_107_22_pad_groupi_n_1092 ,csa_tree_add_107_22_pad_groupi_n_775 ,csa_tree_add_107_22_pad_groupi_n_937);
  xnor csa_tree_add_107_22_pad_groupi_g4644(csa_tree_add_107_22_pad_groupi_n_1089 ,csa_tree_add_107_22_pad_groupi_n_827 ,csa_tree_add_107_22_pad_groupi_n_973);
  xnor csa_tree_add_107_22_pad_groupi_g4645(csa_tree_add_107_22_pad_groupi_n_1088 ,csa_tree_add_107_22_pad_groupi_n_777 ,csa_tree_add_107_22_pad_groupi_n_940);
  xnor csa_tree_add_107_22_pad_groupi_g4646(csa_tree_add_107_22_pad_groupi_n_1087 ,csa_tree_add_107_22_pad_groupi_n_774 ,csa_tree_add_107_22_pad_groupi_n_954);
  xnor csa_tree_add_107_22_pad_groupi_g4647(csa_tree_add_107_22_pad_groupi_n_1086 ,csa_tree_add_107_22_pad_groupi_n_893 ,csa_tree_add_107_22_pad_groupi_n_959);
  xnor csa_tree_add_107_22_pad_groupi_g4648(csa_tree_add_107_22_pad_groupi_n_1084 ,csa_tree_add_107_22_pad_groupi_n_785 ,csa_tree_add_107_22_pad_groupi_n_956);
  xnor csa_tree_add_107_22_pad_groupi_g4649(csa_tree_add_107_22_pad_groupi_n_1082 ,csa_tree_add_107_22_pad_groupi_n_839 ,csa_tree_add_107_22_pad_groupi_n_958);
  xnor csa_tree_add_107_22_pad_groupi_g4650(csa_tree_add_107_22_pad_groupi_n_1080 ,csa_tree_add_107_22_pad_groupi_n_936 ,csa_tree_add_107_22_pad_groupi_n_953);
  not csa_tree_add_107_22_pad_groupi_g4651(csa_tree_add_107_22_pad_groupi_n_1071 ,csa_tree_add_107_22_pad_groupi_n_1070);
  not csa_tree_add_107_22_pad_groupi_g4652(csa_tree_add_107_22_pad_groupi_n_1069 ,csa_tree_add_107_22_pad_groupi_n_1068);
  not csa_tree_add_107_22_pad_groupi_g4653(csa_tree_add_107_22_pad_groupi_n_1065 ,csa_tree_add_107_22_pad_groupi_n_1066);
  not csa_tree_add_107_22_pad_groupi_g4654(csa_tree_add_107_22_pad_groupi_n_1063 ,csa_tree_add_107_22_pad_groupi_n_1064);
  not csa_tree_add_107_22_pad_groupi_g4655(csa_tree_add_107_22_pad_groupi_n_1060 ,csa_tree_add_107_22_pad_groupi_n_1061);
  not csa_tree_add_107_22_pad_groupi_g4656(csa_tree_add_107_22_pad_groupi_n_1057 ,csa_tree_add_107_22_pad_groupi_n_1058);
  or csa_tree_add_107_22_pad_groupi_g4657(csa_tree_add_107_22_pad_groupi_n_1054 ,csa_tree_add_107_22_pad_groupi_n_276 ,csa_tree_add_107_22_pad_groupi_n_975);
  and csa_tree_add_107_22_pad_groupi_g4658(csa_tree_add_107_22_pad_groupi_n_1053 ,csa_tree_add_107_22_pad_groupi_n_934 ,csa_tree_add_107_22_pad_groupi_n_975);
  and csa_tree_add_107_22_pad_groupi_g4659(csa_tree_add_107_22_pad_groupi_n_1052 ,csa_tree_add_107_22_pad_groupi_n_998 ,csa_tree_add_107_22_pad_groupi_n_1020);
  and csa_tree_add_107_22_pad_groupi_g4660(csa_tree_add_107_22_pad_groupi_n_1051 ,csa_tree_add_107_22_pad_groupi_n_933 ,csa_tree_add_107_22_pad_groupi_n_1012);
  or csa_tree_add_107_22_pad_groupi_g4661(csa_tree_add_107_22_pad_groupi_n_1050 ,csa_tree_add_107_22_pad_groupi_n_933 ,csa_tree_add_107_22_pad_groupi_n_1012);
  and csa_tree_add_107_22_pad_groupi_g4662(csa_tree_add_107_22_pad_groupi_n_1049 ,csa_tree_add_107_22_pad_groupi_n_797 ,csa_tree_add_107_22_pad_groupi_n_4);
  and csa_tree_add_107_22_pad_groupi_g4663(csa_tree_add_107_22_pad_groupi_n_1074 ,csa_tree_add_107_22_pad_groupi_n_913 ,csa_tree_add_107_22_pad_groupi_n_1007);
  or csa_tree_add_107_22_pad_groupi_g4664(csa_tree_add_107_22_pad_groupi_n_1073 ,csa_tree_add_107_22_pad_groupi_n_910 ,csa_tree_add_107_22_pad_groupi_n_999);
  and csa_tree_add_107_22_pad_groupi_g4665(csa_tree_add_107_22_pad_groupi_n_1072 ,csa_tree_add_107_22_pad_groupi_n_915 ,csa_tree_add_107_22_pad_groupi_n_996);
  or csa_tree_add_107_22_pad_groupi_g4666(csa_tree_add_107_22_pad_groupi_n_1070 ,csa_tree_add_107_22_pad_groupi_n_890 ,csa_tree_add_107_22_pad_groupi_n_1005);
  or csa_tree_add_107_22_pad_groupi_g4667(csa_tree_add_107_22_pad_groupi_n_1068 ,csa_tree_add_107_22_pad_groupi_n_905 ,csa_tree_add_107_22_pad_groupi_n_1003);
  and csa_tree_add_107_22_pad_groupi_g4668(csa_tree_add_107_22_pad_groupi_n_1067 ,csa_tree_add_107_22_pad_groupi_n_912 ,csa_tree_add_107_22_pad_groupi_n_1002);
  or csa_tree_add_107_22_pad_groupi_g4669(csa_tree_add_107_22_pad_groupi_n_1066 ,csa_tree_add_107_22_pad_groupi_n_903 ,csa_tree_add_107_22_pad_groupi_n_1004);
  or csa_tree_add_107_22_pad_groupi_g4670(csa_tree_add_107_22_pad_groupi_n_1064 ,csa_tree_add_107_22_pad_groupi_n_925 ,csa_tree_add_107_22_pad_groupi_n_1006);
  or csa_tree_add_107_22_pad_groupi_g4671(csa_tree_add_107_22_pad_groupi_n_1062 ,csa_tree_add_107_22_pad_groupi_n_874 ,csa_tree_add_107_22_pad_groupi_n_987);
  or csa_tree_add_107_22_pad_groupi_g4672(csa_tree_add_107_22_pad_groupi_n_1061 ,csa_tree_add_107_22_pad_groupi_n_929 ,csa_tree_add_107_22_pad_groupi_n_979);
  or csa_tree_add_107_22_pad_groupi_g4673(csa_tree_add_107_22_pad_groupi_n_1059 ,csa_tree_add_107_22_pad_groupi_n_889 ,csa_tree_add_107_22_pad_groupi_n_995);
  or csa_tree_add_107_22_pad_groupi_g4674(csa_tree_add_107_22_pad_groupi_n_1058 ,csa_tree_add_107_22_pad_groupi_n_911 ,csa_tree_add_107_22_pad_groupi_n_1008);
  or csa_tree_add_107_22_pad_groupi_g4675(csa_tree_add_107_22_pad_groupi_n_1056 ,csa_tree_add_107_22_pad_groupi_n_869 ,csa_tree_add_107_22_pad_groupi_n_1001);
  or csa_tree_add_107_22_pad_groupi_g4676(csa_tree_add_107_22_pad_groupi_n_1055 ,csa_tree_add_107_22_pad_groupi_n_886 ,csa_tree_add_107_22_pad_groupi_n_993);
  not csa_tree_add_107_22_pad_groupi_g4677(csa_tree_add_107_22_pad_groupi_n_1048 ,csa_tree_add_107_22_pad_groupi_n_1047);
  not csa_tree_add_107_22_pad_groupi_g4678(csa_tree_add_107_22_pad_groupi_n_1037 ,csa_tree_add_107_22_pad_groupi_n_1036);
  not csa_tree_add_107_22_pad_groupi_g4679(csa_tree_add_107_22_pad_groupi_n_1033 ,csa_tree_add_107_22_pad_groupi_n_1034);
  or csa_tree_add_107_22_pad_groupi_g4680(csa_tree_add_107_22_pad_groupi_n_1032 ,csa_tree_add_107_22_pad_groupi_n_876 ,csa_tree_add_107_22_pad_groupi_n_977);
  nor csa_tree_add_107_22_pad_groupi_g4681(csa_tree_add_107_22_pad_groupi_n_1031 ,csa_tree_add_107_22_pad_groupi_n_646 ,csa_tree_add_107_22_pad_groupi_n_1024);
  or csa_tree_add_107_22_pad_groupi_g4682(csa_tree_add_107_22_pad_groupi_n_1030 ,csa_tree_add_107_22_pad_groupi_n_745 ,csa_tree_add_107_22_pad_groupi_n_1014);
  or csa_tree_add_107_22_pad_groupi_g4683(csa_tree_add_107_22_pad_groupi_n_1029 ,csa_tree_add_107_22_pad_groupi_n_797 ,csa_tree_add_107_22_pad_groupi_n_4);
  nor csa_tree_add_107_22_pad_groupi_g4684(csa_tree_add_107_22_pad_groupi_n_1028 ,csa_tree_add_107_22_pad_groupi_n_746 ,csa_tree_add_107_22_pad_groupi_n_1013);
  and csa_tree_add_107_22_pad_groupi_g4685(csa_tree_add_107_22_pad_groupi_n_1027 ,csa_tree_add_107_22_pad_groupi_n_865 ,csa_tree_add_107_22_pad_groupi_n_1021);
  and csa_tree_add_107_22_pad_groupi_g4686(csa_tree_add_107_22_pad_groupi_n_1026 ,csa_tree_add_107_22_pad_groupi_n_646 ,csa_tree_add_107_22_pad_groupi_n_1024);
  and csa_tree_add_107_22_pad_groupi_g4687(csa_tree_add_107_22_pad_groupi_n_1047 ,csa_tree_add_107_22_pad_groupi_n_895 ,csa_tree_add_107_22_pad_groupi_n_994);
  xnor csa_tree_add_107_22_pad_groupi_g4688(csa_tree_add_107_22_pad_groupi_n_1025 ,csa_tree_add_107_22_pad_groupi_n_935 ,csa_tree_add_107_22_pad_groupi_n_820);
  and csa_tree_add_107_22_pad_groupi_g4689(csa_tree_add_107_22_pad_groupi_n_1046 ,csa_tree_add_107_22_pad_groupi_n_853 ,csa_tree_add_107_22_pad_groupi_n_982);
  or csa_tree_add_107_22_pad_groupi_g4690(csa_tree_add_107_22_pad_groupi_n_1045 ,csa_tree_add_107_22_pad_groupi_n_906 ,csa_tree_add_107_22_pad_groupi_n_997);
  or csa_tree_add_107_22_pad_groupi_g4691(csa_tree_add_107_22_pad_groupi_n_1044 ,csa_tree_add_107_22_pad_groupi_n_887 ,csa_tree_add_107_22_pad_groupi_n_992);
  or csa_tree_add_107_22_pad_groupi_g4692(csa_tree_add_107_22_pad_groupi_n_1043 ,csa_tree_add_107_22_pad_groupi_n_926 ,csa_tree_add_107_22_pad_groupi_n_991);
  and csa_tree_add_107_22_pad_groupi_g4693(csa_tree_add_107_22_pad_groupi_n_1042 ,csa_tree_add_107_22_pad_groupi_n_864 ,csa_tree_add_107_22_pad_groupi_n_985);
  or csa_tree_add_107_22_pad_groupi_g4694(csa_tree_add_107_22_pad_groupi_n_1041 ,csa_tree_add_107_22_pad_groupi_n_879 ,csa_tree_add_107_22_pad_groupi_n_984);
  or csa_tree_add_107_22_pad_groupi_g4695(csa_tree_add_107_22_pad_groupi_n_1040 ,csa_tree_add_107_22_pad_groupi_n_870 ,csa_tree_add_107_22_pad_groupi_n_988);
  and csa_tree_add_107_22_pad_groupi_g4696(csa_tree_add_107_22_pad_groupi_n_1039 ,csa_tree_add_107_22_pad_groupi_n_852 ,csa_tree_add_107_22_pad_groupi_n_981);
  and csa_tree_add_107_22_pad_groupi_g4697(csa_tree_add_107_22_pad_groupi_n_1038 ,csa_tree_add_107_22_pad_groupi_n_878 ,csa_tree_add_107_22_pad_groupi_n_989);
  or csa_tree_add_107_22_pad_groupi_g4698(csa_tree_add_107_22_pad_groupi_n_1036 ,csa_tree_add_107_22_pad_groupi_n_897 ,csa_tree_add_107_22_pad_groupi_n_983);
  or csa_tree_add_107_22_pad_groupi_g4699(csa_tree_add_107_22_pad_groupi_n_1035 ,csa_tree_add_107_22_pad_groupi_n_907 ,csa_tree_add_107_22_pad_groupi_n_990);
  or csa_tree_add_107_22_pad_groupi_g4700(csa_tree_add_107_22_pad_groupi_n_1034 ,csa_tree_add_107_22_pad_groupi_n_866 ,csa_tree_add_107_22_pad_groupi_n_986);
  not csa_tree_add_107_22_pad_groupi_g4701(csa_tree_add_107_22_pad_groupi_n_1023 ,csa_tree_add_107_22_pad_groupi_n_1022);
  not csa_tree_add_107_22_pad_groupi_g4702(csa_tree_add_107_22_pad_groupi_n_1018 ,csa_tree_add_107_22_pad_groupi_n_1017);
  not csa_tree_add_107_22_pad_groupi_g4703(csa_tree_add_107_22_pad_groupi_n_1016 ,csa_tree_add_107_22_pad_groupi_n_1015);
  not csa_tree_add_107_22_pad_groupi_g4704(csa_tree_add_107_22_pad_groupi_n_1014 ,csa_tree_add_107_22_pad_groupi_n_1013);
  not csa_tree_add_107_22_pad_groupi_g4705(csa_tree_add_107_22_pad_groupi_n_1010 ,csa_tree_add_107_22_pad_groupi_n_1009);
  nor csa_tree_add_107_22_pad_groupi_g4706(csa_tree_add_107_22_pad_groupi_n_1008 ,csa_tree_add_107_22_pad_groupi_n_841 ,csa_tree_add_107_22_pad_groupi_n_930);
  or csa_tree_add_107_22_pad_groupi_g4707(csa_tree_add_107_22_pad_groupi_n_1007 ,csa_tree_add_107_22_pad_groupi_n_843 ,csa_tree_add_107_22_pad_groupi_n_917);
  nor csa_tree_add_107_22_pad_groupi_g4708(csa_tree_add_107_22_pad_groupi_n_1006 ,csa_tree_add_107_22_pad_groupi_n_824 ,csa_tree_add_107_22_pad_groupi_n_872);
  and csa_tree_add_107_22_pad_groupi_g4709(csa_tree_add_107_22_pad_groupi_n_1005 ,csa_tree_add_107_22_pad_groupi_n_840 ,csa_tree_add_107_22_pad_groupi_n_922);
  and csa_tree_add_107_22_pad_groupi_g4710(csa_tree_add_107_22_pad_groupi_n_1004 ,csa_tree_add_107_22_pad_groupi_n_839 ,csa_tree_add_107_22_pad_groupi_n_909);
  and csa_tree_add_107_22_pad_groupi_g4711(csa_tree_add_107_22_pad_groupi_n_1003 ,csa_tree_add_107_22_pad_groupi_n_770 ,csa_tree_add_107_22_pad_groupi_n_916);
  or csa_tree_add_107_22_pad_groupi_g4712(csa_tree_add_107_22_pad_groupi_n_1002 ,csa_tree_add_107_22_pad_groupi_n_779 ,csa_tree_add_107_22_pad_groupi_n_902);
  and csa_tree_add_107_22_pad_groupi_g4713(csa_tree_add_107_22_pad_groupi_n_1001 ,csa_tree_add_107_22_pad_groupi_n_769 ,csa_tree_add_107_22_pad_groupi_n_904);
  and csa_tree_add_107_22_pad_groupi_g4714(csa_tree_add_107_22_pad_groupi_n_1000 ,csa_tree_add_107_22_pad_groupi_n_820 ,csa_tree_add_107_22_pad_groupi_n_935);
  nor csa_tree_add_107_22_pad_groupi_g4715(csa_tree_add_107_22_pad_groupi_n_999 ,csa_tree_add_107_22_pad_groupi_n_834 ,csa_tree_add_107_22_pad_groupi_n_896);
  or csa_tree_add_107_22_pad_groupi_g4716(csa_tree_add_107_22_pad_groupi_n_998 ,csa_tree_add_107_22_pad_groupi_n_820 ,csa_tree_add_107_22_pad_groupi_n_935);
  and csa_tree_add_107_22_pad_groupi_g4717(csa_tree_add_107_22_pad_groupi_n_997 ,csa_tree_add_107_22_pad_groupi_n_830 ,csa_tree_add_107_22_pad_groupi_n_856);
  or csa_tree_add_107_22_pad_groupi_g4718(csa_tree_add_107_22_pad_groupi_n_996 ,csa_tree_add_107_22_pad_groupi_n_936 ,csa_tree_add_107_22_pad_groupi_n_919);
  and csa_tree_add_107_22_pad_groupi_g4719(csa_tree_add_107_22_pad_groupi_n_995 ,csa_tree_add_107_22_pad_groupi_n_775 ,csa_tree_add_107_22_pad_groupi_n_891);
  or csa_tree_add_107_22_pad_groupi_g4720(csa_tree_add_107_22_pad_groupi_n_994 ,csa_tree_add_107_22_pad_groupi_n_892 ,csa_tree_add_107_22_pad_groupi_n_894);
  and csa_tree_add_107_22_pad_groupi_g4721(csa_tree_add_107_22_pad_groupi_n_993 ,csa_tree_add_107_22_pad_groupi_n_768 ,csa_tree_add_107_22_pad_groupi_n_924);
  and csa_tree_add_107_22_pad_groupi_g4722(csa_tree_add_107_22_pad_groupi_n_992 ,csa_tree_add_107_22_pad_groupi_n_780 ,csa_tree_add_107_22_pad_groupi_n_885);
  nor csa_tree_add_107_22_pad_groupi_g4723(csa_tree_add_107_22_pad_groupi_n_991 ,csa_tree_add_107_22_pad_groupi_n_837 ,csa_tree_add_107_22_pad_groupi_n_877);
  and csa_tree_add_107_22_pad_groupi_g4724(csa_tree_add_107_22_pad_groupi_n_990 ,csa_tree_add_107_22_pad_groupi_n_777 ,csa_tree_add_107_22_pad_groupi_n_928);
  or csa_tree_add_107_22_pad_groupi_g4725(csa_tree_add_107_22_pad_groupi_n_989 ,csa_tree_add_107_22_pad_groupi_n_838 ,csa_tree_add_107_22_pad_groupi_n_875);
  nor csa_tree_add_107_22_pad_groupi_g4726(csa_tree_add_107_22_pad_groupi_n_988 ,csa_tree_add_107_22_pad_groupi_n_774 ,csa_tree_add_107_22_pad_groupi_n_855);
  nor csa_tree_add_107_22_pad_groupi_g4727(csa_tree_add_107_22_pad_groupi_n_987 ,csa_tree_add_107_22_pad_groupi_n_776 ,csa_tree_add_107_22_pad_groupi_n_883);
  and csa_tree_add_107_22_pad_groupi_g4728(csa_tree_add_107_22_pad_groupi_n_986 ,csa_tree_add_107_22_pad_groupi_n_773 ,csa_tree_add_107_22_pad_groupi_n_863);
  or csa_tree_add_107_22_pad_groupi_g4729(csa_tree_add_107_22_pad_groupi_n_985 ,csa_tree_add_107_22_pad_groupi_n_823 ,csa_tree_add_107_22_pad_groupi_n_862);
  nor csa_tree_add_107_22_pad_groupi_g4730(csa_tree_add_107_22_pad_groupi_n_984 ,csa_tree_add_107_22_pad_groupi_n_772 ,csa_tree_add_107_22_pad_groupi_n_859);
  nor csa_tree_add_107_22_pad_groupi_g4731(csa_tree_add_107_22_pad_groupi_n_983 ,csa_tree_add_107_22_pad_groupi_n_771 ,csa_tree_add_107_22_pad_groupi_n_900);
  or csa_tree_add_107_22_pad_groupi_g4732(csa_tree_add_107_22_pad_groupi_n_982 ,csa_tree_add_107_22_pad_groupi_n_835 ,csa_tree_add_107_22_pad_groupi_n_851);
  or csa_tree_add_107_22_pad_groupi_g4733(csa_tree_add_107_22_pad_groupi_n_981 ,csa_tree_add_107_22_pad_groupi_n_893 ,csa_tree_add_107_22_pad_groupi_n_920);
  xnor csa_tree_add_107_22_pad_groupi_g4734(csa_tree_add_107_22_pad_groupi_n_980 ,csa_tree_add_107_22_pad_groupi_n_846 ,csa_tree_add_107_22_pad_groupi_n_848);
  and csa_tree_add_107_22_pad_groupi_g4735(csa_tree_add_107_22_pad_groupi_n_979 ,csa_tree_add_107_22_pad_groupi_n_827 ,csa_tree_add_107_22_pad_groupi_n_927);
  or csa_tree_add_107_22_pad_groupi_g4736(csa_tree_add_107_22_pad_groupi_n_1024 ,csa_tree_add_107_22_pad_groupi_n_19 ,csa_tree_add_107_22_pad_groupi_n_898);
  xnor csa_tree_add_107_22_pad_groupi_g4737(csa_tree_add_107_22_pad_groupi_n_1022 ,csa_tree_add_107_22_pad_groupi_n_706 ,csa_tree_add_107_22_pad_groupi_n_844);
  xnor csa_tree_add_107_22_pad_groupi_g4739(csa_tree_add_107_22_pad_groupi_n_1021 ,csa_tree_add_107_22_pad_groupi_n_711 ,in25[9]);
  xnor csa_tree_add_107_22_pad_groupi_g4740(csa_tree_add_107_22_pad_groupi_n_1020 ,csa_tree_add_107_22_pad_groupi_n_645 ,csa_tree_add_107_22_pad_groupi_n_832);
  and csa_tree_add_107_22_pad_groupi_g4741(csa_tree_add_107_22_pad_groupi_n_1019 ,csa_tree_add_107_22_pad_groupi_n_899 ,csa_tree_add_107_22_pad_groupi_n_359);
  and csa_tree_add_107_22_pad_groupi_g4742(csa_tree_add_107_22_pad_groupi_n_1017 ,csa_tree_add_107_22_pad_groupi_n_656 ,csa_tree_add_107_22_pad_groupi_n_923);
  or csa_tree_add_107_22_pad_groupi_g4743(csa_tree_add_107_22_pad_groupi_n_1015 ,csa_tree_add_107_22_pad_groupi_n_682 ,csa_tree_add_107_22_pad_groupi_n_881);
  or csa_tree_add_107_22_pad_groupi_g4744(csa_tree_add_107_22_pad_groupi_n_1013 ,csa_tree_add_107_22_pad_groupi_n_666 ,csa_tree_add_107_22_pad_groupi_n_861);
  xnor csa_tree_add_107_22_pad_groupi_g4745(csa_tree_add_107_22_pad_groupi_n_1012 ,csa_tree_add_107_22_pad_groupi_n_704 ,csa_tree_add_107_22_pad_groupi_n_767);
  xnor csa_tree_add_107_22_pad_groupi_g4746(csa_tree_add_107_22_pad_groupi_n_1011 ,csa_tree_add_107_22_pad_groupi_n_831 ,csa_tree_add_107_22_pad_groupi_n_1);
  or csa_tree_add_107_22_pad_groupi_g4747(csa_tree_add_107_22_pad_groupi_n_1009 ,csa_tree_add_107_22_pad_groupi_n_702 ,csa_tree_add_107_22_pad_groupi_n_931);
  xnor csa_tree_add_107_22_pad_groupi_g4748(csa_tree_add_107_22_pad_groupi_n_974 ,csa_tree_add_107_22_pad_groupi_n_726 ,csa_tree_add_107_22_pad_groupi_n_821);
  xnor csa_tree_add_107_22_pad_groupi_g4749(csa_tree_add_107_22_pad_groupi_n_973 ,csa_tree_add_107_22_pad_groupi_n_802 ,csa_tree_add_107_22_pad_groupi_n_795);
  xnor csa_tree_add_107_22_pad_groupi_g4750(csa_tree_add_107_22_pad_groupi_n_972 ,csa_tree_add_107_22_pad_groupi_n_837 ,csa_tree_add_107_22_pad_groupi_n_766);
  xnor csa_tree_add_107_22_pad_groupi_g4751(csa_tree_add_107_22_pad_groupi_n_971 ,csa_tree_add_107_22_pad_groupi_n_829 ,in25[12]);
  xnor csa_tree_add_107_22_pad_groupi_g4752(csa_tree_add_107_22_pad_groupi_n_970 ,csa_tree_add_107_22_pad_groupi_n_739 ,csa_tree_add_107_22_pad_groupi_n_728);
  xnor csa_tree_add_107_22_pad_groupi_g4753(csa_tree_add_107_22_pad_groupi_n_969 ,csa_tree_add_107_22_pad_groupi_n_758 ,csa_tree_add_107_22_pad_groupi_n_757);
  xor csa_tree_add_107_22_pad_groupi_g4754(csa_tree_add_107_22_pad_groupi_n_968 ,csa_tree_add_107_22_pad_groupi_n_824 ,csa_tree_add_107_22_pad_groupi_n_809);
  xor csa_tree_add_107_22_pad_groupi_g4755(csa_tree_add_107_22_pad_groupi_n_967 ,csa_tree_add_107_22_pad_groupi_n_834 ,in25[8]);
  xnor csa_tree_add_107_22_pad_groupi_g4756(csa_tree_add_107_22_pad_groupi_n_966 ,csa_tree_add_107_22_pad_groupi_n_733 ,csa_tree_add_107_22_pad_groupi_n_755);
  xnor csa_tree_add_107_22_pad_groupi_g4757(csa_tree_add_107_22_pad_groupi_n_965 ,csa_tree_add_107_22_pad_groupi_n_800 ,csa_tree_add_107_22_pad_groupi_n_799);
  xor csa_tree_add_107_22_pad_groupi_g4758(csa_tree_add_107_22_pad_groupi_n_964 ,csa_tree_add_107_22_pad_groupi_n_776 ,csa_tree_add_107_22_pad_groupi_n_721);
  xor csa_tree_add_107_22_pad_groupi_g4759(csa_tree_add_107_22_pad_groupi_n_963 ,csa_tree_add_107_22_pad_groupi_n_772 ,in25[1]);
  xnor csa_tree_add_107_22_pad_groupi_g4760(csa_tree_add_107_22_pad_groupi_n_962 ,csa_tree_add_107_22_pad_groupi_n_765 ,csa_tree_add_107_22_pad_groupi_n_751);
  xnor csa_tree_add_107_22_pad_groupi_g4761(csa_tree_add_107_22_pad_groupi_n_961 ,csa_tree_add_107_22_pad_groupi_n_735 ,csa_tree_add_107_22_pad_groupi_n_792);
  xor csa_tree_add_107_22_pad_groupi_g4762(csa_tree_add_107_22_pad_groupi_n_960 ,csa_tree_add_107_22_pad_groupi_n_771 ,csa_tree_add_107_22_pad_groupi_n_729);
  xnor csa_tree_add_107_22_pad_groupi_g4763(csa_tree_add_107_22_pad_groupi_n_959 ,csa_tree_add_107_22_pad_groupi_n_725 ,csa_tree_add_107_22_pad_groupi_n_723);
  xnor csa_tree_add_107_22_pad_groupi_g4764(csa_tree_add_107_22_pad_groupi_n_958 ,csa_tree_add_107_22_pad_groupi_n_814 ,csa_tree_add_107_22_pad_groupi_n_796);
  xnor csa_tree_add_107_22_pad_groupi_g4765(csa_tree_add_107_22_pad_groupi_n_957 ,csa_tree_add_107_22_pad_groupi_n_784 ,csa_tree_add_107_22_pad_groupi_n_747);
  xor csa_tree_add_107_22_pad_groupi_g4766(csa_tree_add_107_22_pad_groupi_n_956 ,csa_tree_add_107_22_pad_groupi_n_841 ,csa_tree_add_107_22_pad_groupi_n_748);
  xnor csa_tree_add_107_22_pad_groupi_g4767(csa_tree_add_107_22_pad_groupi_n_955 ,csa_tree_add_107_22_pad_groupi_n_760 ,csa_tree_add_107_22_pad_groupi_n_737);
  xnor csa_tree_add_107_22_pad_groupi_g4768(csa_tree_add_107_22_pad_groupi_n_954 ,csa_tree_add_107_22_pad_groupi_n_756 ,in25[2]);
  xnor csa_tree_add_107_22_pad_groupi_g4769(csa_tree_add_107_22_pad_groupi_n_953 ,csa_tree_add_107_22_pad_groupi_n_763 ,csa_tree_add_107_22_pad_groupi_n_817);
  xor csa_tree_add_107_22_pad_groupi_g4770(csa_tree_add_107_22_pad_groupi_n_952 ,csa_tree_add_107_22_pad_groupi_n_823 ,csa_tree_add_107_22_pad_groupi_n_742);
  xnor csa_tree_add_107_22_pad_groupi_g4771(csa_tree_add_107_22_pad_groupi_n_951 ,csa_tree_add_107_22_pad_groupi_n_806 ,csa_tree_add_107_22_pad_groupi_n_753);
  xnor csa_tree_add_107_22_pad_groupi_g4772(csa_tree_add_107_22_pad_groupi_n_950 ,csa_tree_add_107_22_pad_groupi_n_790 ,csa_tree_add_107_22_pad_groupi_n_819);
  xnor csa_tree_add_107_22_pad_groupi_g4773(csa_tree_add_107_22_pad_groupi_n_949 ,csa_tree_add_107_22_pad_groupi_n_813 ,csa_tree_add_107_22_pad_groupi_n_716);
  xnor csa_tree_add_107_22_pad_groupi_g4774(csa_tree_add_107_22_pad_groupi_n_948 ,csa_tree_add_107_22_pad_groupi_n_731 ,in25[6]);
  xnor csa_tree_add_107_22_pad_groupi_g4775(csa_tree_add_107_22_pad_groupi_n_947 ,csa_tree_add_107_22_pad_groupi_n_787 ,in25[5]);
  xnor csa_tree_add_107_22_pad_groupi_g4776(csa_tree_add_107_22_pad_groupi_n_946 ,csa_tree_add_107_22_pad_groupi_n_713 ,in25[7]);
  xnor csa_tree_add_107_22_pad_groupi_g4777(csa_tree_add_107_22_pad_groupi_n_945 ,csa_tree_add_107_22_pad_groupi_n_808 ,csa_tree_add_107_22_pad_groupi_n_788);
  xnor csa_tree_add_107_22_pad_groupi_g4778(csa_tree_add_107_22_pad_groupi_n_944 ,csa_tree_add_107_22_pad_groupi_n_761 ,csa_tree_add_107_22_pad_groupi_n_786);
  xnor csa_tree_add_107_22_pad_groupi_g4779(csa_tree_add_107_22_pad_groupi_n_943 ,csa_tree_add_107_22_pad_groupi_n_798 ,in25[4]);
  xnor csa_tree_add_107_22_pad_groupi_g4780(csa_tree_add_107_22_pad_groupi_n_942 ,csa_tree_add_107_22_pad_groupi_n_719 ,csa_tree_add_107_22_pad_groupi_n_720);
  xnor csa_tree_add_107_22_pad_groupi_g4781(csa_tree_add_107_22_pad_groupi_n_941 ,csa_tree_add_107_22_pad_groupi_n_815 ,csa_tree_add_107_22_pad_groupi_n_717);
  xnor csa_tree_add_107_22_pad_groupi_g4782(csa_tree_add_107_22_pad_groupi_n_940 ,csa_tree_add_107_22_pad_groupi_n_807 ,csa_tree_add_107_22_pad_groupi_n_714);
  xnor csa_tree_add_107_22_pad_groupi_g4783(csa_tree_add_107_22_pad_groupi_n_939 ,csa_tree_add_107_22_pad_groupi_n_810 ,csa_tree_add_107_22_pad_groupi_n_811);
  xnor csa_tree_add_107_22_pad_groupi_g4784(csa_tree_add_107_22_pad_groupi_n_938 ,csa_tree_add_107_22_pad_groupi_n_804 ,in25[3]);
  xnor csa_tree_add_107_22_pad_groupi_g4785(csa_tree_add_107_22_pad_groupi_n_937 ,csa_tree_add_107_22_pad_groupi_n_718 ,csa_tree_add_107_22_pad_groupi_n_793);
  xnor csa_tree_add_107_22_pad_groupi_g4786(csa_tree_add_107_22_pad_groupi_n_977 ,csa_tree_add_107_22_pad_groupi_n_822 ,csa_tree_add_107_22_pad_groupi_n_709);
  xnor csa_tree_add_107_22_pad_groupi_g4787(csa_tree_add_107_22_pad_groupi_n_976 ,csa_tree_add_107_22_pad_groupi_n_828 ,csa_tree_add_107_22_pad_groupi_n_710);
  xnor csa_tree_add_107_22_pad_groupi_g4788(csa_tree_add_107_22_pad_groupi_n_975 ,csa_tree_add_107_22_pad_groupi_n_825 ,in25[0]);
  or csa_tree_add_107_22_pad_groupi_g4791(csa_tree_add_107_22_pad_groupi_n_932 ,csa_tree_add_107_22_pad_groupi_n_815 ,csa_tree_add_107_22_pad_groupi_n_717);
  nor csa_tree_add_107_22_pad_groupi_g4792(csa_tree_add_107_22_pad_groupi_n_931 ,csa_tree_add_107_22_pad_groupi_n_673 ,csa_tree_add_107_22_pad_groupi_n_831);
  nor csa_tree_add_107_22_pad_groupi_g4793(csa_tree_add_107_22_pad_groupi_n_930 ,csa_tree_add_107_22_pad_groupi_n_748 ,csa_tree_add_107_22_pad_groupi_n_785);
  nor csa_tree_add_107_22_pad_groupi_g4794(csa_tree_add_107_22_pad_groupi_n_929 ,csa_tree_add_107_22_pad_groupi_n_802 ,csa_tree_add_107_22_pad_groupi_n_794);
  or csa_tree_add_107_22_pad_groupi_g4795(csa_tree_add_107_22_pad_groupi_n_928 ,csa_tree_add_107_22_pad_groupi_n_807 ,csa_tree_add_107_22_pad_groupi_n_714);
  or csa_tree_add_107_22_pad_groupi_g4796(csa_tree_add_107_22_pad_groupi_n_927 ,csa_tree_add_107_22_pad_groupi_n_801 ,csa_tree_add_107_22_pad_groupi_n_795);
  nor csa_tree_add_107_22_pad_groupi_g4797(csa_tree_add_107_22_pad_groupi_n_926 ,csa_tree_add_107_22_pad_groupi_n_766 ,csa_tree_add_107_22_pad_groupi_n_744);
  and csa_tree_add_107_22_pad_groupi_g4798(csa_tree_add_107_22_pad_groupi_n_925 ,csa_tree_add_107_22_pad_groupi_n_764 ,csa_tree_add_107_22_pad_groupi_n_809);
  or csa_tree_add_107_22_pad_groupi_g4799(csa_tree_add_107_22_pad_groupi_n_924 ,csa_tree_add_107_22_pad_groupi_n_719 ,csa_tree_add_107_22_pad_groupi_n_720);
  or csa_tree_add_107_22_pad_groupi_g4800(csa_tree_add_107_22_pad_groupi_n_923 ,csa_tree_add_107_22_pad_groupi_n_593 ,csa_tree_add_107_22_pad_groupi_n_836);
  or csa_tree_add_107_22_pad_groupi_g4801(csa_tree_add_107_22_pad_groupi_n_922 ,csa_tree_add_107_22_pad_groupi_n_800 ,csa_tree_add_107_22_pad_groupi_n_799);
  or csa_tree_add_107_22_pad_groupi_g4802(csa_tree_add_107_22_pad_groupi_n_921 ,csa_tree_add_107_22_pad_groupi_n_789 ,csa_tree_add_107_22_pad_groupi_n_818);
  nor csa_tree_add_107_22_pad_groupi_g4803(csa_tree_add_107_22_pad_groupi_n_920 ,csa_tree_add_107_22_pad_groupi_n_725 ,csa_tree_add_107_22_pad_groupi_n_723);
  nor csa_tree_add_107_22_pad_groupi_g4804(csa_tree_add_107_22_pad_groupi_n_919 ,csa_tree_add_107_22_pad_groupi_n_763 ,csa_tree_add_107_22_pad_groupi_n_817);
  nor csa_tree_add_107_22_pad_groupi_g4805(csa_tree_add_107_22_pad_groupi_n_918 ,csa_tree_add_107_22_pad_groupi_n_790 ,csa_tree_add_107_22_pad_groupi_n_819);
  nor csa_tree_add_107_22_pad_groupi_g4806(csa_tree_add_107_22_pad_groupi_n_917 ,csa_tree_add_107_22_pad_groupi_n_806 ,csa_tree_add_107_22_pad_groupi_n_753);
  or csa_tree_add_107_22_pad_groupi_g4807(csa_tree_add_107_22_pad_groupi_n_916 ,in25[5] ,csa_tree_add_107_22_pad_groupi_n_787);
  or csa_tree_add_107_22_pad_groupi_g4808(csa_tree_add_107_22_pad_groupi_n_915 ,csa_tree_add_107_22_pad_groupi_n_762 ,csa_tree_add_107_22_pad_groupi_n_816);
  and csa_tree_add_107_22_pad_groupi_g4809(csa_tree_add_107_22_pad_groupi_n_914 ,csa_tree_add_107_22_pad_groupi_n_815 ,csa_tree_add_107_22_pad_groupi_n_717);
  or csa_tree_add_107_22_pad_groupi_g4810(csa_tree_add_107_22_pad_groupi_n_913 ,csa_tree_add_107_22_pad_groupi_n_805 ,csa_tree_add_107_22_pad_groupi_n_752);
  or csa_tree_add_107_22_pad_groupi_g4811(csa_tree_add_107_22_pad_groupi_n_912 ,csa_tree_add_107_22_pad_groupi_n_812 ,csa_tree_add_107_22_pad_groupi_n_715);
  and csa_tree_add_107_22_pad_groupi_g4812(csa_tree_add_107_22_pad_groupi_n_911 ,csa_tree_add_107_22_pad_groupi_n_748 ,csa_tree_add_107_22_pad_groupi_n_785);
  nor csa_tree_add_107_22_pad_groupi_g4813(csa_tree_add_107_22_pad_groupi_n_910 ,csa_tree_add_107_22_pad_groupi_n_372 ,csa_tree_add_107_22_pad_groupi_n_782);
  or csa_tree_add_107_22_pad_groupi_g4814(csa_tree_add_107_22_pad_groupi_n_909 ,csa_tree_add_107_22_pad_groupi_n_814 ,csa_tree_add_107_22_pad_groupi_n_796);
  and csa_tree_add_107_22_pad_groupi_g4815(csa_tree_add_107_22_pad_groupi_n_908 ,csa_tree_add_107_22_pad_groupi_n_810 ,csa_tree_add_107_22_pad_groupi_n_811);
  and csa_tree_add_107_22_pad_groupi_g4816(csa_tree_add_107_22_pad_groupi_n_907 ,csa_tree_add_107_22_pad_groupi_n_807 ,csa_tree_add_107_22_pad_groupi_n_714);
  and csa_tree_add_107_22_pad_groupi_g4817(csa_tree_add_107_22_pad_groupi_n_906 ,in25[4] ,csa_tree_add_107_22_pad_groupi_n_798);
  and csa_tree_add_107_22_pad_groupi_g4818(csa_tree_add_107_22_pad_groupi_n_905 ,in25[5] ,csa_tree_add_107_22_pad_groupi_n_787);
  or csa_tree_add_107_22_pad_groupi_g4819(csa_tree_add_107_22_pad_groupi_n_904 ,csa_tree_add_107_22_pad_groupi_n_808 ,csa_tree_add_107_22_pad_groupi_n_788);
  and csa_tree_add_107_22_pad_groupi_g4820(csa_tree_add_107_22_pad_groupi_n_903 ,csa_tree_add_107_22_pad_groupi_n_814 ,csa_tree_add_107_22_pad_groupi_n_796);
  nor csa_tree_add_107_22_pad_groupi_g4821(csa_tree_add_107_22_pad_groupi_n_902 ,csa_tree_add_107_22_pad_groupi_n_813 ,csa_tree_add_107_22_pad_groupi_n_716);
  and csa_tree_add_107_22_pad_groupi_g4822(csa_tree_add_107_22_pad_groupi_n_901 ,csa_tree_add_107_22_pad_groupi_n_761 ,csa_tree_add_107_22_pad_groupi_n_786);
  nor csa_tree_add_107_22_pad_groupi_g4823(csa_tree_add_107_22_pad_groupi_n_900 ,csa_tree_add_107_22_pad_groupi_n_783 ,csa_tree_add_107_22_pad_groupi_n_729);
  or csa_tree_add_107_22_pad_groupi_g4824(csa_tree_add_107_22_pad_groupi_n_899 ,csa_tree_add_107_22_pad_groupi_n_708 ,csa_tree_add_107_22_pad_groupi_n_845);
  or csa_tree_add_107_22_pad_groupi_g4825(csa_tree_add_107_22_pad_groupi_n_898 ,csa_tree_add_107_22_pad_groupi_n_112 ,csa_tree_add_107_22_pad_groupi_n_781);
  and csa_tree_add_107_22_pad_groupi_g4826(csa_tree_add_107_22_pad_groupi_n_897 ,csa_tree_add_107_22_pad_groupi_n_783 ,csa_tree_add_107_22_pad_groupi_n_729);
  and csa_tree_add_107_22_pad_groupi_g4827(csa_tree_add_107_22_pad_groupi_n_896 ,csa_tree_add_107_22_pad_groupi_n_372 ,csa_tree_add_107_22_pad_groupi_n_782);
  or csa_tree_add_107_22_pad_groupi_g4828(csa_tree_add_107_22_pad_groupi_n_895 ,csa_tree_add_107_22_pad_groupi_n_734 ,csa_tree_add_107_22_pad_groupi_n_791);
  nor csa_tree_add_107_22_pad_groupi_g4829(csa_tree_add_107_22_pad_groupi_n_894 ,csa_tree_add_107_22_pad_groupi_n_735 ,csa_tree_add_107_22_pad_groupi_n_792);
  or csa_tree_add_107_22_pad_groupi_g4830(csa_tree_add_107_22_pad_groupi_n_936 ,csa_tree_add_107_22_pad_groupi_n_645 ,csa_tree_add_107_22_pad_groupi_n_833);
  and csa_tree_add_107_22_pad_groupi_g4831(csa_tree_add_107_22_pad_groupi_n_935 ,csa_tree_add_107_22_pad_groupi_n_705 ,csa_tree_add_107_22_pad_groupi_n_767);
  and csa_tree_add_107_22_pad_groupi_g4832(csa_tree_add_107_22_pad_groupi_n_934 ,csa_tree_add_107_22_pad_groupi_n_708 ,csa_tree_add_107_22_pad_groupi_n_845);
  and csa_tree_add_107_22_pad_groupi_g4833(csa_tree_add_107_22_pad_groupi_n_933 ,csa_tree_add_107_22_pad_groupi_n_707 ,csa_tree_add_107_22_pad_groupi_n_844);
  or csa_tree_add_107_22_pad_groupi_g4834(csa_tree_add_107_22_pad_groupi_n_891 ,csa_tree_add_107_22_pad_groupi_n_718 ,csa_tree_add_107_22_pad_groupi_n_793);
  and csa_tree_add_107_22_pad_groupi_g4835(csa_tree_add_107_22_pad_groupi_n_890 ,csa_tree_add_107_22_pad_groupi_n_800 ,csa_tree_add_107_22_pad_groupi_n_799);
  and csa_tree_add_107_22_pad_groupi_g4836(csa_tree_add_107_22_pad_groupi_n_889 ,csa_tree_add_107_22_pad_groupi_n_718 ,csa_tree_add_107_22_pad_groupi_n_793);
  or csa_tree_add_107_22_pad_groupi_g4837(csa_tree_add_107_22_pad_groupi_n_888 ,csa_tree_add_107_22_pad_groupi_n_732 ,csa_tree_add_107_22_pad_groupi_n_754);
  and csa_tree_add_107_22_pad_groupi_g4838(csa_tree_add_107_22_pad_groupi_n_887 ,in25[3] ,csa_tree_add_107_22_pad_groupi_n_804);
  and csa_tree_add_107_22_pad_groupi_g4839(csa_tree_add_107_22_pad_groupi_n_886 ,csa_tree_add_107_22_pad_groupi_n_719 ,csa_tree_add_107_22_pad_groupi_n_720);
  or csa_tree_add_107_22_pad_groupi_g4840(csa_tree_add_107_22_pad_groupi_n_885 ,in25[3] ,csa_tree_add_107_22_pad_groupi_n_804);
  or csa_tree_add_107_22_pad_groupi_g4841(csa_tree_add_107_22_pad_groupi_n_884 ,csa_tree_add_107_22_pad_groupi_n_738 ,csa_tree_add_107_22_pad_groupi_n_727);
  nor csa_tree_add_107_22_pad_groupi_g4842(csa_tree_add_107_22_pad_groupi_n_883 ,csa_tree_add_107_22_pad_groupi_n_803 ,csa_tree_add_107_22_pad_groupi_n_721);
  nor csa_tree_add_107_22_pad_groupi_g4843(csa_tree_add_107_22_pad_groupi_n_882 ,csa_tree_add_107_22_pad_groupi_n_739 ,csa_tree_add_107_22_pad_groupi_n_728);
  nor csa_tree_add_107_22_pad_groupi_g4844(csa_tree_add_107_22_pad_groupi_n_881 ,csa_tree_add_107_22_pad_groupi_n_700 ,csa_tree_add_107_22_pad_groupi_n_828);
  or csa_tree_add_107_22_pad_groupi_g4845(csa_tree_add_107_22_pad_groupi_n_880 ,csa_tree_add_107_22_pad_groupi_n_761 ,csa_tree_add_107_22_pad_groupi_n_786);
  nor csa_tree_add_107_22_pad_groupi_g4846(csa_tree_add_107_22_pad_groupi_n_879 ,csa_tree_add_107_22_pad_groupi_n_371 ,csa_tree_add_107_22_pad_groupi_n_740);
  or csa_tree_add_107_22_pad_groupi_g4847(csa_tree_add_107_22_pad_groupi_n_878 ,csa_tree_add_107_22_pad_groupi_n_387 ,csa_tree_add_107_22_pad_groupi_n_712);
  and csa_tree_add_107_22_pad_groupi_g4848(csa_tree_add_107_22_pad_groupi_n_877 ,csa_tree_add_107_22_pad_groupi_n_766 ,csa_tree_add_107_22_pad_groupi_n_744);
  nor csa_tree_add_107_22_pad_groupi_g4849(csa_tree_add_107_22_pad_groupi_n_876 ,csa_tree_add_107_22_pad_groupi_n_733 ,csa_tree_add_107_22_pad_groupi_n_755);
  nor csa_tree_add_107_22_pad_groupi_g4850(csa_tree_add_107_22_pad_groupi_n_875 ,in25[7] ,csa_tree_add_107_22_pad_groupi_n_713);
  and csa_tree_add_107_22_pad_groupi_g4851(csa_tree_add_107_22_pad_groupi_n_874 ,csa_tree_add_107_22_pad_groupi_n_803 ,csa_tree_add_107_22_pad_groupi_n_721);
  and csa_tree_add_107_22_pad_groupi_g4852(csa_tree_add_107_22_pad_groupi_n_873 ,csa_tree_add_107_22_pad_groupi_n_758 ,csa_tree_add_107_22_pad_groupi_n_757);
  nor csa_tree_add_107_22_pad_groupi_g4853(csa_tree_add_107_22_pad_groupi_n_872 ,csa_tree_add_107_22_pad_groupi_n_764 ,csa_tree_add_107_22_pad_groupi_n_809);
  or csa_tree_add_107_22_pad_groupi_g4854(csa_tree_add_107_22_pad_groupi_n_871 ,csa_tree_add_107_22_pad_groupi_n_758 ,csa_tree_add_107_22_pad_groupi_n_757);
  and csa_tree_add_107_22_pad_groupi_g4855(csa_tree_add_107_22_pad_groupi_n_870 ,in25[2] ,csa_tree_add_107_22_pad_groupi_n_756);
  and csa_tree_add_107_22_pad_groupi_g4856(csa_tree_add_107_22_pad_groupi_n_869 ,csa_tree_add_107_22_pad_groupi_n_808 ,csa_tree_add_107_22_pad_groupi_n_788);
  and csa_tree_add_107_22_pad_groupi_g4857(csa_tree_add_107_22_pad_groupi_n_868 ,csa_tree_add_107_22_pad_groupi_n_784 ,csa_tree_add_107_22_pad_groupi_n_747);
  or csa_tree_add_107_22_pad_groupi_g4858(csa_tree_add_107_22_pad_groupi_n_867 ,csa_tree_add_107_22_pad_groupi_n_810 ,csa_tree_add_107_22_pad_groupi_n_811);
  and csa_tree_add_107_22_pad_groupi_g4859(csa_tree_add_107_22_pad_groupi_n_866 ,csa_tree_add_107_22_pad_groupi_n_765 ,csa_tree_add_107_22_pad_groupi_n_751);
  or csa_tree_add_107_22_pad_groupi_g4860(csa_tree_add_107_22_pad_groupi_n_865 ,csa_tree_add_107_22_pad_groupi_n_784 ,csa_tree_add_107_22_pad_groupi_n_747);
  or csa_tree_add_107_22_pad_groupi_g4861(csa_tree_add_107_22_pad_groupi_n_864 ,csa_tree_add_107_22_pad_groupi_n_749 ,csa_tree_add_107_22_pad_groupi_n_741);
  or csa_tree_add_107_22_pad_groupi_g4862(csa_tree_add_107_22_pad_groupi_n_863 ,csa_tree_add_107_22_pad_groupi_n_765 ,csa_tree_add_107_22_pad_groupi_n_751);
  nor csa_tree_add_107_22_pad_groupi_g4863(csa_tree_add_107_22_pad_groupi_n_862 ,csa_tree_add_107_22_pad_groupi_n_750 ,csa_tree_add_107_22_pad_groupi_n_742);
  nor csa_tree_add_107_22_pad_groupi_g4864(csa_tree_add_107_22_pad_groupi_n_861 ,csa_tree_add_107_22_pad_groupi_n_600 ,csa_tree_add_107_22_pad_groupi_n_822);
  or csa_tree_add_107_22_pad_groupi_g4865(csa_tree_add_107_22_pad_groupi_n_860 ,csa_tree_add_107_22_pad_groupi_n_726 ,csa_tree_add_107_22_pad_groupi_n_821);
  and csa_tree_add_107_22_pad_groupi_g4866(csa_tree_add_107_22_pad_groupi_n_859 ,csa_tree_add_107_22_pad_groupi_n_371 ,csa_tree_add_107_22_pad_groupi_n_740);
  and csa_tree_add_107_22_pad_groupi_g4867(csa_tree_add_107_22_pad_groupi_n_858 ,csa_tree_add_107_22_pad_groupi_n_726 ,csa_tree_add_107_22_pad_groupi_n_821);
  or csa_tree_add_107_22_pad_groupi_g4868(csa_tree_add_107_22_pad_groupi_n_857 ,csa_tree_add_107_22_pad_groupi_n_759 ,csa_tree_add_107_22_pad_groupi_n_736);
  or csa_tree_add_107_22_pad_groupi_g4869(csa_tree_add_107_22_pad_groupi_n_856 ,in25[4] ,csa_tree_add_107_22_pad_groupi_n_798);
  nor csa_tree_add_107_22_pad_groupi_g4870(csa_tree_add_107_22_pad_groupi_n_855 ,in25[2] ,csa_tree_add_107_22_pad_groupi_n_756);
  nor csa_tree_add_107_22_pad_groupi_g4871(csa_tree_add_107_22_pad_groupi_n_854 ,csa_tree_add_107_22_pad_groupi_n_760 ,csa_tree_add_107_22_pad_groupi_n_737);
  or csa_tree_add_107_22_pad_groupi_g4872(csa_tree_add_107_22_pad_groupi_n_853 ,csa_tree_add_107_22_pad_groupi_n_370 ,csa_tree_add_107_22_pad_groupi_n_730);
  or csa_tree_add_107_22_pad_groupi_g4873(csa_tree_add_107_22_pad_groupi_n_852 ,csa_tree_add_107_22_pad_groupi_n_724 ,csa_tree_add_107_22_pad_groupi_n_722);
  nor csa_tree_add_107_22_pad_groupi_g4874(csa_tree_add_107_22_pad_groupi_n_851 ,in25[6] ,csa_tree_add_107_22_pad_groupi_n_731);
  or csa_tree_add_107_22_pad_groupi_g4876(csa_tree_add_107_22_pad_groupi_n_893 ,csa_tree_add_107_22_pad_groupi_n_374 ,csa_tree_add_107_22_pad_groupi_n_826);
  or csa_tree_add_107_22_pad_groupi_g4877(csa_tree_add_107_22_pad_groupi_n_892 ,csa_tree_add_107_22_pad_groupi_n_847 ,csa_tree_add_107_22_pad_groupi_n_849);
  not csa_tree_add_107_22_pad_groupi_g4878(csa_tree_add_107_22_pad_groupi_n_849 ,csa_tree_add_107_22_pad_groupi_n_848);
  not csa_tree_add_107_22_pad_groupi_g4879(csa_tree_add_107_22_pad_groupi_n_847 ,csa_tree_add_107_22_pad_groupi_n_846);
  not csa_tree_add_107_22_pad_groupi_g4880(csa_tree_add_107_22_pad_groupi_n_843 ,csa_tree_add_107_22_pad_groupi_n_842);
  not csa_tree_add_107_22_pad_groupi_g4883(csa_tree_add_107_22_pad_groupi_n_833 ,csa_tree_add_107_22_pad_groupi_n_832);
  not csa_tree_add_107_22_pad_groupi_g4884(csa_tree_add_107_22_pad_groupi_n_826 ,csa_tree_add_107_22_pad_groupi_n_825);
  not csa_tree_add_107_22_pad_groupi_g4885(csa_tree_add_107_22_pad_groupi_n_818 ,csa_tree_add_107_22_pad_groupi_n_819);
  not csa_tree_add_107_22_pad_groupi_g4886(csa_tree_add_107_22_pad_groupi_n_816 ,csa_tree_add_107_22_pad_groupi_n_817);
  not csa_tree_add_107_22_pad_groupi_g4887(csa_tree_add_107_22_pad_groupi_n_812 ,csa_tree_add_107_22_pad_groupi_n_813);
  not csa_tree_add_107_22_pad_groupi_g4888(csa_tree_add_107_22_pad_groupi_n_805 ,csa_tree_add_107_22_pad_groupi_n_806);
  not csa_tree_add_107_22_pad_groupi_g4889(csa_tree_add_107_22_pad_groupi_n_801 ,csa_tree_add_107_22_pad_groupi_n_802);
  not csa_tree_add_107_22_pad_groupi_g4890(csa_tree_add_107_22_pad_groupi_n_794 ,csa_tree_add_107_22_pad_groupi_n_795);
  not csa_tree_add_107_22_pad_groupi_g4891(csa_tree_add_107_22_pad_groupi_n_791 ,csa_tree_add_107_22_pad_groupi_n_792);
  not csa_tree_add_107_22_pad_groupi_g4892(csa_tree_add_107_22_pad_groupi_n_789 ,csa_tree_add_107_22_pad_groupi_n_790);
  and csa_tree_add_107_22_pad_groupi_g4893(csa_tree_add_107_22_pad_groupi_n_781 ,csa_tree_add_107_22_pad_groupi_n_459 ,csa_tree_add_107_22_pad_groupi_n_612);
  or csa_tree_add_107_22_pad_groupi_g4894(csa_tree_add_107_22_pad_groupi_n_848 ,csa_tree_add_107_22_pad_groupi_n_466 ,csa_tree_add_107_22_pad_groupi_n_621);
  or csa_tree_add_107_22_pad_groupi_g4895(csa_tree_add_107_22_pad_groupi_n_846 ,csa_tree_add_107_22_pad_groupi_n_576 ,csa_tree_add_107_22_pad_groupi_n_703);
  and csa_tree_add_107_22_pad_groupi_g4896(csa_tree_add_107_22_pad_groupi_n_845 ,csa_tree_add_107_22_pad_groupi_n_531 ,csa_tree_add_107_22_pad_groupi_n_685);
  or csa_tree_add_107_22_pad_groupi_g4897(csa_tree_add_107_22_pad_groupi_n_844 ,csa_tree_add_107_22_pad_groupi_n_526 ,csa_tree_add_107_22_pad_groupi_n_652);
  or csa_tree_add_107_22_pad_groupi_g4898(csa_tree_add_107_22_pad_groupi_n_842 ,csa_tree_add_107_22_pad_groupi_n_533 ,csa_tree_add_107_22_pad_groupi_n_618);
  and csa_tree_add_107_22_pad_groupi_g4899(csa_tree_add_107_22_pad_groupi_n_841 ,csa_tree_add_107_22_pad_groupi_n_472 ,csa_tree_add_107_22_pad_groupi_n_642);
  or csa_tree_add_107_22_pad_groupi_g4900(csa_tree_add_107_22_pad_groupi_n_840 ,csa_tree_add_107_22_pad_groupi_n_557 ,csa_tree_add_107_22_pad_groupi_n_598);
  or csa_tree_add_107_22_pad_groupi_g4901(csa_tree_add_107_22_pad_groupi_n_839 ,csa_tree_add_107_22_pad_groupi_n_574 ,csa_tree_add_107_22_pad_groupi_n_588);
  and csa_tree_add_107_22_pad_groupi_g4903(csa_tree_add_107_22_pad_groupi_n_837 ,csa_tree_add_107_22_pad_groupi_n_483 ,csa_tree_add_107_22_pad_groupi_n_587);
  and csa_tree_add_107_22_pad_groupi_g4906(csa_tree_add_107_22_pad_groupi_n_834 ,csa_tree_add_107_22_pad_groupi_n_460 ,csa_tree_add_107_22_pad_groupi_n_586);
  or csa_tree_add_107_22_pad_groupi_g4907(csa_tree_add_107_22_pad_groupi_n_832 ,csa_tree_add_107_22_pad_groupi_n_548 ,csa_tree_add_107_22_pad_groupi_n_699);
  or csa_tree_add_107_22_pad_groupi_g4912(csa_tree_add_107_22_pad_groupi_n_827 ,csa_tree_add_107_22_pad_groupi_n_487 ,csa_tree_add_107_22_pad_groupi_n_647);
  or csa_tree_add_107_22_pad_groupi_g4913(csa_tree_add_107_22_pad_groupi_n_825 ,csa_tree_add_107_22_pad_groupi_n_462 ,csa_tree_add_107_22_pad_groupi_n_662);
  and csa_tree_add_107_22_pad_groupi_g4914(csa_tree_add_107_22_pad_groupi_n_824 ,csa_tree_add_107_22_pad_groupi_n_485 ,csa_tree_add_107_22_pad_groupi_n_683);
  and csa_tree_add_107_22_pad_groupi_g4915(csa_tree_add_107_22_pad_groupi_n_823 ,csa_tree_add_107_22_pad_groupi_n_518 ,csa_tree_add_107_22_pad_groupi_n_595);
  or csa_tree_add_107_22_pad_groupi_g4917(csa_tree_add_107_22_pad_groupi_n_821 ,csa_tree_add_107_22_pad_groupi_n_551 ,csa_tree_add_107_22_pad_groupi_n_665);
  or csa_tree_add_107_22_pad_groupi_g4918(csa_tree_add_107_22_pad_groupi_n_820 ,csa_tree_add_107_22_pad_groupi_n_556 ,csa_tree_add_107_22_pad_groupi_n_677);
  or csa_tree_add_107_22_pad_groupi_g4919(csa_tree_add_107_22_pad_groupi_n_819 ,csa_tree_add_107_22_pad_groupi_n_516 ,csa_tree_add_107_22_pad_groupi_n_681);
  or csa_tree_add_107_22_pad_groupi_g4920(csa_tree_add_107_22_pad_groupi_n_817 ,csa_tree_add_107_22_pad_groupi_n_527 ,csa_tree_add_107_22_pad_groupi_n_674);
  or csa_tree_add_107_22_pad_groupi_g4921(csa_tree_add_107_22_pad_groupi_n_815 ,csa_tree_add_107_22_pad_groupi_n_491 ,csa_tree_add_107_22_pad_groupi_n_649);
  or csa_tree_add_107_22_pad_groupi_g4922(csa_tree_add_107_22_pad_groupi_n_814 ,csa_tree_add_107_22_pad_groupi_n_475 ,csa_tree_add_107_22_pad_groupi_n_633);
  or csa_tree_add_107_22_pad_groupi_g4923(csa_tree_add_107_22_pad_groupi_n_813 ,csa_tree_add_107_22_pad_groupi_n_525 ,csa_tree_add_107_22_pad_groupi_n_695);
  or csa_tree_add_107_22_pad_groupi_g4924(csa_tree_add_107_22_pad_groupi_n_811 ,csa_tree_add_107_22_pad_groupi_n_476 ,csa_tree_add_107_22_pad_groupi_n_599);
  or csa_tree_add_107_22_pad_groupi_g4925(csa_tree_add_107_22_pad_groupi_n_810 ,csa_tree_add_107_22_pad_groupi_n_470 ,csa_tree_add_107_22_pad_groupi_n_627);
  or csa_tree_add_107_22_pad_groupi_g4926(csa_tree_add_107_22_pad_groupi_n_809 ,csa_tree_add_107_22_pad_groupi_n_528 ,csa_tree_add_107_22_pad_groupi_n_651);
  or csa_tree_add_107_22_pad_groupi_g4927(csa_tree_add_107_22_pad_groupi_n_808 ,csa_tree_add_107_22_pad_groupi_n_541 ,csa_tree_add_107_22_pad_groupi_n_635);
  or csa_tree_add_107_22_pad_groupi_g4928(csa_tree_add_107_22_pad_groupi_n_807 ,csa_tree_add_107_22_pad_groupi_n_512 ,csa_tree_add_107_22_pad_groupi_n_625);
  or csa_tree_add_107_22_pad_groupi_g4929(csa_tree_add_107_22_pad_groupi_n_806 ,csa_tree_add_107_22_pad_groupi_n_523 ,csa_tree_add_107_22_pad_groupi_n_623);
  or csa_tree_add_107_22_pad_groupi_g4930(csa_tree_add_107_22_pad_groupi_n_804 ,csa_tree_add_107_22_pad_groupi_n_461 ,csa_tree_add_107_22_pad_groupi_n_694);
  or csa_tree_add_107_22_pad_groupi_g4931(csa_tree_add_107_22_pad_groupi_n_803 ,csa_tree_add_107_22_pad_groupi_n_529 ,csa_tree_add_107_22_pad_groupi_n_653);
  or csa_tree_add_107_22_pad_groupi_g4933(csa_tree_add_107_22_pad_groupi_n_800 ,csa_tree_add_107_22_pad_groupi_n_477 ,csa_tree_add_107_22_pad_groupi_n_658);
  or csa_tree_add_107_22_pad_groupi_g4934(csa_tree_add_107_22_pad_groupi_n_799 ,csa_tree_add_107_22_pad_groupi_n_467 ,csa_tree_add_107_22_pad_groupi_n_680);
  or csa_tree_add_107_22_pad_groupi_g4935(csa_tree_add_107_22_pad_groupi_n_798 ,csa_tree_add_107_22_pad_groupi_n_468 ,csa_tree_add_107_22_pad_groupi_n_607);
  or csa_tree_add_107_22_pad_groupi_g4936(csa_tree_add_107_22_pad_groupi_n_797 ,csa_tree_add_107_22_pad_groupi_n_394 ,csa_tree_add_107_22_pad_groupi_n_663);
  or csa_tree_add_107_22_pad_groupi_g4937(csa_tree_add_107_22_pad_groupi_n_796 ,csa_tree_add_107_22_pad_groupi_n_555 ,csa_tree_add_107_22_pad_groupi_n_669);
  or csa_tree_add_107_22_pad_groupi_g4938(csa_tree_add_107_22_pad_groupi_n_795 ,csa_tree_add_107_22_pad_groupi_n_547 ,csa_tree_add_107_22_pad_groupi_n_696);
  or csa_tree_add_107_22_pad_groupi_g4939(csa_tree_add_107_22_pad_groupi_n_793 ,csa_tree_add_107_22_pad_groupi_n_540 ,csa_tree_add_107_22_pad_groupi_n_697);
  or csa_tree_add_107_22_pad_groupi_g4940(csa_tree_add_107_22_pad_groupi_n_792 ,csa_tree_add_107_22_pad_groupi_n_456 ,csa_tree_add_107_22_pad_groupi_n_638);
  or csa_tree_add_107_22_pad_groupi_g4941(csa_tree_add_107_22_pad_groupi_n_790 ,csa_tree_add_107_22_pad_groupi_n_524 ,csa_tree_add_107_22_pad_groupi_n_661);
  or csa_tree_add_107_22_pad_groupi_g4942(csa_tree_add_107_22_pad_groupi_n_788 ,csa_tree_add_107_22_pad_groupi_n_537 ,csa_tree_add_107_22_pad_groupi_n_616);
  or csa_tree_add_107_22_pad_groupi_g4943(csa_tree_add_107_22_pad_groupi_n_787 ,csa_tree_add_107_22_pad_groupi_n_469 ,csa_tree_add_107_22_pad_groupi_n_672);
  or csa_tree_add_107_22_pad_groupi_g4944(csa_tree_add_107_22_pad_groupi_n_786 ,csa_tree_add_107_22_pad_groupi_n_473 ,csa_tree_add_107_22_pad_groupi_n_589);
  or csa_tree_add_107_22_pad_groupi_g4945(csa_tree_add_107_22_pad_groupi_n_785 ,csa_tree_add_107_22_pad_groupi_n_484 ,csa_tree_add_107_22_pad_groupi_n_698);
  or csa_tree_add_107_22_pad_groupi_g4946(csa_tree_add_107_22_pad_groupi_n_784 ,csa_tree_add_107_22_pad_groupi_n_488 ,csa_tree_add_107_22_pad_groupi_n_608);
  or csa_tree_add_107_22_pad_groupi_g4947(csa_tree_add_107_22_pad_groupi_n_783 ,csa_tree_add_107_22_pad_groupi_n_546 ,csa_tree_add_107_22_pad_groupi_n_648);
  not csa_tree_add_107_22_pad_groupi_g4949(csa_tree_add_107_22_pad_groupi_n_779 ,csa_tree_add_107_22_pad_groupi_n_778);
  not csa_tree_add_107_22_pad_groupi_g4950(csa_tree_add_107_22_pad_groupi_n_762 ,csa_tree_add_107_22_pad_groupi_n_763);
  not csa_tree_add_107_22_pad_groupi_g4951(csa_tree_add_107_22_pad_groupi_n_759 ,csa_tree_add_107_22_pad_groupi_n_760);
  not csa_tree_add_107_22_pad_groupi_g4952(csa_tree_add_107_22_pad_groupi_n_754 ,csa_tree_add_107_22_pad_groupi_n_755);
  not csa_tree_add_107_22_pad_groupi_g4953(csa_tree_add_107_22_pad_groupi_n_752 ,csa_tree_add_107_22_pad_groupi_n_753);
  not csa_tree_add_107_22_pad_groupi_g4954(csa_tree_add_107_22_pad_groupi_n_749 ,csa_tree_add_107_22_pad_groupi_n_750);
  not csa_tree_add_107_22_pad_groupi_g4955(csa_tree_add_107_22_pad_groupi_n_745 ,csa_tree_add_107_22_pad_groupi_n_746);
  not csa_tree_add_107_22_pad_groupi_g4956(csa_tree_add_107_22_pad_groupi_n_744 ,csa_tree_add_107_22_pad_groupi_n_743);
  not csa_tree_add_107_22_pad_groupi_g4957(csa_tree_add_107_22_pad_groupi_n_741 ,csa_tree_add_107_22_pad_groupi_n_742);
  not csa_tree_add_107_22_pad_groupi_g4958(csa_tree_add_107_22_pad_groupi_n_738 ,csa_tree_add_107_22_pad_groupi_n_739);
  not csa_tree_add_107_22_pad_groupi_g4959(csa_tree_add_107_22_pad_groupi_n_736 ,csa_tree_add_107_22_pad_groupi_n_737);
  not csa_tree_add_107_22_pad_groupi_g4960(csa_tree_add_107_22_pad_groupi_n_734 ,csa_tree_add_107_22_pad_groupi_n_735);
  not csa_tree_add_107_22_pad_groupi_g4961(csa_tree_add_107_22_pad_groupi_n_732 ,csa_tree_add_107_22_pad_groupi_n_733);
  not csa_tree_add_107_22_pad_groupi_g4962(csa_tree_add_107_22_pad_groupi_n_730 ,csa_tree_add_107_22_pad_groupi_n_731);
  not csa_tree_add_107_22_pad_groupi_g4963(csa_tree_add_107_22_pad_groupi_n_727 ,csa_tree_add_107_22_pad_groupi_n_728);
  not csa_tree_add_107_22_pad_groupi_g4964(csa_tree_add_107_22_pad_groupi_n_724 ,csa_tree_add_107_22_pad_groupi_n_725);
  not csa_tree_add_107_22_pad_groupi_g4965(csa_tree_add_107_22_pad_groupi_n_722 ,csa_tree_add_107_22_pad_groupi_n_723);
  not csa_tree_add_107_22_pad_groupi_g4966(csa_tree_add_107_22_pad_groupi_n_715 ,csa_tree_add_107_22_pad_groupi_n_716);
  not csa_tree_add_107_22_pad_groupi_g4967(csa_tree_add_107_22_pad_groupi_n_712 ,csa_tree_add_107_22_pad_groupi_n_713);
  xnor csa_tree_add_107_22_pad_groupi_g4968(csa_tree_add_107_22_pad_groupi_n_711 ,csa_tree_add_107_22_pad_groupi_n_583 ,in25[10]);
  xnor csa_tree_add_107_22_pad_groupi_g4970(csa_tree_add_107_22_pad_groupi_n_710 ,csa_tree_add_107_22_pad_groupi_n_282 ,in25[12]);
  xnor csa_tree_add_107_22_pad_groupi_g4972(csa_tree_add_107_22_pad_groupi_n_709 ,csa_tree_add_107_22_pad_groupi_n_582 ,in25[12]);
  or csa_tree_add_107_22_pad_groupi_g4975(csa_tree_add_107_22_pad_groupi_n_778 ,csa_tree_add_107_22_pad_groupi_n_539 ,csa_tree_add_107_22_pad_groupi_n_626);
  or csa_tree_add_107_22_pad_groupi_g4976(csa_tree_add_107_22_pad_groupi_n_777 ,csa_tree_add_107_22_pad_groupi_n_550 ,csa_tree_add_107_22_pad_groupi_n_624);
  and csa_tree_add_107_22_pad_groupi_g4977(csa_tree_add_107_22_pad_groupi_n_776 ,csa_tree_add_107_22_pad_groupi_n_464 ,csa_tree_add_107_22_pad_groupi_n_655);
  or csa_tree_add_107_22_pad_groupi_g4978(csa_tree_add_107_22_pad_groupi_n_775 ,csa_tree_add_107_22_pad_groupi_n_482 ,csa_tree_add_107_22_pad_groupi_n_637);
  or csa_tree_add_107_22_pad_groupi_g4980(csa_tree_add_107_22_pad_groupi_n_773 ,csa_tree_add_107_22_pad_groupi_n_519 ,csa_tree_add_107_22_pad_groupi_n_605);
  and csa_tree_add_107_22_pad_groupi_g4981(csa_tree_add_107_22_pad_groupi_n_772 ,csa_tree_add_107_22_pad_groupi_n_457 ,csa_tree_add_107_22_pad_groupi_n_594);
  and csa_tree_add_107_22_pad_groupi_g4982(csa_tree_add_107_22_pad_groupi_n_771 ,csa_tree_add_107_22_pad_groupi_n_492 ,csa_tree_add_107_22_pad_groupi_n_606);
  or csa_tree_add_107_22_pad_groupi_g4984(csa_tree_add_107_22_pad_groupi_n_769 ,csa_tree_add_107_22_pad_groupi_n_490 ,csa_tree_add_107_22_pad_groupi_n_689);
  or csa_tree_add_107_22_pad_groupi_g4985(csa_tree_add_107_22_pad_groupi_n_768 ,csa_tree_add_107_22_pad_groupi_n_545 ,csa_tree_add_107_22_pad_groupi_n_640);
  or csa_tree_add_107_22_pad_groupi_g4986(csa_tree_add_107_22_pad_groupi_n_767 ,csa_tree_add_107_22_pad_groupi_n_552 ,csa_tree_add_107_22_pad_groupi_n_659);
  or csa_tree_add_107_22_pad_groupi_g4988(csa_tree_add_107_22_pad_groupi_n_765 ,csa_tree_add_107_22_pad_groupi_n_517 ,csa_tree_add_107_22_pad_groupi_n_688);
  or csa_tree_add_107_22_pad_groupi_g4989(csa_tree_add_107_22_pad_groupi_n_764 ,csa_tree_add_107_22_pad_groupi_n_554 ,csa_tree_add_107_22_pad_groupi_n_654);
  or csa_tree_add_107_22_pad_groupi_g4990(csa_tree_add_107_22_pad_groupi_n_763 ,csa_tree_add_107_22_pad_groupi_n_480 ,csa_tree_add_107_22_pad_groupi_n_602);
  or csa_tree_add_107_22_pad_groupi_g4991(csa_tree_add_107_22_pad_groupi_n_761 ,csa_tree_add_107_22_pad_groupi_n_577 ,csa_tree_add_107_22_pad_groupi_n_693);
  or csa_tree_add_107_22_pad_groupi_g4992(csa_tree_add_107_22_pad_groupi_n_760 ,csa_tree_add_107_22_pad_groupi_n_478 ,csa_tree_add_107_22_pad_groupi_n_591);
  or csa_tree_add_107_22_pad_groupi_g4993(csa_tree_add_107_22_pad_groupi_n_758 ,csa_tree_add_107_22_pad_groupi_n_514 ,csa_tree_add_107_22_pad_groupi_n_604);
  or csa_tree_add_107_22_pad_groupi_g4994(csa_tree_add_107_22_pad_groupi_n_757 ,csa_tree_add_107_22_pad_groupi_n_532 ,csa_tree_add_107_22_pad_groupi_n_617);
  or csa_tree_add_107_22_pad_groupi_g4995(csa_tree_add_107_22_pad_groupi_n_756 ,csa_tree_add_107_22_pad_groupi_n_455 ,csa_tree_add_107_22_pad_groupi_n_670);
  or csa_tree_add_107_22_pad_groupi_g4996(csa_tree_add_107_22_pad_groupi_n_755 ,csa_tree_add_107_22_pad_groupi_n_544 ,csa_tree_add_107_22_pad_groupi_n_660);
  or csa_tree_add_107_22_pad_groupi_g4997(csa_tree_add_107_22_pad_groupi_n_753 ,csa_tree_add_107_22_pad_groupi_n_486 ,csa_tree_add_107_22_pad_groupi_n_679);
  or csa_tree_add_107_22_pad_groupi_g4998(csa_tree_add_107_22_pad_groupi_n_751 ,csa_tree_add_107_22_pad_groupi_n_575 ,csa_tree_add_107_22_pad_groupi_n_619);
  or csa_tree_add_107_22_pad_groupi_g4999(csa_tree_add_107_22_pad_groupi_n_750 ,csa_tree_add_107_22_pad_groupi_n_522 ,csa_tree_add_107_22_pad_groupi_n_671);
  or csa_tree_add_107_22_pad_groupi_g5000(csa_tree_add_107_22_pad_groupi_n_748 ,csa_tree_add_107_22_pad_groupi_n_515 ,csa_tree_add_107_22_pad_groupi_n_631);
  or csa_tree_add_107_22_pad_groupi_g5001(csa_tree_add_107_22_pad_groupi_n_747 ,csa_tree_add_107_22_pad_groupi_n_573 ,csa_tree_add_107_22_pad_groupi_n_620);
  or csa_tree_add_107_22_pad_groupi_g5002(csa_tree_add_107_22_pad_groupi_n_746 ,csa_tree_add_107_22_pad_groupi_n_534 ,csa_tree_add_107_22_pad_groupi_n_643);
  or csa_tree_add_107_22_pad_groupi_g5003(csa_tree_add_107_22_pad_groupi_n_743 ,csa_tree_add_107_22_pad_groupi_n_481 ,csa_tree_add_107_22_pad_groupi_n_629);
  or csa_tree_add_107_22_pad_groupi_g5004(csa_tree_add_107_22_pad_groupi_n_742 ,csa_tree_add_107_22_pad_groupi_n_536 ,csa_tree_add_107_22_pad_groupi_n_650);
  or csa_tree_add_107_22_pad_groupi_g5006(csa_tree_add_107_22_pad_groupi_n_739 ,csa_tree_add_107_22_pad_groupi_n_564 ,csa_tree_add_107_22_pad_groupi_n_628);
  or csa_tree_add_107_22_pad_groupi_g5007(csa_tree_add_107_22_pad_groupi_n_737 ,csa_tree_add_107_22_pad_groupi_n_513 ,csa_tree_add_107_22_pad_groupi_n_603);
  or csa_tree_add_107_22_pad_groupi_g5008(csa_tree_add_107_22_pad_groupi_n_735 ,csa_tree_add_107_22_pad_groupi_n_553 ,csa_tree_add_107_22_pad_groupi_n_691);
  or csa_tree_add_107_22_pad_groupi_g5009(csa_tree_add_107_22_pad_groupi_n_733 ,csa_tree_add_107_22_pad_groupi_n_530 ,csa_tree_add_107_22_pad_groupi_n_622);
  or csa_tree_add_107_22_pad_groupi_g5010(csa_tree_add_107_22_pad_groupi_n_731 ,csa_tree_add_107_22_pad_groupi_n_463 ,csa_tree_add_107_22_pad_groupi_n_590);
  or csa_tree_add_107_22_pad_groupi_g5011(csa_tree_add_107_22_pad_groupi_n_729 ,csa_tree_add_107_22_pad_groupi_n_471 ,csa_tree_add_107_22_pad_groupi_n_610);
  or csa_tree_add_107_22_pad_groupi_g5012(csa_tree_add_107_22_pad_groupi_n_728 ,csa_tree_add_107_22_pad_groupi_n_520 ,csa_tree_add_107_22_pad_groupi_n_639);
  or csa_tree_add_107_22_pad_groupi_g5013(csa_tree_add_107_22_pad_groupi_n_726 ,csa_tree_add_107_22_pad_groupi_n_535 ,csa_tree_add_107_22_pad_groupi_n_690);
  or csa_tree_add_107_22_pad_groupi_g5014(csa_tree_add_107_22_pad_groupi_n_725 ,csa_tree_add_107_22_pad_groupi_n_538 ,csa_tree_add_107_22_pad_groupi_n_675);
  or csa_tree_add_107_22_pad_groupi_g5015(csa_tree_add_107_22_pad_groupi_n_723 ,csa_tree_add_107_22_pad_groupi_n_543 ,csa_tree_add_107_22_pad_groupi_n_676);
  or csa_tree_add_107_22_pad_groupi_g5016(csa_tree_add_107_22_pad_groupi_n_721 ,csa_tree_add_107_22_pad_groupi_n_542 ,csa_tree_add_107_22_pad_groupi_n_634);
  or csa_tree_add_107_22_pad_groupi_g5017(csa_tree_add_107_22_pad_groupi_n_720 ,csa_tree_add_107_22_pad_groupi_n_479 ,csa_tree_add_107_22_pad_groupi_n_644);
  or csa_tree_add_107_22_pad_groupi_g5018(csa_tree_add_107_22_pad_groupi_n_719 ,csa_tree_add_107_22_pad_groupi_n_521 ,csa_tree_add_107_22_pad_groupi_n_611);
  or csa_tree_add_107_22_pad_groupi_g5019(csa_tree_add_107_22_pad_groupi_n_718 ,csa_tree_add_107_22_pad_groupi_n_489 ,csa_tree_add_107_22_pad_groupi_n_609);
  or csa_tree_add_107_22_pad_groupi_g5020(csa_tree_add_107_22_pad_groupi_n_717 ,csa_tree_add_107_22_pad_groupi_n_549 ,csa_tree_add_107_22_pad_groupi_n_692);
  or csa_tree_add_107_22_pad_groupi_g5021(csa_tree_add_107_22_pad_groupi_n_716 ,csa_tree_add_107_22_pad_groupi_n_465 ,csa_tree_add_107_22_pad_groupi_n_613);
  or csa_tree_add_107_22_pad_groupi_g5022(csa_tree_add_107_22_pad_groupi_n_714 ,csa_tree_add_107_22_pad_groupi_n_474 ,csa_tree_add_107_22_pad_groupi_n_657);
  or csa_tree_add_107_22_pad_groupi_g5023(csa_tree_add_107_22_pad_groupi_n_713 ,csa_tree_add_107_22_pad_groupi_n_458 ,csa_tree_add_107_22_pad_groupi_n_667);
  not csa_tree_add_107_22_pad_groupi_g5024(csa_tree_add_107_22_pad_groupi_n_707 ,csa_tree_add_107_22_pad_groupi_n_706);
  not csa_tree_add_107_22_pad_groupi_g5025(csa_tree_add_107_22_pad_groupi_n_705 ,csa_tree_add_107_22_pad_groupi_n_704);
  nor csa_tree_add_107_22_pad_groupi_g5026(csa_tree_add_107_22_pad_groupi_n_703 ,csa_tree_add_107_22_pad_groupi_n_113 ,csa_tree_add_107_22_pad_groupi_n_218);
  nor csa_tree_add_107_22_pad_groupi_g5027(csa_tree_add_107_22_pad_groupi_n_702 ,in25[9] ,csa_tree_add_107_22_pad_groupi_n_358);
  nor csa_tree_add_107_22_pad_groupi_g5029(csa_tree_add_107_22_pad_groupi_n_700 ,in25[12] ,csa_tree_add_107_22_pad_groupi_n_579);
  nor csa_tree_add_107_22_pad_groupi_g5030(csa_tree_add_107_22_pad_groupi_n_699 ,csa_tree_add_107_22_pad_groupi_n_115 ,csa_tree_add_107_22_pad_groupi_n_189);
  and csa_tree_add_107_22_pad_groupi_g5031(csa_tree_add_107_22_pad_groupi_n_698 ,in9[5] ,csa_tree_add_107_22_pad_groupi_n_172);
  nor csa_tree_add_107_22_pad_groupi_g5032(csa_tree_add_107_22_pad_groupi_n_697 ,csa_tree_add_107_22_pad_groupi_n_119 ,csa_tree_add_107_22_pad_groupi_n_38);
  nor csa_tree_add_107_22_pad_groupi_g5033(csa_tree_add_107_22_pad_groupi_n_696 ,csa_tree_add_107_22_pad_groupi_n_93 ,csa_tree_add_107_22_pad_groupi_n_66);
  and csa_tree_add_107_22_pad_groupi_g5034(csa_tree_add_107_22_pad_groupi_n_695 ,in9[2] ,csa_tree_add_107_22_pad_groupi_n_133);
  and csa_tree_add_107_22_pad_groupi_g5035(csa_tree_add_107_22_pad_groupi_n_694 ,in9[10] ,csa_tree_add_107_22_pad_groupi_n_433);
  and csa_tree_add_107_22_pad_groupi_g5036(csa_tree_add_107_22_pad_groupi_n_693 ,in9[8] ,csa_tree_add_107_22_pad_groupi_n_287);
  and csa_tree_add_107_22_pad_groupi_g5037(csa_tree_add_107_22_pad_groupi_n_692 ,in9[14] ,csa_tree_add_107_22_pad_groupi_n_169);
  and csa_tree_add_107_22_pad_groupi_g5038(csa_tree_add_107_22_pad_groupi_n_691 ,in9[1] ,csa_tree_add_107_22_pad_groupi_n_168);
  and csa_tree_add_107_22_pad_groupi_g5039(csa_tree_add_107_22_pad_groupi_n_690 ,in9[5] ,csa_tree_add_107_22_pad_groupi_n_142);
  and csa_tree_add_107_22_pad_groupi_g5040(csa_tree_add_107_22_pad_groupi_n_689 ,in9[7] ,csa_tree_add_107_22_pad_groupi_n_126);
  and csa_tree_add_107_22_pad_groupi_g5041(csa_tree_add_107_22_pad_groupi_n_688 ,in9[11] ,csa_tree_add_107_22_pad_groupi_n_285);
  or csa_tree_add_107_22_pad_groupi_g5044(csa_tree_add_107_22_pad_groupi_n_685 ,csa_tree_add_107_22_pad_groupi_n_17 ,csa_tree_add_107_22_pad_groupi_n_118);
  or csa_tree_add_107_22_pad_groupi_g5046(csa_tree_add_107_22_pad_groupi_n_683 ,csa_tree_add_107_22_pad_groupi_n_149 ,csa_tree_add_107_22_pad_groupi_n_583);
  and csa_tree_add_107_22_pad_groupi_g5047(csa_tree_add_107_22_pad_groupi_n_682 ,in25[12] ,csa_tree_add_107_22_pad_groupi_n_579);
  and csa_tree_add_107_22_pad_groupi_g5048(csa_tree_add_107_22_pad_groupi_n_681 ,in9[11] ,csa_tree_add_107_22_pad_groupi_n_135);
  and csa_tree_add_107_22_pad_groupi_g5049(csa_tree_add_107_22_pad_groupi_n_680 ,in9[6] ,csa_tree_add_107_22_pad_groupi_n_445);
  nor csa_tree_add_107_22_pad_groupi_g5050(csa_tree_add_107_22_pad_groupi_n_679 ,csa_tree_add_107_22_pad_groupi_n_252 ,csa_tree_add_107_22_pad_groupi_n_223);
  and csa_tree_add_107_22_pad_groupi_g5052(csa_tree_add_107_22_pad_groupi_n_677 ,in9[3] ,csa_tree_add_107_22_pad_groupi_n_139);
  and csa_tree_add_107_22_pad_groupi_g5053(csa_tree_add_107_22_pad_groupi_n_676 ,in9[6] ,csa_tree_add_107_22_pad_groupi_n_136);
  and csa_tree_add_107_22_pad_groupi_g5054(csa_tree_add_107_22_pad_groupi_n_675 ,in9[4] ,csa_tree_add_107_22_pad_groupi_n_144);
  and csa_tree_add_107_22_pad_groupi_g5055(csa_tree_add_107_22_pad_groupi_n_674 ,in9[4] ,csa_tree_add_107_22_pad_groupi_n_138);
  nor csa_tree_add_107_22_pad_groupi_g5056(csa_tree_add_107_22_pad_groupi_n_673 ,csa_tree_add_107_22_pad_groupi_n_369 ,csa_tree_add_107_22_pad_groupi_n_581);
  and csa_tree_add_107_22_pad_groupi_g5057(csa_tree_add_107_22_pad_groupi_n_672 ,in9[12] ,csa_tree_add_107_22_pad_groupi_n_428);
  and csa_tree_add_107_22_pad_groupi_g5058(csa_tree_add_107_22_pad_groupi_n_671 ,in9[4] ,csa_tree_add_107_22_pad_groupi_n_124);
  and csa_tree_add_107_22_pad_groupi_g5059(csa_tree_add_107_22_pad_groupi_n_670 ,in9[9] ,csa_tree_add_107_22_pad_groupi_n_439);
  and csa_tree_add_107_22_pad_groupi_g5060(csa_tree_add_107_22_pad_groupi_n_669 ,in9[14] ,csa_tree_add_107_22_pad_groupi_n_288);
  and csa_tree_add_107_22_pad_groupi_g5062(csa_tree_add_107_22_pad_groupi_n_667 ,in9[14] ,csa_tree_add_107_22_pad_groupi_n_425);
  and csa_tree_add_107_22_pad_groupi_g5063(csa_tree_add_107_22_pad_groupi_n_666 ,in25[12] ,csa_tree_add_107_22_pad_groupi_n_280);
  and csa_tree_add_107_22_pad_groupi_g5064(csa_tree_add_107_22_pad_groupi_n_665 ,in9[7] ,csa_tree_add_107_22_pad_groupi_n_171);
  and csa_tree_add_107_22_pad_groupi_g5066(csa_tree_add_107_22_pad_groupi_n_663 ,csa_tree_add_107_22_pad_groupi_n_406 ,csa_tree_add_107_22_pad_groupi_n_583);
  and csa_tree_add_107_22_pad_groupi_g5067(csa_tree_add_107_22_pad_groupi_n_662 ,in9[7] ,csa_tree_add_107_22_pad_groupi_n_429);
  and csa_tree_add_107_22_pad_groupi_g5068(csa_tree_add_107_22_pad_groupi_n_661 ,in9[9] ,csa_tree_add_107_22_pad_groupi_n_145);
  and csa_tree_add_107_22_pad_groupi_g5069(csa_tree_add_107_22_pad_groupi_n_660 ,in9[14] ,csa_tree_add_107_22_pad_groupi_n_127);
  nor csa_tree_add_107_22_pad_groupi_g5070(csa_tree_add_107_22_pad_groupi_n_659 ,csa_tree_add_107_22_pad_groupi_n_112 ,csa_tree_add_107_22_pad_groupi_n_202);
  and csa_tree_add_107_22_pad_groupi_g5071(csa_tree_add_107_22_pad_groupi_n_658 ,in9[3] ,csa_tree_add_107_22_pad_groupi_n_133);
  nor csa_tree_add_107_22_pad_groupi_g5072(csa_tree_add_107_22_pad_groupi_n_657 ,csa_tree_add_107_22_pad_groupi_n_118 ,csa_tree_add_107_22_pad_groupi_n_215);
  or csa_tree_add_107_22_pad_groupi_g5073(csa_tree_add_107_22_pad_groupi_n_656 ,csa_tree_add_107_22_pad_groupi_n_373 ,csa_tree_add_107_22_pad_groupi_n_357);
  or csa_tree_add_107_22_pad_groupi_g5074(csa_tree_add_107_22_pad_groupi_n_655 ,csa_tree_add_107_22_pad_groupi_n_27 ,csa_tree_add_107_22_pad_groupi_n_427);
  and csa_tree_add_107_22_pad_groupi_g5075(csa_tree_add_107_22_pad_groupi_n_654 ,in9[11] ,csa_tree_add_107_22_pad_groupi_n_130);
  and csa_tree_add_107_22_pad_groupi_g5076(csa_tree_add_107_22_pad_groupi_n_653 ,in9[1] ,csa_tree_add_107_22_pad_groupi_n_147);
  nor csa_tree_add_107_22_pad_groupi_g5077(csa_tree_add_107_22_pad_groupi_n_652 ,csa_tree_add_107_22_pad_groupi_n_93 ,csa_tree_add_107_22_pad_groupi_n_74);
  and csa_tree_add_107_22_pad_groupi_g5078(csa_tree_add_107_22_pad_groupi_n_651 ,in9[13] ,csa_tree_add_107_22_pad_groupi_n_148);
  and csa_tree_add_107_22_pad_groupi_g5079(csa_tree_add_107_22_pad_groupi_n_650 ,in9[6] ,csa_tree_add_107_22_pad_groupi_n_148);
  and csa_tree_add_107_22_pad_groupi_g5080(csa_tree_add_107_22_pad_groupi_n_649 ,in9[12] ,csa_tree_add_107_22_pad_groupi_n_142);
  and csa_tree_add_107_22_pad_groupi_g5081(csa_tree_add_107_22_pad_groupi_n_648 ,in9[3] ,csa_tree_add_107_22_pad_groupi_n_129);
  and csa_tree_add_107_22_pad_groupi_g5082(csa_tree_add_107_22_pad_groupi_n_647 ,in9[4] ,csa_tree_add_107_22_pad_groupi_n_284);
  or csa_tree_add_107_22_pad_groupi_g5084(csa_tree_add_107_22_pad_groupi_n_706 ,csa_tree_add_107_22_pad_groupi_n_24 ,csa_tree_add_107_22_pad_groupi_n_502);
  or csa_tree_add_107_22_pad_groupi_g5085(csa_tree_add_107_22_pad_groupi_n_704 ,csa_tree_add_107_22_pad_groupi_n_24 ,csa_tree_add_107_22_pad_groupi_n_257);
  nor csa_tree_add_107_22_pad_groupi_g5086(csa_tree_add_107_22_pad_groupi_n_644 ,csa_tree_add_107_22_pad_groupi_n_113 ,csa_tree_add_107_22_pad_groupi_n_178);
  nor csa_tree_add_107_22_pad_groupi_g5087(csa_tree_add_107_22_pad_groupi_n_643 ,csa_tree_add_107_22_pad_groupi_n_160 ,csa_tree_add_107_22_pad_groupi_n_578);
  or csa_tree_add_107_22_pad_groupi_g5088(csa_tree_add_107_22_pad_groupi_n_642 ,csa_tree_add_107_22_pad_groupi_n_47 ,csa_tree_add_107_22_pad_groupi_n_497);
  and csa_tree_add_107_22_pad_groupi_g5090(csa_tree_add_107_22_pad_groupi_n_640 ,in9[6] ,csa_tree_add_107_22_pad_groupi_n_130);
  and csa_tree_add_107_22_pad_groupi_g5091(csa_tree_add_107_22_pad_groupi_n_639 ,in9[13] ,csa_tree_add_107_22_pad_groupi_n_171);
  nor csa_tree_add_107_22_pad_groupi_g5092(csa_tree_add_107_22_pad_groupi_n_638 ,csa_tree_add_107_22_pad_groupi_n_87 ,csa_tree_add_107_22_pad_groupi_n_434);
  and csa_tree_add_107_22_pad_groupi_g5093(csa_tree_add_107_22_pad_groupi_n_637 ,in9[10] ,csa_tree_add_107_22_pad_groupi_n_166);
  nor csa_tree_add_107_22_pad_groupi_g5095(csa_tree_add_107_22_pad_groupi_n_635 ,csa_tree_add_107_22_pad_groupi_n_96 ,csa_tree_add_107_22_pad_groupi_n_255);
  and csa_tree_add_107_22_pad_groupi_g5096(csa_tree_add_107_22_pad_groupi_n_634 ,in9[2] ,csa_tree_add_107_22_pad_groupi_n_168);
  and csa_tree_add_107_22_pad_groupi_g5097(csa_tree_add_107_22_pad_groupi_n_633 ,in9[13] ,csa_tree_add_107_22_pad_groupi_n_124);
  nor csa_tree_add_107_22_pad_groupi_g5099(csa_tree_add_107_22_pad_groupi_n_631 ,csa_tree_add_107_22_pad_groupi_n_231 ,csa_tree_add_107_22_pad_groupi_n_257);
  and csa_tree_add_107_22_pad_groupi_g5101(csa_tree_add_107_22_pad_groupi_n_629 ,in9[13] ,csa_tree_add_107_22_pad_groupi_n_287);
  and csa_tree_add_107_22_pad_groupi_g5102(csa_tree_add_107_22_pad_groupi_n_628 ,in9[11] ,csa_tree_add_107_22_pad_groupi_n_145);
  and csa_tree_add_107_22_pad_groupi_g5103(csa_tree_add_107_22_pad_groupi_n_627 ,in9[7] ,csa_tree_add_107_22_pad_groupi_n_141);
  nor csa_tree_add_107_22_pad_groupi_g5104(csa_tree_add_107_22_pad_groupi_n_626 ,csa_tree_add_107_22_pad_groupi_n_71 ,csa_tree_add_107_22_pad_groupi_n_507);
  and csa_tree_add_107_22_pad_groupi_g5105(csa_tree_add_107_22_pad_groupi_n_625 ,in9[7] ,csa_tree_add_107_22_pad_groupi_n_285);
  and csa_tree_add_107_22_pad_groupi_g5106(csa_tree_add_107_22_pad_groupi_n_624 ,in9[5] ,csa_tree_add_107_22_pad_groupi_n_165);
  and csa_tree_add_107_22_pad_groupi_g5107(csa_tree_add_107_22_pad_groupi_n_623 ,in9[10] ,csa_tree_add_107_22_pad_groupi_n_132);
  nor csa_tree_add_107_22_pad_groupi_g5108(csa_tree_add_107_22_pad_groupi_n_622 ,csa_tree_add_107_22_pad_groupi_n_159 ,csa_tree_add_107_22_pad_groupi_n_282);
  nor csa_tree_add_107_22_pad_groupi_g5109(csa_tree_add_107_22_pad_groupi_n_621 ,csa_tree_add_107_22_pad_groupi_n_98 ,csa_tree_add_107_22_pad_groupi_n_430);
  nor csa_tree_add_107_22_pad_groupi_g5110(csa_tree_add_107_22_pad_groupi_n_620 ,csa_tree_add_107_22_pad_groupi_n_194 ,csa_tree_add_107_22_pad_groupi_n_502);
  nor csa_tree_add_107_22_pad_groupi_g5111(csa_tree_add_107_22_pad_groupi_n_619 ,csa_tree_add_107_22_pad_groupi_n_116 ,csa_tree_add_107_22_pad_groupi_n_187);
  and csa_tree_add_107_22_pad_groupi_g5112(csa_tree_add_107_22_pad_groupi_n_618 ,in9[8] ,csa_tree_add_107_22_pad_groupi_n_165);
  and csa_tree_add_107_22_pad_groupi_g5113(csa_tree_add_107_22_pad_groupi_n_617 ,in9[8] ,csa_tree_add_107_22_pad_groupi_n_136);
  nor csa_tree_add_107_22_pad_groupi_g5114(csa_tree_add_107_22_pad_groupi_n_616 ,csa_tree_add_107_22_pad_groupi_n_119 ,csa_tree_add_107_22_pad_groupi_n_181);
  nor csa_tree_add_107_22_pad_groupi_g5117(csa_tree_add_107_22_pad_groupi_n_613 ,csa_tree_add_107_22_pad_groupi_n_204 ,csa_tree_add_107_22_pad_groupi_n_432);
  or csa_tree_add_107_22_pad_groupi_g5118(csa_tree_add_107_22_pad_groupi_n_612 ,csa_tree_add_107_22_pad_groupi_n_64 ,csa_tree_add_107_22_pad_groupi_n_438);
  and csa_tree_add_107_22_pad_groupi_g5119(csa_tree_add_107_22_pad_groupi_n_611 ,in9[8] ,csa_tree_add_107_22_pad_groupi_n_284);
  nor csa_tree_add_107_22_pad_groupi_g5120(csa_tree_add_107_22_pad_groupi_n_610 ,csa_tree_add_107_22_pad_groupi_n_116 ,csa_tree_add_107_22_pad_groupi_n_184);
  nor csa_tree_add_107_22_pad_groupi_g5121(csa_tree_add_107_22_pad_groupi_n_609 ,csa_tree_add_107_22_pad_groupi_n_91 ,csa_tree_add_107_22_pad_groupi_n_501);
  and csa_tree_add_107_22_pad_groupi_g5122(csa_tree_add_107_22_pad_groupi_n_608 ,in9[12] ,csa_tree_add_107_22_pad_groupi_n_166);
  and csa_tree_add_107_22_pad_groupi_g5123(csa_tree_add_107_22_pad_groupi_n_607 ,in9[11] ,csa_tree_add_107_22_pad_groupi_n_431);
  or csa_tree_add_107_22_pad_groupi_g5124(csa_tree_add_107_22_pad_groupi_n_606 ,csa_tree_add_107_22_pad_groupi_n_17 ,csa_tree_add_107_22_pad_groupi_n_255);
  and csa_tree_add_107_22_pad_groupi_g5125(csa_tree_add_107_22_pad_groupi_n_605 ,in9[9] ,csa_tree_add_107_22_pad_groupi_n_127);
  nor csa_tree_add_107_22_pad_groupi_g5126(csa_tree_add_107_22_pad_groupi_n_604 ,csa_tree_add_107_22_pad_groupi_n_211 ,csa_tree_add_107_22_pad_groupi_n_508);
  and csa_tree_add_107_22_pad_groupi_g5127(csa_tree_add_107_22_pad_groupi_n_603 ,in9[12] ,csa_tree_add_107_22_pad_groupi_n_169);
  and csa_tree_add_107_22_pad_groupi_g5128(csa_tree_add_107_22_pad_groupi_n_602 ,in9[1] ,csa_tree_add_107_22_pad_groupi_n_123);
  nor csa_tree_add_107_22_pad_groupi_g5130(csa_tree_add_107_22_pad_groupi_n_600 ,in25[12] ,csa_tree_add_107_22_pad_groupi_n_582);
  and csa_tree_add_107_22_pad_groupi_g5131(csa_tree_add_107_22_pad_groupi_n_599 ,in9[9] ,csa_tree_add_107_22_pad_groupi_n_139);
  nor csa_tree_add_107_22_pad_groupi_g5132(csa_tree_add_107_22_pad_groupi_n_598 ,csa_tree_add_107_22_pad_groupi_n_101 ,csa_tree_add_107_22_pad_groupi_n_508);
  or csa_tree_add_107_22_pad_groupi_g5135(csa_tree_add_107_22_pad_groupi_n_595 ,csa_tree_add_107_22_pad_groupi_n_55 ,csa_tree_add_107_22_pad_groupi_n_115);
  or csa_tree_add_107_22_pad_groupi_g5136(csa_tree_add_107_22_pad_groupi_n_594 ,csa_tree_add_107_22_pad_groupi_n_50 ,csa_tree_add_107_22_pad_groupi_n_426);
  nor csa_tree_add_107_22_pad_groupi_g5137(csa_tree_add_107_22_pad_groupi_n_593 ,in25[11] ,csa_tree_add_107_22_pad_groupi_n_580);
  and csa_tree_add_107_22_pad_groupi_g5139(csa_tree_add_107_22_pad_groupi_n_591 ,in9[10] ,csa_tree_add_107_22_pad_groupi_n_288);
  and csa_tree_add_107_22_pad_groupi_g5140(csa_tree_add_107_22_pad_groupi_n_590 ,in9[13] ,csa_tree_add_107_22_pad_groupi_n_435);
  and csa_tree_add_107_22_pad_groupi_g5141(csa_tree_add_107_22_pad_groupi_n_589 ,in9[10] ,csa_tree_add_107_22_pad_groupi_n_172);
  nor csa_tree_add_107_22_pad_groupi_g5142(csa_tree_add_107_22_pad_groupi_n_588 ,csa_tree_add_107_22_pad_groupi_n_158 ,csa_tree_add_107_22_pad_groupi_n_280);
  or csa_tree_add_107_22_pad_groupi_g5143(csa_tree_add_107_22_pad_groupi_n_587 ,csa_tree_add_107_22_pad_groupi_n_151 ,csa_tree_add_107_22_pad_groupi_n_580);
  or csa_tree_add_107_22_pad_groupi_g5144(csa_tree_add_107_22_pad_groupi_n_586 ,csa_tree_add_107_22_pad_groupi_n_15 ,csa_tree_add_107_22_pad_groupi_n_581);
  or csa_tree_add_107_22_pad_groupi_g5145(csa_tree_add_107_22_pad_groupi_n_646 ,csa_tree_add_107_22_pad_groupi_n_57 ,csa_tree_add_107_22_pad_groupi_n_493);
  or csa_tree_add_107_22_pad_groupi_g5146(csa_tree_add_107_22_pad_groupi_n_645 ,csa_tree_add_107_22_pad_groupi_n_42 ,csa_tree_add_107_22_pad_groupi_n_278);
  nor csa_tree_add_107_22_pad_groupi_g5150(csa_tree_add_107_22_pad_groupi_n_577 ,csa_tree_add_107_22_pad_groupi_n_183 ,csa_tree_add_107_22_pad_groupi_n_332);
  nor csa_tree_add_107_22_pad_groupi_g5151(csa_tree_add_107_22_pad_groupi_n_576 ,csa_tree_add_107_22_pad_groupi_n_42 ,csa_tree_add_107_22_pad_groupi_n_302);
  nor csa_tree_add_107_22_pad_groupi_g5152(csa_tree_add_107_22_pad_groupi_n_575 ,csa_tree_add_107_22_pad_groupi_n_233 ,csa_tree_add_107_22_pad_groupi_n_306);
  nor csa_tree_add_107_22_pad_groupi_g5153(csa_tree_add_107_22_pad_groupi_n_574 ,csa_tree_add_107_22_pad_groupi_n_193 ,csa_tree_add_107_22_pad_groupi_n_341);
  nor csa_tree_add_107_22_pad_groupi_g5154(csa_tree_add_107_22_pad_groupi_n_573 ,csa_tree_add_107_22_pad_groupi_n_84 ,csa_tree_add_107_22_pad_groupi_n_312);
  nor csa_tree_add_107_22_pad_groupi_g5163(csa_tree_add_107_22_pad_groupi_n_564 ,csa_tree_add_107_22_pad_groupi_n_78 ,csa_tree_add_107_22_pad_groupi_n_330);
  nor csa_tree_add_107_22_pad_groupi_g5170(csa_tree_add_107_22_pad_groupi_n_557 ,csa_tree_add_107_22_pad_groupi_n_71 ,csa_tree_add_107_22_pad_groupi_n_335);
  nor csa_tree_add_107_22_pad_groupi_g5171(csa_tree_add_107_22_pad_groupi_n_556 ,csa_tree_add_107_22_pad_groupi_n_101 ,csa_tree_add_107_22_pad_groupi_n_315);
  nor csa_tree_add_107_22_pad_groupi_g5172(csa_tree_add_107_22_pad_groupi_n_555 ,csa_tree_add_107_22_pad_groupi_n_186 ,csa_tree_add_107_22_pad_groupi_n_336);
  nor csa_tree_add_107_22_pad_groupi_g5173(csa_tree_add_107_22_pad_groupi_n_554 ,csa_tree_add_107_22_pad_groupi_n_177 ,csa_tree_add_107_22_pad_groupi_n_309);
  nor csa_tree_add_107_22_pad_groupi_g5174(csa_tree_add_107_22_pad_groupi_n_553 ,csa_tree_add_107_22_pad_groupi_n_244 ,csa_tree_add_107_22_pad_groupi_n_320);
  nor csa_tree_add_107_22_pad_groupi_g5175(csa_tree_add_107_22_pad_groupi_n_552 ,csa_tree_add_107_22_pad_groupi_n_247 ,csa_tree_add_107_22_pad_groupi_n_323);
  nor csa_tree_add_107_22_pad_groupi_g5176(csa_tree_add_107_22_pad_groupi_n_551 ,csa_tree_add_107_22_pad_groupi_n_67 ,csa_tree_add_107_22_pad_groupi_n_317);
  nor csa_tree_add_107_22_pad_groupi_g5177(csa_tree_add_107_22_pad_groupi_n_550 ,csa_tree_add_107_22_pad_groupi_n_175 ,csa_tree_add_107_22_pad_groupi_n_339);
  nor csa_tree_add_107_22_pad_groupi_g5178(csa_tree_add_107_22_pad_groupi_n_549 ,csa_tree_add_107_22_pad_groupi_n_85 ,csa_tree_add_107_22_pad_groupi_n_321);
  nor csa_tree_add_107_22_pad_groupi_g5179(csa_tree_add_107_22_pad_groupi_n_548 ,csa_tree_add_107_22_pad_groupi_n_88 ,csa_tree_add_107_22_pad_groupi_n_305);
  nor csa_tree_add_107_22_pad_groupi_g5180(csa_tree_add_107_22_pad_groupi_n_547 ,csa_tree_add_107_22_pad_groupi_n_197 ,csa_tree_add_107_22_pad_groupi_n_323);
  nor csa_tree_add_107_22_pad_groupi_g5181(csa_tree_add_107_22_pad_groupi_n_546 ,csa_tree_add_107_22_pad_groupi_n_100 ,csa_tree_add_107_22_pad_groupi_n_326);
  nor csa_tree_add_107_22_pad_groupi_g5182(csa_tree_add_107_22_pad_groupi_n_545 ,csa_tree_add_107_22_pad_groupi_n_53 ,csa_tree_add_107_22_pad_groupi_n_327);
  nor csa_tree_add_107_22_pad_groupi_g5183(csa_tree_add_107_22_pad_groupi_n_544 ,csa_tree_add_107_22_pad_groupi_n_187 ,csa_tree_add_107_22_pad_groupi_n_326);
  nor csa_tree_add_107_22_pad_groupi_g5184(csa_tree_add_107_22_pad_groupi_n_543 ,csa_tree_add_107_22_pad_groupi_n_196 ,csa_tree_add_107_22_pad_groupi_n_317);
  nor csa_tree_add_107_22_pad_groupi_g5185(csa_tree_add_107_22_pad_groupi_n_542 ,csa_tree_add_107_22_pad_groupi_n_217 ,csa_tree_add_107_22_pad_groupi_n_318);
  nor csa_tree_add_107_22_pad_groupi_g5186(csa_tree_add_107_22_pad_groupi_n_541 ,csa_tree_add_107_22_pad_groupi_n_209 ,csa_tree_add_107_22_pad_groupi_n_344);
  nor csa_tree_add_107_22_pad_groupi_g5187(csa_tree_add_107_22_pad_groupi_n_540 ,csa_tree_add_107_22_pad_groupi_n_229 ,csa_tree_add_107_22_pad_groupi_n_324);
  nor csa_tree_add_107_22_pad_groupi_g5188(csa_tree_add_107_22_pad_groupi_n_539 ,csa_tree_add_107_22_pad_groupi_n_41 ,csa_tree_add_107_22_pad_groupi_n_335);
  nor csa_tree_add_107_22_pad_groupi_g5189(csa_tree_add_107_22_pad_groupi_n_538 ,csa_tree_add_107_22_pad_groupi_n_36 ,csa_tree_add_107_22_pad_groupi_n_336);
  nor csa_tree_add_107_22_pad_groupi_g5190(csa_tree_add_107_22_pad_groupi_n_537 ,csa_tree_add_107_22_pad_groupi_n_79 ,csa_tree_add_107_22_pad_groupi_n_324);
  nor csa_tree_add_107_22_pad_groupi_g5191(csa_tree_add_107_22_pad_groupi_n_536 ,csa_tree_add_107_22_pad_groupi_n_204 ,csa_tree_add_107_22_pad_groupi_n_345);
  nor csa_tree_add_107_22_pad_groupi_g5192(csa_tree_add_107_22_pad_groupi_n_535 ,csa_tree_add_107_22_pad_groupi_n_28 ,csa_tree_add_107_22_pad_groupi_n_329);
  nor csa_tree_add_107_22_pad_groupi_g5193(csa_tree_add_107_22_pad_groupi_n_534 ,csa_tree_add_107_22_pad_groupi_n_194 ,csa_tree_add_107_22_pad_groupi_n_327);
  nor csa_tree_add_107_22_pad_groupi_g5194(csa_tree_add_107_22_pad_groupi_n_533 ,csa_tree_add_107_22_pad_groupi_n_191 ,csa_tree_add_107_22_pad_groupi_n_338);
  nor csa_tree_add_107_22_pad_groupi_g5195(csa_tree_add_107_22_pad_groupi_n_532 ,csa_tree_add_107_22_pad_groupi_n_184 ,csa_tree_add_107_22_pad_groupi_n_318);
  or csa_tree_add_107_22_pad_groupi_g5196(csa_tree_add_107_22_pad_groupi_n_531 ,csa_tree_add_107_22_pad_groupi_n_174 ,csa_tree_add_107_22_pad_groupi_n_305);
  nor csa_tree_add_107_22_pad_groupi_g5197(csa_tree_add_107_22_pad_groupi_n_530 ,csa_tree_add_107_22_pad_groupi_n_39 ,csa_tree_add_107_22_pad_groupi_n_330);
  nor csa_tree_add_107_22_pad_groupi_g5198(csa_tree_add_107_22_pad_groupi_n_529 ,csa_tree_add_107_22_pad_groupi_n_243 ,csa_tree_add_107_22_pad_groupi_n_344);
  nor csa_tree_add_107_22_pad_groupi_g5199(csa_tree_add_107_22_pad_groupi_n_528 ,csa_tree_add_107_22_pad_groupi_n_91 ,csa_tree_add_107_22_pad_groupi_n_345);
  nor csa_tree_add_107_22_pad_groupi_g5200(csa_tree_add_107_22_pad_groupi_n_527 ,csa_tree_add_107_22_pad_groupi_n_231 ,csa_tree_add_107_22_pad_groupi_n_321);
  nor csa_tree_add_107_22_pad_groupi_g5201(csa_tree_add_107_22_pad_groupi_n_526 ,csa_tree_add_107_22_pad_groupi_n_217 ,csa_tree_add_107_22_pad_groupi_n_265);
  nor csa_tree_add_107_22_pad_groupi_g5202(csa_tree_add_107_22_pad_groupi_n_525 ,csa_tree_add_107_22_pad_groupi_n_64 ,csa_tree_add_107_22_pad_groupi_n_311);
  nor csa_tree_add_107_22_pad_groupi_g5203(csa_tree_add_107_22_pad_groupi_n_524 ,csa_tree_add_107_22_pad_groupi_n_55 ,csa_tree_add_107_22_pad_groupi_n_269);
  nor csa_tree_add_107_22_pad_groupi_g5204(csa_tree_add_107_22_pad_groupi_n_523 ,csa_tree_add_107_22_pad_groupi_n_76 ,csa_tree_add_107_22_pad_groupi_n_312);
  nor csa_tree_add_107_22_pad_groupi_g5205(csa_tree_add_107_22_pad_groupi_n_522 ,csa_tree_add_107_22_pad_groupi_n_201 ,csa_tree_add_107_22_pad_groupi_n_339);
  nor csa_tree_add_107_22_pad_groupi_g5206(csa_tree_add_107_22_pad_groupi_n_521 ,csa_tree_add_107_22_pad_groupi_n_22 ,csa_tree_add_107_22_pad_groupi_n_275);
  nor csa_tree_add_107_22_pad_groupi_g5207(csa_tree_add_107_22_pad_groupi_n_520 ,csa_tree_add_107_22_pad_groupi_n_222 ,csa_tree_add_107_22_pad_groupi_n_262);
  nor csa_tree_add_107_22_pad_groupi_g5208(csa_tree_add_107_22_pad_groupi_n_519 ,csa_tree_add_107_22_pad_groupi_n_50 ,csa_tree_add_107_22_pad_groupi_n_272);
  or csa_tree_add_107_22_pad_groupi_g5209(csa_tree_add_107_22_pad_groupi_n_518 ,csa_tree_add_107_22_pad_groupi_n_21 ,csa_tree_add_107_22_pad_groupi_n_266);
  nor csa_tree_add_107_22_pad_groupi_g5210(csa_tree_add_107_22_pad_groupi_n_517 ,csa_tree_add_107_22_pad_groupi_n_178 ,csa_tree_add_107_22_pad_groupi_n_274);
  nor csa_tree_add_107_22_pad_groupi_g5211(csa_tree_add_107_22_pad_groupi_n_516 ,csa_tree_add_107_22_pad_groupi_n_225 ,csa_tree_add_107_22_pad_groupi_n_263);
  nor csa_tree_add_107_22_pad_groupi_g5212(csa_tree_add_107_22_pad_groupi_n_515 ,csa_tree_add_107_22_pad_groupi_n_47 ,csa_tree_add_107_22_pad_groupi_n_268);
  nor csa_tree_add_107_22_pad_groupi_g5213(csa_tree_add_107_22_pad_groupi_n_514 ,csa_tree_add_107_22_pad_groupi_n_197 ,csa_tree_add_107_22_pad_groupi_n_333);
  nor csa_tree_add_107_22_pad_groupi_g5214(csa_tree_add_107_22_pad_groupi_n_513 ,csa_tree_add_107_22_pad_groupi_n_227 ,csa_tree_add_107_22_pad_groupi_n_320);
  nor csa_tree_add_107_22_pad_groupi_g5215(csa_tree_add_107_22_pad_groupi_n_512 ,csa_tree_add_107_22_pad_groupi_n_59 ,csa_tree_add_107_22_pad_groupi_n_342);
  or csa_tree_add_107_22_pad_groupi_g5217(csa_tree_add_107_22_pad_groupi_n_583 ,csa_tree_add_107_22_pad_groupi_n_121 ,csa_tree_add_107_22_pad_groupi_n_424);
  or csa_tree_add_107_22_pad_groupi_g5218(csa_tree_add_107_22_pad_groupi_n_582 ,csa_tree_add_107_22_pad_groupi_n_162 ,csa_tree_add_107_22_pad_groupi_n_402);
  or csa_tree_add_107_22_pad_groupi_g5219(csa_tree_add_107_22_pad_groupi_n_581 ,csa_tree_add_107_22_pad_groupi_n_121 ,csa_tree_add_107_22_pad_groupi_n_109);
  or csa_tree_add_107_22_pad_groupi_g5220(csa_tree_add_107_22_pad_groupi_n_580 ,csa_tree_add_107_22_pad_groupi_n_162 ,csa_tree_add_107_22_pad_groupi_n_404);
  or csa_tree_add_107_22_pad_groupi_g5221(csa_tree_add_107_22_pad_groupi_n_579 ,csa_tree_add_107_22_pad_groupi_n_163 ,csa_tree_add_107_22_pad_groupi_n_403);
  not csa_tree_add_107_22_pad_groupi_g5223(csa_tree_add_107_22_pad_groupi_n_510 ,csa_tree_add_107_22_pad_groupi_n_505);
  not csa_tree_add_107_22_pad_groupi_g5224(csa_tree_add_107_22_pad_groupi_n_509 ,csa_tree_add_107_22_pad_groupi_n_505);
  not csa_tree_add_107_22_pad_groupi_g5225(csa_tree_add_107_22_pad_groupi_n_508 ,csa_tree_add_107_22_pad_groupi_n_506);
  not csa_tree_add_107_22_pad_groupi_g5226(csa_tree_add_107_22_pad_groupi_n_507 ,csa_tree_add_107_22_pad_groupi_n_506);
  not csa_tree_add_107_22_pad_groupi_g5227(csa_tree_add_107_22_pad_groupi_n_506 ,csa_tree_add_107_22_pad_groupi_n_505);
  not csa_tree_add_107_22_pad_groupi_g5228(csa_tree_add_107_22_pad_groupi_n_504 ,csa_tree_add_107_22_pad_groupi_n_499);
  not csa_tree_add_107_22_pad_groupi_g5229(csa_tree_add_107_22_pad_groupi_n_503 ,csa_tree_add_107_22_pad_groupi_n_499);
  not csa_tree_add_107_22_pad_groupi_g5230(csa_tree_add_107_22_pad_groupi_n_502 ,csa_tree_add_107_22_pad_groupi_n_500);
  not csa_tree_add_107_22_pad_groupi_g5231(csa_tree_add_107_22_pad_groupi_n_501 ,csa_tree_add_107_22_pad_groupi_n_500);
  not csa_tree_add_107_22_pad_groupi_g5232(csa_tree_add_107_22_pad_groupi_n_500 ,csa_tree_add_107_22_pad_groupi_n_499);
  not csa_tree_add_107_22_pad_groupi_g5233(csa_tree_add_107_22_pad_groupi_n_498 ,csa_tree_add_107_22_pad_groupi_n_278);
  not csa_tree_add_107_22_pad_groupi_g5234(csa_tree_add_107_22_pad_groupi_n_496 ,csa_tree_add_107_22_pad_groupi_n_497);
  not csa_tree_add_107_22_pad_groupi_g5235(csa_tree_add_107_22_pad_groupi_n_495 ,csa_tree_add_107_22_pad_groupi_n_493);
  not csa_tree_add_107_22_pad_groupi_g5236(csa_tree_add_107_22_pad_groupi_n_494 ,csa_tree_add_107_22_pad_groupi_n_493);
  or csa_tree_add_107_22_pad_groupi_g5237(csa_tree_add_107_22_pad_groupi_n_492 ,csa_tree_add_107_22_pad_groupi_n_27 ,csa_tree_add_107_22_pad_groupi_n_311);
  nor csa_tree_add_107_22_pad_groupi_g5238(csa_tree_add_107_22_pad_groupi_n_491 ,csa_tree_add_107_22_pad_groupi_n_180 ,csa_tree_add_107_22_pad_groupi_n_329);
  nor csa_tree_add_107_22_pad_groupi_g5239(csa_tree_add_107_22_pad_groupi_n_490 ,csa_tree_add_107_22_pad_groupi_n_220 ,csa_tree_add_107_22_pad_groupi_n_271);
  nor csa_tree_add_107_22_pad_groupi_g5240(csa_tree_add_107_22_pad_groupi_n_489 ,csa_tree_add_107_22_pad_groupi_n_82 ,csa_tree_add_107_22_pad_groupi_n_275);
  nor csa_tree_add_107_22_pad_groupi_g5241(csa_tree_add_107_22_pad_groupi_n_488 ,csa_tree_add_107_22_pad_groupi_n_181 ,csa_tree_add_107_22_pad_groupi_n_309);
  nor csa_tree_add_107_22_pad_groupi_g5242(csa_tree_add_107_22_pad_groupi_n_487 ,csa_tree_add_107_22_pad_groupi_n_88 ,csa_tree_add_107_22_pad_groupi_n_341);
  nor csa_tree_add_107_22_pad_groupi_g5243(csa_tree_add_107_22_pad_groupi_n_486 ,csa_tree_add_107_22_pad_groupi_n_227 ,csa_tree_add_107_22_pad_groupi_n_306);
  or csa_tree_add_107_22_pad_groupi_g5244(csa_tree_add_107_22_pad_groupi_n_485 ,csa_tree_add_107_22_pad_groupi_n_30 ,csa_tree_add_107_22_pad_groupi_n_302);
  nor csa_tree_add_107_22_pad_groupi_g5245(csa_tree_add_107_22_pad_groupi_n_484 ,csa_tree_add_107_22_pad_groupi_n_174 ,csa_tree_add_107_22_pad_groupi_n_315);
  or csa_tree_add_107_22_pad_groupi_g5246(csa_tree_add_107_22_pad_groupi_n_483 ,csa_tree_add_107_22_pad_groupi_n_30 ,csa_tree_add_107_22_pad_groupi_n_263);
  nor csa_tree_add_107_22_pad_groupi_g5247(csa_tree_add_107_22_pad_groupi_n_482 ,csa_tree_add_107_22_pad_groupi_n_96 ,csa_tree_add_107_22_pad_groupi_n_338);
  nor csa_tree_add_107_22_pad_groupi_g5248(csa_tree_add_107_22_pad_groupi_n_481 ,csa_tree_add_107_22_pad_groupi_n_233 ,csa_tree_add_107_22_pad_groupi_n_269);
  nor csa_tree_add_107_22_pad_groupi_g5249(csa_tree_add_107_22_pad_groupi_n_480 ,csa_tree_add_107_22_pad_groupi_n_25 ,csa_tree_add_107_22_pad_groupi_n_272);
  nor csa_tree_add_107_22_pad_groupi_g5250(csa_tree_add_107_22_pad_groupi_n_479 ,csa_tree_add_107_22_pad_groupi_n_214 ,csa_tree_add_107_22_pad_groupi_n_266);
  nor csa_tree_add_107_22_pad_groupi_g5251(csa_tree_add_107_22_pad_groupi_n_478 ,csa_tree_add_107_22_pad_groupi_n_235 ,csa_tree_add_107_22_pad_groupi_n_332);
  nor csa_tree_add_107_22_pad_groupi_g5252(csa_tree_add_107_22_pad_groupi_n_477 ,csa_tree_add_107_22_pad_groupi_n_73 ,csa_tree_add_107_22_pad_groupi_n_342);
  nor csa_tree_add_107_22_pad_groupi_g5253(csa_tree_add_107_22_pad_groupi_n_476 ,csa_tree_add_107_22_pad_groupi_n_206 ,csa_tree_add_107_22_pad_groupi_n_314);
  nor csa_tree_add_107_22_pad_groupi_g5254(csa_tree_add_107_22_pad_groupi_n_475 ,csa_tree_add_107_22_pad_groupi_n_69 ,csa_tree_add_107_22_pad_groupi_n_308);
  nor csa_tree_add_107_22_pad_groupi_g5255(csa_tree_add_107_22_pad_groupi_n_474 ,csa_tree_add_107_22_pad_groupi_n_209 ,csa_tree_add_107_22_pad_groupi_n_303);
  nor csa_tree_add_107_22_pad_groupi_g5256(csa_tree_add_107_22_pad_groupi_n_473 ,csa_tree_add_107_22_pad_groupi_n_76 ,csa_tree_add_107_22_pad_groupi_n_314);
  or csa_tree_add_107_22_pad_groupi_g5257(csa_tree_add_107_22_pad_groupi_n_472 ,csa_tree_add_107_22_pad_groupi_n_45 ,csa_tree_add_107_22_pad_groupi_n_308);
  nor csa_tree_add_107_22_pad_groupi_g5258(csa_tree_add_107_22_pad_groupi_n_471 ,csa_tree_add_107_22_pad_groupi_n_211 ,csa_tree_add_107_22_pad_groupi_n_303);
  nor csa_tree_add_107_22_pad_groupi_g5259(csa_tree_add_107_22_pad_groupi_n_470 ,csa_tree_add_107_22_pad_groupi_n_67 ,csa_tree_add_107_22_pad_groupi_n_333);
  nor csa_tree_add_107_22_pad_groupi_g5260(csa_tree_add_107_22_pad_groupi_n_469 ,csa_tree_add_107_22_pad_groupi_n_180 ,csa_tree_add_107_22_pad_groupi_n_300);
  nor csa_tree_add_107_22_pad_groupi_g5261(csa_tree_add_107_22_pad_groupi_n_468 ,csa_tree_add_107_22_pad_groupi_n_177 ,csa_tree_add_107_22_pad_groupi_n_399);
  nor csa_tree_add_107_22_pad_groupi_g5262(csa_tree_add_107_22_pad_groupi_n_467 ,csa_tree_add_107_22_pad_groupi_n_52 ,csa_tree_add_107_22_pad_groupi_n_291);
  nor csa_tree_add_107_22_pad_groupi_g5263(csa_tree_add_107_22_pad_groupi_n_466 ,csa_tree_add_107_22_pad_groupi_n_45 ,csa_tree_add_107_22_pad_groupi_n_290);
  nor csa_tree_add_107_22_pad_groupi_g5264(csa_tree_add_107_22_pad_groupi_n_465 ,csa_tree_add_107_22_pad_groupi_n_175 ,csa_tree_add_107_22_pad_groupi_n_297);
  or csa_tree_add_107_22_pad_groupi_g5265(csa_tree_add_107_22_pad_groupi_n_464 ,csa_tree_add_107_22_pad_groupi_n_36 ,csa_tree_add_107_22_pad_groupi_n_296);
  nor csa_tree_add_107_22_pad_groupi_g5266(csa_tree_add_107_22_pad_groupi_n_463 ,csa_tree_add_107_22_pad_groupi_n_90 ,csa_tree_add_107_22_pad_groupi_n_260);
  nor csa_tree_add_107_22_pad_groupi_g5267(csa_tree_add_107_22_pad_groupi_n_462 ,csa_tree_add_107_22_pad_groupi_n_212 ,csa_tree_add_107_22_pad_groupi_n_299);
  nor csa_tree_add_107_22_pad_groupi_g5268(csa_tree_add_107_22_pad_groupi_n_461 ,csa_tree_add_107_22_pad_groupi_n_95 ,csa_tree_add_107_22_pad_groupi_n_299);
  or csa_tree_add_107_22_pad_groupi_g5269(csa_tree_add_107_22_pad_groupi_n_460 ,csa_tree_add_107_22_pad_groupi_n_39 ,csa_tree_add_107_22_pad_groupi_n_290);
  nor csa_tree_add_107_22_pad_groupi_g5271(csa_tree_add_107_22_pad_groupi_n_458 ,csa_tree_add_107_22_pad_groupi_n_186 ,csa_tree_add_107_22_pad_groupi_n_300);
  or csa_tree_add_107_22_pad_groupi_g5272(csa_tree_add_107_22_pad_groupi_n_457 ,csa_tree_add_107_22_pad_groupi_n_21 ,csa_tree_add_107_22_pad_groupi_n_291);
  nor csa_tree_add_107_22_pad_groupi_g5273(csa_tree_add_107_22_pad_groupi_n_456 ,csa_tree_add_107_22_pad_groupi_n_98 ,csa_tree_add_107_22_pad_groupi_n_296);
  nor csa_tree_add_107_22_pad_groupi_g5274(csa_tree_add_107_22_pad_groupi_n_455 ,csa_tree_add_107_22_pad_groupi_n_207 ,csa_tree_add_107_22_pad_groupi_n_297);
  nor csa_tree_add_107_22_pad_groupi_g5284(csa_tree_add_107_22_pad_groupi_n_445 ,csa_tree_add_107_22_pad_groupi_n_106 ,csa_tree_add_107_22_pad_groupi_n_294);
  nor csa_tree_add_107_22_pad_groupi_g5290(csa_tree_add_107_22_pad_groupi_n_439 ,csa_tree_add_107_22_pad_groupi_n_109 ,csa_tree_add_107_22_pad_groupi_n_241);
  or csa_tree_add_107_22_pad_groupi_g5291(csa_tree_add_107_22_pad_groupi_n_438 ,csa_tree_add_107_22_pad_groupi_n_32 ,csa_tree_add_107_22_pad_groupi_n_103);
  nor csa_tree_add_107_22_pad_groupi_g5294(csa_tree_add_107_22_pad_groupi_n_435 ,csa_tree_add_107_22_pad_groupi_n_107 ,csa_tree_add_107_22_pad_groupi_n_240);
  or csa_tree_add_107_22_pad_groupi_g5295(csa_tree_add_107_22_pad_groupi_n_434 ,csa_tree_add_107_22_pad_groupi_n_293 ,csa_tree_add_107_22_pad_groupi_n_110);
  nor csa_tree_add_107_22_pad_groupi_g5296(csa_tree_add_107_22_pad_groupi_n_433 ,csa_tree_add_107_22_pad_groupi_n_103 ,csa_tree_add_107_22_pad_groupi_n_294);
  or csa_tree_add_107_22_pad_groupi_g5297(csa_tree_add_107_22_pad_groupi_n_432 ,csa_tree_add_107_22_pad_groupi_n_13 ,csa_tree_add_107_22_pad_groupi_n_61);
  nor csa_tree_add_107_22_pad_groupi_g5298(csa_tree_add_107_22_pad_groupi_n_431 ,csa_tree_add_107_22_pad_groupi_n_110 ,csa_tree_add_107_22_pad_groupi_n_238);
  or csa_tree_add_107_22_pad_groupi_g5299(csa_tree_add_107_22_pad_groupi_n_430 ,csa_tree_add_107_22_pad_groupi_n_13 ,csa_tree_add_107_22_pad_groupi_n_104);
  nor csa_tree_add_107_22_pad_groupi_g5300(csa_tree_add_107_22_pad_groupi_n_429 ,csa_tree_add_107_22_pad_groupi_n_61 ,csa_tree_add_107_22_pad_groupi_n_32);
  nor csa_tree_add_107_22_pad_groupi_g5301(csa_tree_add_107_22_pad_groupi_n_428 ,csa_tree_add_107_22_pad_groupi_n_249 ,csa_tree_add_107_22_pad_groupi_n_34);
  or csa_tree_add_107_22_pad_groupi_g5302(csa_tree_add_107_22_pad_groupi_n_427 ,csa_tree_add_107_22_pad_groupi_n_15 ,csa_tree_add_107_22_pad_groupi_n_106);
  or csa_tree_add_107_22_pad_groupi_g5303(csa_tree_add_107_22_pad_groupi_n_426 ,csa_tree_add_107_22_pad_groupi_n_34 ,csa_tree_add_107_22_pad_groupi_n_107);
  nor csa_tree_add_107_22_pad_groupi_g5304(csa_tree_add_107_22_pad_groupi_n_425 ,csa_tree_add_107_22_pad_groupi_n_104 ,csa_tree_add_107_22_pad_groupi_n_237);
  or csa_tree_add_107_22_pad_groupi_g5305(csa_tree_add_107_22_pad_groupi_n_511 ,csa_tree_add_107_22_pad_groupi_n_154 ,csa_tree_add_107_22_pad_groupi_n_424);
  or csa_tree_add_107_22_pad_groupi_g5306(csa_tree_add_107_22_pad_groupi_n_505 ,csa_tree_add_107_22_pad_groupi_n_150 ,csa_tree_add_107_22_pad_groupi_n_403);
  or csa_tree_add_107_22_pad_groupi_g5307(csa_tree_add_107_22_pad_groupi_n_499 ,csa_tree_add_107_22_pad_groupi_n_155 ,csa_tree_add_107_22_pad_groupi_n_402);
  or csa_tree_add_107_22_pad_groupi_g5309(csa_tree_add_107_22_pad_groupi_n_493 ,csa_tree_add_107_22_pad_groupi_n_152 ,csa_tree_add_107_22_pad_groupi_n_404);
  not csa_tree_add_107_22_pad_groupi_g5311(csa_tree_add_107_22_pad_groupi_n_423 ,csa_tree_add_107_22_pad_groupi_n_158);
  not csa_tree_add_107_22_pad_groupi_g5312(csa_tree_add_107_22_pad_groupi_n_422 ,csa_tree_add_107_22_pad_groupi_n_155);
  not csa_tree_add_107_22_pad_groupi_g5315(csa_tree_add_107_22_pad_groupi_n_419 ,csa_tree_add_107_22_pad_groupi_n_154);
  not csa_tree_add_107_22_pad_groupi_g5317(csa_tree_add_107_22_pad_groupi_n_418 ,csa_tree_add_107_22_pad_groupi_n_149);
  not csa_tree_add_107_22_pad_groupi_g5319(csa_tree_add_107_22_pad_groupi_n_416 ,csa_tree_add_107_22_pad_groupi_n_152);
  not csa_tree_add_107_22_pad_groupi_g5321(csa_tree_add_107_22_pad_groupi_n_415 ,csa_tree_add_107_22_pad_groupi_n_151);
  not csa_tree_add_107_22_pad_groupi_g5323(csa_tree_add_107_22_pad_groupi_n_414 ,csa_tree_add_107_22_pad_groupi_n_160);
  not csa_tree_add_107_22_pad_groupi_g5324(csa_tree_add_107_22_pad_groupi_n_413 ,csa_tree_add_107_22_pad_groupi_n_153);
  not csa_tree_add_107_22_pad_groupi_g5327(csa_tree_add_107_22_pad_groupi_n_411 ,csa_tree_add_107_22_pad_groupi_n_159);
  not csa_tree_add_107_22_pad_groupi_g5328(csa_tree_add_107_22_pad_groupi_n_410 ,csa_tree_add_107_22_pad_groupi_n_150);
  or csa_tree_add_107_22_pad_groupi_g5331(csa_tree_add_107_22_pad_groupi_n_406 ,in25[10] ,in25[9]);
  and csa_tree_add_107_22_pad_groupi_g5332(csa_tree_add_107_22_pad_groupi_n_424 ,csa_tree_add_107_22_pad_groupi_n_375 ,csa_tree_add_107_22_pad_groupi_n_388);
  and csa_tree_add_107_22_pad_groupi_g5333(csa_tree_add_107_22_pad_groupi_n_421 ,n_581 ,n_588);
  and csa_tree_add_107_22_pad_groupi_g5334(csa_tree_add_107_22_pad_groupi_n_420 ,in26[0] ,n_590);
  and csa_tree_add_107_22_pad_groupi_g5335(csa_tree_add_107_22_pad_groupi_n_417 ,n_582 ,n_589);
  and csa_tree_add_107_22_pad_groupi_g5337(csa_tree_add_107_22_pad_groupi_n_409 ,n_580 ,n_587);
  not csa_tree_add_107_22_pad_groupi_g5339(csa_tree_add_107_22_pad_groupi_n_399 ,csa_tree_add_107_22_pad_groupi_n_293);
  not csa_tree_add_107_22_pad_groupi_g5340(csa_tree_add_107_22_pad_groupi_n_398 ,csa_tree_add_107_22_pad_groupi_n_395);
  not csa_tree_add_107_22_pad_groupi_g5341(csa_tree_add_107_22_pad_groupi_n_397 ,csa_tree_add_107_22_pad_groupi_n_258);
  not csa_tree_add_107_22_pad_groupi_g5345(csa_tree_add_107_22_pad_groupi_n_396 ,csa_tree_add_107_22_pad_groupi_n_395);
  and csa_tree_add_107_22_pad_groupi_g5346(csa_tree_add_107_22_pad_groupi_n_394 ,in25[10] ,in25[9]);
  and csa_tree_add_107_22_pad_groupi_g5348(csa_tree_add_107_22_pad_groupi_n_404 ,csa_tree_add_107_22_pad_groupi_n_391 ,csa_tree_add_107_22_pad_groupi_n_393);
  and csa_tree_add_107_22_pad_groupi_g5349(csa_tree_add_107_22_pad_groupi_n_403 ,csa_tree_add_107_22_pad_groupi_n_378 ,csa_tree_add_107_22_pad_groupi_n_377);
  and csa_tree_add_107_22_pad_groupi_g5350(csa_tree_add_107_22_pad_groupi_n_402 ,csa_tree_add_107_22_pad_groupi_n_392 ,csa_tree_add_107_22_pad_groupi_n_376);
  and csa_tree_add_107_22_pad_groupi_g5351(csa_tree_add_107_22_pad_groupi_n_401 ,csa_tree_add_107_22_pad_groupi_n_390 ,csa_tree_add_107_22_pad_groupi_n_389);
  or csa_tree_add_107_22_pad_groupi_g5353(csa_tree_add_107_22_pad_groupi_n_395 ,csa_tree_add_107_22_pad_groupi_n_390 ,csa_tree_add_107_22_pad_groupi_n_389);
  not csa_tree_add_107_22_pad_groupi_g5354(csa_tree_add_107_22_pad_groupi_n_393 ,n_589);
  not csa_tree_add_107_22_pad_groupi_g5355(csa_tree_add_107_22_pad_groupi_n_392 ,n_581);
  not csa_tree_add_107_22_pad_groupi_g5356(csa_tree_add_107_22_pad_groupi_n_391 ,n_582);
  not csa_tree_add_107_22_pad_groupi_g5357(csa_tree_add_107_22_pad_groupi_n_390 ,n_584);
  not csa_tree_add_107_22_pad_groupi_g5358(csa_tree_add_107_22_pad_groupi_n_389 ,n_591);
  not csa_tree_add_107_22_pad_groupi_g5359(csa_tree_add_107_22_pad_groupi_n_388 ,n_590);
  not csa_tree_add_107_22_pad_groupi_g5360(csa_tree_add_107_22_pad_groupi_n_387 ,in25[7]);
  not csa_tree_add_107_22_pad_groupi_g5361(csa_tree_add_107_22_pad_groupi_n_386 ,in9[15]);
  not csa_tree_add_107_22_pad_groupi_g5362(csa_tree_add_107_22_pad_groupi_n_385 ,in9[2]);
  not csa_tree_add_107_22_pad_groupi_g5363(csa_tree_add_107_22_pad_groupi_n_384 ,in9[5]);
  not csa_tree_add_107_22_pad_groupi_g5364(csa_tree_add_107_22_pad_groupi_n_383 ,in9[13]);
  not csa_tree_add_107_22_pad_groupi_g5365(csa_tree_add_107_22_pad_groupi_n_382 ,in9[3]);
  not csa_tree_add_107_22_pad_groupi_g5366(csa_tree_add_107_22_pad_groupi_n_381 ,in9[9]);
  not csa_tree_add_107_22_pad_groupi_g5367(csa_tree_add_107_22_pad_groupi_n_380 ,in9[1]);
  not csa_tree_add_107_22_pad_groupi_g5368(csa_tree_add_107_22_pad_groupi_n_379 ,in9[8]);
  not csa_tree_add_107_22_pad_groupi_g5369(csa_tree_add_107_22_pad_groupi_n_378 ,n_580);
  not csa_tree_add_107_22_pad_groupi_g5370(csa_tree_add_107_22_pad_groupi_n_377 ,n_587);
  not csa_tree_add_107_22_pad_groupi_g5371(csa_tree_add_107_22_pad_groupi_n_376 ,n_588);
  not csa_tree_add_107_22_pad_groupi_g5372(csa_tree_add_107_22_pad_groupi_n_375 ,in26[0]);
  not csa_tree_add_107_22_pad_groupi_g5373(csa_tree_add_107_22_pad_groupi_n_374 ,in25[0]);
  not csa_tree_add_107_22_pad_groupi_g5374(csa_tree_add_107_22_pad_groupi_n_373 ,in25[11]);
  not csa_tree_add_107_22_pad_groupi_g5375(csa_tree_add_107_22_pad_groupi_n_372 ,in25[8]);
  not csa_tree_add_107_22_pad_groupi_g5376(csa_tree_add_107_22_pad_groupi_n_371 ,in25[1]);
  not csa_tree_add_107_22_pad_groupi_g5377(csa_tree_add_107_22_pad_groupi_n_370 ,in25[6]);
  not csa_tree_add_107_22_pad_groupi_g5378(csa_tree_add_107_22_pad_groupi_n_369 ,in25[9]);
  not csa_tree_add_107_22_pad_groupi_g5379(csa_tree_add_107_22_pad_groupi_n_368 ,in9[0]);
  not csa_tree_add_107_22_pad_groupi_g5380(csa_tree_add_107_22_pad_groupi_n_367 ,in9[4]);
  not csa_tree_add_107_22_pad_groupi_g5381(csa_tree_add_107_22_pad_groupi_n_366 ,in9[12]);
  not csa_tree_add_107_22_pad_groupi_g5382(csa_tree_add_107_22_pad_groupi_n_365 ,in9[11]);
  not csa_tree_add_107_22_pad_groupi_g5383(csa_tree_add_107_22_pad_groupi_n_364 ,in9[7]);
  not csa_tree_add_107_22_pad_groupi_g5384(csa_tree_add_107_22_pad_groupi_n_363 ,in9[10]);
  not csa_tree_add_107_22_pad_groupi_g5385(csa_tree_add_107_22_pad_groupi_n_362 ,in9[6]);
  not csa_tree_add_107_22_pad_groupi_g5386(csa_tree_add_107_22_pad_groupi_n_361 ,in9[14]);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5534(csa_tree_add_107_22_pad_groupi_n_345 ,csa_tree_add_107_22_pad_groupi_n_343);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5535(csa_tree_add_107_22_pad_groupi_n_344 ,csa_tree_add_107_22_pad_groupi_n_343);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5536(csa_tree_add_107_22_pad_groupi_n_343 ,csa_tree_add_107_22_pad_groupi_n_356);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5538(csa_tree_add_107_22_pad_groupi_n_342 ,csa_tree_add_107_22_pad_groupi_n_340);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5539(csa_tree_add_107_22_pad_groupi_n_341 ,csa_tree_add_107_22_pad_groupi_n_340);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5540(csa_tree_add_107_22_pad_groupi_n_340 ,csa_tree_add_107_22_pad_groupi_n_422);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5542(csa_tree_add_107_22_pad_groupi_n_339 ,csa_tree_add_107_22_pad_groupi_n_337);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5543(csa_tree_add_107_22_pad_groupi_n_338 ,csa_tree_add_107_22_pad_groupi_n_337);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5544(csa_tree_add_107_22_pad_groupi_n_337 ,csa_tree_add_107_22_pad_groupi_n_413);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5546(csa_tree_add_107_22_pad_groupi_n_336 ,csa_tree_add_107_22_pad_groupi_n_334);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5547(csa_tree_add_107_22_pad_groupi_n_335 ,csa_tree_add_107_22_pad_groupi_n_334);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5548(csa_tree_add_107_22_pad_groupi_n_334 ,csa_tree_add_107_22_pad_groupi_n_348);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5550(csa_tree_add_107_22_pad_groupi_n_333 ,csa_tree_add_107_22_pad_groupi_n_331);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5551(csa_tree_add_107_22_pad_groupi_n_332 ,csa_tree_add_107_22_pad_groupi_n_331);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5552(csa_tree_add_107_22_pad_groupi_n_331 ,csa_tree_add_107_22_pad_groupi_n_411);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5554(csa_tree_add_107_22_pad_groupi_n_330 ,csa_tree_add_107_22_pad_groupi_n_328);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5555(csa_tree_add_107_22_pad_groupi_n_329 ,csa_tree_add_107_22_pad_groupi_n_328);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5556(csa_tree_add_107_22_pad_groupi_n_328 ,csa_tree_add_107_22_pad_groupi_n_410);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5558(csa_tree_add_107_22_pad_groupi_n_327 ,csa_tree_add_107_22_pad_groupi_n_325);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5559(csa_tree_add_107_22_pad_groupi_n_326 ,csa_tree_add_107_22_pad_groupi_n_325);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5560(csa_tree_add_107_22_pad_groupi_n_325 ,csa_tree_add_107_22_pad_groupi_n_350);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5562(csa_tree_add_107_22_pad_groupi_n_324 ,csa_tree_add_107_22_pad_groupi_n_322);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5563(csa_tree_add_107_22_pad_groupi_n_323 ,csa_tree_add_107_22_pad_groupi_n_322);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5564(csa_tree_add_107_22_pad_groupi_n_322 ,csa_tree_add_107_22_pad_groupi_n_419);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5566(csa_tree_add_107_22_pad_groupi_n_321 ,csa_tree_add_107_22_pad_groupi_n_319);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5567(csa_tree_add_107_22_pad_groupi_n_320 ,csa_tree_add_107_22_pad_groupi_n_319);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5568(csa_tree_add_107_22_pad_groupi_n_319 ,csa_tree_add_107_22_pad_groupi_n_416);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5570(csa_tree_add_107_22_pad_groupi_n_318 ,csa_tree_add_107_22_pad_groupi_n_316);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5571(csa_tree_add_107_22_pad_groupi_n_317 ,csa_tree_add_107_22_pad_groupi_n_316);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5572(csa_tree_add_107_22_pad_groupi_n_316 ,csa_tree_add_107_22_pad_groupi_n_351);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5574(csa_tree_add_107_22_pad_groupi_n_315 ,csa_tree_add_107_22_pad_groupi_n_313);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5575(csa_tree_add_107_22_pad_groupi_n_314 ,csa_tree_add_107_22_pad_groupi_n_313);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5576(csa_tree_add_107_22_pad_groupi_n_313 ,csa_tree_add_107_22_pad_groupi_n_415);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5578(csa_tree_add_107_22_pad_groupi_n_312 ,csa_tree_add_107_22_pad_groupi_n_310);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5579(csa_tree_add_107_22_pad_groupi_n_311 ,csa_tree_add_107_22_pad_groupi_n_310);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5580(csa_tree_add_107_22_pad_groupi_n_310 ,csa_tree_add_107_22_pad_groupi_n_423);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5582(csa_tree_add_107_22_pad_groupi_n_309 ,csa_tree_add_107_22_pad_groupi_n_307);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5583(csa_tree_add_107_22_pad_groupi_n_308 ,csa_tree_add_107_22_pad_groupi_n_307);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5584(csa_tree_add_107_22_pad_groupi_n_307 ,csa_tree_add_107_22_pad_groupi_n_414);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5586(csa_tree_add_107_22_pad_groupi_n_306 ,csa_tree_add_107_22_pad_groupi_n_304);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5587(csa_tree_add_107_22_pad_groupi_n_305 ,csa_tree_add_107_22_pad_groupi_n_304);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5588(csa_tree_add_107_22_pad_groupi_n_304 ,csa_tree_add_107_22_pad_groupi_n_353);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5590(csa_tree_add_107_22_pad_groupi_n_303 ,csa_tree_add_107_22_pad_groupi_n_301);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5591(csa_tree_add_107_22_pad_groupi_n_302 ,csa_tree_add_107_22_pad_groupi_n_301);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5592(csa_tree_add_107_22_pad_groupi_n_301 ,csa_tree_add_107_22_pad_groupi_n_418);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5594(csa_tree_add_107_22_pad_groupi_n_300 ,csa_tree_add_107_22_pad_groupi_n_298);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5595(csa_tree_add_107_22_pad_groupi_n_299 ,csa_tree_add_107_22_pad_groupi_n_298);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5596(csa_tree_add_107_22_pad_groupi_n_298 ,csa_tree_add_107_22_pad_groupi_n_397);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5598(csa_tree_add_107_22_pad_groupi_n_297 ,csa_tree_add_107_22_pad_groupi_n_295);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5599(csa_tree_add_107_22_pad_groupi_n_296 ,csa_tree_add_107_22_pad_groupi_n_295);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5600(csa_tree_add_107_22_pad_groupi_n_295 ,csa_tree_add_107_22_pad_groupi_n_346);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5602(csa_tree_add_107_22_pad_groupi_n_294 ,csa_tree_add_107_22_pad_groupi_n_292);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5603(csa_tree_add_107_22_pad_groupi_n_293 ,csa_tree_add_107_22_pad_groupi_n_292);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5604(csa_tree_add_107_22_pad_groupi_n_292 ,csa_tree_add_107_22_pad_groupi_n_398);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5606(csa_tree_add_107_22_pad_groupi_n_291 ,csa_tree_add_107_22_pad_groupi_n_289);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5607(csa_tree_add_107_22_pad_groupi_n_290 ,csa_tree_add_107_22_pad_groupi_n_289);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5608(csa_tree_add_107_22_pad_groupi_n_289 ,csa_tree_add_107_22_pad_groupi_n_397);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5610(csa_tree_add_107_22_pad_groupi_n_288 ,csa_tree_add_107_22_pad_groupi_n_286);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5611(csa_tree_add_107_22_pad_groupi_n_287 ,csa_tree_add_107_22_pad_groupi_n_286);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5612(csa_tree_add_107_22_pad_groupi_n_286 ,csa_tree_add_107_22_pad_groupi_n_509);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5614(csa_tree_add_107_22_pad_groupi_n_285 ,csa_tree_add_107_22_pad_groupi_n_283);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5615(csa_tree_add_107_22_pad_groupi_n_284 ,csa_tree_add_107_22_pad_groupi_n_283);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5616(csa_tree_add_107_22_pad_groupi_n_283 ,csa_tree_add_107_22_pad_groupi_n_503);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5620(csa_tree_add_107_22_pad_groupi_n_358 ,csa_tree_add_107_22_pad_groupi_n_581);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5623(csa_tree_add_107_22_pad_groupi_n_282 ,csa_tree_add_107_22_pad_groupi_n_281);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5624(csa_tree_add_107_22_pad_groupi_n_281 ,csa_tree_add_107_22_pad_groupi_n_579);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5627(csa_tree_add_107_22_pad_groupi_n_280 ,csa_tree_add_107_22_pad_groupi_n_279);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5628(csa_tree_add_107_22_pad_groupi_n_279 ,csa_tree_add_107_22_pad_groupi_n_582);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5632(csa_tree_add_107_22_pad_groupi_n_357 ,csa_tree_add_107_22_pad_groupi_n_580);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5635(csa_tree_add_107_22_pad_groupi_n_278 ,csa_tree_add_107_22_pad_groupi_n_277);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5636(csa_tree_add_107_22_pad_groupi_n_277 ,csa_tree_add_107_22_pad_groupi_n_497);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5639(csa_tree_add_107_22_pad_groupi_n_276 ,csa_tree_add_107_22_pad_groupi_n_359);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5640(csa_tree_add_107_22_pad_groupi_n_359 ,csa_tree_add_107_22_pad_groupi_n_934);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5642(csa_tree_add_107_22_pad_groupi_n_275 ,csa_tree_add_107_22_pad_groupi_n_273);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5643(csa_tree_add_107_22_pad_groupi_n_274 ,csa_tree_add_107_22_pad_groupi_n_273);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5644(csa_tree_add_107_22_pad_groupi_n_273 ,csa_tree_add_107_22_pad_groupi_n_355);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5646(csa_tree_add_107_22_pad_groupi_n_272 ,csa_tree_add_107_22_pad_groupi_n_270);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5647(csa_tree_add_107_22_pad_groupi_n_271 ,csa_tree_add_107_22_pad_groupi_n_270);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5648(csa_tree_add_107_22_pad_groupi_n_270 ,csa_tree_add_107_22_pad_groupi_n_349);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5650(csa_tree_add_107_22_pad_groupi_n_269 ,csa_tree_add_107_22_pad_groupi_n_267);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5651(csa_tree_add_107_22_pad_groupi_n_268 ,csa_tree_add_107_22_pad_groupi_n_267);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5652(csa_tree_add_107_22_pad_groupi_n_267 ,csa_tree_add_107_22_pad_groupi_n_347);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5654(csa_tree_add_107_22_pad_groupi_n_266 ,csa_tree_add_107_22_pad_groupi_n_264);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5655(csa_tree_add_107_22_pad_groupi_n_265 ,csa_tree_add_107_22_pad_groupi_n_264);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5656(csa_tree_add_107_22_pad_groupi_n_264 ,csa_tree_add_107_22_pad_groupi_n_354);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5658(csa_tree_add_107_22_pad_groupi_n_263 ,csa_tree_add_107_22_pad_groupi_n_261);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5659(csa_tree_add_107_22_pad_groupi_n_262 ,csa_tree_add_107_22_pad_groupi_n_261);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5660(csa_tree_add_107_22_pad_groupi_n_261 ,csa_tree_add_107_22_pad_groupi_n_352);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5662(csa_tree_add_107_22_pad_groupi_n_260 ,csa_tree_add_107_22_pad_groupi_n_259);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5664(csa_tree_add_107_22_pad_groupi_n_259 ,csa_tree_add_107_22_pad_groupi_n_399);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5686(csa_tree_add_107_22_pad_groupi_n_258 ,csa_tree_add_107_22_pad_groupi_n_346);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5688(csa_tree_add_107_22_pad_groupi_n_346 ,csa_tree_add_107_22_pad_groupi_n_398);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5690(csa_tree_add_107_22_pad_groupi_n_257 ,csa_tree_add_107_22_pad_groupi_n_256);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5692(csa_tree_add_107_22_pad_groupi_n_256 ,csa_tree_add_107_22_pad_groupi_n_507);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5694(csa_tree_add_107_22_pad_groupi_n_255 ,csa_tree_add_107_22_pad_groupi_n_254);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5696(csa_tree_add_107_22_pad_groupi_n_254 ,csa_tree_add_107_22_pad_groupi_n_501);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5709(csa_tree_add_107_22_pad_groupi_n_253 ,csa_tree_add_107_22_pad_groupi_n_251);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5710(csa_tree_add_107_22_pad_groupi_n_252 ,csa_tree_add_107_22_pad_groupi_n_251);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5711(csa_tree_add_107_22_pad_groupi_n_251 ,csa_tree_add_107_22_pad_groupi_n_511);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5713(csa_tree_add_107_22_pad_groupi_n_250 ,csa_tree_add_107_22_pad_groupi_n_248);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5714(csa_tree_add_107_22_pad_groupi_n_249 ,csa_tree_add_107_22_pad_groupi_n_248);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5715(csa_tree_add_107_22_pad_groupi_n_248 ,csa_tree_add_107_22_pad_groupi_n_401);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5721(csa_tree_add_107_22_pad_groupi_n_247 ,csa_tree_add_107_22_pad_groupi_n_245);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5722(csa_tree_add_107_22_pad_groupi_n_246 ,csa_tree_add_107_22_pad_groupi_n_245);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5723(csa_tree_add_107_22_pad_groupi_n_245 ,csa_tree_add_107_22_pad_groupi_n_385);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5733(csa_tree_add_107_22_pad_groupi_n_244 ,csa_tree_add_107_22_pad_groupi_n_242);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5734(csa_tree_add_107_22_pad_groupi_n_243 ,csa_tree_add_107_22_pad_groupi_n_242);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5735(csa_tree_add_107_22_pad_groupi_n_242 ,csa_tree_add_107_22_pad_groupi_n_368);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5737(csa_tree_add_107_22_pad_groupi_n_241 ,csa_tree_add_107_22_pad_groupi_n_239);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5738(csa_tree_add_107_22_pad_groupi_n_240 ,csa_tree_add_107_22_pad_groupi_n_239);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5739(csa_tree_add_107_22_pad_groupi_n_239 ,csa_tree_add_107_22_pad_groupi_n_396);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5741(csa_tree_add_107_22_pad_groupi_n_238 ,csa_tree_add_107_22_pad_groupi_n_236);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5742(csa_tree_add_107_22_pad_groupi_n_237 ,csa_tree_add_107_22_pad_groupi_n_236);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5743(csa_tree_add_107_22_pad_groupi_n_236 ,csa_tree_add_107_22_pad_groupi_n_396);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5746(csa_tree_add_107_22_pad_groupi_n_235 ,csa_tree_add_107_22_pad_groupi_n_234);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5747(csa_tree_add_107_22_pad_groupi_n_234 ,csa_tree_add_107_22_pad_groupi_n_381);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5750(csa_tree_add_107_22_pad_groupi_n_233 ,csa_tree_add_107_22_pad_groupi_n_232);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5751(csa_tree_add_107_22_pad_groupi_n_232 ,csa_tree_add_107_22_pad_groupi_n_366);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5754(csa_tree_add_107_22_pad_groupi_n_231 ,csa_tree_add_107_22_pad_groupi_n_230);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5755(csa_tree_add_107_22_pad_groupi_n_230 ,csa_tree_add_107_22_pad_groupi_n_382);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5758(csa_tree_add_107_22_pad_groupi_n_229 ,csa_tree_add_107_22_pad_groupi_n_228);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5759(csa_tree_add_107_22_pad_groupi_n_228 ,csa_tree_add_107_22_pad_groupi_n_383);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5762(csa_tree_add_107_22_pad_groupi_n_227 ,csa_tree_add_107_22_pad_groupi_n_226);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5763(csa_tree_add_107_22_pad_groupi_n_226 ,csa_tree_add_107_22_pad_groupi_n_365);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5766(csa_tree_add_107_22_pad_groupi_n_225 ,csa_tree_add_107_22_pad_groupi_n_224);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5767(csa_tree_add_107_22_pad_groupi_n_224 ,csa_tree_add_107_22_pad_groupi_n_363);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5769(csa_tree_add_107_22_pad_groupi_n_223 ,csa_tree_add_107_22_pad_groupi_n_221);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5770(csa_tree_add_107_22_pad_groupi_n_222 ,csa_tree_add_107_22_pad_groupi_n_221);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5771(csa_tree_add_107_22_pad_groupi_n_221 ,csa_tree_add_107_22_pad_groupi_n_366);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5774(csa_tree_add_107_22_pad_groupi_n_220 ,csa_tree_add_107_22_pad_groupi_n_219);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5775(csa_tree_add_107_22_pad_groupi_n_219 ,csa_tree_add_107_22_pad_groupi_n_362);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5777(csa_tree_add_107_22_pad_groupi_n_218 ,csa_tree_add_107_22_pad_groupi_n_216);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5778(csa_tree_add_107_22_pad_groupi_n_217 ,csa_tree_add_107_22_pad_groupi_n_216);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5779(csa_tree_add_107_22_pad_groupi_n_216 ,csa_tree_add_107_22_pad_groupi_n_380);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5781(csa_tree_add_107_22_pad_groupi_n_215 ,csa_tree_add_107_22_pad_groupi_n_213);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5782(csa_tree_add_107_22_pad_groupi_n_214 ,csa_tree_add_107_22_pad_groupi_n_213);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5783(csa_tree_add_107_22_pad_groupi_n_213 ,csa_tree_add_107_22_pad_groupi_n_381);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5785(csa_tree_add_107_22_pad_groupi_n_212 ,csa_tree_add_107_22_pad_groupi_n_210);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5786(csa_tree_add_107_22_pad_groupi_n_211 ,csa_tree_add_107_22_pad_groupi_n_210);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5787(csa_tree_add_107_22_pad_groupi_n_210 ,csa_tree_add_107_22_pad_groupi_n_362);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5790(csa_tree_add_107_22_pad_groupi_n_209 ,csa_tree_add_107_22_pad_groupi_n_208);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5791(csa_tree_add_107_22_pad_groupi_n_208 ,csa_tree_add_107_22_pad_groupi_n_379);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5793(csa_tree_add_107_22_pad_groupi_n_207 ,csa_tree_add_107_22_pad_groupi_n_205);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5794(csa_tree_add_107_22_pad_groupi_n_206 ,csa_tree_add_107_22_pad_groupi_n_205);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5795(csa_tree_add_107_22_pad_groupi_n_205 ,csa_tree_add_107_22_pad_groupi_n_379);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5798(csa_tree_add_107_22_pad_groupi_n_204 ,csa_tree_add_107_22_pad_groupi_n_203);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5799(csa_tree_add_107_22_pad_groupi_n_203 ,csa_tree_add_107_22_pad_groupi_n_384);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5801(csa_tree_add_107_22_pad_groupi_n_202 ,csa_tree_add_107_22_pad_groupi_n_200);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5802(csa_tree_add_107_22_pad_groupi_n_201 ,csa_tree_add_107_22_pad_groupi_n_200);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5803(csa_tree_add_107_22_pad_groupi_n_200 ,csa_tree_add_107_22_pad_groupi_n_382);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5807(csa_tree_add_107_22_pad_groupi_n_198 ,csa_tree_add_107_22_pad_groupi_n_361);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5809(csa_tree_add_107_22_pad_groupi_n_197 ,csa_tree_add_107_22_pad_groupi_n_195);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5810(csa_tree_add_107_22_pad_groupi_n_196 ,csa_tree_add_107_22_pad_groupi_n_195);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5811(csa_tree_add_107_22_pad_groupi_n_195 ,csa_tree_add_107_22_pad_groupi_n_384);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5813(csa_tree_add_107_22_pad_groupi_n_194 ,csa_tree_add_107_22_pad_groupi_n_192);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5814(csa_tree_add_107_22_pad_groupi_n_193 ,csa_tree_add_107_22_pad_groupi_n_192);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5815(csa_tree_add_107_22_pad_groupi_n_192 ,csa_tree_add_107_22_pad_groupi_n_361);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5817(csa_tree_add_107_22_pad_groupi_n_191 ,csa_tree_add_107_22_pad_groupi_n_190);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5819(csa_tree_add_107_22_pad_groupi_n_190 ,csa_tree_add_107_22_pad_groupi_n_364);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5822(csa_tree_add_107_22_pad_groupi_n_189 ,csa_tree_add_107_22_pad_groupi_n_188);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5823(csa_tree_add_107_22_pad_groupi_n_188 ,csa_tree_add_107_22_pad_groupi_n_367);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5825(csa_tree_add_107_22_pad_groupi_n_187 ,csa_tree_add_107_22_pad_groupi_n_185);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5826(csa_tree_add_107_22_pad_groupi_n_186 ,csa_tree_add_107_22_pad_groupi_n_185);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5827(csa_tree_add_107_22_pad_groupi_n_185 ,csa_tree_add_107_22_pad_groupi_n_383);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5829(csa_tree_add_107_22_pad_groupi_n_184 ,csa_tree_add_107_22_pad_groupi_n_182);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5830(csa_tree_add_107_22_pad_groupi_n_183 ,csa_tree_add_107_22_pad_groupi_n_182);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5831(csa_tree_add_107_22_pad_groupi_n_182 ,csa_tree_add_107_22_pad_groupi_n_364);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5833(csa_tree_add_107_22_pad_groupi_n_181 ,csa_tree_add_107_22_pad_groupi_n_179);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5834(csa_tree_add_107_22_pad_groupi_n_180 ,csa_tree_add_107_22_pad_groupi_n_179);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5835(csa_tree_add_107_22_pad_groupi_n_179 ,csa_tree_add_107_22_pad_groupi_n_365);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5837(csa_tree_add_107_22_pad_groupi_n_178 ,csa_tree_add_107_22_pad_groupi_n_176);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5838(csa_tree_add_107_22_pad_groupi_n_177 ,csa_tree_add_107_22_pad_groupi_n_176);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5839(csa_tree_add_107_22_pad_groupi_n_176 ,csa_tree_add_107_22_pad_groupi_n_363);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5841(csa_tree_add_107_22_pad_groupi_n_175 ,csa_tree_add_107_22_pad_groupi_n_173);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5842(csa_tree_add_107_22_pad_groupi_n_174 ,csa_tree_add_107_22_pad_groupi_n_173);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5843(csa_tree_add_107_22_pad_groupi_n_173 ,csa_tree_add_107_22_pad_groupi_n_367);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5845(csa_tree_add_107_22_pad_groupi_n_172 ,csa_tree_add_107_22_pad_groupi_n_170);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5846(csa_tree_add_107_22_pad_groupi_n_171 ,csa_tree_add_107_22_pad_groupi_n_170);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5847(csa_tree_add_107_22_pad_groupi_n_170 ,csa_tree_add_107_22_pad_groupi_n_495);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5849(csa_tree_add_107_22_pad_groupi_n_169 ,csa_tree_add_107_22_pad_groupi_n_167);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5850(csa_tree_add_107_22_pad_groupi_n_168 ,csa_tree_add_107_22_pad_groupi_n_167);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5851(csa_tree_add_107_22_pad_groupi_n_167 ,csa_tree_add_107_22_pad_groupi_n_495);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5853(csa_tree_add_107_22_pad_groupi_n_166 ,csa_tree_add_107_22_pad_groupi_n_164);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5854(csa_tree_add_107_22_pad_groupi_n_165 ,csa_tree_add_107_22_pad_groupi_n_164);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5855(csa_tree_add_107_22_pad_groupi_n_164 ,csa_tree_add_107_22_pad_groupi_n_498);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5857(csa_tree_add_107_22_pad_groupi_n_163 ,csa_tree_add_107_22_pad_groupi_n_161);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5858(csa_tree_add_107_22_pad_groupi_n_162 ,csa_tree_add_107_22_pad_groupi_n_161);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5859(csa_tree_add_107_22_pad_groupi_n_161 ,csa_tree_add_107_22_pad_groupi_n_386);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5861(csa_tree_add_107_22_pad_groupi_n_160 ,csa_tree_add_107_22_pad_groupi_n_350);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5863(csa_tree_add_107_22_pad_groupi_n_350 ,csa_tree_add_107_22_pad_groupi_n_412);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5865(csa_tree_add_107_22_pad_groupi_n_159 ,csa_tree_add_107_22_pad_groupi_n_348);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5867(csa_tree_add_107_22_pad_groupi_n_348 ,csa_tree_add_107_22_pad_groupi_n_409);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5869(csa_tree_add_107_22_pad_groupi_n_158 ,csa_tree_add_107_22_pad_groupi_n_356);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5871(csa_tree_add_107_22_pad_groupi_n_356 ,csa_tree_add_107_22_pad_groupi_n_421);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5877(csa_tree_add_107_22_pad_groupi_n_155 ,csa_tree_add_107_22_pad_groupi_n_355);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5879(csa_tree_add_107_22_pad_groupi_n_355 ,csa_tree_add_107_22_pad_groupi_n_421);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5881(csa_tree_add_107_22_pad_groupi_n_154 ,csa_tree_add_107_22_pad_groupi_n_353);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5883(csa_tree_add_107_22_pad_groupi_n_353 ,csa_tree_add_107_22_pad_groupi_n_420);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5885(csa_tree_add_107_22_pad_groupi_n_153 ,csa_tree_add_107_22_pad_groupi_n_349);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5887(csa_tree_add_107_22_pad_groupi_n_349 ,csa_tree_add_107_22_pad_groupi_n_412);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5889(csa_tree_add_107_22_pad_groupi_n_152 ,csa_tree_add_107_22_pad_groupi_n_351);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5891(csa_tree_add_107_22_pad_groupi_n_351 ,csa_tree_add_107_22_pad_groupi_n_417);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5893(csa_tree_add_107_22_pad_groupi_n_151 ,csa_tree_add_107_22_pad_groupi_n_352);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5895(csa_tree_add_107_22_pad_groupi_n_352 ,csa_tree_add_107_22_pad_groupi_n_417);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5897(csa_tree_add_107_22_pad_groupi_n_150 ,csa_tree_add_107_22_pad_groupi_n_347);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5899(csa_tree_add_107_22_pad_groupi_n_347 ,csa_tree_add_107_22_pad_groupi_n_409);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5901(csa_tree_add_107_22_pad_groupi_n_149 ,csa_tree_add_107_22_pad_groupi_n_354);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5903(csa_tree_add_107_22_pad_groupi_n_354 ,csa_tree_add_107_22_pad_groupi_n_420);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5905(csa_tree_add_107_22_pad_groupi_n_148 ,csa_tree_add_107_22_pad_groupi_n_146);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5906(csa_tree_add_107_22_pad_groupi_n_147 ,csa_tree_add_107_22_pad_groupi_n_146);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5907(csa_tree_add_107_22_pad_groupi_n_146 ,csa_tree_add_107_22_pad_groupi_n_504);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5909(csa_tree_add_107_22_pad_groupi_n_145 ,csa_tree_add_107_22_pad_groupi_n_143);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5910(csa_tree_add_107_22_pad_groupi_n_144 ,csa_tree_add_107_22_pad_groupi_n_143);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5911(csa_tree_add_107_22_pad_groupi_n_143 ,csa_tree_add_107_22_pad_groupi_n_510);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5913(csa_tree_add_107_22_pad_groupi_n_142 ,csa_tree_add_107_22_pad_groupi_n_140);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5914(csa_tree_add_107_22_pad_groupi_n_141 ,csa_tree_add_107_22_pad_groupi_n_140);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5915(csa_tree_add_107_22_pad_groupi_n_140 ,csa_tree_add_107_22_pad_groupi_n_510);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5917(csa_tree_add_107_22_pad_groupi_n_139 ,csa_tree_add_107_22_pad_groupi_n_137);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5918(csa_tree_add_107_22_pad_groupi_n_138 ,csa_tree_add_107_22_pad_groupi_n_137);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5919(csa_tree_add_107_22_pad_groupi_n_137 ,csa_tree_add_107_22_pad_groupi_n_494);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5921(csa_tree_add_107_22_pad_groupi_n_136 ,csa_tree_add_107_22_pad_groupi_n_134);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5922(csa_tree_add_107_22_pad_groupi_n_135 ,csa_tree_add_107_22_pad_groupi_n_134);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5923(csa_tree_add_107_22_pad_groupi_n_134 ,csa_tree_add_107_22_pad_groupi_n_494);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5925(csa_tree_add_107_22_pad_groupi_n_133 ,csa_tree_add_107_22_pad_groupi_n_131);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5926(csa_tree_add_107_22_pad_groupi_n_132 ,csa_tree_add_107_22_pad_groupi_n_131);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5927(csa_tree_add_107_22_pad_groupi_n_131 ,csa_tree_add_107_22_pad_groupi_n_504);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5929(csa_tree_add_107_22_pad_groupi_n_130 ,csa_tree_add_107_22_pad_groupi_n_128);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5930(csa_tree_add_107_22_pad_groupi_n_129 ,csa_tree_add_107_22_pad_groupi_n_128);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5931(csa_tree_add_107_22_pad_groupi_n_128 ,csa_tree_add_107_22_pad_groupi_n_498);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5933(csa_tree_add_107_22_pad_groupi_n_127 ,csa_tree_add_107_22_pad_groupi_n_125);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5934(csa_tree_add_107_22_pad_groupi_n_126 ,csa_tree_add_107_22_pad_groupi_n_125);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5935(csa_tree_add_107_22_pad_groupi_n_125 ,csa_tree_add_107_22_pad_groupi_n_496);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5937(csa_tree_add_107_22_pad_groupi_n_124 ,csa_tree_add_107_22_pad_groupi_n_122);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5938(csa_tree_add_107_22_pad_groupi_n_123 ,csa_tree_add_107_22_pad_groupi_n_122);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5939(csa_tree_add_107_22_pad_groupi_n_122 ,csa_tree_add_107_22_pad_groupi_n_496);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5941(csa_tree_add_107_22_pad_groupi_n_121 ,csa_tree_add_107_22_pad_groupi_n_120);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5943(csa_tree_add_107_22_pad_groupi_n_120 ,csa_tree_add_107_22_pad_groupi_n_386);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5945(csa_tree_add_107_22_pad_groupi_n_119 ,csa_tree_add_107_22_pad_groupi_n_117);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5946(csa_tree_add_107_22_pad_groupi_n_118 ,csa_tree_add_107_22_pad_groupi_n_117);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5947(csa_tree_add_107_22_pad_groupi_n_117 ,csa_tree_add_107_22_pad_groupi_n_511);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5949(csa_tree_add_107_22_pad_groupi_n_116 ,csa_tree_add_107_22_pad_groupi_n_114);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5950(csa_tree_add_107_22_pad_groupi_n_115 ,csa_tree_add_107_22_pad_groupi_n_114);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5951(csa_tree_add_107_22_pad_groupi_n_114 ,csa_tree_add_107_22_pad_groupi_n_511);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5953(csa_tree_add_107_22_pad_groupi_n_113 ,csa_tree_add_107_22_pad_groupi_n_111);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5954(csa_tree_add_107_22_pad_groupi_n_112 ,csa_tree_add_107_22_pad_groupi_n_111);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5955(csa_tree_add_107_22_pad_groupi_n_111 ,csa_tree_add_107_22_pad_groupi_n_253);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5957(csa_tree_add_107_22_pad_groupi_n_110 ,csa_tree_add_107_22_pad_groupi_n_108);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5958(csa_tree_add_107_22_pad_groupi_n_109 ,csa_tree_add_107_22_pad_groupi_n_108);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5959(csa_tree_add_107_22_pad_groupi_n_108 ,csa_tree_add_107_22_pad_groupi_n_401);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5961(csa_tree_add_107_22_pad_groupi_n_107 ,csa_tree_add_107_22_pad_groupi_n_105);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5962(csa_tree_add_107_22_pad_groupi_n_106 ,csa_tree_add_107_22_pad_groupi_n_105);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5963(csa_tree_add_107_22_pad_groupi_n_105 ,csa_tree_add_107_22_pad_groupi_n_401);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5965(csa_tree_add_107_22_pad_groupi_n_104 ,csa_tree_add_107_22_pad_groupi_n_102);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5966(csa_tree_add_107_22_pad_groupi_n_103 ,csa_tree_add_107_22_pad_groupi_n_102);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5967(csa_tree_add_107_22_pad_groupi_n_102 ,csa_tree_add_107_22_pad_groupi_n_250);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5969(csa_tree_add_107_22_pad_groupi_n_101 ,csa_tree_add_107_22_pad_groupi_n_99);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5970(csa_tree_add_107_22_pad_groupi_n_100 ,csa_tree_add_107_22_pad_groupi_n_99);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5971(csa_tree_add_107_22_pad_groupi_n_99 ,csa_tree_add_107_22_pad_groupi_n_385);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5973(csa_tree_add_107_22_pad_groupi_n_98 ,csa_tree_add_107_22_pad_groupi_n_97);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5975(csa_tree_add_107_22_pad_groupi_n_97 ,csa_tree_add_107_22_pad_groupi_n_247);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5977(csa_tree_add_107_22_pad_groupi_n_96 ,csa_tree_add_107_22_pad_groupi_n_94);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5978(csa_tree_add_107_22_pad_groupi_n_95 ,csa_tree_add_107_22_pad_groupi_n_94);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5979(csa_tree_add_107_22_pad_groupi_n_94 ,csa_tree_add_107_22_pad_groupi_n_381);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5981(csa_tree_add_107_22_pad_groupi_n_93 ,csa_tree_add_107_22_pad_groupi_n_92);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5983(csa_tree_add_107_22_pad_groupi_n_92 ,csa_tree_add_107_22_pad_groupi_n_252);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5985(csa_tree_add_107_22_pad_groupi_n_91 ,csa_tree_add_107_22_pad_groupi_n_89);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5986(csa_tree_add_107_22_pad_groupi_n_90 ,csa_tree_add_107_22_pad_groupi_n_89);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5987(csa_tree_add_107_22_pad_groupi_n_89 ,csa_tree_add_107_22_pad_groupi_n_366);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5989(csa_tree_add_107_22_pad_groupi_n_88 ,csa_tree_add_107_22_pad_groupi_n_86);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5990(csa_tree_add_107_22_pad_groupi_n_87 ,csa_tree_add_107_22_pad_groupi_n_86);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5991(csa_tree_add_107_22_pad_groupi_n_86 ,csa_tree_add_107_22_pad_groupi_n_382);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5993(csa_tree_add_107_22_pad_groupi_n_85 ,csa_tree_add_107_22_pad_groupi_n_83);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5994(csa_tree_add_107_22_pad_groupi_n_84 ,csa_tree_add_107_22_pad_groupi_n_83);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5995(csa_tree_add_107_22_pad_groupi_n_83 ,csa_tree_add_107_22_pad_groupi_n_383);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5997(csa_tree_add_107_22_pad_groupi_n_82 ,csa_tree_add_107_22_pad_groupi_n_80);
  not csa_tree_add_107_22_pad_groupi_drc_bufs5999(csa_tree_add_107_22_pad_groupi_n_80 ,csa_tree_add_107_22_pad_groupi_n_365);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6001(csa_tree_add_107_22_pad_groupi_n_79 ,csa_tree_add_107_22_pad_groupi_n_77);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6002(csa_tree_add_107_22_pad_groupi_n_78 ,csa_tree_add_107_22_pad_groupi_n_77);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6003(csa_tree_add_107_22_pad_groupi_n_77 ,csa_tree_add_107_22_pad_groupi_n_363);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6005(csa_tree_add_107_22_pad_groupi_n_76 ,csa_tree_add_107_22_pad_groupi_n_75);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6007(csa_tree_add_107_22_pad_groupi_n_75 ,csa_tree_add_107_22_pad_groupi_n_215);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6009(csa_tree_add_107_22_pad_groupi_n_74 ,csa_tree_add_107_22_pad_groupi_n_72);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6010(csa_tree_add_107_22_pad_groupi_n_73 ,csa_tree_add_107_22_pad_groupi_n_72);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6011(csa_tree_add_107_22_pad_groupi_n_72 ,csa_tree_add_107_22_pad_groupi_n_385);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6013(csa_tree_add_107_22_pad_groupi_n_71 ,csa_tree_add_107_22_pad_groupi_n_70);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6015(csa_tree_add_107_22_pad_groupi_n_70 ,csa_tree_add_107_22_pad_groupi_n_218);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6017(csa_tree_add_107_22_pad_groupi_n_69 ,csa_tree_add_107_22_pad_groupi_n_68);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6019(csa_tree_add_107_22_pad_groupi_n_68 ,csa_tree_add_107_22_pad_groupi_n_223);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6021(csa_tree_add_107_22_pad_groupi_n_67 ,csa_tree_add_107_22_pad_groupi_n_65);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6022(csa_tree_add_107_22_pad_groupi_n_66 ,csa_tree_add_107_22_pad_groupi_n_65);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6023(csa_tree_add_107_22_pad_groupi_n_65 ,csa_tree_add_107_22_pad_groupi_n_362);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6025(csa_tree_add_107_22_pad_groupi_n_64 ,csa_tree_add_107_22_pad_groupi_n_62);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6027(csa_tree_add_107_22_pad_groupi_n_62 ,csa_tree_add_107_22_pad_groupi_n_380);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6029(csa_tree_add_107_22_pad_groupi_n_61 ,csa_tree_add_107_22_pad_groupi_n_60);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6031(csa_tree_add_107_22_pad_groupi_n_60 ,csa_tree_add_107_22_pad_groupi_n_249);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6033(csa_tree_add_107_22_pad_groupi_n_59 ,csa_tree_add_107_22_pad_groupi_n_58);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6035(csa_tree_add_107_22_pad_groupi_n_58 ,csa_tree_add_107_22_pad_groupi_n_212);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6037(csa_tree_add_107_22_pad_groupi_n_57 ,csa_tree_add_107_22_pad_groupi_n_56);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6039(csa_tree_add_107_22_pad_groupi_n_56 ,csa_tree_add_107_22_pad_groupi_n_244);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6041(csa_tree_add_107_22_pad_groupi_n_55 ,csa_tree_add_107_22_pad_groupi_n_54);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6043(csa_tree_add_107_22_pad_groupi_n_54 ,csa_tree_add_107_22_pad_groupi_n_207);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6045(csa_tree_add_107_22_pad_groupi_n_53 ,csa_tree_add_107_22_pad_groupi_n_51);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6046(csa_tree_add_107_22_pad_groupi_n_52 ,csa_tree_add_107_22_pad_groupi_n_51);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6047(csa_tree_add_107_22_pad_groupi_n_51 ,csa_tree_add_107_22_pad_groupi_n_384);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6049(csa_tree_add_107_22_pad_groupi_n_50 ,csa_tree_add_107_22_pad_groupi_n_48);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6051(csa_tree_add_107_22_pad_groupi_n_48 ,csa_tree_add_107_22_pad_groupi_n_379);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6053(csa_tree_add_107_22_pad_groupi_n_47 ,csa_tree_add_107_22_pad_groupi_n_46);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6055(csa_tree_add_107_22_pad_groupi_n_46 ,csa_tree_add_107_22_pad_groupi_n_246);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6057(csa_tree_add_107_22_pad_groupi_n_45 ,csa_tree_add_107_22_pad_groupi_n_43);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6059(csa_tree_add_107_22_pad_groupi_n_43 ,csa_tree_add_107_22_pad_groupi_n_380);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6061(csa_tree_add_107_22_pad_groupi_n_42 ,csa_tree_add_107_22_pad_groupi_n_40);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6062(csa_tree_add_107_22_pad_groupi_n_41 ,csa_tree_add_107_22_pad_groupi_n_40);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6063(csa_tree_add_107_22_pad_groupi_n_40 ,csa_tree_add_107_22_pad_groupi_n_368);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6065(csa_tree_add_107_22_pad_groupi_n_39 ,csa_tree_add_107_22_pad_groupi_n_37);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6066(csa_tree_add_107_22_pad_groupi_n_38 ,csa_tree_add_107_22_pad_groupi_n_37);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6067(csa_tree_add_107_22_pad_groupi_n_37 ,csa_tree_add_107_22_pad_groupi_n_361);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6069(csa_tree_add_107_22_pad_groupi_n_36 ,csa_tree_add_107_22_pad_groupi_n_35);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6071(csa_tree_add_107_22_pad_groupi_n_35 ,csa_tree_add_107_22_pad_groupi_n_202);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6073(csa_tree_add_107_22_pad_groupi_n_34 ,csa_tree_add_107_22_pad_groupi_n_33);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6075(csa_tree_add_107_22_pad_groupi_n_33 ,csa_tree_add_107_22_pad_groupi_n_238);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6077(csa_tree_add_107_22_pad_groupi_n_32 ,csa_tree_add_107_22_pad_groupi_n_31);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6079(csa_tree_add_107_22_pad_groupi_n_31 ,csa_tree_add_107_22_pad_groupi_n_241);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6082(csa_tree_add_107_22_pad_groupi_n_30 ,csa_tree_add_107_22_pad_groupi_n_29);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6083(csa_tree_add_107_22_pad_groupi_n_29 ,csa_tree_add_107_22_pad_groupi_n_193);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6085(csa_tree_add_107_22_pad_groupi_n_28 ,csa_tree_add_107_22_pad_groupi_n_26);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6086(csa_tree_add_107_22_pad_groupi_n_27 ,csa_tree_add_107_22_pad_groupi_n_26);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6087(csa_tree_add_107_22_pad_groupi_n_26 ,csa_tree_add_107_22_pad_groupi_n_367);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6089(csa_tree_add_107_22_pad_groupi_n_25 ,csa_tree_add_107_22_pad_groupi_n_23);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6090(csa_tree_add_107_22_pad_groupi_n_24 ,csa_tree_add_107_22_pad_groupi_n_23);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6091(csa_tree_add_107_22_pad_groupi_n_23 ,csa_tree_add_107_22_pad_groupi_n_368);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6093(csa_tree_add_107_22_pad_groupi_n_22 ,csa_tree_add_107_22_pad_groupi_n_20);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6094(csa_tree_add_107_22_pad_groupi_n_21 ,csa_tree_add_107_22_pad_groupi_n_20);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6095(csa_tree_add_107_22_pad_groupi_n_20 ,csa_tree_add_107_22_pad_groupi_n_364);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6098(csa_tree_add_107_22_pad_groupi_n_19 ,csa_tree_add_107_22_pad_groupi_n_18);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6099(csa_tree_add_107_22_pad_groupi_n_18 ,csa_tree_add_107_22_pad_groupi_n_243);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6102(csa_tree_add_107_22_pad_groupi_n_17 ,csa_tree_add_107_22_pad_groupi_n_16);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6103(csa_tree_add_107_22_pad_groupi_n_16 ,csa_tree_add_107_22_pad_groupi_n_196);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6106(csa_tree_add_107_22_pad_groupi_n_15 ,csa_tree_add_107_22_pad_groupi_n_14);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6107(csa_tree_add_107_22_pad_groupi_n_14 ,csa_tree_add_107_22_pad_groupi_n_237);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6110(csa_tree_add_107_22_pad_groupi_n_13 ,csa_tree_add_107_22_pad_groupi_n_12);
  not csa_tree_add_107_22_pad_groupi_drc_bufs6111(csa_tree_add_107_22_pad_groupi_n_12 ,csa_tree_add_107_22_pad_groupi_n_240);
  xor csa_tree_add_107_22_pad_groupi_g2(n_263 ,csa_tree_add_107_22_pad_groupi_n_1537 ,csa_tree_add_107_22_pad_groupi_n_1520);
  xor csa_tree_add_107_22_pad_groupi_g6113(n_261 ,csa_tree_add_107_22_pad_groupi_n_1532 ,csa_tree_add_107_22_pad_groupi_n_1518);
  xor csa_tree_add_107_22_pad_groupi_g6114(n_258 ,csa_tree_add_107_22_pad_groupi_n_1524 ,csa_tree_add_107_22_pad_groupi_n_1482);
  xor csa_tree_add_107_22_pad_groupi_g6115(n_257 ,csa_tree_add_107_22_pad_groupi_n_1522 ,csa_tree_add_107_22_pad_groupi_n_1502);
  xor csa_tree_add_107_22_pad_groupi_g6116(n_256 ,csa_tree_add_107_22_pad_groupi_n_1515 ,csa_tree_add_107_22_pad_groupi_n_1461);
  xor csa_tree_add_107_22_pad_groupi_g6117(csa_tree_add_107_22_pad_groupi_n_6 ,csa_tree_add_107_22_pad_groupi_n_1368 ,csa_tree_add_107_22_pad_groupi_n_1406);
  xor csa_tree_add_107_22_pad_groupi_g6118(csa_tree_add_107_22_pad_groupi_n_5 ,csa_tree_add_107_22_pad_groupi_n_1332 ,csa_tree_add_107_22_pad_groupi_n_1350);
  xor csa_tree_add_107_22_pad_groupi_g6119(csa_tree_add_107_22_pad_groupi_n_4 ,csa_tree_add_107_22_pad_groupi_n_836 ,csa_tree_add_107_22_pad_groupi_n_0);
  xor csa_tree_add_107_22_pad_groupi_g6120(csa_tree_add_107_22_pad_groupi_n_3 ,csa_tree_add_107_22_pad_groupi_n_835 ,csa_tree_add_107_22_pad_groupi_n_948);
  xor csa_tree_add_107_22_pad_groupi_g6122(csa_tree_add_107_22_pad_groupi_n_1 ,csa_tree_add_107_22_pad_groupi_n_358 ,in25[9]);
  xor csa_tree_add_107_22_pad_groupi_g6123(csa_tree_add_107_22_pad_groupi_n_0 ,csa_tree_add_107_22_pad_groupi_n_357 ,in25[11]);
  xnor csa_tree_add_110_49_pad_groupi_g4238(n_142 ,csa_tree_add_110_49_pad_groupi_n_1555 ,csa_tree_add_110_49_pad_groupi_n_1482);
  nor csa_tree_add_110_49_pad_groupi_g4239(csa_tree_add_110_49_pad_groupi_n_1555 ,csa_tree_add_110_49_pad_groupi_n_1553 ,csa_tree_add_110_49_pad_groupi_n_1504);
  xnor csa_tree_add_110_49_pad_groupi_g4240(n_141 ,csa_tree_add_110_49_pad_groupi_n_1552 ,csa_tree_add_110_49_pad_groupi_n_1511);
  nor csa_tree_add_110_49_pad_groupi_g4241(csa_tree_add_110_49_pad_groupi_n_1553 ,csa_tree_add_110_49_pad_groupi_n_1552 ,csa_tree_add_110_49_pad_groupi_n_1505);
  and csa_tree_add_110_49_pad_groupi_g4242(csa_tree_add_110_49_pad_groupi_n_1552 ,csa_tree_add_110_49_pad_groupi_n_1485 ,csa_tree_add_110_49_pad_groupi_n_1551);
  or csa_tree_add_110_49_pad_groupi_g4244(csa_tree_add_110_49_pad_groupi_n_1551 ,csa_tree_add_110_49_pad_groupi_n_1550 ,csa_tree_add_110_49_pad_groupi_n_1491);
  and csa_tree_add_110_49_pad_groupi_g4246(csa_tree_add_110_49_pad_groupi_n_1550 ,csa_tree_add_110_49_pad_groupi_n_1549 ,csa_tree_add_110_49_pad_groupi_n_1513);
  or csa_tree_add_110_49_pad_groupi_g4248(csa_tree_add_110_49_pad_groupi_n_1549 ,csa_tree_add_110_49_pad_groupi_n_1512 ,csa_tree_add_110_49_pad_groupi_n_1548);
  and csa_tree_add_110_49_pad_groupi_g4250(csa_tree_add_110_49_pad_groupi_n_1548 ,csa_tree_add_110_49_pad_groupi_n_1546 ,csa_tree_add_110_49_pad_groupi_n_1506);
  xnor csa_tree_add_110_49_pad_groupi_g4251(n_138 ,csa_tree_add_110_49_pad_groupi_n_1545 ,csa_tree_add_110_49_pad_groupi_n_1510);
  or csa_tree_add_110_49_pad_groupi_g4252(csa_tree_add_110_49_pad_groupi_n_1546 ,csa_tree_add_110_49_pad_groupi_n_1545 ,csa_tree_add_110_49_pad_groupi_n_1507);
  and csa_tree_add_110_49_pad_groupi_g4253(csa_tree_add_110_49_pad_groupi_n_1545 ,csa_tree_add_110_49_pad_groupi_n_1543 ,csa_tree_add_110_49_pad_groupi_n_1515);
  xnor csa_tree_add_110_49_pad_groupi_g4254(n_137 ,csa_tree_add_110_49_pad_groupi_n_1542 ,csa_tree_add_110_49_pad_groupi_n_1517);
  or csa_tree_add_110_49_pad_groupi_g4255(csa_tree_add_110_49_pad_groupi_n_1543 ,csa_tree_add_110_49_pad_groupi_n_1542 ,csa_tree_add_110_49_pad_groupi_n_1516);
  and csa_tree_add_110_49_pad_groupi_g4256(csa_tree_add_110_49_pad_groupi_n_1542 ,csa_tree_add_110_49_pad_groupi_n_1540 ,csa_tree_add_110_49_pad_groupi_n_1492);
  xnor csa_tree_add_110_49_pad_groupi_g4257(n_136 ,csa_tree_add_110_49_pad_groupi_n_1539 ,csa_tree_add_110_49_pad_groupi_n_1500);
  or csa_tree_add_110_49_pad_groupi_g4258(csa_tree_add_110_49_pad_groupi_n_1540 ,csa_tree_add_110_49_pad_groupi_n_1493 ,csa_tree_add_110_49_pad_groupi_n_1539);
  and csa_tree_add_110_49_pad_groupi_g4259(csa_tree_add_110_49_pad_groupi_n_1539 ,csa_tree_add_110_49_pad_groupi_n_1494 ,csa_tree_add_110_49_pad_groupi_n_1537);
  xnor csa_tree_add_110_49_pad_groupi_g4260(n_135 ,csa_tree_add_110_49_pad_groupi_n_1536 ,csa_tree_add_110_49_pad_groupi_n_1499);
  or csa_tree_add_110_49_pad_groupi_g4261(csa_tree_add_110_49_pad_groupi_n_1537 ,csa_tree_add_110_49_pad_groupi_n_1536 ,csa_tree_add_110_49_pad_groupi_n_1495);
  and csa_tree_add_110_49_pad_groupi_g4262(csa_tree_add_110_49_pad_groupi_n_1536 ,csa_tree_add_110_49_pad_groupi_n_1534 ,csa_tree_add_110_49_pad_groupi_n_1472);
  xnor csa_tree_add_110_49_pad_groupi_g4263(n_134 ,csa_tree_add_110_49_pad_groupi_n_1533 ,csa_tree_add_110_49_pad_groupi_n_1483);
  or csa_tree_add_110_49_pad_groupi_g4264(csa_tree_add_110_49_pad_groupi_n_1534 ,csa_tree_add_110_49_pad_groupi_n_1533 ,csa_tree_add_110_49_pad_groupi_n_1473);
  and csa_tree_add_110_49_pad_groupi_g4265(csa_tree_add_110_49_pad_groupi_n_1533 ,csa_tree_add_110_49_pad_groupi_n_1474 ,csa_tree_add_110_49_pad_groupi_n_1531);
  xnor csa_tree_add_110_49_pad_groupi_g4266(n_133 ,csa_tree_add_110_49_pad_groupi_n_1530 ,csa_tree_add_110_49_pad_groupi_n_1484);
  or csa_tree_add_110_49_pad_groupi_g4267(csa_tree_add_110_49_pad_groupi_n_1531 ,csa_tree_add_110_49_pad_groupi_n_1530 ,csa_tree_add_110_49_pad_groupi_n_1471);
  and csa_tree_add_110_49_pad_groupi_g4268(csa_tree_add_110_49_pad_groupi_n_1530 ,csa_tree_add_110_49_pad_groupi_n_1528 ,csa_tree_add_110_49_pad_groupi_n_1454);
  xnor csa_tree_add_110_49_pad_groupi_g4269(n_132 ,csa_tree_add_110_49_pad_groupi_n_1527 ,csa_tree_add_110_49_pad_groupi_n_1464);
  or csa_tree_add_110_49_pad_groupi_g4270(csa_tree_add_110_49_pad_groupi_n_1528 ,csa_tree_add_110_49_pad_groupi_n_1452 ,csa_tree_add_110_49_pad_groupi_n_1527);
  and csa_tree_add_110_49_pad_groupi_g4271(csa_tree_add_110_49_pad_groupi_n_1527 ,csa_tree_add_110_49_pad_groupi_n_1525 ,csa_tree_add_110_49_pad_groupi_n_1453);
  xnor csa_tree_add_110_49_pad_groupi_g4272(n_131 ,csa_tree_add_110_49_pad_groupi_n_1524 ,csa_tree_add_110_49_pad_groupi_n_1463);
  or csa_tree_add_110_49_pad_groupi_g4273(csa_tree_add_110_49_pad_groupi_n_1525 ,csa_tree_add_110_49_pad_groupi_n_1449 ,csa_tree_add_110_49_pad_groupi_n_1524);
  and csa_tree_add_110_49_pad_groupi_g4274(csa_tree_add_110_49_pad_groupi_n_1524 ,csa_tree_add_110_49_pad_groupi_n_1522 ,csa_tree_add_110_49_pad_groupi_n_1450);
  xnor csa_tree_add_110_49_pad_groupi_g4275(n_130 ,csa_tree_add_110_49_pad_groupi_n_1521 ,csa_tree_add_110_49_pad_groupi_n_1461);
  or csa_tree_add_110_49_pad_groupi_g4276(csa_tree_add_110_49_pad_groupi_n_1522 ,csa_tree_add_110_49_pad_groupi_n_1451 ,csa_tree_add_110_49_pad_groupi_n_1521);
  and csa_tree_add_110_49_pad_groupi_g4277(csa_tree_add_110_49_pad_groupi_n_1521 ,csa_tree_add_110_49_pad_groupi_n_1419 ,csa_tree_add_110_49_pad_groupi_n_1519);
  xnor csa_tree_add_110_49_pad_groupi_g4278(n_129 ,csa_tree_add_110_49_pad_groupi_n_1514 ,csa_tree_add_110_49_pad_groupi_n_1437);
  or csa_tree_add_110_49_pad_groupi_g4279(csa_tree_add_110_49_pad_groupi_n_1519 ,csa_tree_add_110_49_pad_groupi_n_1421 ,csa_tree_add_110_49_pad_groupi_n_1514);
  xnor csa_tree_add_110_49_pad_groupi_g4280(csa_tree_add_110_49_pad_groupi_n_1518 ,csa_tree_add_110_49_pad_groupi_n_1481 ,csa_tree_add_110_49_pad_groupi_n_1498);
  xnor csa_tree_add_110_49_pad_groupi_g4281(csa_tree_add_110_49_pad_groupi_n_1517 ,csa_tree_add_110_49_pad_groupi_n_1457 ,csa_tree_add_110_49_pad_groupi_n_1503);
  nor csa_tree_add_110_49_pad_groupi_g4282(csa_tree_add_110_49_pad_groupi_n_1516 ,csa_tree_add_110_49_pad_groupi_n_1457 ,csa_tree_add_110_49_pad_groupi_n_1502);
  or csa_tree_add_110_49_pad_groupi_g4283(csa_tree_add_110_49_pad_groupi_n_1515 ,csa_tree_add_110_49_pad_groupi_n_1456 ,csa_tree_add_110_49_pad_groupi_n_1503);
  and csa_tree_add_110_49_pad_groupi_g4284(csa_tree_add_110_49_pad_groupi_n_1514 ,csa_tree_add_110_49_pad_groupi_n_1422 ,csa_tree_add_110_49_pad_groupi_n_1508);
  or csa_tree_add_110_49_pad_groupi_g4285(csa_tree_add_110_49_pad_groupi_n_1513 ,csa_tree_add_110_49_pad_groupi_n_1480 ,csa_tree_add_110_49_pad_groupi_n_1497);
  nor csa_tree_add_110_49_pad_groupi_g4286(csa_tree_add_110_49_pad_groupi_n_1512 ,csa_tree_add_110_49_pad_groupi_n_1481 ,csa_tree_add_110_49_pad_groupi_n_1498);
  xnor csa_tree_add_110_49_pad_groupi_g4287(csa_tree_add_110_49_pad_groupi_n_1511 ,csa_tree_add_110_49_pad_groupi_n_1448 ,csa_tree_add_110_49_pad_groupi_n_1489);
  xnor csa_tree_add_110_49_pad_groupi_g4288(csa_tree_add_110_49_pad_groupi_n_1510 ,csa_tree_add_110_49_pad_groupi_n_1477 ,csa_tree_add_110_49_pad_groupi_n_1488);
  xnor csa_tree_add_110_49_pad_groupi_g4289(n_128 ,csa_tree_add_110_49_pad_groupi_n_1496 ,csa_tree_add_110_49_pad_groupi_n_1436);
  or csa_tree_add_110_49_pad_groupi_g4290(csa_tree_add_110_49_pad_groupi_n_1508 ,csa_tree_add_110_49_pad_groupi_n_1423 ,csa_tree_add_110_49_pad_groupi_n_1496);
  nor csa_tree_add_110_49_pad_groupi_g4291(csa_tree_add_110_49_pad_groupi_n_1507 ,csa_tree_add_110_49_pad_groupi_n_1476 ,csa_tree_add_110_49_pad_groupi_n_1488);
  or csa_tree_add_110_49_pad_groupi_g4292(csa_tree_add_110_49_pad_groupi_n_1506 ,csa_tree_add_110_49_pad_groupi_n_1477 ,csa_tree_add_110_49_pad_groupi_n_1487);
  and csa_tree_add_110_49_pad_groupi_g4293(csa_tree_add_110_49_pad_groupi_n_1505 ,csa_tree_add_110_49_pad_groupi_n_1448 ,csa_tree_add_110_49_pad_groupi_n_1490);
  nor csa_tree_add_110_49_pad_groupi_g4294(csa_tree_add_110_49_pad_groupi_n_1504 ,csa_tree_add_110_49_pad_groupi_n_1448 ,csa_tree_add_110_49_pad_groupi_n_1490);
  not csa_tree_add_110_49_pad_groupi_g4295(csa_tree_add_110_49_pad_groupi_n_1503 ,csa_tree_add_110_49_pad_groupi_n_1502);
  xnor csa_tree_add_110_49_pad_groupi_g4296(csa_tree_add_110_49_pad_groupi_n_1502 ,csa_tree_add_110_49_pad_groupi_n_1365 ,csa_tree_add_110_49_pad_groupi_n_1462);
  xnor csa_tree_add_110_49_pad_groupi_g4297(csa_tree_add_110_49_pad_groupi_n_1501 ,csa_tree_add_110_49_pad_groupi_n_1479 ,csa_tree_add_110_49_pad_groupi_n_1466);
  xnor csa_tree_add_110_49_pad_groupi_g4298(csa_tree_add_110_49_pad_groupi_n_1500 ,csa_tree_add_110_49_pad_groupi_n_1459 ,csa_tree_add_110_49_pad_groupi_n_1468);
  xnor csa_tree_add_110_49_pad_groupi_g4299(csa_tree_add_110_49_pad_groupi_n_1499 ,csa_tree_add_110_49_pad_groupi_n_1429 ,csa_tree_add_110_49_pad_groupi_n_1470);
  not csa_tree_add_110_49_pad_groupi_g4300(csa_tree_add_110_49_pad_groupi_n_1498 ,csa_tree_add_110_49_pad_groupi_n_1497);
  xnor csa_tree_add_110_49_pad_groupi_g4301(csa_tree_add_110_49_pad_groupi_n_1497 ,csa_tree_add_110_49_pad_groupi_n_1366 ,csa_tree_add_110_49_pad_groupi_n_1);
  nor csa_tree_add_110_49_pad_groupi_g4302(csa_tree_add_110_49_pad_groupi_n_1495 ,csa_tree_add_110_49_pad_groupi_n_1428 ,csa_tree_add_110_49_pad_groupi_n_1470);
  or csa_tree_add_110_49_pad_groupi_g4303(csa_tree_add_110_49_pad_groupi_n_1494 ,csa_tree_add_110_49_pad_groupi_n_1429 ,csa_tree_add_110_49_pad_groupi_n_1469);
  nor csa_tree_add_110_49_pad_groupi_g4304(csa_tree_add_110_49_pad_groupi_n_1493 ,csa_tree_add_110_49_pad_groupi_n_1458 ,csa_tree_add_110_49_pad_groupi_n_1468);
  or csa_tree_add_110_49_pad_groupi_g4305(csa_tree_add_110_49_pad_groupi_n_1492 ,csa_tree_add_110_49_pad_groupi_n_1459 ,csa_tree_add_110_49_pad_groupi_n_1467);
  nor csa_tree_add_110_49_pad_groupi_g4306(csa_tree_add_110_49_pad_groupi_n_1491 ,csa_tree_add_110_49_pad_groupi_n_1479 ,csa_tree_add_110_49_pad_groupi_n_1466);
  and csa_tree_add_110_49_pad_groupi_g4307(csa_tree_add_110_49_pad_groupi_n_1496 ,csa_tree_add_110_49_pad_groupi_n_1295 ,csa_tree_add_110_49_pad_groupi_n_1475);
  not csa_tree_add_110_49_pad_groupi_g4308(csa_tree_add_110_49_pad_groupi_n_1490 ,csa_tree_add_110_49_pad_groupi_n_1489);
  not csa_tree_add_110_49_pad_groupi_g4309(csa_tree_add_110_49_pad_groupi_n_1488 ,csa_tree_add_110_49_pad_groupi_n_1487);
  xnor csa_tree_add_110_49_pad_groupi_g4310(n_127 ,csa_tree_add_110_49_pad_groupi_n_1460 ,csa_tree_add_110_49_pad_groupi_n_1310);
  or csa_tree_add_110_49_pad_groupi_g4311(csa_tree_add_110_49_pad_groupi_n_1485 ,csa_tree_add_110_49_pad_groupi_n_1478 ,csa_tree_add_110_49_pad_groupi_n_1465);
  xnor csa_tree_add_110_49_pad_groupi_g4312(csa_tree_add_110_49_pad_groupi_n_1484 ,csa_tree_add_110_49_pad_groupi_n_1427 ,csa_tree_add_110_49_pad_groupi_n_1445);
  xnor csa_tree_add_110_49_pad_groupi_g4313(csa_tree_add_110_49_pad_groupi_n_1483 ,csa_tree_add_110_49_pad_groupi_n_1431 ,csa_tree_add_110_49_pad_groupi_n_1447);
  xnor csa_tree_add_110_49_pad_groupi_g4314(csa_tree_add_110_49_pad_groupi_n_1482 ,csa_tree_add_110_49_pad_groupi_n_1439 ,csa_tree_add_110_49_pad_groupi_n_1438);
  xnor csa_tree_add_110_49_pad_groupi_g4315(csa_tree_add_110_49_pad_groupi_n_1489 ,csa_tree_add_110_49_pad_groupi_n_1333 ,csa_tree_add_110_49_pad_groupi_n_1441);
  xnor csa_tree_add_110_49_pad_groupi_g4316(csa_tree_add_110_49_pad_groupi_n_1487 ,csa_tree_add_110_49_pad_groupi_n_1400 ,csa_tree_add_110_49_pad_groupi_n_1440);
  not csa_tree_add_110_49_pad_groupi_g4317(csa_tree_add_110_49_pad_groupi_n_1481 ,csa_tree_add_110_49_pad_groupi_n_1480);
  not csa_tree_add_110_49_pad_groupi_g4318(csa_tree_add_110_49_pad_groupi_n_1479 ,csa_tree_add_110_49_pad_groupi_n_1478);
  not csa_tree_add_110_49_pad_groupi_g4319(csa_tree_add_110_49_pad_groupi_n_1477 ,csa_tree_add_110_49_pad_groupi_n_1476);
  or csa_tree_add_110_49_pad_groupi_g4320(csa_tree_add_110_49_pad_groupi_n_1475 ,csa_tree_add_110_49_pad_groupi_n_1272 ,csa_tree_add_110_49_pad_groupi_n_1460);
  or csa_tree_add_110_49_pad_groupi_g4321(csa_tree_add_110_49_pad_groupi_n_1474 ,csa_tree_add_110_49_pad_groupi_n_1427 ,csa_tree_add_110_49_pad_groupi_n_1444);
  nor csa_tree_add_110_49_pad_groupi_g4322(csa_tree_add_110_49_pad_groupi_n_1473 ,csa_tree_add_110_49_pad_groupi_n_1431 ,csa_tree_add_110_49_pad_groupi_n_1446);
  or csa_tree_add_110_49_pad_groupi_g4323(csa_tree_add_110_49_pad_groupi_n_1472 ,csa_tree_add_110_49_pad_groupi_n_1430 ,csa_tree_add_110_49_pad_groupi_n_1447);
  nor csa_tree_add_110_49_pad_groupi_g4324(csa_tree_add_110_49_pad_groupi_n_1471 ,csa_tree_add_110_49_pad_groupi_n_1426 ,csa_tree_add_110_49_pad_groupi_n_1445);
  and csa_tree_add_110_49_pad_groupi_g4325(csa_tree_add_110_49_pad_groupi_n_1480 ,csa_tree_add_110_49_pad_groupi_n_1407 ,csa_tree_add_110_49_pad_groupi_n_1443);
  and csa_tree_add_110_49_pad_groupi_g4326(csa_tree_add_110_49_pad_groupi_n_1478 ,csa_tree_add_110_49_pad_groupi_n_1390 ,csa_tree_add_110_49_pad_groupi_n_1442);
  or csa_tree_add_110_49_pad_groupi_g4327(csa_tree_add_110_49_pad_groupi_n_1476 ,csa_tree_add_110_49_pad_groupi_n_1378 ,csa_tree_add_110_49_pad_groupi_n_1455);
  not csa_tree_add_110_49_pad_groupi_g4328(csa_tree_add_110_49_pad_groupi_n_1470 ,csa_tree_add_110_49_pad_groupi_n_1469);
  not csa_tree_add_110_49_pad_groupi_g4329(csa_tree_add_110_49_pad_groupi_n_1468 ,csa_tree_add_110_49_pad_groupi_n_1467);
  not csa_tree_add_110_49_pad_groupi_g4330(csa_tree_add_110_49_pad_groupi_n_1466 ,csa_tree_add_110_49_pad_groupi_n_1465);
  xnor csa_tree_add_110_49_pad_groupi_g4331(csa_tree_add_110_49_pad_groupi_n_1464 ,csa_tree_add_110_49_pad_groupi_n_1435 ,csa_tree_add_110_49_pad_groupi_n_1414);
  xnor csa_tree_add_110_49_pad_groupi_g4332(csa_tree_add_110_49_pad_groupi_n_1463 ,csa_tree_add_110_49_pad_groupi_n_1433 ,csa_tree_add_110_49_pad_groupi_n_1412);
  xnor csa_tree_add_110_49_pad_groupi_g4333(csa_tree_add_110_49_pad_groupi_n_1462 ,csa_tree_add_110_49_pad_groupi_n_1239 ,csa_tree_add_110_49_pad_groupi_n_1417);
  xnor csa_tree_add_110_49_pad_groupi_g4334(csa_tree_add_110_49_pad_groupi_n_1461 ,csa_tree_add_110_49_pad_groupi_n_1397 ,csa_tree_add_110_49_pad_groupi_n_1416);
  xnor csa_tree_add_110_49_pad_groupi_g4336(csa_tree_add_110_49_pad_groupi_n_1469 ,csa_tree_add_110_49_pad_groupi_n_1369 ,csa_tree_add_110_49_pad_groupi_n_1404);
  xnor csa_tree_add_110_49_pad_groupi_g4337(csa_tree_add_110_49_pad_groupi_n_1467 ,csa_tree_add_110_49_pad_groupi_n_1350 ,csa_tree_add_110_49_pad_groupi_n_1405);
  xnor csa_tree_add_110_49_pad_groupi_g4338(csa_tree_add_110_49_pad_groupi_n_1465 ,csa_tree_add_110_49_pad_groupi_n_1402 ,csa_tree_add_110_49_pad_groupi_n_1406);
  not csa_tree_add_110_49_pad_groupi_g4339(csa_tree_add_110_49_pad_groupi_n_1459 ,csa_tree_add_110_49_pad_groupi_n_1458);
  not csa_tree_add_110_49_pad_groupi_g4340(csa_tree_add_110_49_pad_groupi_n_1456 ,csa_tree_add_110_49_pad_groupi_n_1457);
  and csa_tree_add_110_49_pad_groupi_g4341(csa_tree_add_110_49_pad_groupi_n_1455 ,csa_tree_add_110_49_pad_groupi_n_1374 ,csa_tree_add_110_49_pad_groupi_n_1417);
  or csa_tree_add_110_49_pad_groupi_g4342(csa_tree_add_110_49_pad_groupi_n_1454 ,csa_tree_add_110_49_pad_groupi_n_1435 ,csa_tree_add_110_49_pad_groupi_n_1413);
  or csa_tree_add_110_49_pad_groupi_g4343(csa_tree_add_110_49_pad_groupi_n_1453 ,csa_tree_add_110_49_pad_groupi_n_1432 ,csa_tree_add_110_49_pad_groupi_n_1412);
  nor csa_tree_add_110_49_pad_groupi_g4344(csa_tree_add_110_49_pad_groupi_n_1452 ,csa_tree_add_110_49_pad_groupi_n_1434 ,csa_tree_add_110_49_pad_groupi_n_1414);
  nor csa_tree_add_110_49_pad_groupi_g4345(csa_tree_add_110_49_pad_groupi_n_1451 ,csa_tree_add_110_49_pad_groupi_n_1396 ,csa_tree_add_110_49_pad_groupi_n_1416);
  or csa_tree_add_110_49_pad_groupi_g4346(csa_tree_add_110_49_pad_groupi_n_1450 ,csa_tree_add_110_49_pad_groupi_n_1397 ,csa_tree_add_110_49_pad_groupi_n_1415);
  nor csa_tree_add_110_49_pad_groupi_g4347(csa_tree_add_110_49_pad_groupi_n_1449 ,csa_tree_add_110_49_pad_groupi_n_1433 ,csa_tree_add_110_49_pad_groupi_n_1411);
  and csa_tree_add_110_49_pad_groupi_g4348(csa_tree_add_110_49_pad_groupi_n_1460 ,csa_tree_add_110_49_pad_groupi_n_1208 ,csa_tree_add_110_49_pad_groupi_n_1420);
  or csa_tree_add_110_49_pad_groupi_g4349(csa_tree_add_110_49_pad_groupi_n_1458 ,csa_tree_add_110_49_pad_groupi_n_1391 ,csa_tree_add_110_49_pad_groupi_n_1425);
  or csa_tree_add_110_49_pad_groupi_g4350(csa_tree_add_110_49_pad_groupi_n_1457 ,csa_tree_add_110_49_pad_groupi_n_1393 ,csa_tree_add_110_49_pad_groupi_n_1424);
  not csa_tree_add_110_49_pad_groupi_g4351(csa_tree_add_110_49_pad_groupi_n_1447 ,csa_tree_add_110_49_pad_groupi_n_1446);
  not csa_tree_add_110_49_pad_groupi_g4352(csa_tree_add_110_49_pad_groupi_n_1445 ,csa_tree_add_110_49_pad_groupi_n_1444);
  or csa_tree_add_110_49_pad_groupi_g4353(csa_tree_add_110_49_pad_groupi_n_1443 ,csa_tree_add_110_49_pad_groupi_n_1401 ,csa_tree_add_110_49_pad_groupi_n_1409);
  or csa_tree_add_110_49_pad_groupi_g4354(csa_tree_add_110_49_pad_groupi_n_1442 ,csa_tree_add_110_49_pad_groupi_n_1379 ,csa_tree_add_110_49_pad_groupi_n_1418);
  xnor csa_tree_add_110_49_pad_groupi_g4355(csa_tree_add_110_49_pad_groupi_n_1441 ,csa_tree_add_110_49_pad_groupi_n_1336 ,csa_tree_add_110_49_pad_groupi_n_1386);
  xnor csa_tree_add_110_49_pad_groupi_g4356(csa_tree_add_110_49_pad_groupi_n_1440 ,csa_tree_add_110_49_pad_groupi_n_1279 ,csa_tree_add_110_49_pad_groupi_n_1381);
  nor csa_tree_add_110_49_pad_groupi_g4357(csa_tree_add_110_49_pad_groupi_n_1439 ,csa_tree_add_110_49_pad_groupi_n_1342 ,csa_tree_add_110_49_pad_groupi_n_1408);
  xnor csa_tree_add_110_49_pad_groupi_g4358(csa_tree_add_110_49_pad_groupi_n_1438 ,csa_tree_add_110_49_pad_groupi_n_1354 ,csa_tree_add_110_49_pad_groupi_n_1371);
  xnor csa_tree_add_110_49_pad_groupi_g4359(csa_tree_add_110_49_pad_groupi_n_1437 ,csa_tree_add_110_49_pad_groupi_n_1399 ,csa_tree_add_110_49_pad_groupi_n_1385);
  xnor csa_tree_add_110_49_pad_groupi_g4360(csa_tree_add_110_49_pad_groupi_n_1436 ,csa_tree_add_110_49_pad_groupi_n_1261 ,csa_tree_add_110_49_pad_groupi_n_1383);
  and csa_tree_add_110_49_pad_groupi_g4361(csa_tree_add_110_49_pad_groupi_n_1448 ,csa_tree_add_110_49_pad_groupi_n_1377 ,csa_tree_add_110_49_pad_groupi_n_1410);
  xnor csa_tree_add_110_49_pad_groupi_g4362(csa_tree_add_110_49_pad_groupi_n_1446 ,csa_tree_add_110_49_pad_groupi_n_1351 ,csa_tree_add_110_49_pad_groupi_n_1372);
  xnor csa_tree_add_110_49_pad_groupi_g4363(csa_tree_add_110_49_pad_groupi_n_1444 ,csa_tree_add_110_49_pad_groupi_n_1316 ,csa_tree_add_110_49_pad_groupi_n_1370);
  not csa_tree_add_110_49_pad_groupi_g4364(csa_tree_add_110_49_pad_groupi_n_1434 ,csa_tree_add_110_49_pad_groupi_n_1435);
  not csa_tree_add_110_49_pad_groupi_g4365(csa_tree_add_110_49_pad_groupi_n_1432 ,csa_tree_add_110_49_pad_groupi_n_1433);
  not csa_tree_add_110_49_pad_groupi_g4366(csa_tree_add_110_49_pad_groupi_n_1430 ,csa_tree_add_110_49_pad_groupi_n_1431);
  not csa_tree_add_110_49_pad_groupi_g4367(csa_tree_add_110_49_pad_groupi_n_1429 ,csa_tree_add_110_49_pad_groupi_n_1428);
  not csa_tree_add_110_49_pad_groupi_g4368(csa_tree_add_110_49_pad_groupi_n_1426 ,csa_tree_add_110_49_pad_groupi_n_1427);
  and csa_tree_add_110_49_pad_groupi_g4369(csa_tree_add_110_49_pad_groupi_n_1425 ,csa_tree_add_110_49_pad_groupi_n_1369 ,csa_tree_add_110_49_pad_groupi_n_1373);
  nor csa_tree_add_110_49_pad_groupi_g4370(csa_tree_add_110_49_pad_groupi_n_1424 ,csa_tree_add_110_49_pad_groupi_n_1368 ,csa_tree_add_110_49_pad_groupi_n_1392);
  nor csa_tree_add_110_49_pad_groupi_g4371(csa_tree_add_110_49_pad_groupi_n_1423 ,csa_tree_add_110_49_pad_groupi_n_1260 ,csa_tree_add_110_49_pad_groupi_n_1383);
  or csa_tree_add_110_49_pad_groupi_g4372(csa_tree_add_110_49_pad_groupi_n_1422 ,csa_tree_add_110_49_pad_groupi_n_1261 ,csa_tree_add_110_49_pad_groupi_n_1382);
  nor csa_tree_add_110_49_pad_groupi_g4373(csa_tree_add_110_49_pad_groupi_n_1421 ,csa_tree_add_110_49_pad_groupi_n_1398 ,csa_tree_add_110_49_pad_groupi_n_1385);
  or csa_tree_add_110_49_pad_groupi_g4374(csa_tree_add_110_49_pad_groupi_n_1420 ,csa_tree_add_110_49_pad_groupi_n_1213 ,csa_tree_add_110_49_pad_groupi_n_1389);
  or csa_tree_add_110_49_pad_groupi_g4375(csa_tree_add_110_49_pad_groupi_n_1419 ,csa_tree_add_110_49_pad_groupi_n_1399 ,csa_tree_add_110_49_pad_groupi_n_1384);
  and csa_tree_add_110_49_pad_groupi_g4376(csa_tree_add_110_49_pad_groupi_n_1435 ,csa_tree_add_110_49_pad_groupi_n_1357 ,csa_tree_add_110_49_pad_groupi_n_1388);
  or csa_tree_add_110_49_pad_groupi_g4377(csa_tree_add_110_49_pad_groupi_n_1433 ,csa_tree_add_110_49_pad_groupi_n_1270 ,csa_tree_add_110_49_pad_groupi_n_1387);
  or csa_tree_add_110_49_pad_groupi_g4378(csa_tree_add_110_49_pad_groupi_n_1431 ,csa_tree_add_110_49_pad_groupi_n_1362 ,csa_tree_add_110_49_pad_groupi_n_1394);
  or csa_tree_add_110_49_pad_groupi_g4379(csa_tree_add_110_49_pad_groupi_n_1428 ,csa_tree_add_110_49_pad_groupi_n_1345 ,csa_tree_add_110_49_pad_groupi_n_1375);
  and csa_tree_add_110_49_pad_groupi_g4380(csa_tree_add_110_49_pad_groupi_n_1427 ,csa_tree_add_110_49_pad_groupi_n_1313 ,csa_tree_add_110_49_pad_groupi_n_1395);
  not csa_tree_add_110_49_pad_groupi_g4382(csa_tree_add_110_49_pad_groupi_n_1416 ,csa_tree_add_110_49_pad_groupi_n_1415);
  not csa_tree_add_110_49_pad_groupi_g4383(csa_tree_add_110_49_pad_groupi_n_1414 ,csa_tree_add_110_49_pad_groupi_n_1413);
  not csa_tree_add_110_49_pad_groupi_g4384(csa_tree_add_110_49_pad_groupi_n_1412 ,csa_tree_add_110_49_pad_groupi_n_1411);
  or csa_tree_add_110_49_pad_groupi_g4385(csa_tree_add_110_49_pad_groupi_n_1410 ,csa_tree_add_110_49_pad_groupi_n_1403 ,csa_tree_add_110_49_pad_groupi_n_1376);
  nor csa_tree_add_110_49_pad_groupi_g4386(csa_tree_add_110_49_pad_groupi_n_1409 ,csa_tree_add_110_49_pad_groupi_n_1278 ,csa_tree_add_110_49_pad_groupi_n_1381);
  and csa_tree_add_110_49_pad_groupi_g4387(csa_tree_add_110_49_pad_groupi_n_1408 ,csa_tree_add_110_49_pad_groupi_n_1343 ,csa_tree_add_110_49_pad_groupi_n_1386);
  or csa_tree_add_110_49_pad_groupi_g4388(csa_tree_add_110_49_pad_groupi_n_1407 ,csa_tree_add_110_49_pad_groupi_n_1279 ,csa_tree_add_110_49_pad_groupi_n_1380);
  xnor csa_tree_add_110_49_pad_groupi_g4389(csa_tree_add_110_49_pad_groupi_n_1406 ,csa_tree_add_110_49_pad_groupi_n_1318 ,csa_tree_add_110_49_pad_groupi_n_1349);
  xor csa_tree_add_110_49_pad_groupi_g4390(csa_tree_add_110_49_pad_groupi_n_1405 ,csa_tree_add_110_49_pad_groupi_n_1368 ,csa_tree_add_110_49_pad_groupi_n_1296);
  xnor csa_tree_add_110_49_pad_groupi_g4391(csa_tree_add_110_49_pad_groupi_n_1404 ,csa_tree_add_110_49_pad_groupi_n_1284 ,csa_tree_add_110_49_pad_groupi_n_1347);
  xnor csa_tree_add_110_49_pad_groupi_g4392(csa_tree_add_110_49_pad_groupi_n_1418 ,csa_tree_add_110_49_pad_groupi_n_1302 ,csa_tree_add_110_49_pad_groupi_n_1340);
  xnor csa_tree_add_110_49_pad_groupi_g4393(csa_tree_add_110_49_pad_groupi_n_1417 ,csa_tree_add_110_49_pad_groupi_n_1240 ,csa_tree_add_110_49_pad_groupi_n_1339);
  xnor csa_tree_add_110_49_pad_groupi_g4394(csa_tree_add_110_49_pad_groupi_n_1415 ,csa_tree_add_110_49_pad_groupi_n_1353 ,csa_tree_add_110_49_pad_groupi_n_1307);
  xnor csa_tree_add_110_49_pad_groupi_g4395(csa_tree_add_110_49_pad_groupi_n_1413 ,csa_tree_add_110_49_pad_groupi_n_1352 ,csa_tree_add_110_49_pad_groupi_n_1341);
  xnor csa_tree_add_110_49_pad_groupi_g4396(csa_tree_add_110_49_pad_groupi_n_1411 ,csa_tree_add_110_49_pad_groupi_n_1320 ,csa_tree_add_110_49_pad_groupi_n_1338);
  not csa_tree_add_110_49_pad_groupi_g4397(csa_tree_add_110_49_pad_groupi_n_1403 ,csa_tree_add_110_49_pad_groupi_n_1402);
  not csa_tree_add_110_49_pad_groupi_g4398(csa_tree_add_110_49_pad_groupi_n_1401 ,csa_tree_add_110_49_pad_groupi_n_1400);
  not csa_tree_add_110_49_pad_groupi_g4399(csa_tree_add_110_49_pad_groupi_n_1398 ,csa_tree_add_110_49_pad_groupi_n_1399);
  not csa_tree_add_110_49_pad_groupi_g4400(csa_tree_add_110_49_pad_groupi_n_1397 ,csa_tree_add_110_49_pad_groupi_n_1396);
  or csa_tree_add_110_49_pad_groupi_g4401(csa_tree_add_110_49_pad_groupi_n_1395 ,csa_tree_add_110_49_pad_groupi_n_1314 ,csa_tree_add_110_49_pad_groupi_n_1352);
  and csa_tree_add_110_49_pad_groupi_g4402(csa_tree_add_110_49_pad_groupi_n_1394 ,csa_tree_add_110_49_pad_groupi_n_1337 ,csa_tree_add_110_49_pad_groupi_n_1363);
  nor csa_tree_add_110_49_pad_groupi_g4403(csa_tree_add_110_49_pad_groupi_n_1393 ,csa_tree_add_110_49_pad_groupi_n_1297 ,csa_tree_add_110_49_pad_groupi_n_1350);
  and csa_tree_add_110_49_pad_groupi_g4404(csa_tree_add_110_49_pad_groupi_n_1392 ,csa_tree_add_110_49_pad_groupi_n_1297 ,csa_tree_add_110_49_pad_groupi_n_1350);
  nor csa_tree_add_110_49_pad_groupi_g4405(csa_tree_add_110_49_pad_groupi_n_1391 ,csa_tree_add_110_49_pad_groupi_n_1284 ,csa_tree_add_110_49_pad_groupi_n_1346);
  or csa_tree_add_110_49_pad_groupi_g4406(csa_tree_add_110_49_pad_groupi_n_1390 ,csa_tree_add_110_49_pad_groupi_n_1237 ,csa_tree_add_110_49_pad_groupi_n_1367);
  nor csa_tree_add_110_49_pad_groupi_g4407(csa_tree_add_110_49_pad_groupi_n_1389 ,csa_tree_add_110_49_pad_groupi_n_1123 ,csa_tree_add_110_49_pad_groupi_n_1355);
  or csa_tree_add_110_49_pad_groupi_g4408(csa_tree_add_110_49_pad_groupi_n_1388 ,csa_tree_add_110_49_pad_groupi_n_1300 ,csa_tree_add_110_49_pad_groupi_n_1358);
  and csa_tree_add_110_49_pad_groupi_g4409(csa_tree_add_110_49_pad_groupi_n_1387 ,csa_tree_add_110_49_pad_groupi_n_1271 ,csa_tree_add_110_49_pad_groupi_n_1353);
  or csa_tree_add_110_49_pad_groupi_g4410(csa_tree_add_110_49_pad_groupi_n_1402 ,csa_tree_add_110_49_pad_groupi_n_1329 ,csa_tree_add_110_49_pad_groupi_n_1360);
  or csa_tree_add_110_49_pad_groupi_g4411(csa_tree_add_110_49_pad_groupi_n_1400 ,csa_tree_add_110_49_pad_groupi_n_1324 ,csa_tree_add_110_49_pad_groupi_n_1356);
  and csa_tree_add_110_49_pad_groupi_g4412(csa_tree_add_110_49_pad_groupi_n_1399 ,csa_tree_add_110_49_pad_groupi_n_1255 ,csa_tree_add_110_49_pad_groupi_n_1361);
  or csa_tree_add_110_49_pad_groupi_g4413(csa_tree_add_110_49_pad_groupi_n_1396 ,csa_tree_add_110_49_pad_groupi_n_1311 ,csa_tree_add_110_49_pad_groupi_n_1359);
  not csa_tree_add_110_49_pad_groupi_g4414(csa_tree_add_110_49_pad_groupi_n_1385 ,csa_tree_add_110_49_pad_groupi_n_1384);
  not csa_tree_add_110_49_pad_groupi_g4415(csa_tree_add_110_49_pad_groupi_n_1383 ,csa_tree_add_110_49_pad_groupi_n_1382);
  not csa_tree_add_110_49_pad_groupi_g4416(csa_tree_add_110_49_pad_groupi_n_1381 ,csa_tree_add_110_49_pad_groupi_n_1380);
  and csa_tree_add_110_49_pad_groupi_g4417(csa_tree_add_110_49_pad_groupi_n_1379 ,csa_tree_add_110_49_pad_groupi_n_1237 ,csa_tree_add_110_49_pad_groupi_n_1367);
  nor csa_tree_add_110_49_pad_groupi_g4418(csa_tree_add_110_49_pad_groupi_n_1378 ,csa_tree_add_110_49_pad_groupi_n_1239 ,csa_tree_add_110_49_pad_groupi_n_1365);
  or csa_tree_add_110_49_pad_groupi_g4419(csa_tree_add_110_49_pad_groupi_n_1377 ,csa_tree_add_110_49_pad_groupi_n_1318 ,csa_tree_add_110_49_pad_groupi_n_1348);
  nor csa_tree_add_110_49_pad_groupi_g4420(csa_tree_add_110_49_pad_groupi_n_1376 ,csa_tree_add_110_49_pad_groupi_n_1317 ,csa_tree_add_110_49_pad_groupi_n_1349);
  nor csa_tree_add_110_49_pad_groupi_g4421(csa_tree_add_110_49_pad_groupi_n_1375 ,csa_tree_add_110_49_pad_groupi_n_1351 ,csa_tree_add_110_49_pad_groupi_n_1344);
  or csa_tree_add_110_49_pad_groupi_g4422(csa_tree_add_110_49_pad_groupi_n_1374 ,csa_tree_add_110_49_pad_groupi_n_1238 ,csa_tree_add_110_49_pad_groupi_n_1364);
  or csa_tree_add_110_49_pad_groupi_g4423(csa_tree_add_110_49_pad_groupi_n_1373 ,csa_tree_add_110_49_pad_groupi_n_1283 ,csa_tree_add_110_49_pad_groupi_n_1347);
  xnor csa_tree_add_110_49_pad_groupi_g4424(csa_tree_add_110_49_pad_groupi_n_1372 ,csa_tree_add_110_49_pad_groupi_n_1334 ,csa_tree_add_110_49_pad_groupi_n_1276);
  xnor csa_tree_add_110_49_pad_groupi_g4425(csa_tree_add_110_49_pad_groupi_n_1371 ,csa_tree_add_110_49_pad_groupi_n_1244 ,csa_tree_add_110_49_pad_groupi_n_1309);
  xnor csa_tree_add_110_49_pad_groupi_g4426(csa_tree_add_110_49_pad_groupi_n_1370 ,csa_tree_add_110_49_pad_groupi_n_1337 ,csa_tree_add_110_49_pad_groupi_n_1275);
  xnor csa_tree_add_110_49_pad_groupi_g4427(csa_tree_add_110_49_pad_groupi_n_1386 ,csa_tree_add_110_49_pad_groupi_n_1242 ,csa_tree_add_110_49_pad_groupi_n_1306);
  xnor csa_tree_add_110_49_pad_groupi_g4428(csa_tree_add_110_49_pad_groupi_n_1384 ,csa_tree_add_110_49_pad_groupi_n_1280 ,csa_tree_add_110_49_pad_groupi_n_1305);
  xnor csa_tree_add_110_49_pad_groupi_g4429(csa_tree_add_110_49_pad_groupi_n_1382 ,csa_tree_add_110_49_pad_groupi_n_1321 ,csa_tree_add_110_49_pad_groupi_n_1268);
  xnor csa_tree_add_110_49_pad_groupi_g4430(csa_tree_add_110_49_pad_groupi_n_1380 ,csa_tree_add_110_49_pad_groupi_n_1243 ,csa_tree_add_110_49_pad_groupi_n_1308);
  not csa_tree_add_110_49_pad_groupi_g4431(csa_tree_add_110_49_pad_groupi_n_1367 ,csa_tree_add_110_49_pad_groupi_n_1366);
  not csa_tree_add_110_49_pad_groupi_g4432(csa_tree_add_110_49_pad_groupi_n_1365 ,csa_tree_add_110_49_pad_groupi_n_1364);
  or csa_tree_add_110_49_pad_groupi_g4433(csa_tree_add_110_49_pad_groupi_n_1363 ,csa_tree_add_110_49_pad_groupi_n_287 ,csa_tree_add_110_49_pad_groupi_n_1316);
  nor csa_tree_add_110_49_pad_groupi_g4434(csa_tree_add_110_49_pad_groupi_n_1362 ,csa_tree_add_110_49_pad_groupi_n_187 ,csa_tree_add_110_49_pad_groupi_n_1315);
  or csa_tree_add_110_49_pad_groupi_g4435(csa_tree_add_110_49_pad_groupi_n_1361 ,csa_tree_add_110_49_pad_groupi_n_1254 ,csa_tree_add_110_49_pad_groupi_n_1321);
  and csa_tree_add_110_49_pad_groupi_g4436(csa_tree_add_110_49_pad_groupi_n_1360 ,csa_tree_add_110_49_pad_groupi_n_1328 ,csa_tree_add_110_49_pad_groupi_n_1302);
  nor csa_tree_add_110_49_pad_groupi_g4437(csa_tree_add_110_49_pad_groupi_n_1359 ,csa_tree_add_110_49_pad_groupi_n_1262 ,csa_tree_add_110_49_pad_groupi_n_1312);
  nor csa_tree_add_110_49_pad_groupi_g4438(csa_tree_add_110_49_pad_groupi_n_1358 ,csa_tree_add_110_49_pad_groupi_n_1227 ,csa_tree_add_110_49_pad_groupi_n_1320);
  or csa_tree_add_110_49_pad_groupi_g4439(csa_tree_add_110_49_pad_groupi_n_1357 ,csa_tree_add_110_49_pad_groupi_n_1228 ,csa_tree_add_110_49_pad_groupi_n_1319);
  and csa_tree_add_110_49_pad_groupi_g4440(csa_tree_add_110_49_pad_groupi_n_1356 ,csa_tree_add_110_49_pad_groupi_n_1331 ,csa_tree_add_110_49_pad_groupi_n_1240);
  nor csa_tree_add_110_49_pad_groupi_g4441(csa_tree_add_110_49_pad_groupi_n_1355 ,csa_tree_add_110_49_pad_groupi_n_1122 ,csa_tree_add_110_49_pad_groupi_n_1326);
  nor csa_tree_add_110_49_pad_groupi_g4442(csa_tree_add_110_49_pad_groupi_n_1354 ,csa_tree_add_110_49_pad_groupi_n_1292 ,csa_tree_add_110_49_pad_groupi_n_1322);
  or csa_tree_add_110_49_pad_groupi_g4443(csa_tree_add_110_49_pad_groupi_n_1369 ,csa_tree_add_110_49_pad_groupi_n_1212 ,csa_tree_add_110_49_pad_groupi_n_1327);
  and csa_tree_add_110_49_pad_groupi_g4444(csa_tree_add_110_49_pad_groupi_n_1368 ,csa_tree_add_110_49_pad_groupi_n_1249 ,csa_tree_add_110_49_pad_groupi_n_1325);
  or csa_tree_add_110_49_pad_groupi_g4445(csa_tree_add_110_49_pad_groupi_n_1366 ,csa_tree_add_110_49_pad_groupi_n_1293 ,csa_tree_add_110_49_pad_groupi_n_1330);
  or csa_tree_add_110_49_pad_groupi_g4446(csa_tree_add_110_49_pad_groupi_n_1364 ,csa_tree_add_110_49_pad_groupi_n_1206 ,csa_tree_add_110_49_pad_groupi_n_1323);
  not csa_tree_add_110_49_pad_groupi_g4447(csa_tree_add_110_49_pad_groupi_n_1349 ,csa_tree_add_110_49_pad_groupi_n_1348);
  not csa_tree_add_110_49_pad_groupi_g4448(csa_tree_add_110_49_pad_groupi_n_1347 ,csa_tree_add_110_49_pad_groupi_n_1346);
  nor csa_tree_add_110_49_pad_groupi_g4449(csa_tree_add_110_49_pad_groupi_n_1345 ,csa_tree_add_110_49_pad_groupi_n_1334 ,csa_tree_add_110_49_pad_groupi_n_1277);
  and csa_tree_add_110_49_pad_groupi_g4450(csa_tree_add_110_49_pad_groupi_n_1344 ,csa_tree_add_110_49_pad_groupi_n_1334 ,csa_tree_add_110_49_pad_groupi_n_1277);
  or csa_tree_add_110_49_pad_groupi_g4451(csa_tree_add_110_49_pad_groupi_n_1343 ,csa_tree_add_110_49_pad_groupi_n_1332 ,csa_tree_add_110_49_pad_groupi_n_1335);
  nor csa_tree_add_110_49_pad_groupi_g4452(csa_tree_add_110_49_pad_groupi_n_1342 ,csa_tree_add_110_49_pad_groupi_n_1333 ,csa_tree_add_110_49_pad_groupi_n_1336);
  xnor csa_tree_add_110_49_pad_groupi_g4453(csa_tree_add_110_49_pad_groupi_n_1341 ,csa_tree_add_110_49_pad_groupi_n_1230 ,csa_tree_add_110_49_pad_groupi_n_1299);
  xnor csa_tree_add_110_49_pad_groupi_g4454(csa_tree_add_110_49_pad_groupi_n_1340 ,csa_tree_add_110_49_pad_groupi_n_625 ,csa_tree_add_110_49_pad_groupi_n_1274);
  xnor csa_tree_add_110_49_pad_groupi_g4455(csa_tree_add_110_49_pad_groupi_n_1339 ,csa_tree_add_110_49_pad_groupi_n_1282 ,csa_tree_add_110_49_pad_groupi_n_1184);
  xnor csa_tree_add_110_49_pad_groupi_g4456(csa_tree_add_110_49_pad_groupi_n_1338 ,csa_tree_add_110_49_pad_groupi_n_1228 ,csa_tree_add_110_49_pad_groupi_n_1300);
  xnor csa_tree_add_110_49_pad_groupi_g4457(csa_tree_add_110_49_pad_groupi_n_1353 ,csa_tree_add_110_49_pad_groupi_n_1155 ,csa_tree_add_110_49_pad_groupi_n_1267);
  xnor csa_tree_add_110_49_pad_groupi_g4458(csa_tree_add_110_49_pad_groupi_n_1352 ,csa_tree_add_110_49_pad_groupi_n_1218 ,csa_tree_add_110_49_pad_groupi_n_1265);
  xnor csa_tree_add_110_49_pad_groupi_g4459(csa_tree_add_110_49_pad_groupi_n_1351 ,csa_tree_add_110_49_pad_groupi_n_1301 ,csa_tree_add_110_49_pad_groupi_n_1223);
  xnor csa_tree_add_110_49_pad_groupi_g4460(csa_tree_add_110_49_pad_groupi_n_1350 ,csa_tree_add_110_49_pad_groupi_n_1285 ,csa_tree_add_110_49_pad_groupi_n_1221);
  xnor csa_tree_add_110_49_pad_groupi_g4461(csa_tree_add_110_49_pad_groupi_n_1348 ,csa_tree_add_110_49_pad_groupi_n_1217 ,csa_tree_add_110_49_pad_groupi_n_1266);
  xnor csa_tree_add_110_49_pad_groupi_g4462(csa_tree_add_110_49_pad_groupi_n_1346 ,csa_tree_add_110_49_pad_groupi_n_1303 ,csa_tree_add_110_49_pad_groupi_n_1269);
  not csa_tree_add_110_49_pad_groupi_g4463(csa_tree_add_110_49_pad_groupi_n_1336 ,csa_tree_add_110_49_pad_groupi_n_1335);
  not csa_tree_add_110_49_pad_groupi_g4464(csa_tree_add_110_49_pad_groupi_n_1332 ,csa_tree_add_110_49_pad_groupi_n_1333);
  or csa_tree_add_110_49_pad_groupi_g4465(csa_tree_add_110_49_pad_groupi_n_1331 ,csa_tree_add_110_49_pad_groupi_n_286 ,csa_tree_add_110_49_pad_groupi_n_1281);
  and csa_tree_add_110_49_pad_groupi_g4466(csa_tree_add_110_49_pad_groupi_n_1330 ,csa_tree_add_110_49_pad_groupi_n_1291 ,csa_tree_add_110_49_pad_groupi_n_1243);
  nor csa_tree_add_110_49_pad_groupi_g4467(csa_tree_add_110_49_pad_groupi_n_1329 ,csa_tree_add_110_49_pad_groupi_n_624 ,csa_tree_add_110_49_pad_groupi_n_1274);
  or csa_tree_add_110_49_pad_groupi_g4468(csa_tree_add_110_49_pad_groupi_n_1328 ,csa_tree_add_110_49_pad_groupi_n_625 ,csa_tree_add_110_49_pad_groupi_n_1273);
  and csa_tree_add_110_49_pad_groupi_g4469(csa_tree_add_110_49_pad_groupi_n_1327 ,csa_tree_add_110_49_pad_groupi_n_1210 ,csa_tree_add_110_49_pad_groupi_n_1301);
  nor csa_tree_add_110_49_pad_groupi_g4470(csa_tree_add_110_49_pad_groupi_n_1326 ,csa_tree_add_110_49_pad_groupi_n_1139 ,csa_tree_add_110_49_pad_groupi_n_1288);
  or csa_tree_add_110_49_pad_groupi_g4471(csa_tree_add_110_49_pad_groupi_n_1325 ,csa_tree_add_110_49_pad_groupi_n_1248 ,csa_tree_add_110_49_pad_groupi_n_1304);
  nor csa_tree_add_110_49_pad_groupi_g4472(csa_tree_add_110_49_pad_groupi_n_1324 ,csa_tree_add_110_49_pad_groupi_n_188 ,csa_tree_add_110_49_pad_groupi_n_1282);
  nor csa_tree_add_110_49_pad_groupi_g4473(csa_tree_add_110_49_pad_groupi_n_1323 ,csa_tree_add_110_49_pad_groupi_n_1205 ,csa_tree_add_110_49_pad_groupi_n_1285);
  nor csa_tree_add_110_49_pad_groupi_g4474(csa_tree_add_110_49_pad_groupi_n_1322 ,csa_tree_add_110_49_pad_groupi_n_1242 ,csa_tree_add_110_49_pad_groupi_n_1287);
  or csa_tree_add_110_49_pad_groupi_g4475(csa_tree_add_110_49_pad_groupi_n_1337 ,csa_tree_add_110_49_pad_groupi_n_1250 ,csa_tree_add_110_49_pad_groupi_n_1294);
  or csa_tree_add_110_49_pad_groupi_g4476(csa_tree_add_110_49_pad_groupi_n_1335 ,csa_tree_add_110_49_pad_groupi_n_1247 ,csa_tree_add_110_49_pad_groupi_n_1290);
  and csa_tree_add_110_49_pad_groupi_g4477(csa_tree_add_110_49_pad_groupi_n_1334 ,csa_tree_add_110_49_pad_groupi_n_1207 ,csa_tree_add_110_49_pad_groupi_n_1286);
  and csa_tree_add_110_49_pad_groupi_g4478(csa_tree_add_110_49_pad_groupi_n_1333 ,csa_tree_add_110_49_pad_groupi_n_691 ,csa_tree_add_110_49_pad_groupi_n_1289);
  not csa_tree_add_110_49_pad_groupi_g4479(csa_tree_add_110_49_pad_groupi_n_1320 ,csa_tree_add_110_49_pad_groupi_n_1319);
  not csa_tree_add_110_49_pad_groupi_g4480(csa_tree_add_110_49_pad_groupi_n_1318 ,csa_tree_add_110_49_pad_groupi_n_1317);
  not csa_tree_add_110_49_pad_groupi_g4481(csa_tree_add_110_49_pad_groupi_n_1316 ,csa_tree_add_110_49_pad_groupi_n_1315);
  nor csa_tree_add_110_49_pad_groupi_g4482(csa_tree_add_110_49_pad_groupi_n_1314 ,csa_tree_add_110_49_pad_groupi_n_1230 ,csa_tree_add_110_49_pad_groupi_n_1299);
  or csa_tree_add_110_49_pad_groupi_g4483(csa_tree_add_110_49_pad_groupi_n_1313 ,csa_tree_add_110_49_pad_groupi_n_1229 ,csa_tree_add_110_49_pad_groupi_n_1298);
  nor csa_tree_add_110_49_pad_groupi_g4484(csa_tree_add_110_49_pad_groupi_n_1312 ,csa_tree_add_110_49_pad_groupi_n_1225 ,csa_tree_add_110_49_pad_groupi_n_1280);
  and csa_tree_add_110_49_pad_groupi_g4485(csa_tree_add_110_49_pad_groupi_n_1311 ,csa_tree_add_110_49_pad_groupi_n_1225 ,csa_tree_add_110_49_pad_groupi_n_1280);
  xnor csa_tree_add_110_49_pad_groupi_g4486(csa_tree_add_110_49_pad_groupi_n_1310 ,csa_tree_add_110_49_pad_groupi_n_1185 ,csa_tree_add_110_49_pad_groupi_n_1226);
  xnor csa_tree_add_110_49_pad_groupi_g4487(csa_tree_add_110_49_pad_groupi_n_1309 ,csa_tree_add_110_49_pad_groupi_n_1055 ,csa_tree_add_110_49_pad_groupi_n_1222);
  xnor csa_tree_add_110_49_pad_groupi_g4488(csa_tree_add_110_49_pad_groupi_n_1308 ,csa_tree_add_110_49_pad_groupi_n_634 ,csa_tree_add_110_49_pad_groupi_n_1234);
  xnor csa_tree_add_110_49_pad_groupi_g4489(csa_tree_add_110_49_pad_groupi_n_1307 ,csa_tree_add_110_49_pad_groupi_n_1188 ,csa_tree_add_110_49_pad_groupi_n_1232);
  xnor csa_tree_add_110_49_pad_groupi_g4490(csa_tree_add_110_49_pad_groupi_n_1306 ,csa_tree_add_110_49_pad_groupi_n_575 ,csa_tree_add_110_49_pad_groupi_n_1236);
  xnor csa_tree_add_110_49_pad_groupi_g4491(csa_tree_add_110_49_pad_groupi_n_1305 ,csa_tree_add_110_49_pad_groupi_n_1262 ,csa_tree_add_110_49_pad_groupi_n_1225);
  xnor csa_tree_add_110_49_pad_groupi_g4492(csa_tree_add_110_49_pad_groupi_n_1321 ,csa_tree_add_110_49_pad_groupi_n_1014 ,csa_tree_add_110_49_pad_groupi_n_1224);
  xnor csa_tree_add_110_49_pad_groupi_g4493(csa_tree_add_110_49_pad_groupi_n_1319 ,csa_tree_add_110_49_pad_groupi_n_1196 ,csa_tree_add_110_49_pad_groupi_n_1220);
  xnor csa_tree_add_110_49_pad_groupi_g4494(csa_tree_add_110_49_pad_groupi_n_1317 ,csa_tree_add_110_49_pad_groupi_n_1263 ,csa_tree_add_110_49_pad_groupi_n_799);
  xnor csa_tree_add_110_49_pad_groupi_g4495(csa_tree_add_110_49_pad_groupi_n_1315 ,csa_tree_add_110_49_pad_groupi_n_1241 ,csa_tree_add_110_49_pad_groupi_n_1219);
  not csa_tree_add_110_49_pad_groupi_g4496(csa_tree_add_110_49_pad_groupi_n_1304 ,csa_tree_add_110_49_pad_groupi_n_1303);
  not csa_tree_add_110_49_pad_groupi_g4497(csa_tree_add_110_49_pad_groupi_n_1298 ,csa_tree_add_110_49_pad_groupi_n_1299);
  not csa_tree_add_110_49_pad_groupi_g4498(csa_tree_add_110_49_pad_groupi_n_1297 ,csa_tree_add_110_49_pad_groupi_n_1296);
  or csa_tree_add_110_49_pad_groupi_g4499(csa_tree_add_110_49_pad_groupi_n_1295 ,csa_tree_add_110_49_pad_groupi_n_1186 ,csa_tree_add_110_49_pad_groupi_n_1226);
  and csa_tree_add_110_49_pad_groupi_g4500(csa_tree_add_110_49_pad_groupi_n_1294 ,csa_tree_add_110_49_pad_groupi_n_1218 ,csa_tree_add_110_49_pad_groupi_n_1258);
  nor csa_tree_add_110_49_pad_groupi_g4501(csa_tree_add_110_49_pad_groupi_n_1293 ,csa_tree_add_110_49_pad_groupi_n_633 ,csa_tree_add_110_49_pad_groupi_n_1234);
  and csa_tree_add_110_49_pad_groupi_g4502(csa_tree_add_110_49_pad_groupi_n_1292 ,csa_tree_add_110_49_pad_groupi_n_575 ,csa_tree_add_110_49_pad_groupi_n_1235);
  or csa_tree_add_110_49_pad_groupi_g4503(csa_tree_add_110_49_pad_groupi_n_1291 ,csa_tree_add_110_49_pad_groupi_n_634 ,csa_tree_add_110_49_pad_groupi_n_1233);
  and csa_tree_add_110_49_pad_groupi_g4504(csa_tree_add_110_49_pad_groupi_n_1290 ,csa_tree_add_110_49_pad_groupi_n_1217 ,csa_tree_add_110_49_pad_groupi_n_1246);
  or csa_tree_add_110_49_pad_groupi_g4505(csa_tree_add_110_49_pad_groupi_n_1289 ,csa_tree_add_110_49_pad_groupi_n_690 ,csa_tree_add_110_49_pad_groupi_n_1264);
  nor csa_tree_add_110_49_pad_groupi_g4506(csa_tree_add_110_49_pad_groupi_n_1288 ,csa_tree_add_110_49_pad_groupi_n_1146 ,csa_tree_add_110_49_pad_groupi_n_1253);
  and csa_tree_add_110_49_pad_groupi_g4507(csa_tree_add_110_49_pad_groupi_n_1287 ,csa_tree_add_110_49_pad_groupi_n_574 ,csa_tree_add_110_49_pad_groupi_n_1236);
  or csa_tree_add_110_49_pad_groupi_g4508(csa_tree_add_110_49_pad_groupi_n_1286 ,csa_tree_add_110_49_pad_groupi_n_1215 ,csa_tree_add_110_49_pad_groupi_n_1241);
  or csa_tree_add_110_49_pad_groupi_g4509(csa_tree_add_110_49_pad_groupi_n_1303 ,csa_tree_add_110_49_pad_groupi_n_1145 ,csa_tree_add_110_49_pad_groupi_n_1256);
  or csa_tree_add_110_49_pad_groupi_g4510(csa_tree_add_110_49_pad_groupi_n_1302 ,csa_tree_add_110_49_pad_groupi_n_1120 ,csa_tree_add_110_49_pad_groupi_n_1251);
  or csa_tree_add_110_49_pad_groupi_g4511(csa_tree_add_110_49_pad_groupi_n_1301 ,csa_tree_add_110_49_pad_groupi_n_1150 ,csa_tree_add_110_49_pad_groupi_n_1252);
  and csa_tree_add_110_49_pad_groupi_g4512(csa_tree_add_110_49_pad_groupi_n_1300 ,csa_tree_add_110_49_pad_groupi_n_1204 ,csa_tree_add_110_49_pad_groupi_n_1257);
  or csa_tree_add_110_49_pad_groupi_g4513(csa_tree_add_110_49_pad_groupi_n_1299 ,csa_tree_add_110_49_pad_groupi_n_1202 ,csa_tree_add_110_49_pad_groupi_n_1245);
  or csa_tree_add_110_49_pad_groupi_g4514(csa_tree_add_110_49_pad_groupi_n_1296 ,csa_tree_add_110_49_pad_groupi_n_1176 ,csa_tree_add_110_49_pad_groupi_n_1259);
  not csa_tree_add_110_49_pad_groupi_g4515(csa_tree_add_110_49_pad_groupi_n_1284 ,csa_tree_add_110_49_pad_groupi_n_1283);
  not csa_tree_add_110_49_pad_groupi_g4516(csa_tree_add_110_49_pad_groupi_n_1281 ,csa_tree_add_110_49_pad_groupi_n_1282);
  not csa_tree_add_110_49_pad_groupi_g4517(csa_tree_add_110_49_pad_groupi_n_1279 ,csa_tree_add_110_49_pad_groupi_n_1278);
  not csa_tree_add_110_49_pad_groupi_g4518(csa_tree_add_110_49_pad_groupi_n_1277 ,csa_tree_add_110_49_pad_groupi_n_1276);
  not csa_tree_add_110_49_pad_groupi_g4520(csa_tree_add_110_49_pad_groupi_n_1274 ,csa_tree_add_110_49_pad_groupi_n_1273);
  and csa_tree_add_110_49_pad_groupi_g4521(csa_tree_add_110_49_pad_groupi_n_1272 ,csa_tree_add_110_49_pad_groupi_n_1186 ,csa_tree_add_110_49_pad_groupi_n_1226);
  or csa_tree_add_110_49_pad_groupi_g4522(csa_tree_add_110_49_pad_groupi_n_1271 ,csa_tree_add_110_49_pad_groupi_n_1187 ,csa_tree_add_110_49_pad_groupi_n_1232);
  nor csa_tree_add_110_49_pad_groupi_g4523(csa_tree_add_110_49_pad_groupi_n_1270 ,csa_tree_add_110_49_pad_groupi_n_1188 ,csa_tree_add_110_49_pad_groupi_n_1231);
  xnor csa_tree_add_110_49_pad_groupi_g4524(csa_tree_add_110_49_pad_groupi_n_1269 ,csa_tree_add_110_49_pad_groupi_n_1159 ,csa_tree_add_110_49_pad_groupi_n_1192);
  xnor csa_tree_add_110_49_pad_groupi_g4525(csa_tree_add_110_49_pad_groupi_n_1268 ,csa_tree_add_110_49_pad_groupi_n_630 ,csa_tree_add_110_49_pad_groupi_n_1190);
  xnor csa_tree_add_110_49_pad_groupi_g4526(csa_tree_add_110_49_pad_groupi_n_1267 ,csa_tree_add_110_49_pad_groupi_n_621 ,csa_tree_add_110_49_pad_groupi_n_1195);
  xnor csa_tree_add_110_49_pad_groupi_g4527(csa_tree_add_110_49_pad_groupi_n_1266 ,csa_tree_add_110_49_pad_groupi_n_1181 ,n_156);
  xnor csa_tree_add_110_49_pad_groupi_g4528(csa_tree_add_110_49_pad_groupi_n_1265 ,csa_tree_add_110_49_pad_groupi_n_1128 ,csa_tree_add_110_49_pad_groupi_n_1183);
  xnor csa_tree_add_110_49_pad_groupi_g4529(csa_tree_add_110_49_pad_groupi_n_1285 ,csa_tree_add_110_49_pad_groupi_n_1135 ,csa_tree_add_110_49_pad_groupi_n_1174);
  xnor csa_tree_add_110_49_pad_groupi_g4530(csa_tree_add_110_49_pad_groupi_n_1283 ,csa_tree_add_110_49_pad_groupi_n_1126 ,csa_tree_add_110_49_pad_groupi_n_1170);
  xnor csa_tree_add_110_49_pad_groupi_g4531(csa_tree_add_110_49_pad_groupi_n_1282 ,csa_tree_add_110_49_pad_groupi_n_1173 ,n_153);
  xnor csa_tree_add_110_49_pad_groupi_g4532(csa_tree_add_110_49_pad_groupi_n_1280 ,csa_tree_add_110_49_pad_groupi_n_1161 ,csa_tree_add_110_49_pad_groupi_n_1175);
  xnor csa_tree_add_110_49_pad_groupi_g4533(csa_tree_add_110_49_pad_groupi_n_1278 ,csa_tree_add_110_49_pad_groupi_n_1216 ,csa_tree_add_110_49_pad_groupi_n_1171);
  xnor csa_tree_add_110_49_pad_groupi_g4534(csa_tree_add_110_49_pad_groupi_n_1276 ,csa_tree_add_110_49_pad_groupi_n_1194 ,csa_tree_add_110_49_pad_groupi_n_1169);
  xnor csa_tree_add_110_49_pad_groupi_g4535(csa_tree_add_110_49_pad_groupi_n_1275 ,csa_tree_add_110_49_pad_groupi_n_1193 ,csa_tree_add_110_49_pad_groupi_n_1172);
  xnor csa_tree_add_110_49_pad_groupi_g4536(csa_tree_add_110_49_pad_groupi_n_1273 ,csa_tree_add_110_49_pad_groupi_n_1168 ,n_187);
  not csa_tree_add_110_49_pad_groupi_g4537(csa_tree_add_110_49_pad_groupi_n_1264 ,csa_tree_add_110_49_pad_groupi_n_1263);
  not csa_tree_add_110_49_pad_groupi_g4538(csa_tree_add_110_49_pad_groupi_n_1261 ,csa_tree_add_110_49_pad_groupi_n_1260);
  and csa_tree_add_110_49_pad_groupi_g4539(csa_tree_add_110_49_pad_groupi_n_1259 ,csa_tree_add_110_49_pad_groupi_n_1109 ,csa_tree_add_110_49_pad_groupi_n_1177);
  or csa_tree_add_110_49_pad_groupi_g4540(csa_tree_add_110_49_pad_groupi_n_1258 ,csa_tree_add_110_49_pad_groupi_n_1127 ,csa_tree_add_110_49_pad_groupi_n_1183);
  or csa_tree_add_110_49_pad_groupi_g4541(csa_tree_add_110_49_pad_groupi_n_1257 ,csa_tree_add_110_49_pad_groupi_n_1214 ,csa_tree_add_110_49_pad_groupi_n_1195);
  and csa_tree_add_110_49_pad_groupi_g4542(csa_tree_add_110_49_pad_groupi_n_1256 ,csa_tree_add_110_49_pad_groupi_n_1144 ,csa_tree_add_110_49_pad_groupi_n_1194);
  or csa_tree_add_110_49_pad_groupi_g4543(csa_tree_add_110_49_pad_groupi_n_1255 ,csa_tree_add_110_49_pad_groupi_n_629 ,csa_tree_add_110_49_pad_groupi_n_1189);
  nor csa_tree_add_110_49_pad_groupi_g4544(csa_tree_add_110_49_pad_groupi_n_1254 ,csa_tree_add_110_49_pad_groupi_n_630 ,csa_tree_add_110_49_pad_groupi_n_1190);
  nor csa_tree_add_110_49_pad_groupi_g4545(csa_tree_add_110_49_pad_groupi_n_1253 ,csa_tree_add_110_49_pad_groupi_n_1027 ,csa_tree_add_110_49_pad_groupi_n_1199);
  and csa_tree_add_110_49_pad_groupi_g4546(csa_tree_add_110_49_pad_groupi_n_1252 ,csa_tree_add_110_49_pad_groupi_n_1140 ,csa_tree_add_110_49_pad_groupi_n_1193);
  nor csa_tree_add_110_49_pad_groupi_g4547(csa_tree_add_110_49_pad_groupi_n_1251 ,csa_tree_add_110_49_pad_groupi_n_1216 ,csa_tree_add_110_49_pad_groupi_n_1121);
  nor csa_tree_add_110_49_pad_groupi_g4548(csa_tree_add_110_49_pad_groupi_n_1250 ,csa_tree_add_110_49_pad_groupi_n_1128 ,csa_tree_add_110_49_pad_groupi_n_1182);
  or csa_tree_add_110_49_pad_groupi_g4549(csa_tree_add_110_49_pad_groupi_n_1249 ,csa_tree_add_110_49_pad_groupi_n_1159 ,csa_tree_add_110_49_pad_groupi_n_1191);
  nor csa_tree_add_110_49_pad_groupi_g4550(csa_tree_add_110_49_pad_groupi_n_1248 ,csa_tree_add_110_49_pad_groupi_n_1158 ,csa_tree_add_110_49_pad_groupi_n_1192);
  nor csa_tree_add_110_49_pad_groupi_g4551(csa_tree_add_110_49_pad_groupi_n_1247 ,csa_tree_add_110_49_pad_groupi_n_310 ,csa_tree_add_110_49_pad_groupi_n_1181);
  or csa_tree_add_110_49_pad_groupi_g4552(csa_tree_add_110_49_pad_groupi_n_1246 ,n_156 ,csa_tree_add_110_49_pad_groupi_n_1180);
  and csa_tree_add_110_49_pad_groupi_g4553(csa_tree_add_110_49_pad_groupi_n_1245 ,csa_tree_add_110_49_pad_groupi_n_1201 ,csa_tree_add_110_49_pad_groupi_n_1196);
  nor csa_tree_add_110_49_pad_groupi_g4554(csa_tree_add_110_49_pad_groupi_n_1244 ,csa_tree_add_110_49_pad_groupi_n_316 ,csa_tree_add_110_49_pad_groupi_n_1203);
  or csa_tree_add_110_49_pad_groupi_g4555(csa_tree_add_110_49_pad_groupi_n_1263 ,csa_tree_add_110_49_pad_groupi_n_1086 ,csa_tree_add_110_49_pad_groupi_n_1209);
  and csa_tree_add_110_49_pad_groupi_g4556(csa_tree_add_110_49_pad_groupi_n_1262 ,csa_tree_add_110_49_pad_groupi_n_1095 ,csa_tree_add_110_49_pad_groupi_n_1198);
  or csa_tree_add_110_49_pad_groupi_g4557(csa_tree_add_110_49_pad_groupi_n_1260 ,csa_tree_add_110_49_pad_groupi_n_1091 ,csa_tree_add_110_49_pad_groupi_n_1211);
  not csa_tree_add_110_49_pad_groupi_g4558(csa_tree_add_110_49_pad_groupi_n_1239 ,csa_tree_add_110_49_pad_groupi_n_1238);
  not csa_tree_add_110_49_pad_groupi_g4559(csa_tree_add_110_49_pad_groupi_n_1236 ,csa_tree_add_110_49_pad_groupi_n_1235);
  not csa_tree_add_110_49_pad_groupi_g4560(csa_tree_add_110_49_pad_groupi_n_1234 ,csa_tree_add_110_49_pad_groupi_n_1233);
  not csa_tree_add_110_49_pad_groupi_g4561(csa_tree_add_110_49_pad_groupi_n_1232 ,csa_tree_add_110_49_pad_groupi_n_1231);
  not csa_tree_add_110_49_pad_groupi_g4562(csa_tree_add_110_49_pad_groupi_n_1230 ,csa_tree_add_110_49_pad_groupi_n_1229);
  not csa_tree_add_110_49_pad_groupi_g4563(csa_tree_add_110_49_pad_groupi_n_1227 ,csa_tree_add_110_49_pad_groupi_n_1228);
  xnor csa_tree_add_110_49_pad_groupi_g4564(csa_tree_add_110_49_pad_groupi_n_1224 ,csa_tree_add_110_49_pad_groupi_n_581 ,csa_tree_add_110_49_pad_groupi_n_1162);
  xnor csa_tree_add_110_49_pad_groupi_g4565(csa_tree_add_110_49_pad_groupi_n_1223 ,csa_tree_add_110_49_pad_groupi_n_1157 ,csa_tree_add_110_49_pad_groupi_n_1132);
  xnor csa_tree_add_110_49_pad_groupi_g4566(csa_tree_add_110_49_pad_groupi_n_1222 ,csa_tree_add_110_49_pad_groupi_n_1138 ,csa_tree_add_110_49_pad_groupi_n_1110);
  xnor csa_tree_add_110_49_pad_groupi_g4567(csa_tree_add_110_49_pad_groupi_n_1221 ,csa_tree_add_110_49_pad_groupi_n_1130 ,csa_tree_add_110_49_pad_groupi_n_1133);
  xnor csa_tree_add_110_49_pad_groupi_g4568(csa_tree_add_110_49_pad_groupi_n_1220 ,csa_tree_add_110_49_pad_groupi_n_623 ,csa_tree_add_110_49_pad_groupi_n_1152);
  xnor csa_tree_add_110_49_pad_groupi_g4569(csa_tree_add_110_49_pad_groupi_n_1219 ,csa_tree_add_110_49_pad_groupi_n_1129 ,csa_tree_add_110_49_pad_groupi_n_1153);
  or csa_tree_add_110_49_pad_groupi_g4570(csa_tree_add_110_49_pad_groupi_n_1243 ,csa_tree_add_110_49_pad_groupi_n_1063 ,csa_tree_add_110_49_pad_groupi_n_1178);
  xnor csa_tree_add_110_49_pad_groupi_g4571(csa_tree_add_110_49_pad_groupi_n_1242 ,csa_tree_add_110_49_pad_groupi_n_1134 ,csa_tree_add_110_49_pad_groupi_n_369);
  and csa_tree_add_110_49_pad_groupi_g4572(csa_tree_add_110_49_pad_groupi_n_1241 ,csa_tree_add_110_49_pad_groupi_n_1090 ,csa_tree_add_110_49_pad_groupi_n_1197);
  or csa_tree_add_110_49_pad_groupi_g4573(csa_tree_add_110_49_pad_groupi_n_1240 ,csa_tree_add_110_49_pad_groupi_n_1148 ,csa_tree_add_110_49_pad_groupi_n_1200);
  xnor csa_tree_add_110_49_pad_groupi_g4574(csa_tree_add_110_49_pad_groupi_n_1238 ,csa_tree_add_110_49_pad_groupi_n_1166 ,csa_tree_add_110_49_pad_groupi_n_1113);
  xnor csa_tree_add_110_49_pad_groupi_g4575(csa_tree_add_110_49_pad_groupi_n_1237 ,csa_tree_add_110_49_pad_groupi_n_1160 ,csa_tree_add_110_49_pad_groupi_n_1111);
  xnor csa_tree_add_110_49_pad_groupi_g4576(csa_tree_add_110_49_pad_groupi_n_1235 ,csa_tree_add_110_49_pad_groupi_n_1112 ,n_157);
  xnor csa_tree_add_110_49_pad_groupi_g4577(csa_tree_add_110_49_pad_groupi_n_1233 ,csa_tree_add_110_49_pad_groupi_n_1115 ,n_218);
  and csa_tree_add_110_49_pad_groupi_g4578(csa_tree_add_110_49_pad_groupi_n_1231 ,csa_tree_add_110_49_pad_groupi_n_1149 ,csa_tree_add_110_49_pad_groupi_n_1179);
  xnor csa_tree_add_110_49_pad_groupi_g4579(csa_tree_add_110_49_pad_groupi_n_1229 ,csa_tree_add_110_49_pad_groupi_n_1164 ,csa_tree_add_110_49_pad_groupi_n_1117);
  xnor csa_tree_add_110_49_pad_groupi_g4580(csa_tree_add_110_49_pad_groupi_n_1228 ,csa_tree_add_110_49_pad_groupi_n_1076 ,csa_tree_add_110_49_pad_groupi_n_1118);
  xnor csa_tree_add_110_49_pad_groupi_g4581(csa_tree_add_110_49_pad_groupi_n_1226 ,csa_tree_add_110_49_pad_groupi_n_1167 ,csa_tree_add_110_49_pad_groupi_n_1116);
  xnor csa_tree_add_110_49_pad_groupi_g4582(csa_tree_add_110_49_pad_groupi_n_1225 ,csa_tree_add_110_49_pad_groupi_n_583 ,csa_tree_add_110_49_pad_groupi_n_1114);
  and csa_tree_add_110_49_pad_groupi_g4583(csa_tree_add_110_49_pad_groupi_n_1215 ,csa_tree_add_110_49_pad_groupi_n_1153 ,csa_tree_add_110_49_pad_groupi_n_1129);
  nor csa_tree_add_110_49_pad_groupi_g4584(csa_tree_add_110_49_pad_groupi_n_1214 ,csa_tree_add_110_49_pad_groupi_n_621 ,csa_tree_add_110_49_pad_groupi_n_1154);
  nor csa_tree_add_110_49_pad_groupi_g4585(csa_tree_add_110_49_pad_groupi_n_1213 ,csa_tree_add_110_49_pad_groupi_n_1080 ,csa_tree_add_110_49_pad_groupi_n_1137);
  nor csa_tree_add_110_49_pad_groupi_g4586(csa_tree_add_110_49_pad_groupi_n_1212 ,csa_tree_add_110_49_pad_groupi_n_1156 ,csa_tree_add_110_49_pad_groupi_n_1132);
  nor csa_tree_add_110_49_pad_groupi_g4587(csa_tree_add_110_49_pad_groupi_n_1211 ,csa_tree_add_110_49_pad_groupi_n_1089 ,csa_tree_add_110_49_pad_groupi_n_1167);
  or csa_tree_add_110_49_pad_groupi_g4588(csa_tree_add_110_49_pad_groupi_n_1210 ,csa_tree_add_110_49_pad_groupi_n_1157 ,csa_tree_add_110_49_pad_groupi_n_1131);
  and csa_tree_add_110_49_pad_groupi_g4589(csa_tree_add_110_49_pad_groupi_n_1209 ,csa_tree_add_110_49_pad_groupi_n_1085 ,csa_tree_add_110_49_pad_groupi_n_1160);
  or csa_tree_add_110_49_pad_groupi_g4590(csa_tree_add_110_49_pad_groupi_n_1208 ,csa_tree_add_110_49_pad_groupi_n_1081 ,csa_tree_add_110_49_pad_groupi_n_1136);
  or csa_tree_add_110_49_pad_groupi_g4591(csa_tree_add_110_49_pad_groupi_n_1207 ,csa_tree_add_110_49_pad_groupi_n_1153 ,csa_tree_add_110_49_pad_groupi_n_1129);
  nor csa_tree_add_110_49_pad_groupi_g4592(csa_tree_add_110_49_pad_groupi_n_1206 ,csa_tree_add_110_49_pad_groupi_n_1133 ,csa_tree_add_110_49_pad_groupi_n_1130);
  and csa_tree_add_110_49_pad_groupi_g4593(csa_tree_add_110_49_pad_groupi_n_1205 ,csa_tree_add_110_49_pad_groupi_n_1133 ,csa_tree_add_110_49_pad_groupi_n_1130);
  or csa_tree_add_110_49_pad_groupi_g4594(csa_tree_add_110_49_pad_groupi_n_1204 ,csa_tree_add_110_49_pad_groupi_n_620 ,csa_tree_add_110_49_pad_groupi_n_1155);
  nor csa_tree_add_110_49_pad_groupi_g4595(csa_tree_add_110_49_pad_groupi_n_1203 ,csa_tree_add_110_49_pad_groupi_n_358 ,csa_tree_add_110_49_pad_groupi_n_1134);
  nor csa_tree_add_110_49_pad_groupi_g4596(csa_tree_add_110_49_pad_groupi_n_1202 ,csa_tree_add_110_49_pad_groupi_n_622 ,csa_tree_add_110_49_pad_groupi_n_1152);
  or csa_tree_add_110_49_pad_groupi_g4597(csa_tree_add_110_49_pad_groupi_n_1201 ,csa_tree_add_110_49_pad_groupi_n_623 ,csa_tree_add_110_49_pad_groupi_n_1151);
  and csa_tree_add_110_49_pad_groupi_g4598(csa_tree_add_110_49_pad_groupi_n_1200 ,csa_tree_add_110_49_pad_groupi_n_1135 ,csa_tree_add_110_49_pad_groupi_n_1124);
  nor csa_tree_add_110_49_pad_groupi_g4599(csa_tree_add_110_49_pad_groupi_n_1199 ,csa_tree_add_110_49_pad_groupi_n_1031 ,csa_tree_add_110_49_pad_groupi_n_1143);
  or csa_tree_add_110_49_pad_groupi_g4600(csa_tree_add_110_49_pad_groupi_n_1198 ,csa_tree_add_110_49_pad_groupi_n_1094 ,csa_tree_add_110_49_pad_groupi_n_1163);
  or csa_tree_add_110_49_pad_groupi_g4601(csa_tree_add_110_49_pad_groupi_n_1197 ,csa_tree_add_110_49_pad_groupi_n_1088 ,csa_tree_add_110_49_pad_groupi_n_1165);
  or csa_tree_add_110_49_pad_groupi_g4602(csa_tree_add_110_49_pad_groupi_n_1218 ,csa_tree_add_110_49_pad_groupi_n_1066 ,csa_tree_add_110_49_pad_groupi_n_1119);
  or csa_tree_add_110_49_pad_groupi_g4603(csa_tree_add_110_49_pad_groupi_n_1217 ,csa_tree_add_110_49_pad_groupi_n_836 ,csa_tree_add_110_49_pad_groupi_n_1142);
  and csa_tree_add_110_49_pad_groupi_g4604(csa_tree_add_110_49_pad_groupi_n_1216 ,csa_tree_add_110_49_pad_groupi_n_325 ,csa_tree_add_110_49_pad_groupi_n_1141);
  not csa_tree_add_110_49_pad_groupi_g4605(csa_tree_add_110_49_pad_groupi_n_1191 ,csa_tree_add_110_49_pad_groupi_n_1192);
  not csa_tree_add_110_49_pad_groupi_g4606(csa_tree_add_110_49_pad_groupi_n_1190 ,csa_tree_add_110_49_pad_groupi_n_1189);
  not csa_tree_add_110_49_pad_groupi_g4607(csa_tree_add_110_49_pad_groupi_n_1188 ,csa_tree_add_110_49_pad_groupi_n_1187);
  not csa_tree_add_110_49_pad_groupi_g4608(csa_tree_add_110_49_pad_groupi_n_1186 ,csa_tree_add_110_49_pad_groupi_n_1185);
  not csa_tree_add_110_49_pad_groupi_g4610(csa_tree_add_110_49_pad_groupi_n_1182 ,csa_tree_add_110_49_pad_groupi_n_1183);
  not csa_tree_add_110_49_pad_groupi_g4611(csa_tree_add_110_49_pad_groupi_n_1181 ,csa_tree_add_110_49_pad_groupi_n_1180);
  or csa_tree_add_110_49_pad_groupi_g4612(csa_tree_add_110_49_pad_groupi_n_1179 ,csa_tree_add_110_49_pad_groupi_n_1161 ,csa_tree_add_110_49_pad_groupi_n_1147);
  nor csa_tree_add_110_49_pad_groupi_g4613(csa_tree_add_110_49_pad_groupi_n_1178 ,csa_tree_add_110_49_pad_groupi_n_1166 ,csa_tree_add_110_49_pad_groupi_n_1064);
  or csa_tree_add_110_49_pad_groupi_g4614(csa_tree_add_110_49_pad_groupi_n_1177 ,csa_tree_add_110_49_pad_groupi_n_1006 ,csa_tree_add_110_49_pad_groupi_n_1125);
  nor csa_tree_add_110_49_pad_groupi_g4615(csa_tree_add_110_49_pad_groupi_n_1176 ,csa_tree_add_110_49_pad_groupi_n_1007 ,csa_tree_add_110_49_pad_groupi_n_1126);
  xnor csa_tree_add_110_49_pad_groupi_g4616(csa_tree_add_110_49_pad_groupi_n_1175 ,csa_tree_add_110_49_pad_groupi_n_632 ,csa_tree_add_110_49_pad_groupi_n_1073);
  xnor csa_tree_add_110_49_pad_groupi_g4617(csa_tree_add_110_49_pad_groupi_n_1174 ,csa_tree_add_110_49_pad_groupi_n_1105 ,csa_tree_add_110_49_pad_groupi_n_1075);
  xnor csa_tree_add_110_49_pad_groupi_g4618(csa_tree_add_110_49_pad_groupi_n_1173 ,csa_tree_add_110_49_pad_groupi_n_1107 ,n_185);
  xnor csa_tree_add_110_49_pad_groupi_g4619(csa_tree_add_110_49_pad_groupi_n_1172 ,csa_tree_add_110_49_pad_groupi_n_1103 ,csa_tree_add_110_49_pad_groupi_n_1012);
  xnor csa_tree_add_110_49_pad_groupi_g4620(csa_tree_add_110_49_pad_groupi_n_1171 ,csa_tree_add_110_49_pad_groupi_n_1069 ,csa_tree_add_110_49_pad_groupi_n_1070);
  xnor csa_tree_add_110_49_pad_groupi_g4621(csa_tree_add_110_49_pad_groupi_n_1170 ,csa_tree_add_110_49_pad_groupi_n_1109 ,csa_tree_add_110_49_pad_groupi_n_1007);
  xnor csa_tree_add_110_49_pad_groupi_g4622(csa_tree_add_110_49_pad_groupi_n_1169 ,csa_tree_add_110_49_pad_groupi_n_1106 ,csa_tree_add_110_49_pad_groupi_n_1008);
  xnor csa_tree_add_110_49_pad_groupi_g4623(csa_tree_add_110_49_pad_groupi_n_1168 ,csa_tree_add_110_49_pad_groupi_n_1108 ,csa_tree_add_110_49_pad_groupi_n_743);
  xnor csa_tree_add_110_49_pad_groupi_g4624(csa_tree_add_110_49_pad_groupi_n_1196 ,csa_tree_add_110_49_pad_groupi_n_934 ,csa_tree_add_110_49_pad_groupi_n_1061);
  xnor csa_tree_add_110_49_pad_groupi_g4625(csa_tree_add_110_49_pad_groupi_n_1195 ,csa_tree_add_110_49_pad_groupi_n_932 ,csa_tree_add_110_49_pad_groupi_n_1052);
  xnor csa_tree_add_110_49_pad_groupi_g4626(csa_tree_add_110_49_pad_groupi_n_1194 ,csa_tree_add_110_49_pad_groupi_n_1051 ,n_182);
  xnor csa_tree_add_110_49_pad_groupi_g4627(csa_tree_add_110_49_pad_groupi_n_1193 ,csa_tree_add_110_49_pad_groupi_n_1060 ,n_181);
  xnor csa_tree_add_110_49_pad_groupi_g4628(csa_tree_add_110_49_pad_groupi_n_1192 ,csa_tree_add_110_49_pad_groupi_n_1050 ,n_247);
  xnor csa_tree_add_110_49_pad_groupi_g4629(csa_tree_add_110_49_pad_groupi_n_1189 ,csa_tree_add_110_49_pad_groupi_n_943 ,csa_tree_add_110_49_pad_groupi_n_1054);
  xnor csa_tree_add_110_49_pad_groupi_g4630(csa_tree_add_110_49_pad_groupi_n_1187 ,csa_tree_add_110_49_pad_groupi_n_1022 ,csa_tree_add_110_49_pad_groupi_n_1056);
  xnor csa_tree_add_110_49_pad_groupi_g4631(csa_tree_add_110_49_pad_groupi_n_1185 ,csa_tree_add_110_49_pad_groupi_n_989 ,csa_tree_add_110_49_pad_groupi_n_1059);
  xnor csa_tree_add_110_49_pad_groupi_g4632(csa_tree_add_110_49_pad_groupi_n_1184 ,csa_tree_add_110_49_pad_groupi_n_1057 ,n_217);
  xnor csa_tree_add_110_49_pad_groupi_g4633(csa_tree_add_110_49_pad_groupi_n_1183 ,csa_tree_add_110_49_pad_groupi_n_1053 ,n_212);
  xnor csa_tree_add_110_49_pad_groupi_g4634(csa_tree_add_110_49_pad_groupi_n_1180 ,csa_tree_add_110_49_pad_groupi_n_1023 ,csa_tree_add_110_49_pad_groupi_n_1058);
  not csa_tree_add_110_49_pad_groupi_g4635(csa_tree_add_110_49_pad_groupi_n_1165 ,csa_tree_add_110_49_pad_groupi_n_1164);
  not csa_tree_add_110_49_pad_groupi_g4636(csa_tree_add_110_49_pad_groupi_n_1163 ,csa_tree_add_110_49_pad_groupi_n_1162);
  not csa_tree_add_110_49_pad_groupi_g4637(csa_tree_add_110_49_pad_groupi_n_1159 ,csa_tree_add_110_49_pad_groupi_n_1158);
  not csa_tree_add_110_49_pad_groupi_g4638(csa_tree_add_110_49_pad_groupi_n_1156 ,csa_tree_add_110_49_pad_groupi_n_1157);
  not csa_tree_add_110_49_pad_groupi_g4639(csa_tree_add_110_49_pad_groupi_n_1154 ,csa_tree_add_110_49_pad_groupi_n_1155);
  not csa_tree_add_110_49_pad_groupi_g4640(csa_tree_add_110_49_pad_groupi_n_1152 ,csa_tree_add_110_49_pad_groupi_n_1151);
  nor csa_tree_add_110_49_pad_groupi_g4641(csa_tree_add_110_49_pad_groupi_n_1150 ,csa_tree_add_110_49_pad_groupi_n_1102 ,csa_tree_add_110_49_pad_groupi_n_1012);
  or csa_tree_add_110_49_pad_groupi_g4642(csa_tree_add_110_49_pad_groupi_n_1149 ,csa_tree_add_110_49_pad_groupi_n_631 ,csa_tree_add_110_49_pad_groupi_n_1073);
  nor csa_tree_add_110_49_pad_groupi_g4643(csa_tree_add_110_49_pad_groupi_n_1148 ,csa_tree_add_110_49_pad_groupi_n_1104 ,csa_tree_add_110_49_pad_groupi_n_1075);
  nor csa_tree_add_110_49_pad_groupi_g4644(csa_tree_add_110_49_pad_groupi_n_1147 ,csa_tree_add_110_49_pad_groupi_n_632 ,csa_tree_add_110_49_pad_groupi_n_1072);
  and csa_tree_add_110_49_pad_groupi_g4645(csa_tree_add_110_49_pad_groupi_n_1146 ,csa_tree_add_110_49_pad_groupi_n_950 ,csa_tree_add_110_49_pad_groupi_n_1079);
  and csa_tree_add_110_49_pad_groupi_g4646(csa_tree_add_110_49_pad_groupi_n_1145 ,csa_tree_add_110_49_pad_groupi_n_1106 ,csa_tree_add_110_49_pad_groupi_n_1008);
  or csa_tree_add_110_49_pad_groupi_g4647(csa_tree_add_110_49_pad_groupi_n_1144 ,csa_tree_add_110_49_pad_groupi_n_1106 ,csa_tree_add_110_49_pad_groupi_n_1008);
  nor csa_tree_add_110_49_pad_groupi_g4648(csa_tree_add_110_49_pad_groupi_n_1143 ,csa_tree_add_110_49_pad_groupi_n_1030 ,csa_tree_add_110_49_pad_groupi_n_1082);
  and csa_tree_add_110_49_pad_groupi_g4649(csa_tree_add_110_49_pad_groupi_n_1142 ,csa_tree_add_110_49_pad_groupi_n_862 ,csa_tree_add_110_49_pad_groupi_n_1108);
  or csa_tree_add_110_49_pad_groupi_g4650(csa_tree_add_110_49_pad_groupi_n_1141 ,csa_tree_add_110_49_pad_groupi_n_335 ,csa_tree_add_110_49_pad_groupi_n_1107);
  or csa_tree_add_110_49_pad_groupi_g4651(csa_tree_add_110_49_pad_groupi_n_1140 ,csa_tree_add_110_49_pad_groupi_n_1103 ,csa_tree_add_110_49_pad_groupi_n_1011);
  nor csa_tree_add_110_49_pad_groupi_g4652(csa_tree_add_110_49_pad_groupi_n_1139 ,csa_tree_add_110_49_pad_groupi_n_950 ,csa_tree_add_110_49_pad_groupi_n_1079);
  nor csa_tree_add_110_49_pad_groupi_g4653(csa_tree_add_110_49_pad_groupi_n_1138 ,csa_tree_add_110_49_pad_groupi_n_345 ,csa_tree_add_110_49_pad_groupi_n_1098);
  and csa_tree_add_110_49_pad_groupi_g4654(csa_tree_add_110_49_pad_groupi_n_1167 ,csa_tree_add_110_49_pad_groupi_n_999 ,csa_tree_add_110_49_pad_groupi_n_1101);
  and csa_tree_add_110_49_pad_groupi_g4655(csa_tree_add_110_49_pad_groupi_n_1166 ,csa_tree_add_110_49_pad_groupi_n_323 ,csa_tree_add_110_49_pad_groupi_n_1087);
  or csa_tree_add_110_49_pad_groupi_g4656(csa_tree_add_110_49_pad_groupi_n_1164 ,csa_tree_add_110_49_pad_groupi_n_1035 ,csa_tree_add_110_49_pad_groupi_n_1096);
  or csa_tree_add_110_49_pad_groupi_g4657(csa_tree_add_110_49_pad_groupi_n_1162 ,csa_tree_add_110_49_pad_groupi_n_1043 ,csa_tree_add_110_49_pad_groupi_n_1093);
  and csa_tree_add_110_49_pad_groupi_g4658(csa_tree_add_110_49_pad_groupi_n_1161 ,csa_tree_add_110_49_pad_groupi_n_1039 ,csa_tree_add_110_49_pad_groupi_n_1097);
  or csa_tree_add_110_49_pad_groupi_g4659(csa_tree_add_110_49_pad_groupi_n_1160 ,csa_tree_add_110_49_pad_groupi_n_977 ,csa_tree_add_110_49_pad_groupi_n_1084);
  or csa_tree_add_110_49_pad_groupi_g4660(csa_tree_add_110_49_pad_groupi_n_1158 ,csa_tree_add_110_49_pad_groupi_n_341 ,csa_tree_add_110_49_pad_groupi_n_1099);
  or csa_tree_add_110_49_pad_groupi_g4661(csa_tree_add_110_49_pad_groupi_n_1157 ,csa_tree_add_110_49_pad_groupi_n_330 ,csa_tree_add_110_49_pad_groupi_n_1092);
  and csa_tree_add_110_49_pad_groupi_g4662(csa_tree_add_110_49_pad_groupi_n_1155 ,csa_tree_add_110_49_pad_groupi_n_1041 ,csa_tree_add_110_49_pad_groupi_n_1100);
  and csa_tree_add_110_49_pad_groupi_g4663(csa_tree_add_110_49_pad_groupi_n_1153 ,csa_tree_add_110_49_pad_groupi_n_324 ,csa_tree_add_110_49_pad_groupi_n_1083);
  or csa_tree_add_110_49_pad_groupi_g4664(csa_tree_add_110_49_pad_groupi_n_1151 ,csa_tree_add_110_49_pad_groupi_n_1002 ,csa_tree_add_110_49_pad_groupi_n_1068);
  not csa_tree_add_110_49_pad_groupi_g4665(csa_tree_add_110_49_pad_groupi_n_1137 ,csa_tree_add_110_49_pad_groupi_n_1136);
  not csa_tree_add_110_49_pad_groupi_g4666(csa_tree_add_110_49_pad_groupi_n_1131 ,csa_tree_add_110_49_pad_groupi_n_1132);
  not csa_tree_add_110_49_pad_groupi_g4667(csa_tree_add_110_49_pad_groupi_n_1127 ,csa_tree_add_110_49_pad_groupi_n_1128);
  not csa_tree_add_110_49_pad_groupi_g4668(csa_tree_add_110_49_pad_groupi_n_1126 ,csa_tree_add_110_49_pad_groupi_n_1125);
  or csa_tree_add_110_49_pad_groupi_g4669(csa_tree_add_110_49_pad_groupi_n_1124 ,csa_tree_add_110_49_pad_groupi_n_1105 ,csa_tree_add_110_49_pad_groupi_n_1074);
  nor csa_tree_add_110_49_pad_groupi_g4670(csa_tree_add_110_49_pad_groupi_n_1123 ,csa_tree_add_110_49_pad_groupi_n_972 ,csa_tree_add_110_49_pad_groupi_n_1078);
  nor csa_tree_add_110_49_pad_groupi_g4671(csa_tree_add_110_49_pad_groupi_n_1122 ,csa_tree_add_110_49_pad_groupi_n_973 ,csa_tree_add_110_49_pad_groupi_n_1077);
  and csa_tree_add_110_49_pad_groupi_g4672(csa_tree_add_110_49_pad_groupi_n_1121 ,csa_tree_add_110_49_pad_groupi_n_1069 ,csa_tree_add_110_49_pad_groupi_n_1071);
  nor csa_tree_add_110_49_pad_groupi_g4673(csa_tree_add_110_49_pad_groupi_n_1120 ,csa_tree_add_110_49_pad_groupi_n_1069 ,csa_tree_add_110_49_pad_groupi_n_1071);
  and csa_tree_add_110_49_pad_groupi_g4674(csa_tree_add_110_49_pad_groupi_n_1119 ,csa_tree_add_110_49_pad_groupi_n_1065 ,csa_tree_add_110_49_pad_groupi_n_1076);
  xnor csa_tree_add_110_49_pad_groupi_g4675(csa_tree_add_110_49_pad_groupi_n_1118 ,csa_tree_add_110_49_pad_groupi_n_519 ,csa_tree_add_110_49_pad_groupi_n_1010);
  xnor csa_tree_add_110_49_pad_groupi_g4676(csa_tree_add_110_49_pad_groupi_n_1117 ,csa_tree_add_110_49_pad_groupi_n_577 ,csa_tree_add_110_49_pad_groupi_n_1016);
  xnor csa_tree_add_110_49_pad_groupi_g4677(csa_tree_add_110_49_pad_groupi_n_1116 ,csa_tree_add_110_49_pad_groupi_n_626 ,csa_tree_add_110_49_pad_groupi_n_1019);
  xnor csa_tree_add_110_49_pad_groupi_g4678(csa_tree_add_110_49_pad_groupi_n_1115 ,csa_tree_add_110_49_pad_groupi_n_930 ,csa_tree_add_110_49_pad_groupi_n_1045);
  xnor csa_tree_add_110_49_pad_groupi_g4679(csa_tree_add_110_49_pad_groupi_n_1114 ,csa_tree_add_110_49_pad_groupi_n_962 ,csa_tree_add_110_49_pad_groupi_n_1047);
  xnor csa_tree_add_110_49_pad_groupi_g4680(csa_tree_add_110_49_pad_groupi_n_1113 ,csa_tree_add_110_49_pad_groupi_n_1044 ,csa_tree_add_110_49_pad_groupi_n_1017);
  xnor csa_tree_add_110_49_pad_groupi_g4681(csa_tree_add_110_49_pad_groupi_n_1112 ,csa_tree_add_110_49_pad_groupi_n_1020 ,n_253);
  xnor csa_tree_add_110_49_pad_groupi_g4682(csa_tree_add_110_49_pad_groupi_n_1111 ,csa_tree_add_110_49_pad_groupi_n_517 ,csa_tree_add_110_49_pad_groupi_n_1005);
  xnor csa_tree_add_110_49_pad_groupi_g4683(csa_tree_add_110_49_pad_groupi_n_1110 ,csa_tree_add_110_49_pad_groupi_n_377 ,csa_tree_add_110_49_pad_groupi_n_995);
  xnor csa_tree_add_110_49_pad_groupi_g4684(csa_tree_add_110_49_pad_groupi_n_1136 ,csa_tree_add_110_49_pad_groupi_n_954 ,csa_tree_add_110_49_pad_groupi_n_993);
  or csa_tree_add_110_49_pad_groupi_g4685(csa_tree_add_110_49_pad_groupi_n_1135 ,csa_tree_add_110_49_pad_groupi_n_333 ,csa_tree_add_110_49_pad_groupi_n_1067);
  and csa_tree_add_110_49_pad_groupi_g4686(csa_tree_add_110_49_pad_groupi_n_1134 ,csa_tree_add_110_49_pad_groupi_n_1026 ,csa_tree_add_110_49_pad_groupi_n_1062);
  xnor csa_tree_add_110_49_pad_groupi_g4687(csa_tree_add_110_49_pad_groupi_n_1133 ,csa_tree_add_110_49_pad_groupi_n_1021 ,csa_tree_add_110_49_pad_groupi_n_368);
  xnor csa_tree_add_110_49_pad_groupi_g4688(csa_tree_add_110_49_pad_groupi_n_1132 ,csa_tree_add_110_49_pad_groupi_n_1048 ,csa_tree_add_110_49_pad_groupi_n_366);
  xnor csa_tree_add_110_49_pad_groupi_g4689(csa_tree_add_110_49_pad_groupi_n_1130 ,csa_tree_add_110_49_pad_groupi_n_994 ,n_152);
  xnor csa_tree_add_110_49_pad_groupi_g4690(csa_tree_add_110_49_pad_groupi_n_1129 ,csa_tree_add_110_49_pad_groupi_n_1049 ,csa_tree_add_110_49_pad_groupi_n_370);
  xnor csa_tree_add_110_49_pad_groupi_g4691(csa_tree_add_110_49_pad_groupi_n_1128 ,csa_tree_add_110_49_pad_groupi_n_1046 ,csa_tree_add_110_49_pad_groupi_n_381);
  xnor csa_tree_add_110_49_pad_groupi_g4692(csa_tree_add_110_49_pad_groupi_n_1125 ,csa_tree_add_110_49_pad_groupi_n_1024 ,csa_tree_add_110_49_pad_groupi_n_378);
  not csa_tree_add_110_49_pad_groupi_g4693(csa_tree_add_110_49_pad_groupi_n_1104 ,csa_tree_add_110_49_pad_groupi_n_1105);
  not csa_tree_add_110_49_pad_groupi_g4694(csa_tree_add_110_49_pad_groupi_n_1102 ,csa_tree_add_110_49_pad_groupi_n_1103);
  or csa_tree_add_110_49_pad_groupi_g4695(csa_tree_add_110_49_pad_groupi_n_1101 ,csa_tree_add_110_49_pad_groupi_n_945 ,csa_tree_add_110_49_pad_groupi_n_1003);
  or csa_tree_add_110_49_pad_groupi_g4696(csa_tree_add_110_49_pad_groupi_n_1100 ,csa_tree_add_110_49_pad_groupi_n_1047 ,csa_tree_add_110_49_pad_groupi_n_1040);
  nor csa_tree_add_110_49_pad_groupi_g4697(csa_tree_add_110_49_pad_groupi_n_1099 ,csa_tree_add_110_49_pad_groupi_n_314 ,csa_tree_add_110_49_pad_groupi_n_1048);
  and csa_tree_add_110_49_pad_groupi_g4698(csa_tree_add_110_49_pad_groupi_n_1098 ,csa_tree_add_110_49_pad_groupi_n_320 ,csa_tree_add_110_49_pad_groupi_n_1020);
  or csa_tree_add_110_49_pad_groupi_g4699(csa_tree_add_110_49_pad_groupi_n_1097 ,csa_tree_add_110_49_pad_groupi_n_943 ,csa_tree_add_110_49_pad_groupi_n_1037);
  and csa_tree_add_110_49_pad_groupi_g4700(csa_tree_add_110_49_pad_groupi_n_1096 ,csa_tree_add_110_49_pad_groupi_n_934 ,csa_tree_add_110_49_pad_groupi_n_1028);
  or csa_tree_add_110_49_pad_groupi_g4701(csa_tree_add_110_49_pad_groupi_n_1095 ,csa_tree_add_110_49_pad_groupi_n_580 ,csa_tree_add_110_49_pad_groupi_n_1014);
  nor csa_tree_add_110_49_pad_groupi_g4702(csa_tree_add_110_49_pad_groupi_n_1094 ,csa_tree_add_110_49_pad_groupi_n_581 ,csa_tree_add_110_49_pad_groupi_n_1013);
  nor csa_tree_add_110_49_pad_groupi_g4703(csa_tree_add_110_49_pad_groupi_n_1093 ,csa_tree_add_110_49_pad_groupi_n_989 ,csa_tree_add_110_49_pad_groupi_n_1034);
  nor csa_tree_add_110_49_pad_groupi_g4704(csa_tree_add_110_49_pad_groupi_n_1092 ,csa_tree_add_110_49_pad_groupi_n_365 ,csa_tree_add_110_49_pad_groupi_n_1049);
  and csa_tree_add_110_49_pad_groupi_g4705(csa_tree_add_110_49_pad_groupi_n_1091 ,csa_tree_add_110_49_pad_groupi_n_626 ,csa_tree_add_110_49_pad_groupi_n_1019);
  or csa_tree_add_110_49_pad_groupi_g4706(csa_tree_add_110_49_pad_groupi_n_1090 ,csa_tree_add_110_49_pad_groupi_n_576 ,csa_tree_add_110_49_pad_groupi_n_1016);
  nor csa_tree_add_110_49_pad_groupi_g4707(csa_tree_add_110_49_pad_groupi_n_1089 ,csa_tree_add_110_49_pad_groupi_n_626 ,csa_tree_add_110_49_pad_groupi_n_1019);
  nor csa_tree_add_110_49_pad_groupi_g4708(csa_tree_add_110_49_pad_groupi_n_1088 ,csa_tree_add_110_49_pad_groupi_n_577 ,csa_tree_add_110_49_pad_groupi_n_1015);
  or csa_tree_add_110_49_pad_groupi_g4709(csa_tree_add_110_49_pad_groupi_n_1087 ,csa_tree_add_110_49_pad_groupi_n_326 ,csa_tree_add_110_49_pad_groupi_n_1021);
  nor csa_tree_add_110_49_pad_groupi_g4710(csa_tree_add_110_49_pad_groupi_n_1086 ,csa_tree_add_110_49_pad_groupi_n_516 ,csa_tree_add_110_49_pad_groupi_n_1005);
  or csa_tree_add_110_49_pad_groupi_g4711(csa_tree_add_110_49_pad_groupi_n_1085 ,csa_tree_add_110_49_pad_groupi_n_517 ,csa_tree_add_110_49_pad_groupi_n_1004);
  and csa_tree_add_110_49_pad_groupi_g4712(csa_tree_add_110_49_pad_groupi_n_1084 ,csa_tree_add_110_49_pad_groupi_n_988 ,csa_tree_add_110_49_pad_groupi_n_1045);
  or csa_tree_add_110_49_pad_groupi_g4713(csa_tree_add_110_49_pad_groupi_n_1083 ,csa_tree_add_110_49_pad_groupi_n_363 ,csa_tree_add_110_49_pad_groupi_n_1046);
  nor csa_tree_add_110_49_pad_groupi_g4714(csa_tree_add_110_49_pad_groupi_n_1082 ,csa_tree_add_110_49_pad_groupi_n_905 ,csa_tree_add_110_49_pad_groupi_n_1029);
  or csa_tree_add_110_49_pad_groupi_g4715(csa_tree_add_110_49_pad_groupi_n_1109 ,csa_tree_add_110_49_pad_groupi_n_353 ,csa_tree_add_110_49_pad_groupi_n_1042);
  or csa_tree_add_110_49_pad_groupi_g4716(csa_tree_add_110_49_pad_groupi_n_1108 ,csa_tree_add_110_49_pad_groupi_n_814 ,csa_tree_add_110_49_pad_groupi_n_1033);
  and csa_tree_add_110_49_pad_groupi_g4717(csa_tree_add_110_49_pad_groupi_n_1107 ,csa_tree_add_110_49_pad_groupi_n_857 ,csa_tree_add_110_49_pad_groupi_n_1038);
  or csa_tree_add_110_49_pad_groupi_g4718(csa_tree_add_110_49_pad_groupi_n_1106 ,csa_tree_add_110_49_pad_groupi_n_328 ,csa_tree_add_110_49_pad_groupi_n_1036);
  or csa_tree_add_110_49_pad_groupi_g4719(csa_tree_add_110_49_pad_groupi_n_1105 ,csa_tree_add_110_49_pad_groupi_n_346 ,csa_tree_add_110_49_pad_groupi_n_1000);
  or csa_tree_add_110_49_pad_groupi_g4720(csa_tree_add_110_49_pad_groupi_n_1103 ,csa_tree_add_110_49_pad_groupi_n_338 ,csa_tree_add_110_49_pad_groupi_n_1032);
  not csa_tree_add_110_49_pad_groupi_g4721(csa_tree_add_110_49_pad_groupi_n_1081 ,csa_tree_add_110_49_pad_groupi_n_1080);
  not csa_tree_add_110_49_pad_groupi_g4722(csa_tree_add_110_49_pad_groupi_n_1078 ,csa_tree_add_110_49_pad_groupi_n_1077);
  not csa_tree_add_110_49_pad_groupi_g4723(csa_tree_add_110_49_pad_groupi_n_1074 ,csa_tree_add_110_49_pad_groupi_n_1075);
  not csa_tree_add_110_49_pad_groupi_g4724(csa_tree_add_110_49_pad_groupi_n_1072 ,csa_tree_add_110_49_pad_groupi_n_1073);
  not csa_tree_add_110_49_pad_groupi_g4725(csa_tree_add_110_49_pad_groupi_n_1071 ,csa_tree_add_110_49_pad_groupi_n_1070);
  nor csa_tree_add_110_49_pad_groupi_g4726(csa_tree_add_110_49_pad_groupi_n_1068 ,csa_tree_add_110_49_pad_groupi_n_1001 ,csa_tree_add_110_49_pad_groupi_n_1022);
  and csa_tree_add_110_49_pad_groupi_g4727(csa_tree_add_110_49_pad_groupi_n_1067 ,csa_tree_add_110_49_pad_groupi_n_343 ,csa_tree_add_110_49_pad_groupi_n_1024);
  nor csa_tree_add_110_49_pad_groupi_g4728(csa_tree_add_110_49_pad_groupi_n_1066 ,csa_tree_add_110_49_pad_groupi_n_518 ,csa_tree_add_110_49_pad_groupi_n_1010);
  or csa_tree_add_110_49_pad_groupi_g4729(csa_tree_add_110_49_pad_groupi_n_1065 ,csa_tree_add_110_49_pad_groupi_n_519 ,csa_tree_add_110_49_pad_groupi_n_1009);
  and csa_tree_add_110_49_pad_groupi_g4730(csa_tree_add_110_49_pad_groupi_n_1064 ,csa_tree_add_110_49_pad_groupi_n_1044 ,csa_tree_add_110_49_pad_groupi_n_1018);
  nor csa_tree_add_110_49_pad_groupi_g4731(csa_tree_add_110_49_pad_groupi_n_1063 ,csa_tree_add_110_49_pad_groupi_n_1044 ,csa_tree_add_110_49_pad_groupi_n_1018);
  or csa_tree_add_110_49_pad_groupi_g4732(csa_tree_add_110_49_pad_groupi_n_1062 ,csa_tree_add_110_49_pad_groupi_n_1023 ,csa_tree_add_110_49_pad_groupi_n_1025);
  or csa_tree_add_110_49_pad_groupi_g4733(csa_tree_add_110_49_pad_groupi_n_1080 ,csa_tree_add_110_49_pad_groupi_n_917 ,csa_tree_add_110_49_pad_groupi_n_996);
  xnor csa_tree_add_110_49_pad_groupi_g4734(csa_tree_add_110_49_pad_groupi_n_1061 ,csa_tree_add_110_49_pad_groupi_n_958 ,n_179);
  xnor csa_tree_add_110_49_pad_groupi_g4735(csa_tree_add_110_49_pad_groupi_n_1060 ,csa_tree_add_110_49_pad_groupi_n_963 ,n_213);
  xnor csa_tree_add_110_49_pad_groupi_g4736(csa_tree_add_110_49_pad_groupi_n_1059 ,csa_tree_add_110_49_pad_groupi_n_957 ,n_143);
  xnor csa_tree_add_110_49_pad_groupi_g4737(csa_tree_add_110_49_pad_groupi_n_1058 ,csa_tree_add_110_49_pad_groupi_n_960 ,csa_tree_add_110_49_pad_groupi_n_146);
  xnor csa_tree_add_110_49_pad_groupi_g4738(csa_tree_add_110_49_pad_groupi_n_1057 ,csa_tree_add_110_49_pad_groupi_n_967 ,n_249);
  xnor csa_tree_add_110_49_pad_groupi_g4739(csa_tree_add_110_49_pad_groupi_n_1056 ,csa_tree_add_110_49_pad_groupi_n_578 ,csa_tree_add_110_49_pad_groupi_n_953);
  xnor csa_tree_add_110_49_pad_groupi_g4740(csa_tree_add_110_49_pad_groupi_n_1079 ,csa_tree_add_110_49_pad_groupi_n_703 ,csa_tree_add_110_49_pad_groupi_n_951);
  xnor csa_tree_add_110_49_pad_groupi_g4741(csa_tree_add_110_49_pad_groupi_n_1077 ,csa_tree_add_110_49_pad_groupi_n_991 ,csa_tree_add_110_49_pad_groupi_n_926);
  xnor csa_tree_add_110_49_pad_groupi_g4742(csa_tree_add_110_49_pad_groupi_n_1055 ,csa_tree_add_110_49_pad_groupi_n_0 ,csa_tree_add_110_49_pad_groupi_n_375);
  xnor csa_tree_add_110_49_pad_groupi_g4743(csa_tree_add_110_49_pad_groupi_n_1054 ,csa_tree_add_110_49_pad_groupi_n_956 ,n_176);
  xnor csa_tree_add_110_49_pad_groupi_g4744(csa_tree_add_110_49_pad_groupi_n_1053 ,csa_tree_add_110_49_pad_groupi_n_969 ,n_180);
  xnor csa_tree_add_110_49_pad_groupi_g4745(csa_tree_add_110_49_pad_groupi_n_1052 ,csa_tree_add_110_49_pad_groupi_n_965 ,n_242);
  xnor csa_tree_add_110_49_pad_groupi_g4746(csa_tree_add_110_49_pad_groupi_n_1051 ,csa_tree_add_110_49_pad_groupi_n_990 ,n_214);
  xnor csa_tree_add_110_49_pad_groupi_g4747(csa_tree_add_110_49_pad_groupi_n_1050 ,csa_tree_add_110_49_pad_groupi_n_964 ,n_215);
  or csa_tree_add_110_49_pad_groupi_g4748(csa_tree_add_110_49_pad_groupi_n_1076 ,csa_tree_add_110_49_pad_groupi_n_979 ,csa_tree_add_110_49_pad_groupi_n_998);
  xnor csa_tree_add_110_49_pad_groupi_g4749(csa_tree_add_110_49_pad_groupi_n_1075 ,csa_tree_add_110_49_pad_groupi_n_966 ,csa_tree_add_110_49_pad_groupi_n_892);
  xnor csa_tree_add_110_49_pad_groupi_g4750(csa_tree_add_110_49_pad_groupi_n_1073 ,csa_tree_add_110_49_pad_groupi_n_937 ,csa_tree_add_110_49_pad_groupi_n_952);
  xnor csa_tree_add_110_49_pad_groupi_g4751(csa_tree_add_110_49_pad_groupi_n_1070 ,csa_tree_add_110_49_pad_groupi_n_968 ,csa_tree_add_110_49_pad_groupi_n_876);
  and csa_tree_add_110_49_pad_groupi_g4752(csa_tree_add_110_49_pad_groupi_n_1069 ,csa_tree_add_110_49_pad_groupi_n_331 ,csa_tree_add_110_49_pad_groupi_n_997);
  nor csa_tree_add_110_49_pad_groupi_g4753(csa_tree_add_110_49_pad_groupi_n_1043 ,csa_tree_add_110_49_pad_groupi_n_298 ,csa_tree_add_110_49_pad_groupi_n_957);
  and csa_tree_add_110_49_pad_groupi_g4754(csa_tree_add_110_49_pad_groupi_n_1042 ,csa_tree_add_110_49_pad_groupi_n_352 ,csa_tree_add_110_49_pad_groupi_n_990);
  or csa_tree_add_110_49_pad_groupi_g4755(csa_tree_add_110_49_pad_groupi_n_1041 ,csa_tree_add_110_49_pad_groupi_n_582 ,csa_tree_add_110_49_pad_groupi_n_962);
  nor csa_tree_add_110_49_pad_groupi_g4756(csa_tree_add_110_49_pad_groupi_n_1040 ,csa_tree_add_110_49_pad_groupi_n_583 ,csa_tree_add_110_49_pad_groupi_n_961);
  or csa_tree_add_110_49_pad_groupi_g4757(csa_tree_add_110_49_pad_groupi_n_1039 ,csa_tree_add_110_49_pad_groupi_n_307 ,csa_tree_add_110_49_pad_groupi_n_955);
  or csa_tree_add_110_49_pad_groupi_g4758(csa_tree_add_110_49_pad_groupi_n_1038 ,csa_tree_add_110_49_pad_groupi_n_853 ,csa_tree_add_110_49_pad_groupi_n_966);
  nor csa_tree_add_110_49_pad_groupi_g4759(csa_tree_add_110_49_pad_groupi_n_1037 ,n_176 ,csa_tree_add_110_49_pad_groupi_n_956);
  and csa_tree_add_110_49_pad_groupi_g4760(csa_tree_add_110_49_pad_groupi_n_1036 ,csa_tree_add_110_49_pad_groupi_n_339 ,csa_tree_add_110_49_pad_groupi_n_963);
  and csa_tree_add_110_49_pad_groupi_g4761(csa_tree_add_110_49_pad_groupi_n_1035 ,n_179 ,csa_tree_add_110_49_pad_groupi_n_958);
  and csa_tree_add_110_49_pad_groupi_g4762(csa_tree_add_110_49_pad_groupi_n_1034 ,csa_tree_add_110_49_pad_groupi_n_298 ,csa_tree_add_110_49_pad_groupi_n_957);
  and csa_tree_add_110_49_pad_groupi_g4763(csa_tree_add_110_49_pad_groupi_n_1033 ,csa_tree_add_110_49_pad_groupi_n_842 ,csa_tree_add_110_49_pad_groupi_n_968);
  and csa_tree_add_110_49_pad_groupi_g4764(csa_tree_add_110_49_pad_groupi_n_1032 ,csa_tree_add_110_49_pad_groupi_n_357 ,csa_tree_add_110_49_pad_groupi_n_969);
  nor csa_tree_add_110_49_pad_groupi_g4765(csa_tree_add_110_49_pad_groupi_n_1031 ,csa_tree_add_110_49_pad_groupi_n_833 ,csa_tree_add_110_49_pad_groupi_n_971);
  nor csa_tree_add_110_49_pad_groupi_g4766(csa_tree_add_110_49_pad_groupi_n_1030 ,csa_tree_add_110_49_pad_groupi_n_739 ,csa_tree_add_110_49_pad_groupi_n_992);
  and csa_tree_add_110_49_pad_groupi_g4767(csa_tree_add_110_49_pad_groupi_n_1029 ,csa_tree_add_110_49_pad_groupi_n_739 ,csa_tree_add_110_49_pad_groupi_n_992);
  or csa_tree_add_110_49_pad_groupi_g4768(csa_tree_add_110_49_pad_groupi_n_1028 ,n_179 ,csa_tree_add_110_49_pad_groupi_n_958);
  nor csa_tree_add_110_49_pad_groupi_g4769(csa_tree_add_110_49_pad_groupi_n_1027 ,csa_tree_add_110_49_pad_groupi_n_834 ,csa_tree_add_110_49_pad_groupi_n_970);
  or csa_tree_add_110_49_pad_groupi_g4770(csa_tree_add_110_49_pad_groupi_n_1026 ,csa_tree_add_110_49_pad_groupi_n_139 ,csa_tree_add_110_49_pad_groupi_n_959);
  nor csa_tree_add_110_49_pad_groupi_g4771(csa_tree_add_110_49_pad_groupi_n_1025 ,csa_tree_add_110_49_pad_groupi_n_285 ,csa_tree_add_110_49_pad_groupi_n_960);
  and csa_tree_add_110_49_pad_groupi_g4772(csa_tree_add_110_49_pad_groupi_n_1049 ,csa_tree_add_110_49_pad_groupi_n_848 ,csa_tree_add_110_49_pad_groupi_n_982);
  and csa_tree_add_110_49_pad_groupi_g4773(csa_tree_add_110_49_pad_groupi_n_1048 ,csa_tree_add_110_49_pad_groupi_n_863 ,csa_tree_add_110_49_pad_groupi_n_985);
  and csa_tree_add_110_49_pad_groupi_g4774(csa_tree_add_110_49_pad_groupi_n_1047 ,csa_tree_add_110_49_pad_groupi_n_866 ,csa_tree_add_110_49_pad_groupi_n_986);
  and csa_tree_add_110_49_pad_groupi_g4775(csa_tree_add_110_49_pad_groupi_n_1046 ,csa_tree_add_110_49_pad_groupi_n_816 ,csa_tree_add_110_49_pad_groupi_n_976);
  or csa_tree_add_110_49_pad_groupi_g4776(csa_tree_add_110_49_pad_groupi_n_1045 ,csa_tree_add_110_49_pad_groupi_n_826 ,csa_tree_add_110_49_pad_groupi_n_980);
  and csa_tree_add_110_49_pad_groupi_g4777(csa_tree_add_110_49_pad_groupi_n_1044 ,csa_tree_add_110_49_pad_groupi_n_334 ,csa_tree_add_110_49_pad_groupi_n_983);
  not csa_tree_add_110_49_pad_groupi_g4778(csa_tree_add_110_49_pad_groupi_n_1018 ,csa_tree_add_110_49_pad_groupi_n_1017);
  not csa_tree_add_110_49_pad_groupi_g4779(csa_tree_add_110_49_pad_groupi_n_1015 ,csa_tree_add_110_49_pad_groupi_n_1016);
  not csa_tree_add_110_49_pad_groupi_g4780(csa_tree_add_110_49_pad_groupi_n_1013 ,csa_tree_add_110_49_pad_groupi_n_1014);
  not csa_tree_add_110_49_pad_groupi_g4781(csa_tree_add_110_49_pad_groupi_n_1011 ,csa_tree_add_110_49_pad_groupi_n_1012);
  not csa_tree_add_110_49_pad_groupi_g4782(csa_tree_add_110_49_pad_groupi_n_1009 ,csa_tree_add_110_49_pad_groupi_n_1010);
  not csa_tree_add_110_49_pad_groupi_g4783(csa_tree_add_110_49_pad_groupi_n_1007 ,csa_tree_add_110_49_pad_groupi_n_1006);
  not csa_tree_add_110_49_pad_groupi_g4784(csa_tree_add_110_49_pad_groupi_n_1005 ,csa_tree_add_110_49_pad_groupi_n_1004);
  and csa_tree_add_110_49_pad_groupi_g4785(csa_tree_add_110_49_pad_groupi_n_1003 ,csa_tree_add_110_49_pad_groupi_n_705 ,csa_tree_add_110_49_pad_groupi_n_954);
  nor csa_tree_add_110_49_pad_groupi_g4786(csa_tree_add_110_49_pad_groupi_n_1002 ,csa_tree_add_110_49_pad_groupi_n_579 ,csa_tree_add_110_49_pad_groupi_n_953);
  and csa_tree_add_110_49_pad_groupi_g4787(csa_tree_add_110_49_pad_groupi_n_1001 ,csa_tree_add_110_49_pad_groupi_n_579 ,csa_tree_add_110_49_pad_groupi_n_953);
  and csa_tree_add_110_49_pad_groupi_g4788(csa_tree_add_110_49_pad_groupi_n_1000 ,csa_tree_add_110_49_pad_groupi_n_318 ,csa_tree_add_110_49_pad_groupi_n_964);
  or csa_tree_add_110_49_pad_groupi_g4789(csa_tree_add_110_49_pad_groupi_n_999 ,csa_tree_add_110_49_pad_groupi_n_705 ,csa_tree_add_110_49_pad_groupi_n_954);
  and csa_tree_add_110_49_pad_groupi_g4790(csa_tree_add_110_49_pad_groupi_n_998 ,csa_tree_add_110_49_pad_groupi_n_987 ,csa_tree_add_110_49_pad_groupi_n_965);
  or csa_tree_add_110_49_pad_groupi_g4791(csa_tree_add_110_49_pad_groupi_n_997 ,csa_tree_add_110_49_pad_groupi_n_361 ,csa_tree_add_110_49_pad_groupi_n_967);
  nor csa_tree_add_110_49_pad_groupi_g4792(csa_tree_add_110_49_pad_groupi_n_996 ,csa_tree_add_110_49_pad_groupi_n_915 ,csa_tree_add_110_49_pad_groupi_n_991);
  or csa_tree_add_110_49_pad_groupi_g4793(csa_tree_add_110_49_pad_groupi_n_995 ,csa_tree_add_110_49_pad_groupi_n_815 ,csa_tree_add_110_49_pad_groupi_n_978);
  xnor csa_tree_add_110_49_pad_groupi_g4794(csa_tree_add_110_49_pad_groupi_n_994 ,csa_tree_add_110_49_pad_groupi_n_949 ,n_248);
  xnor csa_tree_add_110_49_pad_groupi_g4795(csa_tree_add_110_49_pad_groupi_n_993 ,csa_tree_add_110_49_pad_groupi_n_945 ,csa_tree_add_110_49_pad_groupi_n_705);
  or csa_tree_add_110_49_pad_groupi_g4796(csa_tree_add_110_49_pad_groupi_n_1024 ,csa_tree_add_110_49_pad_groupi_n_810 ,csa_tree_add_110_49_pad_groupi_n_974);
  and csa_tree_add_110_49_pad_groupi_g4797(csa_tree_add_110_49_pad_groupi_n_1023 ,csa_tree_add_110_49_pad_groupi_n_869 ,csa_tree_add_110_49_pad_groupi_n_984);
  and csa_tree_add_110_49_pad_groupi_g4798(csa_tree_add_110_49_pad_groupi_n_1022 ,csa_tree_add_110_49_pad_groupi_n_928 ,csa_tree_add_110_49_pad_groupi_n_975);
  and csa_tree_add_110_49_pad_groupi_g4799(csa_tree_add_110_49_pad_groupi_n_1021 ,csa_tree_add_110_49_pad_groupi_n_822 ,csa_tree_add_110_49_pad_groupi_n_981);
  xnor csa_tree_add_110_49_pad_groupi_g4800(csa_tree_add_110_49_pad_groupi_n_1020 ,csa_tree_add_110_49_pad_groupi_n_936 ,csa_tree_add_110_49_pad_groupi_n_880);
  xnor csa_tree_add_110_49_pad_groupi_g4801(csa_tree_add_110_49_pad_groupi_n_1019 ,csa_tree_add_110_49_pad_groupi_n_707 ,csa_tree_add_110_49_pad_groupi_n_927);
  xnor csa_tree_add_110_49_pad_groupi_g4802(csa_tree_add_110_49_pad_groupi_n_1017 ,csa_tree_add_110_49_pad_groupi_n_933 ,csa_tree_add_110_49_pad_groupi_n_872);
  xnor csa_tree_add_110_49_pad_groupi_g4803(csa_tree_add_110_49_pad_groupi_n_1016 ,csa_tree_add_110_49_pad_groupi_n_946 ,csa_tree_add_110_49_pad_groupi_n_883);
  xnor csa_tree_add_110_49_pad_groupi_g4804(csa_tree_add_110_49_pad_groupi_n_1014 ,csa_tree_add_110_49_pad_groupi_n_947 ,csa_tree_add_110_49_pad_groupi_n_885);
  xnor csa_tree_add_110_49_pad_groupi_g4805(csa_tree_add_110_49_pad_groupi_n_1012 ,csa_tree_add_110_49_pad_groupi_n_944 ,csa_tree_add_110_49_pad_groupi_n_884);
  xnor csa_tree_add_110_49_pad_groupi_g4806(csa_tree_add_110_49_pad_groupi_n_1010 ,csa_tree_add_110_49_pad_groupi_n_942 ,csa_tree_add_110_49_pad_groupi_n_881);
  xnor csa_tree_add_110_49_pad_groupi_g4807(csa_tree_add_110_49_pad_groupi_n_1008 ,csa_tree_add_110_49_pad_groupi_n_935 ,csa_tree_add_110_49_pad_groupi_n_886);
  xnor csa_tree_add_110_49_pad_groupi_g4808(csa_tree_add_110_49_pad_groupi_n_1006 ,csa_tree_add_110_49_pad_groupi_n_948 ,csa_tree_add_110_49_pad_groupi_n_893);
  xnor csa_tree_add_110_49_pad_groupi_g4809(csa_tree_add_110_49_pad_groupi_n_1004 ,csa_tree_add_110_49_pad_groupi_n_938 ,csa_tree_add_110_49_pad_groupi_n_894);
  or csa_tree_add_110_49_pad_groupi_g4810(csa_tree_add_110_49_pad_groupi_n_988 ,n_218 ,csa_tree_add_110_49_pad_groupi_n_930);
  or csa_tree_add_110_49_pad_groupi_g4811(csa_tree_add_110_49_pad_groupi_n_987 ,n_242 ,csa_tree_add_110_49_pad_groupi_n_931);
  or csa_tree_add_110_49_pad_groupi_g4812(csa_tree_add_110_49_pad_groupi_n_986 ,csa_tree_add_110_49_pad_groupi_n_865 ,csa_tree_add_110_49_pad_groupi_n_947);
  or csa_tree_add_110_49_pad_groupi_g4813(csa_tree_add_110_49_pad_groupi_n_985 ,csa_tree_add_110_49_pad_groupi_n_860 ,csa_tree_add_110_49_pad_groupi_n_944);
  or csa_tree_add_110_49_pad_groupi_g4814(csa_tree_add_110_49_pad_groupi_n_984 ,csa_tree_add_110_49_pad_groupi_n_820 ,csa_tree_add_110_49_pad_groupi_n_938);
  or csa_tree_add_110_49_pad_groupi_g4815(csa_tree_add_110_49_pad_groupi_n_983 ,csa_tree_add_110_49_pad_groupi_n_350 ,csa_tree_add_110_49_pad_groupi_n_949);
  or csa_tree_add_110_49_pad_groupi_g4816(csa_tree_add_110_49_pad_groupi_n_982 ,csa_tree_add_110_49_pad_groupi_n_846 ,csa_tree_add_110_49_pad_groupi_n_946);
  or csa_tree_add_110_49_pad_groupi_g4817(csa_tree_add_110_49_pad_groupi_n_981 ,csa_tree_add_110_49_pad_groupi_n_817 ,csa_tree_add_110_49_pad_groupi_n_948);
  and csa_tree_add_110_49_pad_groupi_g4818(csa_tree_add_110_49_pad_groupi_n_980 ,csa_tree_add_110_49_pad_groupi_n_838 ,csa_tree_add_110_49_pad_groupi_n_933);
  nor csa_tree_add_110_49_pad_groupi_g4819(csa_tree_add_110_49_pad_groupi_n_979 ,csa_tree_add_110_49_pad_groupi_n_306 ,csa_tree_add_110_49_pad_groupi_n_932);
  and csa_tree_add_110_49_pad_groupi_g4820(csa_tree_add_110_49_pad_groupi_n_978 ,csa_tree_add_110_49_pad_groupi_n_800 ,csa_tree_add_110_49_pad_groupi_n_936);
  and csa_tree_add_110_49_pad_groupi_g4821(csa_tree_add_110_49_pad_groupi_n_977 ,n_218 ,csa_tree_add_110_49_pad_groupi_n_930);
  or csa_tree_add_110_49_pad_groupi_g4822(csa_tree_add_110_49_pad_groupi_n_976 ,csa_tree_add_110_49_pad_groupi_n_829 ,csa_tree_add_110_49_pad_groupi_n_942);
  or csa_tree_add_110_49_pad_groupi_g4823(csa_tree_add_110_49_pad_groupi_n_975 ,csa_tree_add_110_49_pad_groupi_n_929 ,csa_tree_add_110_49_pad_groupi_n_937);
  and csa_tree_add_110_49_pad_groupi_g4824(csa_tree_add_110_49_pad_groupi_n_974 ,csa_tree_add_110_49_pad_groupi_n_807 ,csa_tree_add_110_49_pad_groupi_n_935);
  and csa_tree_add_110_49_pad_groupi_g4825(csa_tree_add_110_49_pad_groupi_n_992 ,csa_tree_add_110_49_pad_groupi_n_840 ,csa_tree_add_110_49_pad_groupi_n_939);
  and csa_tree_add_110_49_pad_groupi_g4826(csa_tree_add_110_49_pad_groupi_n_991 ,csa_tree_add_110_49_pad_groupi_n_841 ,csa_tree_add_110_49_pad_groupi_n_941);
  xnor csa_tree_add_110_49_pad_groupi_g4827(csa_tree_add_110_49_pad_groupi_n_990 ,csa_tree_add_110_49_pad_groupi_n_732 ,csa_tree_add_110_49_pad_groupi_n_875);
  and csa_tree_add_110_49_pad_groupi_g4828(csa_tree_add_110_49_pad_groupi_n_989 ,csa_tree_add_110_49_pad_groupi_n_852 ,csa_tree_add_110_49_pad_groupi_n_940);
  not csa_tree_add_110_49_pad_groupi_g4829(csa_tree_add_110_49_pad_groupi_n_973 ,csa_tree_add_110_49_pad_groupi_n_972);
  not csa_tree_add_110_49_pad_groupi_g4830(csa_tree_add_110_49_pad_groupi_n_971 ,csa_tree_add_110_49_pad_groupi_n_970);
  not csa_tree_add_110_49_pad_groupi_g4831(csa_tree_add_110_49_pad_groupi_n_961 ,csa_tree_add_110_49_pad_groupi_n_962);
  not csa_tree_add_110_49_pad_groupi_g4832(csa_tree_add_110_49_pad_groupi_n_959 ,csa_tree_add_110_49_pad_groupi_n_960);
  not csa_tree_add_110_49_pad_groupi_g4833(csa_tree_add_110_49_pad_groupi_n_955 ,csa_tree_add_110_49_pad_groupi_n_956);
  xnor csa_tree_add_110_49_pad_groupi_g4835(csa_tree_add_110_49_pad_groupi_n_952 ,csa_tree_add_110_49_pad_groupi_n_897 ,n_209);
  xnor csa_tree_add_110_49_pad_groupi_g4836(csa_tree_add_110_49_pad_groupi_n_972 ,csa_tree_add_110_49_pad_groupi_n_798 ,csa_tree_add_110_49_pad_groupi_n_877);
  xnor csa_tree_add_110_49_pad_groupi_g4837(csa_tree_add_110_49_pad_groupi_n_970 ,csa_tree_add_110_49_pad_groupi_n_702 ,csa_tree_add_110_49_pad_groupi_n_878);
  xnor csa_tree_add_110_49_pad_groupi_g4838(csa_tree_add_110_49_pad_groupi_n_951 ,csa_tree_add_110_49_pad_groupi_n_898 ,csa_tree_add_110_49_pad_groupi_n_764);
  xnor csa_tree_add_110_49_pad_groupi_g4839(csa_tree_add_110_49_pad_groupi_n_969 ,csa_tree_add_110_49_pad_groupi_n_797 ,csa_tree_add_110_49_pad_groupi_n_902);
  xnor csa_tree_add_110_49_pad_groupi_g4840(csa_tree_add_110_49_pad_groupi_n_968 ,csa_tree_add_110_49_pad_groupi_n_737 ,csa_tree_add_110_49_pad_groupi_n_889);
  xnor csa_tree_add_110_49_pad_groupi_g4841(csa_tree_add_110_49_pad_groupi_n_967 ,csa_tree_add_110_49_pad_groupi_n_734 ,csa_tree_add_110_49_pad_groupi_n_890);
  xnor csa_tree_add_110_49_pad_groupi_g4842(csa_tree_add_110_49_pad_groupi_n_966 ,csa_tree_add_110_49_pad_groupi_n_785 ,csa_tree_add_110_49_pad_groupi_n_888);
  xnor csa_tree_add_110_49_pad_groupi_g4843(csa_tree_add_110_49_pad_groupi_n_965 ,csa_tree_add_110_49_pad_groupi_n_793 ,csa_tree_add_110_49_pad_groupi_n_882);
  xnor csa_tree_add_110_49_pad_groupi_g4844(csa_tree_add_110_49_pad_groupi_n_964 ,csa_tree_add_110_49_pad_groupi_n_790 ,csa_tree_add_110_49_pad_groupi_n_901);
  xnor csa_tree_add_110_49_pad_groupi_g4845(csa_tree_add_110_49_pad_groupi_n_963 ,csa_tree_add_110_49_pad_groupi_n_735 ,csa_tree_add_110_49_pad_groupi_n_874);
  xnor csa_tree_add_110_49_pad_groupi_g4846(csa_tree_add_110_49_pad_groupi_n_962 ,csa_tree_add_110_49_pad_groupi_n_719 ,csa_tree_add_110_49_pad_groupi_n_887);
  xnor csa_tree_add_110_49_pad_groupi_g4847(csa_tree_add_110_49_pad_groupi_n_960 ,csa_tree_add_110_49_pad_groupi_n_787 ,csa_tree_add_110_49_pad_groupi_n_891);
  xnor csa_tree_add_110_49_pad_groupi_g4848(csa_tree_add_110_49_pad_groupi_n_958 ,csa_tree_add_110_49_pad_groupi_n_792 ,csa_tree_add_110_49_pad_groupi_n_903);
  xnor csa_tree_add_110_49_pad_groupi_g4849(csa_tree_add_110_49_pad_groupi_n_957 ,csa_tree_add_110_49_pad_groupi_n_768 ,csa_tree_add_110_49_pad_groupi_n_879);
  xnor csa_tree_add_110_49_pad_groupi_g4850(csa_tree_add_110_49_pad_groupi_n_956 ,csa_tree_add_110_49_pad_groupi_n_698 ,csa_tree_add_110_49_pad_groupi_n_900);
  xnor csa_tree_add_110_49_pad_groupi_g4851(csa_tree_add_110_49_pad_groupi_n_954 ,csa_tree_add_110_49_pad_groupi_n_899 ,csa_tree_add_110_49_pad_groupi_n_873);
  xnor csa_tree_add_110_49_pad_groupi_g4852(csa_tree_add_110_49_pad_groupi_n_953 ,csa_tree_add_110_49_pad_groupi_n_835 ,csa_tree_add_110_49_pad_groupi_n_895);
  or csa_tree_add_110_49_pad_groupi_g4853(csa_tree_add_110_49_pad_groupi_n_941 ,csa_tree_add_110_49_pad_groupi_n_839 ,csa_tree_add_110_49_pad_groupi_n_898);
  or csa_tree_add_110_49_pad_groupi_g4854(csa_tree_add_110_49_pad_groupi_n_940 ,csa_tree_add_110_49_pad_groupi_n_849 ,csa_tree_add_110_49_pad_groupi_n_899);
  or csa_tree_add_110_49_pad_groupi_g4855(csa_tree_add_110_49_pad_groupi_n_939 ,csa_tree_add_110_49_pad_groupi_n_914 ,csa_tree_add_110_49_pad_groupi_n_830);
  and csa_tree_add_110_49_pad_groupi_g4856(csa_tree_add_110_49_pad_groupi_n_950 ,csa_tree_add_110_49_pad_groupi_n_851 ,csa_tree_add_110_49_pad_groupi_n_918);
  and csa_tree_add_110_49_pad_groupi_g4857(csa_tree_add_110_49_pad_groupi_n_949 ,csa_tree_add_110_49_pad_groupi_n_847 ,csa_tree_add_110_49_pad_groupi_n_916);
  and csa_tree_add_110_49_pad_groupi_g4858(csa_tree_add_110_49_pad_groupi_n_948 ,csa_tree_add_110_49_pad_groupi_n_823 ,csa_tree_add_110_49_pad_groupi_n_909);
  and csa_tree_add_110_49_pad_groupi_g4859(csa_tree_add_110_49_pad_groupi_n_947 ,csa_tree_add_110_49_pad_groupi_n_858 ,csa_tree_add_110_49_pad_groupi_n_923);
  and csa_tree_add_110_49_pad_groupi_g4860(csa_tree_add_110_49_pad_groupi_n_946 ,csa_tree_add_110_49_pad_groupi_n_844 ,csa_tree_add_110_49_pad_groupi_n_920);
  and csa_tree_add_110_49_pad_groupi_g4861(csa_tree_add_110_49_pad_groupi_n_945 ,csa_tree_add_110_49_pad_groupi_n_827 ,csa_tree_add_110_49_pad_groupi_n_919);
  and csa_tree_add_110_49_pad_groupi_g4862(csa_tree_add_110_49_pad_groupi_n_944 ,csa_tree_add_110_49_pad_groupi_n_859 ,csa_tree_add_110_49_pad_groupi_n_922);
  and csa_tree_add_110_49_pad_groupi_g4863(csa_tree_add_110_49_pad_groupi_n_943 ,csa_tree_add_110_49_pad_groupi_n_856 ,csa_tree_add_110_49_pad_groupi_n_921);
  and csa_tree_add_110_49_pad_groupi_g4864(csa_tree_add_110_49_pad_groupi_n_942 ,csa_tree_add_110_49_pad_groupi_n_861 ,csa_tree_add_110_49_pad_groupi_n_912);
  not csa_tree_add_110_49_pad_groupi_g4865(csa_tree_add_110_49_pad_groupi_n_931 ,csa_tree_add_110_49_pad_groupi_n_932);
  nor csa_tree_add_110_49_pad_groupi_g4866(csa_tree_add_110_49_pad_groupi_n_929 ,n_209 ,csa_tree_add_110_49_pad_groupi_n_897);
  or csa_tree_add_110_49_pad_groupi_g4867(csa_tree_add_110_49_pad_groupi_n_928 ,csa_tree_add_110_49_pad_groupi_n_305 ,csa_tree_add_110_49_pad_groupi_n_896);
  xnor csa_tree_add_110_49_pad_groupi_g4868(csa_tree_add_110_49_pad_groupi_n_927 ,csa_tree_add_110_49_pad_groupi_n_784 ,csa_tree_add_110_49_pad_groupi_n_870);
  xnor csa_tree_add_110_49_pad_groupi_g4869(csa_tree_add_110_49_pad_groupi_n_926 ,csa_tree_add_110_49_pad_groupi_n_704 ,csa_tree_add_110_49_pad_groupi_n_831);
  and csa_tree_add_110_49_pad_groupi_g4870(csa_tree_add_110_49_pad_groupi_n_938 ,csa_tree_add_110_49_pad_groupi_n_811 ,csa_tree_add_110_49_pad_groupi_n_908);
  and csa_tree_add_110_49_pad_groupi_g4871(csa_tree_add_110_49_pad_groupi_n_937 ,csa_tree_add_110_49_pad_groupi_n_812 ,csa_tree_add_110_49_pad_groupi_n_910);
  or csa_tree_add_110_49_pad_groupi_g4872(csa_tree_add_110_49_pad_groupi_n_936 ,csa_tree_add_110_49_pad_groupi_n_867 ,csa_tree_add_110_49_pad_groupi_n_924);
  or csa_tree_add_110_49_pad_groupi_g4873(csa_tree_add_110_49_pad_groupi_n_935 ,csa_tree_add_110_49_pad_groupi_n_806 ,csa_tree_add_110_49_pad_groupi_n_906);
  or csa_tree_add_110_49_pad_groupi_g4874(csa_tree_add_110_49_pad_groupi_n_934 ,csa_tree_add_110_49_pad_groupi_n_825 ,csa_tree_add_110_49_pad_groupi_n_925);
  or csa_tree_add_110_49_pad_groupi_g4875(csa_tree_add_110_49_pad_groupi_n_933 ,csa_tree_add_110_49_pad_groupi_n_843 ,csa_tree_add_110_49_pad_groupi_n_913);
  and csa_tree_add_110_49_pad_groupi_g4876(csa_tree_add_110_49_pad_groupi_n_932 ,csa_tree_add_110_49_pad_groupi_n_804 ,csa_tree_add_110_49_pad_groupi_n_907);
  or csa_tree_add_110_49_pad_groupi_g4877(csa_tree_add_110_49_pad_groupi_n_930 ,csa_tree_add_110_49_pad_groupi_n_805 ,csa_tree_add_110_49_pad_groupi_n_911);
  nor csa_tree_add_110_49_pad_groupi_g4878(csa_tree_add_110_49_pad_groupi_n_925 ,csa_tree_add_110_49_pad_groupi_n_835 ,csa_tree_add_110_49_pad_groupi_n_854);
  and csa_tree_add_110_49_pad_groupi_g4879(csa_tree_add_110_49_pad_groupi_n_924 ,csa_tree_add_110_49_pad_groupi_n_787 ,csa_tree_add_110_49_pad_groupi_n_868);
  or csa_tree_add_110_49_pad_groupi_g4880(csa_tree_add_110_49_pad_groupi_n_923 ,csa_tree_add_110_49_pad_groupi_n_791 ,csa_tree_add_110_49_pad_groupi_n_864);
  or csa_tree_add_110_49_pad_groupi_g4881(csa_tree_add_110_49_pad_groupi_n_922 ,csa_tree_add_110_49_pad_groupi_n_797 ,csa_tree_add_110_49_pad_groupi_n_855);
  or csa_tree_add_110_49_pad_groupi_g4882(csa_tree_add_110_49_pad_groupi_n_921 ,csa_tree_add_110_49_pad_groupi_n_871 ,csa_tree_add_110_49_pad_groupi_n_819);
  or csa_tree_add_110_49_pad_groupi_g4883(csa_tree_add_110_49_pad_groupi_n_920 ,csa_tree_add_110_49_pad_groupi_n_792 ,csa_tree_add_110_49_pad_groupi_n_821);
  or csa_tree_add_110_49_pad_groupi_g4884(csa_tree_add_110_49_pad_groupi_n_919 ,csa_tree_add_110_49_pad_groupi_n_798 ,csa_tree_add_110_49_pad_groupi_n_850);
  or csa_tree_add_110_49_pad_groupi_g4885(csa_tree_add_110_49_pad_groupi_n_918 ,csa_tree_add_110_49_pad_groupi_n_845 ,csa_tree_add_110_49_pad_groupi_n_794);
  nor csa_tree_add_110_49_pad_groupi_g4886(csa_tree_add_110_49_pad_groupi_n_917 ,csa_tree_add_110_49_pad_groupi_n_704 ,csa_tree_add_110_49_pad_groupi_n_832);
  or csa_tree_add_110_49_pad_groupi_g4887(csa_tree_add_110_49_pad_groupi_n_916 ,csa_tree_add_110_49_pad_groupi_n_790 ,csa_tree_add_110_49_pad_groupi_n_837);
  and csa_tree_add_110_49_pad_groupi_g4888(csa_tree_add_110_49_pad_groupi_n_915 ,csa_tree_add_110_49_pad_groupi_n_704 ,csa_tree_add_110_49_pad_groupi_n_832);
  or csa_tree_add_110_49_pad_groupi_g4889(csa_tree_add_110_49_pad_groupi_n_914 ,csa_tree_add_110_49_pad_groupi_n_322 ,csa_tree_add_110_49_pad_groupi_n_818);
  nor csa_tree_add_110_49_pad_groupi_g4890(csa_tree_add_110_49_pad_groupi_n_913 ,csa_tree_add_110_49_pad_groupi_n_828 ,csa_tree_add_110_49_pad_groupi_n_785);
  or csa_tree_add_110_49_pad_groupi_g4891(csa_tree_add_110_49_pad_groupi_n_912 ,csa_tree_add_110_49_pad_groupi_n_793 ,csa_tree_add_110_49_pad_groupi_n_824);
  nor csa_tree_add_110_49_pad_groupi_g4892(csa_tree_add_110_49_pad_groupi_n_911 ,csa_tree_add_110_49_pad_groupi_n_813 ,csa_tree_add_110_49_pad_groupi_n_734);
  or csa_tree_add_110_49_pad_groupi_g4893(csa_tree_add_110_49_pad_groupi_n_910 ,csa_tree_add_110_49_pad_groupi_n_731 ,csa_tree_add_110_49_pad_groupi_n_809);
  or csa_tree_add_110_49_pad_groupi_g4894(csa_tree_add_110_49_pad_groupi_n_909 ,csa_tree_add_110_49_pad_groupi_n_733 ,csa_tree_add_110_49_pad_groupi_n_808);
  or csa_tree_add_110_49_pad_groupi_g4895(csa_tree_add_110_49_pad_groupi_n_908 ,csa_tree_add_110_49_pad_groupi_n_738 ,csa_tree_add_110_49_pad_groupi_n_803);
  or csa_tree_add_110_49_pad_groupi_g4896(csa_tree_add_110_49_pad_groupi_n_907 ,csa_tree_add_110_49_pad_groupi_n_736 ,csa_tree_add_110_49_pad_groupi_n_802);
  and csa_tree_add_110_49_pad_groupi_g4897(csa_tree_add_110_49_pad_groupi_n_906 ,csa_tree_add_110_49_pad_groupi_n_735 ,csa_tree_add_110_49_pad_groupi_n_801);
  xnor csa_tree_add_110_49_pad_groupi_g4898(csa_tree_add_110_49_pad_groupi_n_905 ,csa_tree_add_110_49_pad_groupi_n_639 ,csa_tree_add_110_49_pad_groupi_n_740);
  xnor csa_tree_add_110_49_pad_groupi_g4899(csa_tree_add_110_49_pad_groupi_n_904 ,csa_tree_add_110_49_pad_groupi_n_687 ,csa_tree_add_110_49_pad_groupi_n_688);
  xnor csa_tree_add_110_49_pad_groupi_g4900(csa_tree_add_110_49_pad_groupi_n_903 ,csa_tree_add_110_49_pad_groupi_n_766 ,csa_tree_add_110_49_pad_groupi_n_771);
  xnor csa_tree_add_110_49_pad_groupi_g4901(csa_tree_add_110_49_pad_groupi_n_902 ,csa_tree_add_110_49_pad_groupi_n_761 ,csa_tree_add_110_49_pad_groupi_n_755);
  xnor csa_tree_add_110_49_pad_groupi_g4902(csa_tree_add_110_49_pad_groupi_n_901 ,csa_tree_add_110_49_pad_groupi_n_773 ,csa_tree_add_110_49_pad_groupi_n_745);
  xnor csa_tree_add_110_49_pad_groupi_g4903(csa_tree_add_110_49_pad_groupi_n_900 ,csa_tree_add_110_49_pad_groupi_n_701 ,csa_tree_add_110_49_pad_groupi_n_731);
  not csa_tree_add_110_49_pad_groupi_g4904(csa_tree_add_110_49_pad_groupi_n_896 ,csa_tree_add_110_49_pad_groupi_n_897);
  xnor csa_tree_add_110_49_pad_groupi_g4905(csa_tree_add_110_49_pad_groupi_n_895 ,csa_tree_add_110_49_pad_groupi_n_753 ,csa_tree_add_110_49_pad_groupi_n_710);
  xnor csa_tree_add_110_49_pad_groupi_g4906(csa_tree_add_110_49_pad_groupi_n_894 ,csa_tree_add_110_49_pad_groupi_n_715 ,csa_tree_add_110_49_pad_groupi_n_712);
  xnor csa_tree_add_110_49_pad_groupi_g4907(csa_tree_add_110_49_pad_groupi_n_893 ,csa_tree_add_110_49_pad_groupi_n_727 ,csa_tree_add_110_49_pad_groupi_n_723);
  xnor csa_tree_add_110_49_pad_groupi_g4908(csa_tree_add_110_49_pad_groupi_n_892 ,csa_tree_add_110_49_pad_groupi_n_783 ,csa_tree_add_110_49_pad_groupi_n_756);
  xnor csa_tree_add_110_49_pad_groupi_g4909(csa_tree_add_110_49_pad_groupi_n_891 ,csa_tree_add_110_49_pad_groupi_n_748 ,csa_tree_add_110_49_pad_groupi_n_750);
  xnor csa_tree_add_110_49_pad_groupi_g4910(csa_tree_add_110_49_pad_groupi_n_890 ,csa_tree_add_110_49_pad_groupi_n_774 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g4911(csa_tree_add_110_49_pad_groupi_n_889 ,csa_tree_add_110_49_pad_groupi_n_728 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g4912(csa_tree_add_110_49_pad_groupi_n_888 ,csa_tree_add_110_49_pad_groupi_n_759 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g4913(csa_tree_add_110_49_pad_groupi_n_887 ,csa_tree_add_110_49_pad_groupi_n_736 ,csa_tree_add_110_49_pad_groupi_n_711);
  xnor csa_tree_add_110_49_pad_groupi_g4914(csa_tree_add_110_49_pad_groupi_n_886 ,csa_tree_add_110_49_pad_groupi_n_725 ,csa_tree_add_110_49_pad_groupi_n_696);
  xnor csa_tree_add_110_49_pad_groupi_g4915(csa_tree_add_110_49_pad_groupi_n_885 ,csa_tree_add_110_49_pad_groupi_n_770 ,csa_tree_add_110_49_pad_groupi_n_709);
  xnor csa_tree_add_110_49_pad_groupi_g4916(csa_tree_add_110_49_pad_groupi_n_884 ,csa_tree_add_110_49_pad_groupi_n_765 ,csa_tree_add_110_49_pad_groupi_n_708);
  xnor csa_tree_add_110_49_pad_groupi_g4917(csa_tree_add_110_49_pad_groupi_n_883 ,csa_tree_add_110_49_pad_groupi_n_775 ,csa_tree_add_110_49_pad_groupi_n_706);
  xnor csa_tree_add_110_49_pad_groupi_g4918(csa_tree_add_110_49_pad_groupi_n_882 ,csa_tree_add_110_49_pad_groupi_n_751 ,csa_tree_add_110_49_pad_groupi_n_746);
  xnor csa_tree_add_110_49_pad_groupi_g4919(csa_tree_add_110_49_pad_groupi_n_881 ,csa_tree_add_110_49_pad_groupi_n_780 ,csa_tree_add_110_49_pad_groupi_n_699);
  xnor csa_tree_add_110_49_pad_groupi_g4920(csa_tree_add_110_49_pad_groupi_n_880 ,csa_tree_add_110_49_pad_groupi_n_714 ,csa_tree_add_110_49_pad_groupi_n_692);
  xnor csa_tree_add_110_49_pad_groupi_g4921(csa_tree_add_110_49_pad_groupi_n_879 ,csa_tree_add_110_49_pad_groupi_n_515 ,csa_tree_add_110_49_pad_groupi_n_791);
  xnor csa_tree_add_110_49_pad_groupi_g4922(csa_tree_add_110_49_pad_groupi_n_878 ,csa_tree_add_110_49_pad_groupi_n_521 ,csa_tree_add_110_49_pad_groupi_n_794);
  xnor csa_tree_add_110_49_pad_groupi_g4923(csa_tree_add_110_49_pad_groupi_n_877 ,csa_tree_add_110_49_pad_groupi_n_520 ,csa_tree_add_110_49_pad_groupi_n_769);
  xnor csa_tree_add_110_49_pad_groupi_g4924(csa_tree_add_110_49_pad_groupi_n_876 ,csa_tree_add_110_49_pad_groupi_n_782 ,csa_tree_add_110_49_pad_groupi_n_777);
  xnor csa_tree_add_110_49_pad_groupi_g4925(csa_tree_add_110_49_pad_groupi_n_875 ,csa_tree_add_110_49_pad_groupi_n_718 ,csa_tree_add_110_49_pad_groupi_n_717);
  xnor csa_tree_add_110_49_pad_groupi_g4926(csa_tree_add_110_49_pad_groupi_n_874 ,csa_tree_add_110_49_pad_groupi_n_721 ,csa_tree_add_110_49_pad_groupi_n_763);
  xnor csa_tree_add_110_49_pad_groupi_g4927(csa_tree_add_110_49_pad_groupi_n_873 ,csa_tree_add_110_49_pad_groupi_n_778 ,csa_tree_add_110_49_pad_groupi_n_779);
  xnor csa_tree_add_110_49_pad_groupi_g4928(csa_tree_add_110_49_pad_groupi_n_872 ,csa_tree_add_110_49_pad_groupi_n_758 ,csa_tree_add_110_49_pad_groupi_n_694);
  xnor csa_tree_add_110_49_pad_groupi_g4929(csa_tree_add_110_49_pad_groupi_n_899 ,csa_tree_add_110_49_pad_groupi_n_795 ,csa_tree_add_110_49_pad_groupi_n_635);
  xnor csa_tree_add_110_49_pad_groupi_g4930(csa_tree_add_110_49_pad_groupi_n_898 ,csa_tree_add_110_49_pad_groupi_n_788 ,csa_tree_add_110_49_pad_groupi_n_637);
  xnor csa_tree_add_110_49_pad_groupi_g4931(csa_tree_add_110_49_pad_groupi_n_897 ,csa_tree_add_110_49_pad_groupi_n_729 ,csa_tree_add_110_49_pad_groupi_n_786);
  not csa_tree_add_110_49_pad_groupi_g4932(csa_tree_add_110_49_pad_groupi_n_871 ,csa_tree_add_110_49_pad_groupi_n_870);
  or csa_tree_add_110_49_pad_groupi_g4933(csa_tree_add_110_49_pad_groupi_n_869 ,csa_tree_add_110_49_pad_groupi_n_716 ,csa_tree_add_110_49_pad_groupi_n_712);
  or csa_tree_add_110_49_pad_groupi_g4934(csa_tree_add_110_49_pad_groupi_n_868 ,csa_tree_add_110_49_pad_groupi_n_749 ,csa_tree_add_110_49_pad_groupi_n_747);
  nor csa_tree_add_110_49_pad_groupi_g4935(csa_tree_add_110_49_pad_groupi_n_867 ,csa_tree_add_110_49_pad_groupi_n_750 ,csa_tree_add_110_49_pad_groupi_n_748);
  or csa_tree_add_110_49_pad_groupi_g4936(csa_tree_add_110_49_pad_groupi_n_866 ,csa_tree_add_110_49_pad_groupi_n_709 ,csa_tree_add_110_49_pad_groupi_n_770);
  and csa_tree_add_110_49_pad_groupi_g4937(csa_tree_add_110_49_pad_groupi_n_865 ,csa_tree_add_110_49_pad_groupi_n_709 ,csa_tree_add_110_49_pad_groupi_n_770);
  and csa_tree_add_110_49_pad_groupi_g4938(csa_tree_add_110_49_pad_groupi_n_864 ,csa_tree_add_110_49_pad_groupi_n_515 ,csa_tree_add_110_49_pad_groupi_n_768);
  or csa_tree_add_110_49_pad_groupi_g4939(csa_tree_add_110_49_pad_groupi_n_863 ,csa_tree_add_110_49_pad_groupi_n_708 ,csa_tree_add_110_49_pad_groupi_n_765);
  or csa_tree_add_110_49_pad_groupi_g4940(csa_tree_add_110_49_pad_groupi_n_862 ,n_187 ,csa_tree_add_110_49_pad_groupi_n_146);
  or csa_tree_add_110_49_pad_groupi_g4941(csa_tree_add_110_49_pad_groupi_n_861 ,csa_tree_add_110_49_pad_groupi_n_752 ,csa_tree_add_110_49_pad_groupi_n_746);
  and csa_tree_add_110_49_pad_groupi_g4942(csa_tree_add_110_49_pad_groupi_n_860 ,csa_tree_add_110_49_pad_groupi_n_708 ,csa_tree_add_110_49_pad_groupi_n_765);
  or csa_tree_add_110_49_pad_groupi_g4943(csa_tree_add_110_49_pad_groupi_n_859 ,csa_tree_add_110_49_pad_groupi_n_760 ,csa_tree_add_110_49_pad_groupi_n_755);
  or csa_tree_add_110_49_pad_groupi_g4944(csa_tree_add_110_49_pad_groupi_n_858 ,csa_tree_add_110_49_pad_groupi_n_515 ,csa_tree_add_110_49_pad_groupi_n_768);
  or csa_tree_add_110_49_pad_groupi_g4945(csa_tree_add_110_49_pad_groupi_n_857 ,csa_tree_add_110_49_pad_groupi_n_756 ,csa_tree_add_110_49_pad_groupi_n_783);
  or csa_tree_add_110_49_pad_groupi_g4946(csa_tree_add_110_49_pad_groupi_n_856 ,csa_tree_add_110_49_pad_groupi_n_707 ,csa_tree_add_110_49_pad_groupi_n_784);
  nor csa_tree_add_110_49_pad_groupi_g4947(csa_tree_add_110_49_pad_groupi_n_855 ,csa_tree_add_110_49_pad_groupi_n_761 ,csa_tree_add_110_49_pad_groupi_n_754);
  and csa_tree_add_110_49_pad_groupi_g4948(csa_tree_add_110_49_pad_groupi_n_854 ,csa_tree_add_110_49_pad_groupi_n_710 ,csa_tree_add_110_49_pad_groupi_n_753);
  and csa_tree_add_110_49_pad_groupi_g4949(csa_tree_add_110_49_pad_groupi_n_853 ,csa_tree_add_110_49_pad_groupi_n_756 ,csa_tree_add_110_49_pad_groupi_n_783);
  or csa_tree_add_110_49_pad_groupi_g4950(csa_tree_add_110_49_pad_groupi_n_852 ,csa_tree_add_110_49_pad_groupi_n_779 ,csa_tree_add_110_49_pad_groupi_n_778);
  or csa_tree_add_110_49_pad_groupi_g4951(csa_tree_add_110_49_pad_groupi_n_851 ,csa_tree_add_110_49_pad_groupi_n_521 ,csa_tree_add_110_49_pad_groupi_n_702);
  and csa_tree_add_110_49_pad_groupi_g4952(csa_tree_add_110_49_pad_groupi_n_850 ,csa_tree_add_110_49_pad_groupi_n_520 ,csa_tree_add_110_49_pad_groupi_n_769);
  and csa_tree_add_110_49_pad_groupi_g4953(csa_tree_add_110_49_pad_groupi_n_849 ,csa_tree_add_110_49_pad_groupi_n_779 ,csa_tree_add_110_49_pad_groupi_n_778);
  or csa_tree_add_110_49_pad_groupi_g4954(csa_tree_add_110_49_pad_groupi_n_848 ,csa_tree_add_110_49_pad_groupi_n_706 ,csa_tree_add_110_49_pad_groupi_n_775);
  or csa_tree_add_110_49_pad_groupi_g4955(csa_tree_add_110_49_pad_groupi_n_847 ,csa_tree_add_110_49_pad_groupi_n_772 ,csa_tree_add_110_49_pad_groupi_n_745);
  and csa_tree_add_110_49_pad_groupi_g4956(csa_tree_add_110_49_pad_groupi_n_846 ,csa_tree_add_110_49_pad_groupi_n_706 ,csa_tree_add_110_49_pad_groupi_n_775);
  and csa_tree_add_110_49_pad_groupi_g4957(csa_tree_add_110_49_pad_groupi_n_845 ,csa_tree_add_110_49_pad_groupi_n_521 ,csa_tree_add_110_49_pad_groupi_n_702);
  or csa_tree_add_110_49_pad_groupi_g4958(csa_tree_add_110_49_pad_groupi_n_844 ,csa_tree_add_110_49_pad_groupi_n_767 ,csa_tree_add_110_49_pad_groupi_n_771);
  and csa_tree_add_110_49_pad_groupi_g4959(csa_tree_add_110_49_pad_groupi_n_843 ,in16[1] ,csa_tree_add_110_49_pad_groupi_n_759);
  or csa_tree_add_110_49_pad_groupi_g4960(csa_tree_add_110_49_pad_groupi_n_842 ,csa_tree_add_110_49_pad_groupi_n_776 ,csa_tree_add_110_49_pad_groupi_n_781);
  or csa_tree_add_110_49_pad_groupi_g4961(csa_tree_add_110_49_pad_groupi_n_841 ,csa_tree_add_110_49_pad_groupi_n_703 ,csa_tree_add_110_49_pad_groupi_n_764);
  or csa_tree_add_110_49_pad_groupi_g4962(csa_tree_add_110_49_pad_groupi_n_840 ,csa_tree_add_110_49_pad_groupi_n_524 ,csa_tree_add_110_49_pad_groupi_n_742);
  and csa_tree_add_110_49_pad_groupi_g4963(csa_tree_add_110_49_pad_groupi_n_839 ,csa_tree_add_110_49_pad_groupi_n_703 ,csa_tree_add_110_49_pad_groupi_n_764);
  or csa_tree_add_110_49_pad_groupi_g4964(csa_tree_add_110_49_pad_groupi_n_838 ,csa_tree_add_110_49_pad_groupi_n_693 ,csa_tree_add_110_49_pad_groupi_n_757);
  nor csa_tree_add_110_49_pad_groupi_g4965(csa_tree_add_110_49_pad_groupi_n_837 ,csa_tree_add_110_49_pad_groupi_n_773 ,csa_tree_add_110_49_pad_groupi_n_744);
  and csa_tree_add_110_49_pad_groupi_g4966(csa_tree_add_110_49_pad_groupi_n_836 ,n_187 ,csa_tree_add_110_49_pad_groupi_n_139);
  and csa_tree_add_110_49_pad_groupi_g4967(csa_tree_add_110_49_pad_groupi_n_870 ,csa_tree_add_110_49_pad_groupi_n_636 ,csa_tree_add_110_49_pad_groupi_n_796);
  not csa_tree_add_110_49_pad_groupi_g4968(csa_tree_add_110_49_pad_groupi_n_834 ,csa_tree_add_110_49_pad_groupi_n_833);
  not csa_tree_add_110_49_pad_groupi_g4969(csa_tree_add_110_49_pad_groupi_n_832 ,csa_tree_add_110_49_pad_groupi_n_831);
  and csa_tree_add_110_49_pad_groupi_g4970(csa_tree_add_110_49_pad_groupi_n_830 ,csa_tree_add_110_49_pad_groupi_n_524 ,csa_tree_add_110_49_pad_groupi_n_742);
  and csa_tree_add_110_49_pad_groupi_g4971(csa_tree_add_110_49_pad_groupi_n_829 ,csa_tree_add_110_49_pad_groupi_n_699 ,csa_tree_add_110_49_pad_groupi_n_780);
  nor csa_tree_add_110_49_pad_groupi_g4972(csa_tree_add_110_49_pad_groupi_n_828 ,in16[1] ,csa_tree_add_110_49_pad_groupi_n_759);
  or csa_tree_add_110_49_pad_groupi_g4973(csa_tree_add_110_49_pad_groupi_n_827 ,csa_tree_add_110_49_pad_groupi_n_520 ,csa_tree_add_110_49_pad_groupi_n_769);
  nor csa_tree_add_110_49_pad_groupi_g4974(csa_tree_add_110_49_pad_groupi_n_826 ,csa_tree_add_110_49_pad_groupi_n_694 ,csa_tree_add_110_49_pad_groupi_n_758);
  nor csa_tree_add_110_49_pad_groupi_g4975(csa_tree_add_110_49_pad_groupi_n_825 ,csa_tree_add_110_49_pad_groupi_n_710 ,csa_tree_add_110_49_pad_groupi_n_753);
  and csa_tree_add_110_49_pad_groupi_g4976(csa_tree_add_110_49_pad_groupi_n_824 ,csa_tree_add_110_49_pad_groupi_n_752 ,csa_tree_add_110_49_pad_groupi_n_746);
  or csa_tree_add_110_49_pad_groupi_g4977(csa_tree_add_110_49_pad_groupi_n_823 ,csa_tree_add_110_49_pad_groupi_n_717 ,csa_tree_add_110_49_pad_groupi_n_718);
  or csa_tree_add_110_49_pad_groupi_g4978(csa_tree_add_110_49_pad_groupi_n_822 ,csa_tree_add_110_49_pad_groupi_n_726 ,csa_tree_add_110_49_pad_groupi_n_723);
  and csa_tree_add_110_49_pad_groupi_g4979(csa_tree_add_110_49_pad_groupi_n_821 ,csa_tree_add_110_49_pad_groupi_n_767 ,csa_tree_add_110_49_pad_groupi_n_771);
  and csa_tree_add_110_49_pad_groupi_g4980(csa_tree_add_110_49_pad_groupi_n_820 ,csa_tree_add_110_49_pad_groupi_n_716 ,csa_tree_add_110_49_pad_groupi_n_712);
  and csa_tree_add_110_49_pad_groupi_g4981(csa_tree_add_110_49_pad_groupi_n_819 ,csa_tree_add_110_49_pad_groupi_n_707 ,csa_tree_add_110_49_pad_groupi_n_784);
  or csa_tree_add_110_49_pad_groupi_g4982(csa_tree_add_110_49_pad_groupi_n_818 ,csa_tree_add_110_49_pad_groupi_n_194 ,csa_tree_add_110_49_pad_groupi_n_689);
  nor csa_tree_add_110_49_pad_groupi_g4983(csa_tree_add_110_49_pad_groupi_n_817 ,csa_tree_add_110_49_pad_groupi_n_727 ,csa_tree_add_110_49_pad_groupi_n_722);
  or csa_tree_add_110_49_pad_groupi_g4984(csa_tree_add_110_49_pad_groupi_n_816 ,csa_tree_add_110_49_pad_groupi_n_699 ,csa_tree_add_110_49_pad_groupi_n_780);
  nor csa_tree_add_110_49_pad_groupi_g4985(csa_tree_add_110_49_pad_groupi_n_815 ,csa_tree_add_110_49_pad_groupi_n_692 ,csa_tree_add_110_49_pad_groupi_n_714);
  nor csa_tree_add_110_49_pad_groupi_g4986(csa_tree_add_110_49_pad_groupi_n_814 ,csa_tree_add_110_49_pad_groupi_n_777 ,csa_tree_add_110_49_pad_groupi_n_782);
  nor csa_tree_add_110_49_pad_groupi_g4987(csa_tree_add_110_49_pad_groupi_n_813 ,in16[1] ,csa_tree_add_110_49_pad_groupi_n_774);
  or csa_tree_add_110_49_pad_groupi_g4988(csa_tree_add_110_49_pad_groupi_n_812 ,csa_tree_add_110_49_pad_groupi_n_700 ,csa_tree_add_110_49_pad_groupi_n_698);
  or csa_tree_add_110_49_pad_groupi_g4989(csa_tree_add_110_49_pad_groupi_n_811 ,in16[1] ,csa_tree_add_110_49_pad_groupi_n_728);
  nor csa_tree_add_110_49_pad_groupi_g4990(csa_tree_add_110_49_pad_groupi_n_810 ,csa_tree_add_110_49_pad_groupi_n_696 ,csa_tree_add_110_49_pad_groupi_n_725);
  nor csa_tree_add_110_49_pad_groupi_g4991(csa_tree_add_110_49_pad_groupi_n_809 ,csa_tree_add_110_49_pad_groupi_n_701 ,csa_tree_add_110_49_pad_groupi_n_697);
  and csa_tree_add_110_49_pad_groupi_g4992(csa_tree_add_110_49_pad_groupi_n_808 ,csa_tree_add_110_49_pad_groupi_n_717 ,csa_tree_add_110_49_pad_groupi_n_718);
  or csa_tree_add_110_49_pad_groupi_g4993(csa_tree_add_110_49_pad_groupi_n_807 ,csa_tree_add_110_49_pad_groupi_n_695 ,csa_tree_add_110_49_pad_groupi_n_724);
  nor csa_tree_add_110_49_pad_groupi_g4994(csa_tree_add_110_49_pad_groupi_n_806 ,csa_tree_add_110_49_pad_groupi_n_763 ,csa_tree_add_110_49_pad_groupi_n_721);
  and csa_tree_add_110_49_pad_groupi_g4995(csa_tree_add_110_49_pad_groupi_n_805 ,in16[1] ,csa_tree_add_110_49_pad_groupi_n_774);
  or csa_tree_add_110_49_pad_groupi_g4996(csa_tree_add_110_49_pad_groupi_n_804 ,csa_tree_add_110_49_pad_groupi_n_711 ,csa_tree_add_110_49_pad_groupi_n_719);
  and csa_tree_add_110_49_pad_groupi_g4997(csa_tree_add_110_49_pad_groupi_n_803 ,in16[1] ,csa_tree_add_110_49_pad_groupi_n_728);
  and csa_tree_add_110_49_pad_groupi_g4998(csa_tree_add_110_49_pad_groupi_n_802 ,csa_tree_add_110_49_pad_groupi_n_711 ,csa_tree_add_110_49_pad_groupi_n_719);
  or csa_tree_add_110_49_pad_groupi_g4999(csa_tree_add_110_49_pad_groupi_n_801 ,csa_tree_add_110_49_pad_groupi_n_762 ,csa_tree_add_110_49_pad_groupi_n_720);
  or csa_tree_add_110_49_pad_groupi_g5000(csa_tree_add_110_49_pad_groupi_n_800 ,csa_tree_add_110_49_pad_groupi_n_284 ,csa_tree_add_110_49_pad_groupi_n_713);
  xnor csa_tree_add_110_49_pad_groupi_g5001(csa_tree_add_110_49_pad_groupi_n_799 ,csa_tree_add_110_49_pad_groupi_n_573 ,csa_tree_add_110_49_pad_groupi_n_628);
  or csa_tree_add_110_49_pad_groupi_g5002(csa_tree_add_110_49_pad_groupi_n_835 ,csa_tree_add_110_49_pad_groupi_n_730 ,csa_tree_add_110_49_pad_groupi_n_786);
  and csa_tree_add_110_49_pad_groupi_g5003(csa_tree_add_110_49_pad_groupi_n_833 ,csa_tree_add_110_49_pad_groupi_n_640 ,csa_tree_add_110_49_pad_groupi_n_741);
  and csa_tree_add_110_49_pad_groupi_g5004(csa_tree_add_110_49_pad_groupi_n_831 ,csa_tree_add_110_49_pad_groupi_n_638 ,csa_tree_add_110_49_pad_groupi_n_789);
  not csa_tree_add_110_49_pad_groupi_g5005(csa_tree_add_110_49_pad_groupi_n_796 ,csa_tree_add_110_49_pad_groupi_n_795);
  not csa_tree_add_110_49_pad_groupi_g5006(csa_tree_add_110_49_pad_groupi_n_789 ,csa_tree_add_110_49_pad_groupi_n_788);
  not csa_tree_add_110_49_pad_groupi_g5007(csa_tree_add_110_49_pad_groupi_n_781 ,csa_tree_add_110_49_pad_groupi_n_782);
  not csa_tree_add_110_49_pad_groupi_g5008(csa_tree_add_110_49_pad_groupi_n_776 ,csa_tree_add_110_49_pad_groupi_n_777);
  not csa_tree_add_110_49_pad_groupi_g5009(csa_tree_add_110_49_pad_groupi_n_772 ,csa_tree_add_110_49_pad_groupi_n_773);
  not csa_tree_add_110_49_pad_groupi_g5010(csa_tree_add_110_49_pad_groupi_n_767 ,csa_tree_add_110_49_pad_groupi_n_766);
  not csa_tree_add_110_49_pad_groupi_g5011(csa_tree_add_110_49_pad_groupi_n_762 ,csa_tree_add_110_49_pad_groupi_n_763);
  not csa_tree_add_110_49_pad_groupi_g5012(csa_tree_add_110_49_pad_groupi_n_760 ,csa_tree_add_110_49_pad_groupi_n_761);
  not csa_tree_add_110_49_pad_groupi_g5013(csa_tree_add_110_49_pad_groupi_n_757 ,csa_tree_add_110_49_pad_groupi_n_758);
  not csa_tree_add_110_49_pad_groupi_g5014(csa_tree_add_110_49_pad_groupi_n_754 ,csa_tree_add_110_49_pad_groupi_n_755);
  not csa_tree_add_110_49_pad_groupi_g5015(csa_tree_add_110_49_pad_groupi_n_752 ,csa_tree_add_110_49_pad_groupi_n_751);
  not csa_tree_add_110_49_pad_groupi_g5016(csa_tree_add_110_49_pad_groupi_n_749 ,csa_tree_add_110_49_pad_groupi_n_750);
  not csa_tree_add_110_49_pad_groupi_g5017(csa_tree_add_110_49_pad_groupi_n_747 ,csa_tree_add_110_49_pad_groupi_n_748);
  not csa_tree_add_110_49_pad_groupi_g5018(csa_tree_add_110_49_pad_groupi_n_744 ,csa_tree_add_110_49_pad_groupi_n_745);
  and csa_tree_add_110_49_pad_groupi_g5020(csa_tree_add_110_49_pad_groupi_n_798 ,csa_tree_add_110_49_pad_groupi_n_504 ,csa_tree_add_110_49_pad_groupi_n_617);
  and csa_tree_add_110_49_pad_groupi_g5021(csa_tree_add_110_49_pad_groupi_n_797 ,csa_tree_add_110_49_pad_groupi_n_545 ,csa_tree_add_110_49_pad_groupi_n_647);
  and csa_tree_add_110_49_pad_groupi_g5022(csa_tree_add_110_49_pad_groupi_n_795 ,csa_tree_add_110_49_pad_groupi_n_531 ,csa_tree_add_110_49_pad_groupi_n_671);
  and csa_tree_add_110_49_pad_groupi_g5023(csa_tree_add_110_49_pad_groupi_n_794 ,csa_tree_add_110_49_pad_groupi_n_503 ,csa_tree_add_110_49_pad_groupi_n_615);
  and csa_tree_add_110_49_pad_groupi_g5024(csa_tree_add_110_49_pad_groupi_n_793 ,csa_tree_add_110_49_pad_groupi_n_536 ,csa_tree_add_110_49_pad_groupi_n_669);
  and csa_tree_add_110_49_pad_groupi_g5025(csa_tree_add_110_49_pad_groupi_n_792 ,csa_tree_add_110_49_pad_groupi_n_542 ,csa_tree_add_110_49_pad_groupi_n_641);
  and csa_tree_add_110_49_pad_groupi_g5026(csa_tree_add_110_49_pad_groupi_n_791 ,csa_tree_add_110_49_pad_groupi_n_550 ,csa_tree_add_110_49_pad_groupi_n_664);
  and csa_tree_add_110_49_pad_groupi_g5027(csa_tree_add_110_49_pad_groupi_n_790 ,csa_tree_add_110_49_pad_groupi_n_501 ,csa_tree_add_110_49_pad_groupi_n_611);
  and csa_tree_add_110_49_pad_groupi_g5028(csa_tree_add_110_49_pad_groupi_n_788 ,csa_tree_add_110_49_pad_groupi_n_554 ,csa_tree_add_110_49_pad_groupi_n_613);
  or csa_tree_add_110_49_pad_groupi_g5029(csa_tree_add_110_49_pad_groupi_n_787 ,csa_tree_add_110_49_pad_groupi_n_563 ,csa_tree_add_110_49_pad_groupi_n_683);
  and csa_tree_add_110_49_pad_groupi_g5030(csa_tree_add_110_49_pad_groupi_n_786 ,csa_tree_add_110_49_pad_groupi_n_497 ,csa_tree_add_110_49_pad_groupi_n_659);
  and csa_tree_add_110_49_pad_groupi_g5031(csa_tree_add_110_49_pad_groupi_n_785 ,csa_tree_add_110_49_pad_groupi_n_499 ,csa_tree_add_110_49_pad_groupi_n_661);
  and csa_tree_add_110_49_pad_groupi_g5032(csa_tree_add_110_49_pad_groupi_n_784 ,csa_tree_add_110_49_pad_groupi_n_533 ,csa_tree_add_110_49_pad_groupi_n_646);
  and csa_tree_add_110_49_pad_groupi_g5033(csa_tree_add_110_49_pad_groupi_n_783 ,csa_tree_add_110_49_pad_groupi_n_496 ,csa_tree_add_110_49_pad_groupi_n_645);
  and csa_tree_add_110_49_pad_groupi_g5034(csa_tree_add_110_49_pad_groupi_n_782 ,csa_tree_add_110_49_pad_groupi_n_553 ,csa_tree_add_110_49_pad_groupi_n_653);
  and csa_tree_add_110_49_pad_groupi_g5035(csa_tree_add_110_49_pad_groupi_n_780 ,csa_tree_add_110_49_pad_groupi_n_529 ,csa_tree_add_110_49_pad_groupi_n_665);
  and csa_tree_add_110_49_pad_groupi_g5036(csa_tree_add_110_49_pad_groupi_n_779 ,csa_tree_add_110_49_pad_groupi_n_543 ,csa_tree_add_110_49_pad_groupi_n_612);
  and csa_tree_add_110_49_pad_groupi_g5037(csa_tree_add_110_49_pad_groupi_n_778 ,csa_tree_add_110_49_pad_groupi_n_540 ,csa_tree_add_110_49_pad_groupi_n_644);
  and csa_tree_add_110_49_pad_groupi_g5038(csa_tree_add_110_49_pad_groupi_n_777 ,csa_tree_add_110_49_pad_groupi_n_552 ,csa_tree_add_110_49_pad_groupi_n_672);
  and csa_tree_add_110_49_pad_groupi_g5039(csa_tree_add_110_49_pad_groupi_n_775 ,csa_tree_add_110_49_pad_groupi_n_502 ,csa_tree_add_110_49_pad_groupi_n_670);
  or csa_tree_add_110_49_pad_groupi_g5040(csa_tree_add_110_49_pad_groupi_n_774 ,csa_tree_add_110_49_pad_groupi_n_569 ,csa_tree_add_110_49_pad_groupi_n_679);
  or csa_tree_add_110_49_pad_groupi_g5041(csa_tree_add_110_49_pad_groupi_n_773 ,csa_tree_add_110_49_pad_groupi_n_564 ,csa_tree_add_110_49_pad_groupi_n_682);
  and csa_tree_add_110_49_pad_groupi_g5042(csa_tree_add_110_49_pad_groupi_n_771 ,csa_tree_add_110_49_pad_groupi_n_535 ,csa_tree_add_110_49_pad_groupi_n_642);
  and csa_tree_add_110_49_pad_groupi_g5043(csa_tree_add_110_49_pad_groupi_n_770 ,csa_tree_add_110_49_pad_groupi_n_551 ,csa_tree_add_110_49_pad_groupi_n_652);
  and csa_tree_add_110_49_pad_groupi_g5044(csa_tree_add_110_49_pad_groupi_n_769 ,csa_tree_add_110_49_pad_groupi_n_473 ,csa_tree_add_110_49_pad_groupi_n_618);
  and csa_tree_add_110_49_pad_groupi_g5045(csa_tree_add_110_49_pad_groupi_n_768 ,csa_tree_add_110_49_pad_groupi_n_538 ,csa_tree_add_110_49_pad_groupi_n_651);
  or csa_tree_add_110_49_pad_groupi_g5046(csa_tree_add_110_49_pad_groupi_n_766 ,csa_tree_add_110_49_pad_groupi_n_562 ,csa_tree_add_110_49_pad_groupi_n_675);
  and csa_tree_add_110_49_pad_groupi_g5047(csa_tree_add_110_49_pad_groupi_n_765 ,csa_tree_add_110_49_pad_groupi_n_506 ,csa_tree_add_110_49_pad_groupi_n_650);
  and csa_tree_add_110_49_pad_groupi_g5048(csa_tree_add_110_49_pad_groupi_n_764 ,csa_tree_add_110_49_pad_groupi_n_532 ,csa_tree_add_110_49_pad_groupi_n_616);
  and csa_tree_add_110_49_pad_groupi_g5049(csa_tree_add_110_49_pad_groupi_n_763 ,csa_tree_add_110_49_pad_groupi_n_495 ,csa_tree_add_110_49_pad_groupi_n_660);
  or csa_tree_add_110_49_pad_groupi_g5050(csa_tree_add_110_49_pad_groupi_n_761 ,csa_tree_add_110_49_pad_groupi_n_566 ,csa_tree_add_110_49_pad_groupi_n_681);
  or csa_tree_add_110_49_pad_groupi_g5051(csa_tree_add_110_49_pad_groupi_n_759 ,csa_tree_add_110_49_pad_groupi_n_565 ,csa_tree_add_110_49_pad_groupi_n_684);
  and csa_tree_add_110_49_pad_groupi_g5052(csa_tree_add_110_49_pad_groupi_n_758 ,csa_tree_add_110_49_pad_groupi_n_549 ,csa_tree_add_110_49_pad_groupi_n_643);
  and csa_tree_add_110_49_pad_groupi_g5053(csa_tree_add_110_49_pad_groupi_n_756 ,csa_tree_add_110_49_pad_groupi_n_546 ,csa_tree_add_110_49_pad_groupi_n_649);
  and csa_tree_add_110_49_pad_groupi_g5054(csa_tree_add_110_49_pad_groupi_n_755 ,csa_tree_add_110_49_pad_groupi_n_534 ,csa_tree_add_110_49_pad_groupi_n_596);
  and csa_tree_add_110_49_pad_groupi_g5055(csa_tree_add_110_49_pad_groupi_n_753 ,csa_tree_add_110_49_pad_groupi_n_491 ,csa_tree_add_110_49_pad_groupi_n_610);
  or csa_tree_add_110_49_pad_groupi_g5056(csa_tree_add_110_49_pad_groupi_n_751 ,csa_tree_add_110_49_pad_groupi_n_568 ,csa_tree_add_110_49_pad_groupi_n_677);
  or csa_tree_add_110_49_pad_groupi_g5057(csa_tree_add_110_49_pad_groupi_n_750 ,csa_tree_add_110_49_pad_groupi_n_527 ,csa_tree_add_110_49_pad_groupi_n_584);
  and csa_tree_add_110_49_pad_groupi_g5058(csa_tree_add_110_49_pad_groupi_n_748 ,csa_tree_add_110_49_pad_groupi_n_530 ,csa_tree_add_110_49_pad_groupi_n_662);
  and csa_tree_add_110_49_pad_groupi_g5059(csa_tree_add_110_49_pad_groupi_n_746 ,csa_tree_add_110_49_pad_groupi_n_507 ,csa_tree_add_110_49_pad_groupi_n_655);
  and csa_tree_add_110_49_pad_groupi_g5060(csa_tree_add_110_49_pad_groupi_n_745 ,csa_tree_add_110_49_pad_groupi_n_500 ,csa_tree_add_110_49_pad_groupi_n_666);
  and csa_tree_add_110_49_pad_groupi_g5061(csa_tree_add_110_49_pad_groupi_n_743 ,csa_tree_add_110_49_pad_groupi_n_537 ,csa_tree_add_110_49_pad_groupi_n_668);
  not csa_tree_add_110_49_pad_groupi_g5062(csa_tree_add_110_49_pad_groupi_n_741 ,csa_tree_add_110_49_pad_groupi_n_740);
  not csa_tree_add_110_49_pad_groupi_g5063(csa_tree_add_110_49_pad_groupi_n_738 ,csa_tree_add_110_49_pad_groupi_n_737);
  not csa_tree_add_110_49_pad_groupi_g5064(csa_tree_add_110_49_pad_groupi_n_733 ,csa_tree_add_110_49_pad_groupi_n_732);
  not csa_tree_add_110_49_pad_groupi_g5065(csa_tree_add_110_49_pad_groupi_n_730 ,csa_tree_add_110_49_pad_groupi_n_729);
  not csa_tree_add_110_49_pad_groupi_g5066(csa_tree_add_110_49_pad_groupi_n_726 ,csa_tree_add_110_49_pad_groupi_n_727);
  not csa_tree_add_110_49_pad_groupi_g5067(csa_tree_add_110_49_pad_groupi_n_724 ,csa_tree_add_110_49_pad_groupi_n_725);
  not csa_tree_add_110_49_pad_groupi_g5068(csa_tree_add_110_49_pad_groupi_n_722 ,csa_tree_add_110_49_pad_groupi_n_723);
  not csa_tree_add_110_49_pad_groupi_g5069(csa_tree_add_110_49_pad_groupi_n_720 ,csa_tree_add_110_49_pad_groupi_n_721);
  not csa_tree_add_110_49_pad_groupi_g5070(csa_tree_add_110_49_pad_groupi_n_716 ,csa_tree_add_110_49_pad_groupi_n_715);
  not csa_tree_add_110_49_pad_groupi_g5071(csa_tree_add_110_49_pad_groupi_n_713 ,csa_tree_add_110_49_pad_groupi_n_714);
  not csa_tree_add_110_49_pad_groupi_g5072(csa_tree_add_110_49_pad_groupi_n_700 ,csa_tree_add_110_49_pad_groupi_n_701);
  not csa_tree_add_110_49_pad_groupi_g5073(csa_tree_add_110_49_pad_groupi_n_697 ,csa_tree_add_110_49_pad_groupi_n_698);
  not csa_tree_add_110_49_pad_groupi_g5074(csa_tree_add_110_49_pad_groupi_n_695 ,csa_tree_add_110_49_pad_groupi_n_696);
  not csa_tree_add_110_49_pad_groupi_g5075(csa_tree_add_110_49_pad_groupi_n_693 ,csa_tree_add_110_49_pad_groupi_n_694);
  or csa_tree_add_110_49_pad_groupi_g5077(csa_tree_add_110_49_pad_groupi_n_691 ,csa_tree_add_110_49_pad_groupi_n_572 ,csa_tree_add_110_49_pad_groupi_n_627);
  nor csa_tree_add_110_49_pad_groupi_g5078(csa_tree_add_110_49_pad_groupi_n_690 ,csa_tree_add_110_49_pad_groupi_n_573 ,csa_tree_add_110_49_pad_groupi_n_628);
  nor csa_tree_add_110_49_pad_groupi_g5079(csa_tree_add_110_49_pad_groupi_n_689 ,csa_tree_add_110_49_pad_groupi_n_486 ,csa_tree_add_110_49_pad_groupi_n_594);
  or csa_tree_add_110_49_pad_groupi_g5080(csa_tree_add_110_49_pad_groupi_n_688 ,csa_tree_add_110_49_pad_groupi_n_559 ,csa_tree_add_110_49_pad_groupi_n_678);
  and csa_tree_add_110_49_pad_groupi_g5081(csa_tree_add_110_49_pad_groupi_n_742 ,csa_tree_add_110_49_pad_groupi_n_482 ,csa_tree_add_110_49_pad_groupi_n_602);
  and csa_tree_add_110_49_pad_groupi_g5082(csa_tree_add_110_49_pad_groupi_n_740 ,csa_tree_add_110_49_pad_groupi_n_505 ,csa_tree_add_110_49_pad_groupi_n_614);
  and csa_tree_add_110_49_pad_groupi_g5083(csa_tree_add_110_49_pad_groupi_n_739 ,csa_tree_add_110_49_pad_groupi_n_484 ,csa_tree_add_110_49_pad_groupi_n_591);
  or csa_tree_add_110_49_pad_groupi_g5084(csa_tree_add_110_49_pad_groupi_n_687 ,csa_tree_add_110_49_pad_groupi_n_522 ,csa_tree_add_110_49_pad_groupi_n_586);
  or csa_tree_add_110_49_pad_groupi_g5085(csa_tree_add_110_49_pad_groupi_n_737 ,csa_tree_add_110_49_pad_groupi_n_557 ,csa_tree_add_110_49_pad_groupi_n_673);
  and csa_tree_add_110_49_pad_groupi_g5086(csa_tree_add_110_49_pad_groupi_n_736 ,csa_tree_add_110_49_pad_groupi_n_488 ,csa_tree_add_110_49_pad_groupi_n_603);
  or csa_tree_add_110_49_pad_groupi_g5087(csa_tree_add_110_49_pad_groupi_n_735 ,csa_tree_add_110_49_pad_groupi_n_556 ,csa_tree_add_110_49_pad_groupi_n_680);
  and csa_tree_add_110_49_pad_groupi_g5088(csa_tree_add_110_49_pad_groupi_n_734 ,csa_tree_add_110_49_pad_groupi_n_526 ,csa_tree_add_110_49_pad_groupi_n_648);
  or csa_tree_add_110_49_pad_groupi_g5089(csa_tree_add_110_49_pad_groupi_n_732 ,csa_tree_add_110_49_pad_groupi_n_558 ,csa_tree_add_110_49_pad_groupi_n_674);
  and csa_tree_add_110_49_pad_groupi_g5090(csa_tree_add_110_49_pad_groupi_n_731 ,csa_tree_add_110_49_pad_groupi_n_541 ,csa_tree_add_110_49_pad_groupi_n_658);
  or csa_tree_add_110_49_pad_groupi_g5091(csa_tree_add_110_49_pad_groupi_n_729 ,csa_tree_add_110_49_pad_groupi_n_560 ,csa_tree_add_110_49_pad_groupi_n_676);
  or csa_tree_add_110_49_pad_groupi_g5092(csa_tree_add_110_49_pad_groupi_n_728 ,csa_tree_add_110_49_pad_groupi_n_525 ,csa_tree_add_110_49_pad_groupi_n_585);
  or csa_tree_add_110_49_pad_groupi_g5093(csa_tree_add_110_49_pad_groupi_n_727 ,csa_tree_add_110_49_pad_groupi_n_327 ,csa_tree_add_110_49_pad_groupi_n_592);
  and csa_tree_add_110_49_pad_groupi_g5094(csa_tree_add_110_49_pad_groupi_n_725 ,csa_tree_add_110_49_pad_groupi_n_492 ,csa_tree_add_110_49_pad_groupi_n_606);
  and csa_tree_add_110_49_pad_groupi_g5095(csa_tree_add_110_49_pad_groupi_n_723 ,csa_tree_add_110_49_pad_groupi_n_498 ,csa_tree_add_110_49_pad_groupi_n_609);
  and csa_tree_add_110_49_pad_groupi_g5096(csa_tree_add_110_49_pad_groupi_n_721 ,csa_tree_add_110_49_pad_groupi_n_489 ,csa_tree_add_110_49_pad_groupi_n_605);
  and csa_tree_add_110_49_pad_groupi_g5097(csa_tree_add_110_49_pad_groupi_n_719 ,csa_tree_add_110_49_pad_groupi_n_544 ,csa_tree_add_110_49_pad_groupi_n_604);
  and csa_tree_add_110_49_pad_groupi_g5098(csa_tree_add_110_49_pad_groupi_n_718 ,csa_tree_add_110_49_pad_groupi_n_494 ,csa_tree_add_110_49_pad_groupi_n_608);
  and csa_tree_add_110_49_pad_groupi_g5099(csa_tree_add_110_49_pad_groupi_n_717 ,csa_tree_add_110_49_pad_groupi_n_490 ,csa_tree_add_110_49_pad_groupi_n_667);
  or csa_tree_add_110_49_pad_groupi_g5100(csa_tree_add_110_49_pad_groupi_n_715 ,csa_tree_add_110_49_pad_groupi_n_555 ,csa_tree_add_110_49_pad_groupi_n_663);
  and csa_tree_add_110_49_pad_groupi_g5101(csa_tree_add_110_49_pad_groupi_n_714 ,csa_tree_add_110_49_pad_groupi_n_523 ,csa_tree_add_110_49_pad_groupi_n_686);
  and csa_tree_add_110_49_pad_groupi_g5102(csa_tree_add_110_49_pad_groupi_n_712 ,csa_tree_add_110_49_pad_groupi_n_528 ,csa_tree_add_110_49_pad_groupi_n_654);
  and csa_tree_add_110_49_pad_groupi_g5103(csa_tree_add_110_49_pad_groupi_n_711 ,csa_tree_add_110_49_pad_groupi_n_483 ,csa_tree_add_110_49_pad_groupi_n_587);
  and csa_tree_add_110_49_pad_groupi_g5104(csa_tree_add_110_49_pad_groupi_n_710 ,csa_tree_add_110_49_pad_groupi_n_487 ,csa_tree_add_110_49_pad_groupi_n_590);
  and csa_tree_add_110_49_pad_groupi_g5105(csa_tree_add_110_49_pad_groupi_n_709 ,csa_tree_add_110_49_pad_groupi_n_478 ,csa_tree_add_110_49_pad_groupi_n_601);
  and csa_tree_add_110_49_pad_groupi_g5106(csa_tree_add_110_49_pad_groupi_n_708 ,csa_tree_add_110_49_pad_groupi_n_485 ,csa_tree_add_110_49_pad_groupi_n_600);
  and csa_tree_add_110_49_pad_groupi_g5107(csa_tree_add_110_49_pad_groupi_n_707 ,csa_tree_add_110_49_pad_groupi_n_479 ,csa_tree_add_110_49_pad_groupi_n_599);
  and csa_tree_add_110_49_pad_groupi_g5108(csa_tree_add_110_49_pad_groupi_n_706 ,csa_tree_add_110_49_pad_groupi_n_509 ,csa_tree_add_110_49_pad_groupi_n_598);
  and csa_tree_add_110_49_pad_groupi_g5109(csa_tree_add_110_49_pad_groupi_n_705 ,csa_tree_add_110_49_pad_groupi_n_481 ,csa_tree_add_110_49_pad_groupi_n_597);
  and csa_tree_add_110_49_pad_groupi_g5110(csa_tree_add_110_49_pad_groupi_n_704 ,csa_tree_add_110_49_pad_groupi_n_476 ,csa_tree_add_110_49_pad_groupi_n_619);
  and csa_tree_add_110_49_pad_groupi_g5111(csa_tree_add_110_49_pad_groupi_n_703 ,csa_tree_add_110_49_pad_groupi_n_477 ,csa_tree_add_110_49_pad_groupi_n_595);
  and csa_tree_add_110_49_pad_groupi_g5112(csa_tree_add_110_49_pad_groupi_n_702 ,csa_tree_add_110_49_pad_groupi_n_474 ,csa_tree_add_110_49_pad_groupi_n_589);
  or csa_tree_add_110_49_pad_groupi_g5113(csa_tree_add_110_49_pad_groupi_n_701 ,csa_tree_add_110_49_pad_groupi_n_567 ,csa_tree_add_110_49_pad_groupi_n_656);
  and csa_tree_add_110_49_pad_groupi_g5114(csa_tree_add_110_49_pad_groupi_n_699 ,csa_tree_add_110_49_pad_groupi_n_475 ,csa_tree_add_110_49_pad_groupi_n_593);
  and csa_tree_add_110_49_pad_groupi_g5115(csa_tree_add_110_49_pad_groupi_n_698 ,csa_tree_add_110_49_pad_groupi_n_493 ,csa_tree_add_110_49_pad_groupi_n_607);
  and csa_tree_add_110_49_pad_groupi_g5116(csa_tree_add_110_49_pad_groupi_n_696 ,csa_tree_add_110_49_pad_groupi_n_480 ,csa_tree_add_110_49_pad_groupi_n_588);
  and csa_tree_add_110_49_pad_groupi_g5117(csa_tree_add_110_49_pad_groupi_n_694 ,csa_tree_add_110_49_pad_groupi_n_548 ,csa_tree_add_110_49_pad_groupi_n_657);
  or csa_tree_add_110_49_pad_groupi_g5118(csa_tree_add_110_49_pad_groupi_n_692 ,csa_tree_add_110_49_pad_groupi_n_561 ,csa_tree_add_110_49_pad_groupi_n_685);
  or csa_tree_add_110_49_pad_groupi_g5119(csa_tree_add_110_49_pad_groupi_n_686 ,csa_tree_add_110_49_pad_groupi_n_402 ,csa_tree_add_110_49_pad_groupi_n_25);
  and csa_tree_add_110_49_pad_groupi_g5120(csa_tree_add_110_49_pad_groupi_n_685 ,csa_tree_add_110_49_pad_groupi_n_83 ,csa_tree_add_110_49_pad_groupi_n_155);
  and csa_tree_add_110_49_pad_groupi_g5121(csa_tree_add_110_49_pad_groupi_n_684 ,csa_tree_add_110_49_pad_groupi_n_77 ,csa_tree_add_110_49_pad_groupi_n_152);
  and csa_tree_add_110_49_pad_groupi_g5122(csa_tree_add_110_49_pad_groupi_n_683 ,csa_tree_add_110_49_pad_groupi_n_81 ,csa_tree_add_110_49_pad_groupi_n_151);
  and csa_tree_add_110_49_pad_groupi_g5123(csa_tree_add_110_49_pad_groupi_n_682 ,csa_tree_add_110_49_pad_groupi_n_95 ,csa_tree_add_110_49_pad_groupi_n_136);
  and csa_tree_add_110_49_pad_groupi_g5124(csa_tree_add_110_49_pad_groupi_n_681 ,csa_tree_add_110_49_pad_groupi_n_97 ,csa_tree_add_110_49_pad_groupi_n_134);
  and csa_tree_add_110_49_pad_groupi_g5125(csa_tree_add_110_49_pad_groupi_n_680 ,csa_tree_add_110_49_pad_groupi_n_89 ,csa_tree_add_110_49_pad_groupi_n_137);
  and csa_tree_add_110_49_pad_groupi_g5126(csa_tree_add_110_49_pad_groupi_n_679 ,csa_tree_add_110_49_pad_groupi_n_111 ,csa_tree_add_110_49_pad_groupi_n_133);
  and csa_tree_add_110_49_pad_groupi_g5127(csa_tree_add_110_49_pad_groupi_n_678 ,csa_tree_add_110_49_pad_groupi_n_75 ,csa_tree_add_110_49_pad_groupi_n_154);
  and csa_tree_add_110_49_pad_groupi_g5128(csa_tree_add_110_49_pad_groupi_n_677 ,csa_tree_add_110_49_pad_groupi_n_107 ,csa_tree_add_110_49_pad_groupi_n_154);
  and csa_tree_add_110_49_pad_groupi_g5129(csa_tree_add_110_49_pad_groupi_n_676 ,csa_tree_add_110_49_pad_groupi_n_119 ,csa_tree_add_110_49_pad_groupi_n_151);
  and csa_tree_add_110_49_pad_groupi_g5130(csa_tree_add_110_49_pad_groupi_n_675 ,csa_tree_add_110_49_pad_groupi_n_117 ,csa_tree_add_110_49_pad_groupi_n_137);
  and csa_tree_add_110_49_pad_groupi_g5131(csa_tree_add_110_49_pad_groupi_n_674 ,csa_tree_add_110_49_pad_groupi_n_125 ,csa_tree_add_110_49_pad_groupi_n_152);
  and csa_tree_add_110_49_pad_groupi_g5132(csa_tree_add_110_49_pad_groupi_n_673 ,csa_tree_add_110_49_pad_groupi_n_87 ,csa_tree_add_110_49_pad_groupi_n_134);
  or csa_tree_add_110_49_pad_groupi_g5133(csa_tree_add_110_49_pad_groupi_n_672 ,csa_tree_add_110_49_pad_groupi_n_398 ,csa_tree_add_110_49_pad_groupi_n_46);
  or csa_tree_add_110_49_pad_groupi_g5134(csa_tree_add_110_49_pad_groupi_n_671 ,csa_tree_add_110_49_pad_groupi_n_385 ,csa_tree_add_110_49_pad_groupi_n_28);
  or csa_tree_add_110_49_pad_groupi_g5135(csa_tree_add_110_49_pad_groupi_n_670 ,csa_tree_add_110_49_pad_groupi_n_403 ,csa_tree_add_110_49_pad_groupi_n_45);
  or csa_tree_add_110_49_pad_groupi_g5136(csa_tree_add_110_49_pad_groupi_n_669 ,csa_tree_add_110_49_pad_groupi_n_395 ,csa_tree_add_110_49_pad_groupi_n_66);
  or csa_tree_add_110_49_pad_groupi_g5137(csa_tree_add_110_49_pad_groupi_n_668 ,csa_tree_add_110_49_pad_groupi_n_405 ,csa_tree_add_110_49_pad_groupi_n_27);
  or csa_tree_add_110_49_pad_groupi_g5138(csa_tree_add_110_49_pad_groupi_n_667 ,csa_tree_add_110_49_pad_groupi_n_393 ,csa_tree_add_110_49_pad_groupi_n_25);
  or csa_tree_add_110_49_pad_groupi_g5139(csa_tree_add_110_49_pad_groupi_n_666 ,csa_tree_add_110_49_pad_groupi_n_392 ,csa_tree_add_110_49_pad_groupi_n_24);
  or csa_tree_add_110_49_pad_groupi_g5140(csa_tree_add_110_49_pad_groupi_n_665 ,csa_tree_add_110_49_pad_groupi_n_408 ,csa_tree_add_110_49_pad_groupi_n_24);
  or csa_tree_add_110_49_pad_groupi_g5141(csa_tree_add_110_49_pad_groupi_n_664 ,csa_tree_add_110_49_pad_groupi_n_406 ,csa_tree_add_110_49_pad_groupi_n_28);
  and csa_tree_add_110_49_pad_groupi_g5142(csa_tree_add_110_49_pad_groupi_n_663 ,csa_tree_add_110_49_pad_groupi_n_93 ,csa_tree_add_110_49_pad_groupi_n_155);
  or csa_tree_add_110_49_pad_groupi_g5143(csa_tree_add_110_49_pad_groupi_n_662 ,csa_tree_add_110_49_pad_groupi_n_401 ,csa_tree_add_110_49_pad_groupi_n_45);
  or csa_tree_add_110_49_pad_groupi_g5144(csa_tree_add_110_49_pad_groupi_n_661 ,csa_tree_add_110_49_pad_groupi_n_404 ,csa_tree_add_110_49_pad_groupi_n_66);
  or csa_tree_add_110_49_pad_groupi_g5145(csa_tree_add_110_49_pad_groupi_n_660 ,csa_tree_add_110_49_pad_groupi_n_400 ,csa_tree_add_110_49_pad_groupi_n_27);
  or csa_tree_add_110_49_pad_groupi_g5146(csa_tree_add_110_49_pad_groupi_n_659 ,csa_tree_add_110_49_pad_groupi_n_394 ,csa_tree_add_110_49_pad_groupi_n_7);
  or csa_tree_add_110_49_pad_groupi_g5147(csa_tree_add_110_49_pad_groupi_n_658 ,csa_tree_add_110_49_pad_groupi_n_419 ,csa_tree_add_110_49_pad_groupi_n_7);
  or csa_tree_add_110_49_pad_groupi_g5148(csa_tree_add_110_49_pad_groupi_n_657 ,csa_tree_add_110_49_pad_groupi_n_397 ,csa_tree_add_110_49_pad_groupi_n_67);
  nor csa_tree_add_110_49_pad_groupi_g5149(csa_tree_add_110_49_pad_groupi_n_656 ,csa_tree_add_110_49_pad_groupi_n_176 ,csa_tree_add_110_49_pad_groupi_n_512);
  or csa_tree_add_110_49_pad_groupi_g5150(csa_tree_add_110_49_pad_groupi_n_655 ,csa_tree_add_110_49_pad_groupi_n_417 ,csa_tree_add_110_49_pad_groupi_n_37);
  or csa_tree_add_110_49_pad_groupi_g5151(csa_tree_add_110_49_pad_groupi_n_654 ,csa_tree_add_110_49_pad_groupi_n_457 ,csa_tree_add_110_49_pad_groupi_n_31);
  or csa_tree_add_110_49_pad_groupi_g5152(csa_tree_add_110_49_pad_groupi_n_653 ,csa_tree_add_110_49_pad_groupi_n_413 ,csa_tree_add_110_49_pad_groupi_n_43);
  or csa_tree_add_110_49_pad_groupi_g5153(csa_tree_add_110_49_pad_groupi_n_652 ,csa_tree_add_110_49_pad_groupi_n_451 ,csa_tree_add_110_49_pad_groupi_n_55);
  or csa_tree_add_110_49_pad_groupi_g5154(csa_tree_add_110_49_pad_groupi_n_651 ,csa_tree_add_110_49_pad_groupi_n_453 ,csa_tree_add_110_49_pad_groupi_n_22);
  or csa_tree_add_110_49_pad_groupi_g5155(csa_tree_add_110_49_pad_groupi_n_650 ,csa_tree_add_110_49_pad_groupi_n_416 ,csa_tree_add_110_49_pad_groupi_n_16);
  or csa_tree_add_110_49_pad_groupi_g5156(csa_tree_add_110_49_pad_groupi_n_649 ,csa_tree_add_110_49_pad_groupi_n_458 ,csa_tree_add_110_49_pad_groupi_n_42);
  or csa_tree_add_110_49_pad_groupi_g5157(csa_tree_add_110_49_pad_groupi_n_648 ,csa_tree_add_110_49_pad_groupi_n_449 ,csa_tree_add_110_49_pad_groupi_n_54);
  or csa_tree_add_110_49_pad_groupi_g5158(csa_tree_add_110_49_pad_groupi_n_647 ,csa_tree_add_110_49_pad_groupi_n_415 ,csa_tree_add_110_49_pad_groupi_n_69);
  or csa_tree_add_110_49_pad_groupi_g5159(csa_tree_add_110_49_pad_groupi_n_646 ,csa_tree_add_110_49_pad_groupi_n_452 ,csa_tree_add_110_49_pad_groupi_n_15);
  or csa_tree_add_110_49_pad_groupi_g5160(csa_tree_add_110_49_pad_groupi_n_645 ,csa_tree_add_110_49_pad_groupi_n_443 ,csa_tree_add_110_49_pad_groupi_n_37);
  or csa_tree_add_110_49_pad_groupi_g5161(csa_tree_add_110_49_pad_groupi_n_644 ,csa_tree_add_110_49_pad_groupi_n_447 ,csa_tree_add_110_49_pad_groupi_n_36);
  or csa_tree_add_110_49_pad_groupi_g5162(csa_tree_add_110_49_pad_groupi_n_643 ,csa_tree_add_110_49_pad_groupi_n_445 ,csa_tree_add_110_49_pad_groupi_n_63);
  or csa_tree_add_110_49_pad_groupi_g5163(csa_tree_add_110_49_pad_groupi_n_642 ,csa_tree_add_110_49_pad_groupi_n_418 ,csa_tree_add_110_49_pad_groupi_n_36);
  or csa_tree_add_110_49_pad_groupi_g5164(csa_tree_add_110_49_pad_groupi_n_641 ,csa_tree_add_110_49_pad_groupi_n_459 ,csa_tree_add_110_49_pad_groupi_n_21);
  not csa_tree_add_110_49_pad_groupi_g5165(csa_tree_add_110_49_pad_groupi_n_640 ,csa_tree_add_110_49_pad_groupi_n_639);
  not csa_tree_add_110_49_pad_groupi_g5166(csa_tree_add_110_49_pad_groupi_n_638 ,csa_tree_add_110_49_pad_groupi_n_637);
  not csa_tree_add_110_49_pad_groupi_g5167(csa_tree_add_110_49_pad_groupi_n_636 ,csa_tree_add_110_49_pad_groupi_n_635);
  not csa_tree_add_110_49_pad_groupi_g5168(csa_tree_add_110_49_pad_groupi_n_633 ,csa_tree_add_110_49_pad_groupi_n_634);
  not csa_tree_add_110_49_pad_groupi_g5169(csa_tree_add_110_49_pad_groupi_n_631 ,csa_tree_add_110_49_pad_groupi_n_632);
  not csa_tree_add_110_49_pad_groupi_g5170(csa_tree_add_110_49_pad_groupi_n_629 ,csa_tree_add_110_49_pad_groupi_n_630);
  not csa_tree_add_110_49_pad_groupi_g5171(csa_tree_add_110_49_pad_groupi_n_627 ,csa_tree_add_110_49_pad_groupi_n_628);
  not csa_tree_add_110_49_pad_groupi_g5172(csa_tree_add_110_49_pad_groupi_n_624 ,csa_tree_add_110_49_pad_groupi_n_625);
  not csa_tree_add_110_49_pad_groupi_g5173(csa_tree_add_110_49_pad_groupi_n_622 ,csa_tree_add_110_49_pad_groupi_n_623);
  not csa_tree_add_110_49_pad_groupi_g5174(csa_tree_add_110_49_pad_groupi_n_620 ,csa_tree_add_110_49_pad_groupi_n_621);
  or csa_tree_add_110_49_pad_groupi_g5175(csa_tree_add_110_49_pad_groupi_n_619 ,csa_tree_add_110_49_pad_groupi_n_442 ,csa_tree_add_110_49_pad_groupi_n_58);
  or csa_tree_add_110_49_pad_groupi_g5176(csa_tree_add_110_49_pad_groupi_n_618 ,csa_tree_add_110_49_pad_groupi_n_407 ,csa_tree_add_110_49_pad_groupi_n_31);
  or csa_tree_add_110_49_pad_groupi_g5177(csa_tree_add_110_49_pad_groupi_n_617 ,csa_tree_add_110_49_pad_groupi_n_448 ,csa_tree_add_110_49_pad_groupi_n_16);
  or csa_tree_add_110_49_pad_groupi_g5178(csa_tree_add_110_49_pad_groupi_n_616 ,csa_tree_add_110_49_pad_groupi_n_399 ,csa_tree_add_110_49_pad_groupi_n_54);
  or csa_tree_add_110_49_pad_groupi_g5179(csa_tree_add_110_49_pad_groupi_n_615 ,csa_tree_add_110_49_pad_groupi_n_412 ,csa_tree_add_110_49_pad_groupi_n_69);
  or csa_tree_add_110_49_pad_groupi_g5180(csa_tree_add_110_49_pad_groupi_n_614 ,csa_tree_add_110_49_pad_groupi_n_422 ,csa_tree_add_110_49_pad_groupi_n_15);
  or csa_tree_add_110_49_pad_groupi_g5181(csa_tree_add_110_49_pad_groupi_n_613 ,csa_tree_add_110_49_pad_groupi_n_382 ,csa_tree_add_110_49_pad_groupi_n_30);
  or csa_tree_add_110_49_pad_groupi_g5182(csa_tree_add_110_49_pad_groupi_n_612 ,csa_tree_add_110_49_pad_groupi_n_446 ,csa_tree_add_110_49_pad_groupi_n_30);
  or csa_tree_add_110_49_pad_groupi_g5183(csa_tree_add_110_49_pad_groupi_n_611 ,csa_tree_add_110_49_pad_groupi_n_455 ,csa_tree_add_110_49_pad_groupi_n_5);
  or csa_tree_add_110_49_pad_groupi_g5184(csa_tree_add_110_49_pad_groupi_n_610 ,csa_tree_add_110_49_pad_groupi_n_409 ,csa_tree_add_110_49_pad_groupi_n_22);
  or csa_tree_add_110_49_pad_groupi_g5185(csa_tree_add_110_49_pad_groupi_n_609 ,csa_tree_add_110_49_pad_groupi_n_396 ,csa_tree_add_110_49_pad_groupi_n_42);
  or csa_tree_add_110_49_pad_groupi_g5186(csa_tree_add_110_49_pad_groupi_n_608 ,csa_tree_add_110_49_pad_groupi_n_441 ,csa_tree_add_110_49_pad_groupi_n_63);
  or csa_tree_add_110_49_pad_groupi_g5187(csa_tree_add_110_49_pad_groupi_n_607 ,csa_tree_add_110_49_pad_groupi_n_444 ,csa_tree_add_110_49_pad_groupi_n_21);
  or csa_tree_add_110_49_pad_groupi_g5188(csa_tree_add_110_49_pad_groupi_n_606 ,csa_tree_add_110_49_pad_groupi_n_454 ,csa_tree_add_110_49_pad_groupi_n_5);
  or csa_tree_add_110_49_pad_groupi_g5189(csa_tree_add_110_49_pad_groupi_n_605 ,csa_tree_add_110_49_pad_groupi_n_456 ,csa_tree_add_110_49_pad_groupi_n_9);
  or csa_tree_add_110_49_pad_groupi_g5190(csa_tree_add_110_49_pad_groupi_n_604 ,csa_tree_add_110_49_pad_groupi_n_411 ,csa_tree_add_110_49_pad_groupi_n_9);
  or csa_tree_add_110_49_pad_groupi_g5191(csa_tree_add_110_49_pad_groupi_n_603 ,csa_tree_add_110_49_pad_groupi_n_410 ,csa_tree_add_110_49_pad_groupi_n_70);
  or csa_tree_add_110_49_pad_groupi_g5192(csa_tree_add_110_49_pad_groupi_n_602 ,csa_tree_add_110_49_pad_groupi_n_467 ,csa_tree_add_110_49_pad_groupi_n_33);
  or csa_tree_add_110_49_pad_groupi_g5193(csa_tree_add_110_49_pad_groupi_n_601 ,csa_tree_add_110_49_pad_groupi_n_464 ,csa_tree_add_110_49_pad_groupi_n_19);
  or csa_tree_add_110_49_pad_groupi_g5194(csa_tree_add_110_49_pad_groupi_n_600 ,csa_tree_add_110_49_pad_groupi_n_450 ,csa_tree_add_110_49_pad_groupi_n_34);
  or csa_tree_add_110_49_pad_groupi_g5195(csa_tree_add_110_49_pad_groupi_n_599 ,csa_tree_add_110_49_pad_groupi_n_469 ,csa_tree_add_110_49_pad_groupi_n_18);
  or csa_tree_add_110_49_pad_groupi_g5196(csa_tree_add_110_49_pad_groupi_n_598 ,csa_tree_add_110_49_pad_groupi_n_460 ,csa_tree_add_110_49_pad_groupi_n_57);
  or csa_tree_add_110_49_pad_groupi_g5197(csa_tree_add_110_49_pad_groupi_n_597 ,csa_tree_add_110_49_pad_groupi_n_472 ,csa_tree_add_110_49_pad_groupi_n_39);
  or csa_tree_add_110_49_pad_groupi_g5198(csa_tree_add_110_49_pad_groupi_n_596 ,csa_tree_add_110_49_pad_groupi_n_414 ,csa_tree_add_110_49_pad_groupi_n_64);
  or csa_tree_add_110_49_pad_groupi_g5199(csa_tree_add_110_49_pad_groupi_n_595 ,csa_tree_add_110_49_pad_groupi_n_471 ,csa_tree_add_110_49_pad_groupi_n_19);
  nor csa_tree_add_110_49_pad_groupi_g5200(csa_tree_add_110_49_pad_groupi_n_594 ,csa_tree_add_110_49_pad_groupi_n_40 ,csa_tree_add_110_49_pad_groupi_n_420);
  or csa_tree_add_110_49_pad_groupi_g5201(csa_tree_add_110_49_pad_groupi_n_593 ,csa_tree_add_110_49_pad_groupi_n_470 ,csa_tree_add_110_49_pad_groupi_n_33);
  nor csa_tree_add_110_49_pad_groupi_g5202(csa_tree_add_110_49_pad_groupi_n_592 ,csa_tree_add_110_49_pad_groupi_n_58 ,csa_tree_add_110_49_pad_groupi_n_463);
  or csa_tree_add_110_49_pad_groupi_g5203(csa_tree_add_110_49_pad_groupi_n_591 ,csa_tree_add_110_49_pad_groupi_n_461 ,csa_tree_add_110_49_pad_groupi_n_57);
  or csa_tree_add_110_49_pad_groupi_g5204(csa_tree_add_110_49_pad_groupi_n_590 ,csa_tree_add_110_49_pad_groupi_n_468 ,csa_tree_add_110_49_pad_groupi_n_40);
  or csa_tree_add_110_49_pad_groupi_g5205(csa_tree_add_110_49_pad_groupi_n_589 ,csa_tree_add_110_49_pad_groupi_n_466 ,csa_tree_add_110_49_pad_groupi_n_39);
  or csa_tree_add_110_49_pad_groupi_g5206(csa_tree_add_110_49_pad_groupi_n_588 ,csa_tree_add_110_49_pad_groupi_n_462 ,csa_tree_add_110_49_pad_groupi_n_34);
  or csa_tree_add_110_49_pad_groupi_g5207(csa_tree_add_110_49_pad_groupi_n_587 ,csa_tree_add_110_49_pad_groupi_n_465 ,csa_tree_add_110_49_pad_groupi_n_18);
  nor csa_tree_add_110_49_pad_groupi_g5208(csa_tree_add_110_49_pad_groupi_n_586 ,csa_tree_add_110_49_pad_groupi_n_46 ,csa_tree_add_110_49_pad_groupi_n_292);
  nor csa_tree_add_110_49_pad_groupi_g5209(csa_tree_add_110_49_pad_groupi_n_585 ,csa_tree_add_110_49_pad_groupi_n_55 ,csa_tree_add_110_49_pad_groupi_n_291);
  nor csa_tree_add_110_49_pad_groupi_g5210(csa_tree_add_110_49_pad_groupi_n_584 ,csa_tree_add_110_49_pad_groupi_n_43 ,csa_tree_add_110_49_pad_groupi_n_290);
  or csa_tree_add_110_49_pad_groupi_g5211(csa_tree_add_110_49_pad_groupi_n_639 ,csa_tree_add_110_49_pad_groupi_n_192 ,csa_tree_add_110_49_pad_groupi_n_539);
  or csa_tree_add_110_49_pad_groupi_g5212(csa_tree_add_110_49_pad_groupi_n_637 ,csa_tree_add_110_49_pad_groupi_n_190 ,csa_tree_add_110_49_pad_groupi_n_547);
  or csa_tree_add_110_49_pad_groupi_g5213(csa_tree_add_110_49_pad_groupi_n_635 ,csa_tree_add_110_49_pad_groupi_n_292 ,csa_tree_add_110_49_pad_groupi_n_508);
  xnor csa_tree_add_110_49_pad_groupi_g5214(csa_tree_add_110_49_pad_groupi_n_634 ,csa_tree_add_110_49_pad_groupi_n_371 ,n_186);
  xnor csa_tree_add_110_49_pad_groupi_g5215(csa_tree_add_110_49_pad_groupi_n_632 ,csa_tree_add_110_49_pad_groupi_n_374 ,n_177);
  xnor csa_tree_add_110_49_pad_groupi_g5216(csa_tree_add_110_49_pad_groupi_n_630 ,csa_tree_add_110_49_pad_groupi_n_380 ,n_144);
  xnor csa_tree_add_110_49_pad_groupi_g5217(csa_tree_add_110_49_pad_groupi_n_628 ,csa_tree_add_110_49_pad_groupi_n_376 ,n_252);
  xnor csa_tree_add_110_49_pad_groupi_g5218(csa_tree_add_110_49_pad_groupi_n_626 ,csa_tree_add_110_49_pad_groupi_n_367 ,n_175);
  xnor csa_tree_add_110_49_pad_groupi_g5219(csa_tree_add_110_49_pad_groupi_n_625 ,csa_tree_add_110_49_pad_groupi_n_373 ,n_155);
  xnor csa_tree_add_110_49_pad_groupi_g5220(csa_tree_add_110_49_pad_groupi_n_623 ,csa_tree_add_110_49_pad_groupi_n_379 ,n_243);
  xnor csa_tree_add_110_49_pad_groupi_g5221(csa_tree_add_110_49_pad_groupi_n_621 ,csa_tree_add_110_49_pad_groupi_n_372 ,n_146);
  not csa_tree_add_110_49_pad_groupi_g5222(csa_tree_add_110_49_pad_groupi_n_582 ,csa_tree_add_110_49_pad_groupi_n_583);
  not csa_tree_add_110_49_pad_groupi_g5223(csa_tree_add_110_49_pad_groupi_n_580 ,csa_tree_add_110_49_pad_groupi_n_581);
  not csa_tree_add_110_49_pad_groupi_g5224(csa_tree_add_110_49_pad_groupi_n_579 ,csa_tree_add_110_49_pad_groupi_n_578);
  not csa_tree_add_110_49_pad_groupi_g5225(csa_tree_add_110_49_pad_groupi_n_576 ,csa_tree_add_110_49_pad_groupi_n_577);
  not csa_tree_add_110_49_pad_groupi_g5226(csa_tree_add_110_49_pad_groupi_n_574 ,csa_tree_add_110_49_pad_groupi_n_575);
  not csa_tree_add_110_49_pad_groupi_g5227(csa_tree_add_110_49_pad_groupi_n_572 ,csa_tree_add_110_49_pad_groupi_n_573);
  and csa_tree_add_110_49_pad_groupi_g5228(csa_tree_add_110_49_pad_groupi_n_569 ,csa_tree_add_110_49_pad_groupi_n_87 ,csa_tree_add_110_49_pad_groupi_n_157);
  and csa_tree_add_110_49_pad_groupi_g5229(csa_tree_add_110_49_pad_groupi_n_568 ,csa_tree_add_110_49_pad_groupi_n_117 ,csa_tree_add_110_49_pad_groupi_n_160);
  and csa_tree_add_110_49_pad_groupi_g5230(csa_tree_add_110_49_pad_groupi_n_567 ,csa_tree_add_110_49_pad_groupi_n_119 ,csa_tree_add_110_49_pad_groupi_n_161);
  and csa_tree_add_110_49_pad_groupi_g5231(csa_tree_add_110_49_pad_groupi_n_566 ,csa_tree_add_110_49_pad_groupi_n_89 ,csa_tree_add_110_49_pad_groupi_n_161);
  and csa_tree_add_110_49_pad_groupi_g5232(csa_tree_add_110_49_pad_groupi_n_565 ,csa_tree_add_110_49_pad_groupi_n_111 ,csa_tree_add_110_49_pad_groupi_n_163);
  and csa_tree_add_110_49_pad_groupi_g5233(csa_tree_add_110_49_pad_groupi_n_564 ,csa_tree_add_110_49_pad_groupi_n_77 ,csa_tree_add_110_49_pad_groupi_n_149);
  and csa_tree_add_110_49_pad_groupi_g5234(csa_tree_add_110_49_pad_groupi_n_563 ,csa_tree_add_110_49_pad_groupi_n_83 ,csa_tree_add_110_49_pad_groupi_n_148);
  and csa_tree_add_110_49_pad_groupi_g5235(csa_tree_add_110_49_pad_groupi_n_562 ,csa_tree_add_110_49_pad_groupi_n_97 ,csa_tree_add_110_49_pad_groupi_n_158);
  and csa_tree_add_110_49_pad_groupi_g5236(csa_tree_add_110_49_pad_groupi_n_561 ,csa_tree_add_110_49_pad_groupi_n_75 ,csa_tree_add_110_49_pad_groupi_n_164);
  and csa_tree_add_110_49_pad_groupi_g5237(csa_tree_add_110_49_pad_groupi_n_560 ,csa_tree_add_110_49_pad_groupi_n_107 ,csa_tree_add_110_49_pad_groupi_n_160);
  and csa_tree_add_110_49_pad_groupi_g5238(csa_tree_add_110_49_pad_groupi_n_559 ,csa_tree_add_110_49_pad_groupi_n_233 ,csa_tree_add_110_49_pad_groupi_n_157);
  and csa_tree_add_110_49_pad_groupi_g5239(csa_tree_add_110_49_pad_groupi_n_558 ,csa_tree_add_110_49_pad_groupi_n_95 ,csa_tree_add_110_49_pad_groupi_n_158);
  and csa_tree_add_110_49_pad_groupi_g5240(csa_tree_add_110_49_pad_groupi_n_557 ,csa_tree_add_110_49_pad_groupi_n_93 ,csa_tree_add_110_49_pad_groupi_n_149);
  and csa_tree_add_110_49_pad_groupi_g5241(csa_tree_add_110_49_pad_groupi_n_556 ,csa_tree_add_110_49_pad_groupi_n_125 ,csa_tree_add_110_49_pad_groupi_n_164);
  and csa_tree_add_110_49_pad_groupi_g5242(csa_tree_add_110_49_pad_groupi_n_555 ,csa_tree_add_110_49_pad_groupi_n_81 ,csa_tree_add_110_49_pad_groupi_n_148);
  or csa_tree_add_110_49_pad_groupi_g5243(csa_tree_add_110_49_pad_groupi_n_554 ,csa_tree_add_110_49_pad_groupi_n_407 ,csa_tree_add_110_49_pad_groupi_n_217);
  or csa_tree_add_110_49_pad_groupi_g5244(csa_tree_add_110_49_pad_groupi_n_553 ,csa_tree_add_110_49_pad_groupi_n_457 ,csa_tree_add_110_49_pad_groupi_n_226);
  or csa_tree_add_110_49_pad_groupi_g5245(csa_tree_add_110_49_pad_groupi_n_552 ,csa_tree_add_110_49_pad_groupi_n_405 ,csa_tree_add_110_49_pad_groupi_n_199);
  or csa_tree_add_110_49_pad_groupi_g5246(csa_tree_add_110_49_pad_groupi_n_551 ,csa_tree_add_110_49_pad_groupi_n_410 ,csa_tree_add_110_49_pad_groupi_n_214);
  or csa_tree_add_110_49_pad_groupi_g5247(csa_tree_add_110_49_pad_groupi_n_550 ,csa_tree_add_110_49_pad_groupi_n_419 ,csa_tree_add_110_49_pad_groupi_n_205);
  or csa_tree_add_110_49_pad_groupi_g5248(csa_tree_add_110_49_pad_groupi_n_549 ,csa_tree_add_110_49_pad_groupi_n_413 ,csa_tree_add_110_49_pad_groupi_n_226);
  or csa_tree_add_110_49_pad_groupi_g5249(csa_tree_add_110_49_pad_groupi_n_548 ,csa_tree_add_110_49_pad_groupi_n_398 ,csa_tree_add_110_49_pad_groupi_n_205);
  nor csa_tree_add_110_49_pad_groupi_g5250(csa_tree_add_110_49_pad_groupi_n_547 ,csa_tree_add_110_49_pad_groupi_n_351 ,csa_tree_add_110_49_pad_groupi_n_424);
  or csa_tree_add_110_49_pad_groupi_g5251(csa_tree_add_110_49_pad_groupi_n_546 ,csa_tree_add_110_49_pad_groupi_n_445 ,csa_tree_add_110_49_pad_groupi_n_218);
  or csa_tree_add_110_49_pad_groupi_g5252(csa_tree_add_110_49_pad_groupi_n_545 ,csa_tree_add_110_49_pad_groupi_n_416 ,csa_tree_add_110_49_pad_groupi_n_196);
  or csa_tree_add_110_49_pad_groupi_g5253(csa_tree_add_110_49_pad_groupi_n_544 ,csa_tree_add_110_49_pad_groupi_n_409 ,csa_tree_add_110_49_pad_groupi_n_221);
  or csa_tree_add_110_49_pad_groupi_g5254(csa_tree_add_110_49_pad_groupi_n_543 ,csa_tree_add_110_49_pad_groupi_n_453 ,csa_tree_add_110_49_pad_groupi_n_217);
  or csa_tree_add_110_49_pad_groupi_g5255(csa_tree_add_110_49_pad_groupi_n_542 ,csa_tree_add_110_49_pad_groupi_n_414 ,csa_tree_add_110_49_pad_groupi_n_220);
  or csa_tree_add_110_49_pad_groupi_g5256(csa_tree_add_110_49_pad_groupi_n_541 ,csa_tree_add_110_49_pad_groupi_n_394 ,csa_tree_add_110_49_pad_groupi_n_200);
  or csa_tree_add_110_49_pad_groupi_g5257(csa_tree_add_110_49_pad_groupi_n_540 ,csa_tree_add_110_49_pad_groupi_n_452 ,csa_tree_add_110_49_pad_groupi_n_196);
  nor csa_tree_add_110_49_pad_groupi_g5258(csa_tree_add_110_49_pad_groupi_n_539 ,csa_tree_add_110_49_pad_groupi_n_332 ,csa_tree_add_110_49_pad_groupi_n_426);
  or csa_tree_add_110_49_pad_groupi_g5259(csa_tree_add_110_49_pad_groupi_n_538 ,csa_tree_add_110_49_pad_groupi_n_444 ,csa_tree_add_110_49_pad_groupi_n_223);
  or csa_tree_add_110_49_pad_groupi_g5260(csa_tree_add_110_49_pad_groupi_n_537 ,csa_tree_add_110_49_pad_groupi_n_401 ,csa_tree_add_110_49_pad_groupi_n_203);
  or csa_tree_add_110_49_pad_groupi_g5261(csa_tree_add_110_49_pad_groupi_n_536 ,csa_tree_add_110_49_pad_groupi_n_408 ,csa_tree_add_110_49_pad_groupi_n_199);
  or csa_tree_add_110_49_pad_groupi_g5262(csa_tree_add_110_49_pad_groupi_n_535 ,csa_tree_add_110_49_pad_groupi_n_415 ,csa_tree_add_110_49_pad_groupi_n_215);
  or csa_tree_add_110_49_pad_groupi_g5263(csa_tree_add_110_49_pad_groupi_n_534 ,csa_tree_add_110_49_pad_groupi_n_456 ,csa_tree_add_110_49_pad_groupi_n_223);
  or csa_tree_add_110_49_pad_groupi_g5264(csa_tree_add_110_49_pad_groupi_n_533 ,csa_tree_add_110_49_pad_groupi_n_451 ,csa_tree_add_110_49_pad_groupi_n_209);
  or csa_tree_add_110_49_pad_groupi_g5265(csa_tree_add_110_49_pad_groupi_n_532 ,csa_tree_add_110_49_pad_groupi_n_448 ,csa_tree_add_110_49_pad_groupi_n_214);
  or csa_tree_add_110_49_pad_groupi_g5266(csa_tree_add_110_49_pad_groupi_n_531 ,csa_tree_add_110_49_pad_groupi_n_406 ,csa_tree_add_110_49_pad_groupi_n_202);
  or csa_tree_add_110_49_pad_groupi_g5267(csa_tree_add_110_49_pad_groupi_n_530 ,csa_tree_add_110_49_pad_groupi_n_402 ,csa_tree_add_110_49_pad_groupi_n_229);
  or csa_tree_add_110_49_pad_groupi_g5268(csa_tree_add_110_49_pad_groupi_n_529 ,csa_tree_add_110_49_pad_groupi_n_403 ,csa_tree_add_110_49_pad_groupi_n_229);
  or csa_tree_add_110_49_pad_groupi_g5269(csa_tree_add_110_49_pad_groupi_n_583 ,csa_tree_add_110_49_pad_groupi_n_349 ,csa_tree_add_110_49_pad_groupi_n_432);
  or csa_tree_add_110_49_pad_groupi_g5270(csa_tree_add_110_49_pad_groupi_n_581 ,csa_tree_add_110_49_pad_groupi_n_321 ,csa_tree_add_110_49_pad_groupi_n_433);
  or csa_tree_add_110_49_pad_groupi_g5271(csa_tree_add_110_49_pad_groupi_n_578 ,csa_tree_add_110_49_pad_groupi_n_364 ,csa_tree_add_110_49_pad_groupi_n_431);
  or csa_tree_add_110_49_pad_groupi_g5272(csa_tree_add_110_49_pad_groupi_n_577 ,csa_tree_add_110_49_pad_groupi_n_315 ,csa_tree_add_110_49_pad_groupi_n_428);
  or csa_tree_add_110_49_pad_groupi_g5273(csa_tree_add_110_49_pad_groupi_n_575 ,csa_tree_add_110_49_pad_groupi_n_356 ,csa_tree_add_110_49_pad_groupi_n_429);
  or csa_tree_add_110_49_pad_groupi_g5274(csa_tree_add_110_49_pad_groupi_n_573 ,csa_tree_add_110_49_pad_groupi_n_362 ,csa_tree_add_110_49_pad_groupi_n_423);
  or csa_tree_add_110_49_pad_groupi_g5275(csa_tree_add_110_49_pad_groupi_n_571 ,in16[0] ,csa_tree_add_110_49_pad_groupi_n_421);
  or csa_tree_add_110_49_pad_groupi_g5276(csa_tree_add_110_49_pad_groupi_n_570 ,csa_tree_add_110_49_pad_groupi_n_383 ,csa_tree_add_110_49_pad_groupi_n_141);
  not csa_tree_add_110_49_pad_groupi_g5277(csa_tree_add_110_49_pad_groupi_n_528 ,csa_tree_add_110_49_pad_groupi_n_527);
  not csa_tree_add_110_49_pad_groupi_g5278(csa_tree_add_110_49_pad_groupi_n_526 ,csa_tree_add_110_49_pad_groupi_n_525);
  not csa_tree_add_110_49_pad_groupi_g5279(csa_tree_add_110_49_pad_groupi_n_523 ,csa_tree_add_110_49_pad_groupi_n_522);
  not csa_tree_add_110_49_pad_groupi_g5280(csa_tree_add_110_49_pad_groupi_n_518 ,csa_tree_add_110_49_pad_groupi_n_519);
  not csa_tree_add_110_49_pad_groupi_g5281(csa_tree_add_110_49_pad_groupi_n_516 ,csa_tree_add_110_49_pad_groupi_n_517);
  not csa_tree_add_110_49_pad_groupi_g5282(csa_tree_add_110_49_pad_groupi_n_514 ,csa_tree_add_110_49_pad_groupi_n_512);
  not csa_tree_add_110_49_pad_groupi_g5283(csa_tree_add_110_49_pad_groupi_n_513 ,csa_tree_add_110_49_pad_groupi_n_512);
  or csa_tree_add_110_49_pad_groupi_g5284(csa_tree_add_110_49_pad_groupi_n_509 ,csa_tree_add_110_49_pad_groupi_n_52 ,csa_tree_add_110_49_pad_groupi_n_450);
  nor csa_tree_add_110_49_pad_groupi_g5285(csa_tree_add_110_49_pad_groupi_n_508 ,csa_tree_add_110_49_pad_groupi_n_355 ,csa_tree_add_110_49_pad_groupi_n_425);
  or csa_tree_add_110_49_pad_groupi_g5286(csa_tree_add_110_49_pad_groupi_n_507 ,csa_tree_add_110_49_pad_groupi_n_418 ,csa_tree_add_110_49_pad_groupi_n_208);
  or csa_tree_add_110_49_pad_groupi_g5287(csa_tree_add_110_49_pad_groupi_n_506 ,csa_tree_add_110_49_pad_groupi_n_454 ,csa_tree_add_110_49_pad_groupi_n_211);
  or csa_tree_add_110_49_pad_groupi_g5288(csa_tree_add_110_49_pad_groupi_n_505 ,csa_tree_add_110_49_pad_groupi_n_412 ,csa_tree_add_110_49_pad_groupi_n_211);
  or csa_tree_add_110_49_pad_groupi_g5289(csa_tree_add_110_49_pad_groupi_n_504 ,csa_tree_add_110_49_pad_groupi_n_447 ,csa_tree_add_110_49_pad_groupi_n_208);
  or csa_tree_add_110_49_pad_groupi_g5290(csa_tree_add_110_49_pad_groupi_n_503 ,csa_tree_add_110_49_pad_groupi_n_399 ,csa_tree_add_110_49_pad_groupi_n_197);
  or csa_tree_add_110_49_pad_groupi_g5291(csa_tree_add_110_49_pad_groupi_n_502 ,csa_tree_add_110_49_pad_groupi_n_400 ,csa_tree_add_110_49_pad_groupi_n_202);
  or csa_tree_add_110_49_pad_groupi_g5292(csa_tree_add_110_49_pad_groupi_n_501 ,csa_tree_add_110_49_pad_groupi_n_443 ,csa_tree_add_110_49_pad_groupi_n_209);
  or csa_tree_add_110_49_pad_groupi_g5293(csa_tree_add_110_49_pad_groupi_n_500 ,csa_tree_add_110_49_pad_groupi_n_404 ,csa_tree_add_110_49_pad_groupi_n_206);
  or csa_tree_add_110_49_pad_groupi_g5294(csa_tree_add_110_49_pad_groupi_n_499 ,csa_tree_add_110_49_pad_groupi_n_397 ,csa_tree_add_110_49_pad_groupi_n_203);
  or csa_tree_add_110_49_pad_groupi_g5295(csa_tree_add_110_49_pad_groupi_n_498 ,csa_tree_add_110_49_pad_groupi_n_458 ,csa_tree_add_110_49_pad_groupi_n_220);
  or csa_tree_add_110_49_pad_groupi_g5296(csa_tree_add_110_49_pad_groupi_n_497 ,csa_tree_add_110_49_pad_groupi_n_395 ,csa_tree_add_110_49_pad_groupi_n_230);
  or csa_tree_add_110_49_pad_groupi_g5297(csa_tree_add_110_49_pad_groupi_n_496 ,csa_tree_add_110_49_pad_groupi_n_449 ,csa_tree_add_110_49_pad_groupi_n_212);
  or csa_tree_add_110_49_pad_groupi_g5298(csa_tree_add_110_49_pad_groupi_n_495 ,csa_tree_add_110_49_pad_groupi_n_393 ,csa_tree_add_110_49_pad_groupi_n_200);
  or csa_tree_add_110_49_pad_groupi_g5299(csa_tree_add_110_49_pad_groupi_n_494 ,csa_tree_add_110_49_pad_groupi_n_396 ,csa_tree_add_110_49_pad_groupi_n_227);
  or csa_tree_add_110_49_pad_groupi_g5300(csa_tree_add_110_49_pad_groupi_n_493 ,csa_tree_add_110_49_pad_groupi_n_411 ,csa_tree_add_110_49_pad_groupi_n_221);
  or csa_tree_add_110_49_pad_groupi_g5301(csa_tree_add_110_49_pad_groupi_n_492 ,csa_tree_add_110_49_pad_groupi_n_455 ,csa_tree_add_110_49_pad_groupi_n_215);
  or csa_tree_add_110_49_pad_groupi_g5302(csa_tree_add_110_49_pad_groupi_n_491 ,csa_tree_add_110_49_pad_groupi_n_459 ,csa_tree_add_110_49_pad_groupi_n_224);
  or csa_tree_add_110_49_pad_groupi_g5303(csa_tree_add_110_49_pad_groupi_n_490 ,csa_tree_add_110_49_pad_groupi_n_392 ,csa_tree_add_110_49_pad_groupi_n_206);
  or csa_tree_add_110_49_pad_groupi_g5304(csa_tree_add_110_49_pad_groupi_n_489 ,csa_tree_add_110_49_pad_groupi_n_441 ,csa_tree_add_110_49_pad_groupi_n_218);
  or csa_tree_add_110_49_pad_groupi_g5305(csa_tree_add_110_49_pad_groupi_n_488 ,csa_tree_add_110_49_pad_groupi_n_417 ,csa_tree_add_110_49_pad_groupi_n_197);
  or csa_tree_add_110_49_pad_groupi_g5306(csa_tree_add_110_49_pad_groupi_n_487 ,csa_tree_add_110_49_pad_groupi_n_49 ,csa_tree_add_110_49_pad_groupi_n_470);
  nor csa_tree_add_110_49_pad_groupi_g5307(csa_tree_add_110_49_pad_groupi_n_486 ,csa_tree_add_110_49_pad_groupi_n_61 ,csa_tree_add_110_49_pad_groupi_n_467);
  or csa_tree_add_110_49_pad_groupi_g5308(csa_tree_add_110_49_pad_groupi_n_485 ,csa_tree_add_110_49_pad_groupi_n_72 ,csa_tree_add_110_49_pad_groupi_n_462);
  or csa_tree_add_110_49_pad_groupi_g5309(csa_tree_add_110_49_pad_groupi_n_484 ,csa_tree_add_110_49_pad_groupi_n_48 ,csa_tree_add_110_49_pad_groupi_n_466);
  or csa_tree_add_110_49_pad_groupi_g5310(csa_tree_add_110_49_pad_groupi_n_483 ,csa_tree_add_110_49_pad_groupi_n_51 ,csa_tree_add_110_49_pad_groupi_n_468);
  or csa_tree_add_110_49_pad_groupi_g5311(csa_tree_add_110_49_pad_groupi_n_482 ,csa_tree_add_110_49_pad_groupi_n_60 ,csa_tree_add_110_49_pad_groupi_n_461);
  or csa_tree_add_110_49_pad_groupi_g5312(csa_tree_add_110_49_pad_groupi_n_481 ,csa_tree_add_110_49_pad_groupi_n_11 ,csa_tree_add_110_49_pad_groupi_n_469);
  or csa_tree_add_110_49_pad_groupi_g5313(csa_tree_add_110_49_pad_groupi_n_480 ,csa_tree_add_110_49_pad_groupi_n_48 ,csa_tree_add_110_49_pad_groupi_n_463);
  or csa_tree_add_110_49_pad_groupi_g5314(csa_tree_add_110_49_pad_groupi_n_479 ,csa_tree_add_110_49_pad_groupi_n_51 ,csa_tree_add_110_49_pad_groupi_n_464);
  or csa_tree_add_110_49_pad_groupi_g5315(csa_tree_add_110_49_pad_groupi_n_478 ,csa_tree_add_110_49_pad_groupi_n_60 ,csa_tree_add_110_49_pad_groupi_n_465);
  or csa_tree_add_110_49_pad_groupi_g5316(csa_tree_add_110_49_pad_groupi_n_477 ,csa_tree_add_110_49_pad_groupi_n_72 ,csa_tree_add_110_49_pad_groupi_n_442);
  or csa_tree_add_110_49_pad_groupi_g5317(csa_tree_add_110_49_pad_groupi_n_476 ,csa_tree_add_110_49_pad_groupi_n_11 ,csa_tree_add_110_49_pad_groupi_n_472);
  or csa_tree_add_110_49_pad_groupi_g5318(csa_tree_add_110_49_pad_groupi_n_475 ,csa_tree_add_110_49_pad_groupi_n_61 ,csa_tree_add_110_49_pad_groupi_n_460);
  or csa_tree_add_110_49_pad_groupi_g5319(csa_tree_add_110_49_pad_groupi_n_474 ,csa_tree_add_110_49_pad_groupi_n_73 ,csa_tree_add_110_49_pad_groupi_n_471);
  or csa_tree_add_110_49_pad_groupi_g5320(csa_tree_add_110_49_pad_groupi_n_473 ,csa_tree_add_110_49_pad_groupi_n_446 ,csa_tree_add_110_49_pad_groupi_n_227);
  and csa_tree_add_110_49_pad_groupi_g5321(csa_tree_add_110_49_pad_groupi_n_527 ,in16[5] ,csa_tree_add_110_49_pad_groupi_n_145);
  and csa_tree_add_110_49_pad_groupi_g5322(csa_tree_add_110_49_pad_groupi_n_525 ,in16[3] ,csa_tree_add_110_49_pad_groupi_n_143);
  or csa_tree_add_110_49_pad_groupi_g5323(csa_tree_add_110_49_pad_groupi_n_524 ,csa_tree_add_110_49_pad_groupi_n_167 ,csa_tree_add_110_49_pad_groupi_n_212);
  and csa_tree_add_110_49_pad_groupi_g5324(csa_tree_add_110_49_pad_groupi_n_522 ,in16[7] ,csa_tree_add_110_49_pad_groupi_n_140);
  or csa_tree_add_110_49_pad_groupi_g5325(csa_tree_add_110_49_pad_groupi_n_521 ,csa_tree_add_110_49_pad_groupi_n_176 ,csa_tree_add_110_49_pad_groupi_n_224);
  or csa_tree_add_110_49_pad_groupi_g5326(csa_tree_add_110_49_pad_groupi_n_520 ,csa_tree_add_110_49_pad_groupi_n_166 ,csa_tree_add_110_49_pad_groupi_n_230);
  or csa_tree_add_110_49_pad_groupi_g5327(csa_tree_add_110_49_pad_groupi_n_519 ,csa_tree_add_110_49_pad_groupi_n_337 ,csa_tree_add_110_49_pad_groupi_n_427);
  or csa_tree_add_110_49_pad_groupi_g5328(csa_tree_add_110_49_pad_groupi_n_517 ,csa_tree_add_110_49_pad_groupi_n_340 ,csa_tree_add_110_49_pad_groupi_n_430);
  or csa_tree_add_110_49_pad_groupi_g5329(csa_tree_add_110_49_pad_groupi_n_515 ,csa_tree_add_110_49_pad_groupi_n_175 ,csa_tree_add_110_49_pad_groupi_n_389);
  or csa_tree_add_110_49_pad_groupi_g5330(csa_tree_add_110_49_pad_groupi_n_512 ,csa_tree_add_110_49_pad_groupi_n_300 ,csa_tree_add_110_49_pad_groupi_n_163);
  or csa_tree_add_110_49_pad_groupi_g5331(csa_tree_add_110_49_pad_groupi_n_511 ,csa_tree_add_110_49_pad_groupi_n_384 ,csa_tree_add_110_49_pad_groupi_n_142);
  or csa_tree_add_110_49_pad_groupi_g5332(csa_tree_add_110_49_pad_groupi_n_510 ,csa_tree_add_110_49_pad_groupi_n_434 ,csa_tree_add_110_49_pad_groupi_n_144);
  not csa_tree_add_110_49_pad_groupi_g5333(csa_tree_add_110_49_pad_groupi_n_440 ,csa_tree_add_110_49_pad_groupi_n_145);
  not csa_tree_add_110_49_pad_groupi_g5334(csa_tree_add_110_49_pad_groupi_n_439 ,csa_tree_add_110_49_pad_groupi_n_144);
  not csa_tree_add_110_49_pad_groupi_g5337(csa_tree_add_110_49_pad_groupi_n_437 ,csa_tree_add_110_49_pad_groupi_n_143);
  not csa_tree_add_110_49_pad_groupi_g5338(csa_tree_add_110_49_pad_groupi_n_436 ,csa_tree_add_110_49_pad_groupi_n_142);
  xnor csa_tree_add_110_49_pad_groupi_g5341(csa_tree_add_110_49_pad_groupi_n_434 ,in16[5] ,in16[4]);
  and csa_tree_add_110_49_pad_groupi_g5342(csa_tree_add_110_49_pad_groupi_n_433 ,n_175 ,csa_tree_add_110_49_pad_groupi_n_336);
  and csa_tree_add_110_49_pad_groupi_g5343(csa_tree_add_110_49_pad_groupi_n_432 ,n_144 ,csa_tree_add_110_49_pad_groupi_n_354);
  and csa_tree_add_110_49_pad_groupi_g5344(csa_tree_add_110_49_pad_groupi_n_431 ,n_145 ,csa_tree_add_110_49_pad_groupi_n_360);
  and csa_tree_add_110_49_pad_groupi_g5345(csa_tree_add_110_49_pad_groupi_n_430 ,n_154 ,csa_tree_add_110_49_pad_groupi_n_359);
  and csa_tree_add_110_49_pad_groupi_g5346(csa_tree_add_110_49_pad_groupi_n_429 ,n_188 ,csa_tree_add_110_49_pad_groupi_n_319);
  and csa_tree_add_110_49_pad_groupi_g5347(csa_tree_add_110_49_pad_groupi_n_428 ,n_147 ,csa_tree_add_110_49_pad_groupi_n_317);
  and csa_tree_add_110_49_pad_groupi_g5348(csa_tree_add_110_49_pad_groupi_n_427 ,n_146 ,csa_tree_add_110_49_pad_groupi_n_347);
  and csa_tree_add_110_49_pad_groupi_g5349(csa_tree_add_110_49_pad_groupi_n_426 ,csa_tree_add_110_49_pad_groupi_n_289 ,csa_tree_add_110_49_pad_groupi_n_329);
  and csa_tree_add_110_49_pad_groupi_g5350(csa_tree_add_110_49_pad_groupi_n_425 ,csa_tree_add_110_49_pad_groupi_n_290 ,csa_tree_add_110_49_pad_groupi_n_344);
  and csa_tree_add_110_49_pad_groupi_g5351(csa_tree_add_110_49_pad_groupi_n_424 ,csa_tree_add_110_49_pad_groupi_n_291 ,csa_tree_add_110_49_pad_groupi_n_348);
  and csa_tree_add_110_49_pad_groupi_g5352(csa_tree_add_110_49_pad_groupi_n_423 ,n_155 ,csa_tree_add_110_49_pad_groupi_n_342);
  xnor csa_tree_add_110_49_pad_groupi_g5353(csa_tree_add_110_49_pad_groupi_n_422 ,csa_tree_add_110_49_pad_groupi_n_169 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5356(csa_tree_add_110_49_pad_groupi_n_472 ,csa_tree_add_110_49_pad_groupi_n_259 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5357(csa_tree_add_110_49_pad_groupi_n_471 ,csa_tree_add_110_49_pad_groupi_n_250 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5358(csa_tree_add_110_49_pad_groupi_n_470 ,csa_tree_add_110_49_pad_groupi_n_262 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5359(csa_tree_add_110_49_pad_groupi_n_469 ,csa_tree_add_110_49_pad_groupi_n_265 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5360(csa_tree_add_110_49_pad_groupi_n_468 ,csa_tree_add_110_49_pad_groupi_n_247 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5362(csa_tree_add_110_49_pad_groupi_n_466 ,csa_tree_add_110_49_pad_groupi_n_244 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5363(csa_tree_add_110_49_pad_groupi_n_465 ,csa_tree_add_110_49_pad_groupi_n_238 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5364(csa_tree_add_110_49_pad_groupi_n_464 ,csa_tree_add_110_49_pad_groupi_n_271 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5365(csa_tree_add_110_49_pad_groupi_n_463 ,csa_tree_add_110_49_pad_groupi_n_232 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5366(csa_tree_add_110_49_pad_groupi_n_462 ,csa_tree_add_110_49_pad_groupi_n_274 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5367(csa_tree_add_110_49_pad_groupi_n_461 ,csa_tree_add_110_49_pad_groupi_n_241 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5368(csa_tree_add_110_49_pad_groupi_n_460 ,csa_tree_add_110_49_pad_groupi_n_268 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5369(csa_tree_add_110_49_pad_groupi_n_459 ,csa_tree_add_110_49_pad_groupi_n_266 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5370(csa_tree_add_110_49_pad_groupi_n_458 ,csa_tree_add_110_49_pad_groupi_n_269 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5371(csa_tree_add_110_49_pad_groupi_n_457 ,csa_tree_add_110_49_pad_groupi_n_109 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5372(csa_tree_add_110_49_pad_groupi_n_456 ,csa_tree_add_110_49_pad_groupi_n_239 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5373(csa_tree_add_110_49_pad_groupi_n_455 ,csa_tree_add_110_49_pad_groupi_n_253 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5374(csa_tree_add_110_49_pad_groupi_n_454 ,csa_tree_add_110_49_pad_groupi_n_105 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5375(csa_tree_add_110_49_pad_groupi_n_453 ,csa_tree_add_110_49_pad_groupi_n_245 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5376(csa_tree_add_110_49_pad_groupi_n_452 ,csa_tree_add_110_49_pad_groupi_n_256 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5377(csa_tree_add_110_49_pad_groupi_n_451 ,csa_tree_add_110_49_pad_groupi_n_260 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5378(csa_tree_add_110_49_pad_groupi_n_450 ,csa_tree_add_110_49_pad_groupi_n_254 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5379(csa_tree_add_110_49_pad_groupi_n_449 ,csa_tree_add_110_49_pad_groupi_n_232 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5380(csa_tree_add_110_49_pad_groupi_n_448 ,csa_tree_add_110_49_pad_groupi_n_123 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5381(csa_tree_add_110_49_pad_groupi_n_447 ,csa_tree_add_110_49_pad_groupi_n_251 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5382(csa_tree_add_110_49_pad_groupi_n_446 ,csa_tree_add_110_49_pad_groupi_n_242 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5383(csa_tree_add_110_49_pad_groupi_n_445 ,csa_tree_add_110_49_pad_groupi_n_115 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5384(csa_tree_add_110_49_pad_groupi_n_444 ,csa_tree_add_110_49_pad_groupi_n_99 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5385(csa_tree_add_110_49_pad_groupi_n_443 ,csa_tree_add_110_49_pad_groupi_n_275 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5386(csa_tree_add_110_49_pad_groupi_n_442 ,csa_tree_add_110_49_pad_groupi_n_257 ,in16[1]);
  xnor csa_tree_add_110_49_pad_groupi_g5387(csa_tree_add_110_49_pad_groupi_n_441 ,csa_tree_add_110_49_pad_groupi_n_248 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5388(csa_tree_add_110_49_pad_groupi_n_438 ,csa_tree_add_110_49_pad_groupi_n_192 ,in16[4]);
  xnor csa_tree_add_110_49_pad_groupi_g5389(csa_tree_add_110_49_pad_groupi_n_435 ,csa_tree_add_110_49_pad_groupi_n_194 ,in16[2]);
  not csa_tree_add_110_49_pad_groupi_g5390(csa_tree_add_110_49_pad_groupi_n_391 ,csa_tree_add_110_49_pad_groupi_n_389);
  not csa_tree_add_110_49_pad_groupi_g5391(csa_tree_add_110_49_pad_groupi_n_390 ,csa_tree_add_110_49_pad_groupi_n_389);
  not csa_tree_add_110_49_pad_groupi_g5392(csa_tree_add_110_49_pad_groupi_n_388 ,csa_tree_add_110_49_pad_groupi_n_141);
  not csa_tree_add_110_49_pad_groupi_g5393(csa_tree_add_110_49_pad_groupi_n_387 ,csa_tree_add_110_49_pad_groupi_n_140);
  xnor csa_tree_add_110_49_pad_groupi_g5396(csa_tree_add_110_49_pad_groupi_n_385 ,csa_tree_add_110_49_pad_groupi_n_172 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5397(csa_tree_add_110_49_pad_groupi_n_384 ,in16[3] ,in16[2]);
  xnor csa_tree_add_110_49_pad_groupi_g5398(csa_tree_add_110_49_pad_groupi_n_383 ,in16[7] ,in16[6]);
  xnor csa_tree_add_110_49_pad_groupi_g5399(csa_tree_add_110_49_pad_groupi_n_382 ,csa_tree_add_110_49_pad_groupi_n_170 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5400(csa_tree_add_110_49_pad_groupi_n_419 ,csa_tree_add_110_49_pad_groupi_n_113 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5401(csa_tree_add_110_49_pad_groupi_n_418 ,csa_tree_add_110_49_pad_groupi_n_85 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5402(csa_tree_add_110_49_pad_groupi_n_417 ,csa_tree_add_110_49_pad_groupi_n_272 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5403(csa_tree_add_110_49_pad_groupi_n_416 ,csa_tree_add_110_49_pad_groupi_n_263 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5404(csa_tree_add_110_49_pad_groupi_n_415 ,csa_tree_add_110_49_pad_groupi_n_129 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5405(csa_tree_add_110_49_pad_groupi_n_414 ,csa_tree_add_110_49_pad_groupi_n_79 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5406(csa_tree_add_110_49_pad_groupi_n_413 ,csa_tree_add_110_49_pad_groupi_n_131 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5407(csa_tree_add_110_49_pad_groupi_n_412 ,csa_tree_add_110_49_pad_groupi_n_236 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5408(csa_tree_add_110_49_pad_groupi_n_411 ,csa_tree_add_110_49_pad_groupi_n_101 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5409(csa_tree_add_110_49_pad_groupi_n_410 ,csa_tree_add_110_49_pad_groupi_n_91 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5410(csa_tree_add_110_49_pad_groupi_n_409 ,csa_tree_add_110_49_pad_groupi_n_127 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5411(csa_tree_add_110_49_pad_groupi_n_408 ,csa_tree_add_110_49_pad_groupi_n_101 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5412(csa_tree_add_110_49_pad_groupi_n_407 ,csa_tree_add_110_49_pad_groupi_n_103 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5413(csa_tree_add_110_49_pad_groupi_n_406 ,csa_tree_add_110_49_pad_groupi_n_103 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5414(csa_tree_add_110_49_pad_groupi_n_405 ,csa_tree_add_110_49_pad_groupi_n_115 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5415(csa_tree_add_110_49_pad_groupi_n_404 ,csa_tree_add_110_49_pad_groupi_n_129 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5416(csa_tree_add_110_49_pad_groupi_n_403 ,csa_tree_add_110_49_pad_groupi_n_127 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5417(csa_tree_add_110_49_pad_groupi_n_402 ,csa_tree_add_110_49_pad_groupi_n_109 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5418(csa_tree_add_110_49_pad_groupi_n_401 ,csa_tree_add_110_49_pad_groupi_n_131 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5419(csa_tree_add_110_49_pad_groupi_n_400 ,csa_tree_add_110_49_pad_groupi_n_91 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5420(csa_tree_add_110_49_pad_groupi_n_399 ,csa_tree_add_110_49_pad_groupi_n_113 ,in16[3]);
  xnor csa_tree_add_110_49_pad_groupi_g5421(csa_tree_add_110_49_pad_groupi_n_398 ,csa_tree_add_110_49_pad_groupi_n_105 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5422(csa_tree_add_110_49_pad_groupi_n_397 ,csa_tree_add_110_49_pad_groupi_n_121 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5423(csa_tree_add_110_49_pad_groupi_n_396 ,csa_tree_add_110_49_pad_groupi_n_121 ,in16[5]);
  xnor csa_tree_add_110_49_pad_groupi_g5424(csa_tree_add_110_49_pad_groupi_n_381 ,n_244 ,n_148);
  xnor csa_tree_add_110_49_pad_groupi_g5425(csa_tree_add_110_49_pad_groupi_n_395 ,csa_tree_add_110_49_pad_groupi_n_99 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5426(csa_tree_add_110_49_pad_groupi_n_394 ,csa_tree_add_110_49_pad_groupi_n_123 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5427(csa_tree_add_110_49_pad_groupi_n_393 ,csa_tree_add_110_49_pad_groupi_n_79 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5428(csa_tree_add_110_49_pad_groupi_n_392 ,csa_tree_add_110_49_pad_groupi_n_85 ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5429(csa_tree_add_110_49_pad_groupi_n_380 ,n_240 ,n_208);
  xnor csa_tree_add_110_49_pad_groupi_g5430(csa_tree_add_110_49_pad_groupi_n_379 ,n_211 ,n_147);
  xnor csa_tree_add_110_49_pad_groupi_g5431(csa_tree_add_110_49_pad_groupi_n_378 ,n_183 ,n_151);
  xnor csa_tree_add_110_49_pad_groupi_g5432(csa_tree_add_110_49_pad_groupi_n_377 ,n_254 ,n_222);
  xnor csa_tree_add_110_49_pad_groupi_g5433(csa_tree_add_110_49_pad_groupi_n_376 ,n_220 ,n_188);
  xnor csa_tree_add_110_49_pad_groupi_g5434(csa_tree_add_110_49_pad_groupi_n_375 ,n_190 ,n_158);
  xnor csa_tree_add_110_49_pad_groupi_g5435(csa_tree_add_110_49_pad_groupi_n_374 ,n_241 ,n_145);
  xnor csa_tree_add_110_49_pad_groupi_g5436(csa_tree_add_110_49_pad_groupi_n_373 ,n_251 ,n_219);
  xnor csa_tree_add_110_49_pad_groupi_g5437(csa_tree_add_110_49_pad_groupi_n_372 ,n_210 ,n_178);
  xnor csa_tree_add_110_49_pad_groupi_g5438(csa_tree_add_110_49_pad_groupi_n_371 ,n_250 ,n_154);
  xnor csa_tree_add_110_49_pad_groupi_g5439(csa_tree_add_110_49_pad_groupi_n_370 ,n_245 ,n_149);
  xnor csa_tree_add_110_49_pad_groupi_g5440(csa_tree_add_110_49_pad_groupi_n_369 ,n_221 ,n_189);
  xnor csa_tree_add_110_49_pad_groupi_g5441(csa_tree_add_110_49_pad_groupi_n_368 ,n_216 ,n_184);
  xnor csa_tree_add_110_49_pad_groupi_g5442(csa_tree_add_110_49_pad_groupi_n_367 ,n_239 ,n_207);
  xnor csa_tree_add_110_49_pad_groupi_g5443(csa_tree_add_110_49_pad_groupi_n_366 ,n_246 ,n_150);
  xnor csa_tree_add_110_49_pad_groupi_g5444(csa_tree_add_110_49_pad_groupi_n_389 ,in16[8] ,in16[7]);
  xnor csa_tree_add_110_49_pad_groupi_g5445(csa_tree_add_110_49_pad_groupi_n_386 ,csa_tree_add_110_49_pad_groupi_n_190 ,in16[6]);
  nor csa_tree_add_110_49_pad_groupi_g5446(csa_tree_add_110_49_pad_groupi_n_365 ,n_245 ,n_149);
  and csa_tree_add_110_49_pad_groupi_g5447(csa_tree_add_110_49_pad_groupi_n_364 ,n_241 ,n_177);
  nor csa_tree_add_110_49_pad_groupi_g5448(csa_tree_add_110_49_pad_groupi_n_363 ,n_244 ,n_148);
  and csa_tree_add_110_49_pad_groupi_g5449(csa_tree_add_110_49_pad_groupi_n_362 ,n_251 ,n_219);
  nor csa_tree_add_110_49_pad_groupi_g5450(csa_tree_add_110_49_pad_groupi_n_361 ,n_249 ,n_217);
  or csa_tree_add_110_49_pad_groupi_g5451(csa_tree_add_110_49_pad_groupi_n_360 ,n_241 ,n_177);
  or csa_tree_add_110_49_pad_groupi_g5452(csa_tree_add_110_49_pad_groupi_n_359 ,n_250 ,n_186);
  nor csa_tree_add_110_49_pad_groupi_g5453(csa_tree_add_110_49_pad_groupi_n_358 ,n_221 ,n_189);
  or csa_tree_add_110_49_pad_groupi_g5454(csa_tree_add_110_49_pad_groupi_n_357 ,n_212 ,n_180);
  and csa_tree_add_110_49_pad_groupi_g5455(csa_tree_add_110_49_pad_groupi_n_356 ,n_252 ,n_220);
  nor csa_tree_add_110_49_pad_groupi_g5456(csa_tree_add_110_49_pad_groupi_n_355 ,csa_tree_add_110_49_pad_groupi_n_172 ,in16[6]);
  or csa_tree_add_110_49_pad_groupi_g5457(csa_tree_add_110_49_pad_groupi_n_354 ,n_240 ,n_208);
  and csa_tree_add_110_49_pad_groupi_g5458(csa_tree_add_110_49_pad_groupi_n_353 ,n_214 ,n_182);
  or csa_tree_add_110_49_pad_groupi_g5459(csa_tree_add_110_49_pad_groupi_n_352 ,n_214 ,n_182);
  nor csa_tree_add_110_49_pad_groupi_g5460(csa_tree_add_110_49_pad_groupi_n_351 ,csa_tree_add_110_49_pad_groupi_n_169 ,in16[4]);
  nor csa_tree_add_110_49_pad_groupi_g5461(csa_tree_add_110_49_pad_groupi_n_350 ,n_248 ,n_152);
  and csa_tree_add_110_49_pad_groupi_g5462(csa_tree_add_110_49_pad_groupi_n_349 ,n_240 ,n_208);
  or csa_tree_add_110_49_pad_groupi_g5463(csa_tree_add_110_49_pad_groupi_n_348 ,csa_tree_add_110_49_pad_groupi_n_166 ,csa_tree_add_110_49_pad_groupi_n_302);
  or csa_tree_add_110_49_pad_groupi_g5464(csa_tree_add_110_49_pad_groupi_n_347 ,n_210 ,n_178);
  and csa_tree_add_110_49_pad_groupi_g5465(csa_tree_add_110_49_pad_groupi_n_346 ,n_247 ,n_215);
  and csa_tree_add_110_49_pad_groupi_g5466(csa_tree_add_110_49_pad_groupi_n_345 ,n_253 ,n_157);
  or csa_tree_add_110_49_pad_groupi_g5467(csa_tree_add_110_49_pad_groupi_n_344 ,csa_tree_add_110_49_pad_groupi_n_13 ,csa_tree_add_110_49_pad_groupi_n_303);
  or csa_tree_add_110_49_pad_groupi_g5468(csa_tree_add_110_49_pad_groupi_n_343 ,n_183 ,n_151);
  or csa_tree_add_110_49_pad_groupi_g5469(csa_tree_add_110_49_pad_groupi_n_342 ,n_251 ,n_219);
  and csa_tree_add_110_49_pad_groupi_g5470(csa_tree_add_110_49_pad_groupi_n_341 ,n_246 ,n_150);
  and csa_tree_add_110_49_pad_groupi_g5471(csa_tree_add_110_49_pad_groupi_n_340 ,n_250 ,n_186);
  or csa_tree_add_110_49_pad_groupi_g5472(csa_tree_add_110_49_pad_groupi_n_339 ,n_213 ,n_181);
  and csa_tree_add_110_49_pad_groupi_g5473(csa_tree_add_110_49_pad_groupi_n_338 ,n_212 ,n_180);
  and csa_tree_add_110_49_pad_groupi_g5474(csa_tree_add_110_49_pad_groupi_n_337 ,n_210 ,n_178);
  or csa_tree_add_110_49_pad_groupi_g5475(csa_tree_add_110_49_pad_groupi_n_336 ,n_239 ,n_207);
  nor csa_tree_add_110_49_pad_groupi_g5476(csa_tree_add_110_49_pad_groupi_n_335 ,n_185 ,n_153);
  or csa_tree_add_110_49_pad_groupi_g5477(csa_tree_add_110_49_pad_groupi_n_334 ,csa_tree_add_110_49_pad_groupi_n_296 ,csa_tree_add_110_49_pad_groupi_n_309);
  and csa_tree_add_110_49_pad_groupi_g5478(csa_tree_add_110_49_pad_groupi_n_333 ,n_183 ,n_151);
  nor csa_tree_add_110_49_pad_groupi_g5479(csa_tree_add_110_49_pad_groupi_n_332 ,csa_tree_add_110_49_pad_groupi_n_173 ,in16[2]);
  or csa_tree_add_110_49_pad_groupi_g5480(csa_tree_add_110_49_pad_groupi_n_331 ,csa_tree_add_110_49_pad_groupi_n_295 ,csa_tree_add_110_49_pad_groupi_n_299);
  and csa_tree_add_110_49_pad_groupi_g5481(csa_tree_add_110_49_pad_groupi_n_330 ,n_245 ,n_149);
  or csa_tree_add_110_49_pad_groupi_g5482(csa_tree_add_110_49_pad_groupi_n_329 ,csa_tree_add_110_49_pad_groupi_n_13 ,csa_tree_add_110_49_pad_groupi_n_304);
  and csa_tree_add_110_49_pad_groupi_g5483(csa_tree_add_110_49_pad_groupi_n_328 ,n_213 ,n_181);
  nor csa_tree_add_110_49_pad_groupi_g5484(csa_tree_add_110_49_pad_groupi_n_327 ,csa_tree_add_110_49_pad_groupi_n_52 ,csa_tree_add_110_49_pad_groupi_n_289);
  nor csa_tree_add_110_49_pad_groupi_g5485(csa_tree_add_110_49_pad_groupi_n_326 ,n_216 ,n_184);
  or csa_tree_add_110_49_pad_groupi_g5486(csa_tree_add_110_49_pad_groupi_n_325 ,csa_tree_add_110_49_pad_groupi_n_312 ,csa_tree_add_110_49_pad_groupi_n_294);
  or csa_tree_add_110_49_pad_groupi_g5487(csa_tree_add_110_49_pad_groupi_n_324 ,csa_tree_add_110_49_pad_groupi_n_313 ,csa_tree_add_110_49_pad_groupi_n_311);
  or csa_tree_add_110_49_pad_groupi_g5488(csa_tree_add_110_49_pad_groupi_n_323 ,csa_tree_add_110_49_pad_groupi_n_297 ,csa_tree_add_110_49_pad_groupi_n_308);
  nor csa_tree_add_110_49_pad_groupi_g5489(csa_tree_add_110_49_pad_groupi_n_322 ,csa_tree_add_110_49_pad_groupi_n_49 ,csa_tree_add_110_49_pad_groupi_n_167);
  and csa_tree_add_110_49_pad_groupi_g5490(csa_tree_add_110_49_pad_groupi_n_321 ,n_239 ,n_207);
  or csa_tree_add_110_49_pad_groupi_g5491(csa_tree_add_110_49_pad_groupi_n_320 ,n_253 ,n_157);
  or csa_tree_add_110_49_pad_groupi_g5492(csa_tree_add_110_49_pad_groupi_n_319 ,n_252 ,n_220);
  or csa_tree_add_110_49_pad_groupi_g5493(csa_tree_add_110_49_pad_groupi_n_318 ,n_247 ,n_215);
  or csa_tree_add_110_49_pad_groupi_g5494(csa_tree_add_110_49_pad_groupi_n_317 ,n_243 ,n_211);
  and csa_tree_add_110_49_pad_groupi_g5495(csa_tree_add_110_49_pad_groupi_n_316 ,n_221 ,n_189);
  and csa_tree_add_110_49_pad_groupi_g5496(csa_tree_add_110_49_pad_groupi_n_315 ,n_243 ,n_211);
  nor csa_tree_add_110_49_pad_groupi_g5497(csa_tree_add_110_49_pad_groupi_n_314 ,n_246 ,n_150);
  not csa_tree_add_110_49_pad_groupi_g5498(csa_tree_add_110_49_pad_groupi_n_313 ,n_244);
  not csa_tree_add_110_49_pad_groupi_g5499(csa_tree_add_110_49_pad_groupi_n_312 ,n_185);
  not csa_tree_add_110_49_pad_groupi_g5500(csa_tree_add_110_49_pad_groupi_n_311 ,n_148);
  not csa_tree_add_110_49_pad_groupi_g5501(csa_tree_add_110_49_pad_groupi_n_310 ,n_156);
  not csa_tree_add_110_49_pad_groupi_g5502(csa_tree_add_110_49_pad_groupi_n_309 ,n_152);
  not csa_tree_add_110_49_pad_groupi_g5503(csa_tree_add_110_49_pad_groupi_n_308 ,n_184);
  not csa_tree_add_110_49_pad_groupi_g5504(csa_tree_add_110_49_pad_groupi_n_307 ,n_176);
  not csa_tree_add_110_49_pad_groupi_g5505(csa_tree_add_110_49_pad_groupi_n_306 ,n_242);
  not csa_tree_add_110_49_pad_groupi_g5506(csa_tree_add_110_49_pad_groupi_n_305 ,n_209);
  not csa_tree_add_110_49_pad_groupi_g5507(csa_tree_add_110_49_pad_groupi_n_304 ,in16[2]);
  not csa_tree_add_110_49_pad_groupi_g5508(csa_tree_add_110_49_pad_groupi_n_303 ,in16[6]);
  not csa_tree_add_110_49_pad_groupi_g5509(csa_tree_add_110_49_pad_groupi_n_302 ,in16[4]);
  not csa_tree_add_110_49_pad_groupi_g5510(csa_tree_add_110_49_pad_groupi_n_301 ,csa_tree_add_110_49_pad_groupi_n_170);
  not csa_tree_add_110_49_pad_groupi_g5511(csa_tree_add_110_49_pad_groupi_n_300 ,in16[8]);
  not csa_tree_add_110_49_pad_groupi_g5512(csa_tree_add_110_49_pad_groupi_n_299 ,n_217);
  not csa_tree_add_110_49_pad_groupi_g5513(csa_tree_add_110_49_pad_groupi_n_298 ,n_143);
  not csa_tree_add_110_49_pad_groupi_g5514(csa_tree_add_110_49_pad_groupi_n_297 ,n_216);
  not csa_tree_add_110_49_pad_groupi_g5515(csa_tree_add_110_49_pad_groupi_n_296 ,n_248);
  not csa_tree_add_110_49_pad_groupi_g5516(csa_tree_add_110_49_pad_groupi_n_295 ,n_249);
  not csa_tree_add_110_49_pad_groupi_g5517(csa_tree_add_110_49_pad_groupi_n_294 ,n_153);
  not csa_tree_add_110_49_pad_groupi_g5518(csa_tree_add_110_49_pad_groupi_n_293 ,in16[0]);
  not csa_tree_add_110_49_pad_groupi_g5519(csa_tree_add_110_49_pad_groupi_n_292 ,in16[7]);
  not csa_tree_add_110_49_pad_groupi_g5520(csa_tree_add_110_49_pad_groupi_n_291 ,in16[3]);
  not csa_tree_add_110_49_pad_groupi_g5521(csa_tree_add_110_49_pad_groupi_n_290 ,in16[5]);
  not csa_tree_add_110_49_pad_groupi_g5522(csa_tree_add_110_49_pad_groupi_n_289 ,in16[1]);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5577(csa_tree_add_110_49_pad_groupi_n_277 ,csa_tree_add_110_49_pad_groupi_n_276);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5579(csa_tree_add_110_49_pad_groupi_n_276 ,n_271);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5602(csa_tree_add_110_49_pad_groupi_n_275 ,csa_tree_add_110_49_pad_groupi_n_273);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5603(csa_tree_add_110_49_pad_groupi_n_274 ,csa_tree_add_110_49_pad_groupi_n_273);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5604(csa_tree_add_110_49_pad_groupi_n_273 ,n_285);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5606(csa_tree_add_110_49_pad_groupi_n_272 ,csa_tree_add_110_49_pad_groupi_n_270);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5607(csa_tree_add_110_49_pad_groupi_n_271 ,csa_tree_add_110_49_pad_groupi_n_270);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5608(csa_tree_add_110_49_pad_groupi_n_270 ,n_279);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5610(csa_tree_add_110_49_pad_groupi_n_269 ,csa_tree_add_110_49_pad_groupi_n_267);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5611(csa_tree_add_110_49_pad_groupi_n_268 ,csa_tree_add_110_49_pad_groupi_n_267);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5612(csa_tree_add_110_49_pad_groupi_n_267 ,n_283);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5614(csa_tree_add_110_49_pad_groupi_n_266 ,csa_tree_add_110_49_pad_groupi_n_264);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5615(csa_tree_add_110_49_pad_groupi_n_265 ,csa_tree_add_110_49_pad_groupi_n_264);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5616(csa_tree_add_110_49_pad_groupi_n_264 ,n_278);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5618(csa_tree_add_110_49_pad_groupi_n_263 ,csa_tree_add_110_49_pad_groupi_n_261);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5619(csa_tree_add_110_49_pad_groupi_n_262 ,csa_tree_add_110_49_pad_groupi_n_261);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5620(csa_tree_add_110_49_pad_groupi_n_261 ,n_282);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5622(csa_tree_add_110_49_pad_groupi_n_260 ,csa_tree_add_110_49_pad_groupi_n_258);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5623(csa_tree_add_110_49_pad_groupi_n_259 ,csa_tree_add_110_49_pad_groupi_n_258);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5624(csa_tree_add_110_49_pad_groupi_n_258 ,n_277);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5626(csa_tree_add_110_49_pad_groupi_n_257 ,csa_tree_add_110_49_pad_groupi_n_255);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5627(csa_tree_add_110_49_pad_groupi_n_256 ,csa_tree_add_110_49_pad_groupi_n_255);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5628(csa_tree_add_110_49_pad_groupi_n_255 ,n_276);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5630(csa_tree_add_110_49_pad_groupi_n_254 ,csa_tree_add_110_49_pad_groupi_n_252);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5631(csa_tree_add_110_49_pad_groupi_n_253 ,csa_tree_add_110_49_pad_groupi_n_252);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5632(csa_tree_add_110_49_pad_groupi_n_252 ,n_284);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5634(csa_tree_add_110_49_pad_groupi_n_251 ,csa_tree_add_110_49_pad_groupi_n_249);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5635(csa_tree_add_110_49_pad_groupi_n_250 ,csa_tree_add_110_49_pad_groupi_n_249);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5636(csa_tree_add_110_49_pad_groupi_n_249 ,n_275);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5638(csa_tree_add_110_49_pad_groupi_n_248 ,csa_tree_add_110_49_pad_groupi_n_246);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5639(csa_tree_add_110_49_pad_groupi_n_247 ,csa_tree_add_110_49_pad_groupi_n_246);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5640(csa_tree_add_110_49_pad_groupi_n_246 ,n_281);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5642(csa_tree_add_110_49_pad_groupi_n_245 ,csa_tree_add_110_49_pad_groupi_n_243);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5643(csa_tree_add_110_49_pad_groupi_n_244 ,csa_tree_add_110_49_pad_groupi_n_243);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5644(csa_tree_add_110_49_pad_groupi_n_243 ,n_274);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5646(csa_tree_add_110_49_pad_groupi_n_242 ,csa_tree_add_110_49_pad_groupi_n_240);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5647(csa_tree_add_110_49_pad_groupi_n_241 ,csa_tree_add_110_49_pad_groupi_n_240);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5648(csa_tree_add_110_49_pad_groupi_n_240 ,n_273);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5650(csa_tree_add_110_49_pad_groupi_n_239 ,csa_tree_add_110_49_pad_groupi_n_237);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5651(csa_tree_add_110_49_pad_groupi_n_238 ,csa_tree_add_110_49_pad_groupi_n_237);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5652(csa_tree_add_110_49_pad_groupi_n_237 ,n_280);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5654(csa_tree_add_110_49_pad_groupi_n_236 ,csa_tree_add_110_49_pad_groupi_n_234);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5655(csa_tree_add_110_49_pad_groupi_n_235 ,csa_tree_add_110_49_pad_groupi_n_234);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5656(csa_tree_add_110_49_pad_groupi_n_234 ,n_272);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5658(csa_tree_add_110_49_pad_groupi_n_233 ,csa_tree_add_110_49_pad_groupi_n_231);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5659(csa_tree_add_110_49_pad_groupi_n_232 ,csa_tree_add_110_49_pad_groupi_n_231);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5660(csa_tree_add_110_49_pad_groupi_n_231 ,n_286);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5662(csa_tree_add_110_49_pad_groupi_n_230 ,csa_tree_add_110_49_pad_groupi_n_228);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5663(csa_tree_add_110_49_pad_groupi_n_229 ,csa_tree_add_110_49_pad_groupi_n_228);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5664(csa_tree_add_110_49_pad_groupi_n_228 ,csa_tree_add_110_49_pad_groupi_n_387);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5666(csa_tree_add_110_49_pad_groupi_n_227 ,csa_tree_add_110_49_pad_groupi_n_225);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5667(csa_tree_add_110_49_pad_groupi_n_226 ,csa_tree_add_110_49_pad_groupi_n_225);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5668(csa_tree_add_110_49_pad_groupi_n_225 ,csa_tree_add_110_49_pad_groupi_n_440);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5670(csa_tree_add_110_49_pad_groupi_n_224 ,csa_tree_add_110_49_pad_groupi_n_222);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5671(csa_tree_add_110_49_pad_groupi_n_223 ,csa_tree_add_110_49_pad_groupi_n_222);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5672(csa_tree_add_110_49_pad_groupi_n_222 ,csa_tree_add_110_49_pad_groupi_n_439);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5674(csa_tree_add_110_49_pad_groupi_n_221 ,csa_tree_add_110_49_pad_groupi_n_219);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5675(csa_tree_add_110_49_pad_groupi_n_220 ,csa_tree_add_110_49_pad_groupi_n_219);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5676(csa_tree_add_110_49_pad_groupi_n_219 ,csa_tree_add_110_49_pad_groupi_n_283);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5678(csa_tree_add_110_49_pad_groupi_n_218 ,csa_tree_add_110_49_pad_groupi_n_216);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5679(csa_tree_add_110_49_pad_groupi_n_217 ,csa_tree_add_110_49_pad_groupi_n_216);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5680(csa_tree_add_110_49_pad_groupi_n_216 ,csa_tree_add_110_49_pad_groupi_n_282);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5682(csa_tree_add_110_49_pad_groupi_n_215 ,csa_tree_add_110_49_pad_groupi_n_213);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5683(csa_tree_add_110_49_pad_groupi_n_214 ,csa_tree_add_110_49_pad_groupi_n_213);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5684(csa_tree_add_110_49_pad_groupi_n_213 ,csa_tree_add_110_49_pad_groupi_n_280);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5686(csa_tree_add_110_49_pad_groupi_n_212 ,csa_tree_add_110_49_pad_groupi_n_210);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5687(csa_tree_add_110_49_pad_groupi_n_211 ,csa_tree_add_110_49_pad_groupi_n_210);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5688(csa_tree_add_110_49_pad_groupi_n_210 ,csa_tree_add_110_49_pad_groupi_n_436);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5690(csa_tree_add_110_49_pad_groupi_n_209 ,csa_tree_add_110_49_pad_groupi_n_207);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5691(csa_tree_add_110_49_pad_groupi_n_208 ,csa_tree_add_110_49_pad_groupi_n_207);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5692(csa_tree_add_110_49_pad_groupi_n_207 ,csa_tree_add_110_49_pad_groupi_n_281);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5694(csa_tree_add_110_49_pad_groupi_n_206 ,csa_tree_add_110_49_pad_groupi_n_204);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5695(csa_tree_add_110_49_pad_groupi_n_205 ,csa_tree_add_110_49_pad_groupi_n_204);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5696(csa_tree_add_110_49_pad_groupi_n_204 ,csa_tree_add_110_49_pad_groupi_n_388);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5698(csa_tree_add_110_49_pad_groupi_n_203 ,csa_tree_add_110_49_pad_groupi_n_201);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5699(csa_tree_add_110_49_pad_groupi_n_202 ,csa_tree_add_110_49_pad_groupi_n_201);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5700(csa_tree_add_110_49_pad_groupi_n_201 ,csa_tree_add_110_49_pad_groupi_n_279);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5702(csa_tree_add_110_49_pad_groupi_n_200 ,csa_tree_add_110_49_pad_groupi_n_198);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5703(csa_tree_add_110_49_pad_groupi_n_199 ,csa_tree_add_110_49_pad_groupi_n_198);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5704(csa_tree_add_110_49_pad_groupi_n_198 ,csa_tree_add_110_49_pad_groupi_n_278);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5706(csa_tree_add_110_49_pad_groupi_n_197 ,csa_tree_add_110_49_pad_groupi_n_195);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5707(csa_tree_add_110_49_pad_groupi_n_196 ,csa_tree_add_110_49_pad_groupi_n_195);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5708(csa_tree_add_110_49_pad_groupi_n_195 ,csa_tree_add_110_49_pad_groupi_n_437);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5712(csa_tree_add_110_49_pad_groupi_n_284 ,csa_tree_add_110_49_pad_groupi_n_692);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5715(csa_tree_add_110_49_pad_groupi_n_194 ,csa_tree_add_110_49_pad_groupi_n_193);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5716(csa_tree_add_110_49_pad_groupi_n_193 ,csa_tree_add_110_49_pad_groupi_n_289);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5719(csa_tree_add_110_49_pad_groupi_n_192 ,csa_tree_add_110_49_pad_groupi_n_191);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5720(csa_tree_add_110_49_pad_groupi_n_191 ,csa_tree_add_110_49_pad_groupi_n_291);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5723(csa_tree_add_110_49_pad_groupi_n_190 ,csa_tree_add_110_49_pad_groupi_n_189);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5724(csa_tree_add_110_49_pad_groupi_n_189 ,csa_tree_add_110_49_pad_groupi_n_290);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5735(csa_tree_add_110_49_pad_groupi_n_188 ,csa_tree_add_110_49_pad_groupi_n_286);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5736(csa_tree_add_110_49_pad_groupi_n_286 ,csa_tree_add_110_49_pad_groupi_n_1184);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5739(csa_tree_add_110_49_pad_groupi_n_187 ,csa_tree_add_110_49_pad_groupi_n_287);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5740(csa_tree_add_110_49_pad_groupi_n_287 ,csa_tree_add_110_49_pad_groupi_n_1275);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5762(csa_tree_add_110_49_pad_groupi_n_186 ,csa_tree_add_110_49_pad_groupi_n_185);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5764(csa_tree_add_110_49_pad_groupi_n_185 ,csa_tree_add_110_49_pad_groupi_n_293);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5767(csa_tree_add_110_49_pad_groupi_n_184 ,csa_tree_add_110_49_pad_groupi_n_183);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5769(csa_tree_add_110_49_pad_groupi_n_183 ,csa_tree_add_110_49_pad_groupi_n_570);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5772(csa_tree_add_110_49_pad_groupi_n_182 ,csa_tree_add_110_49_pad_groupi_n_181);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5774(csa_tree_add_110_49_pad_groupi_n_181 ,csa_tree_add_110_49_pad_groupi_n_510);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5782(csa_tree_add_110_49_pad_groupi_n_180 ,csa_tree_add_110_49_pad_groupi_n_179);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5784(csa_tree_add_110_49_pad_groupi_n_179 ,csa_tree_add_110_49_pad_groupi_n_571);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5787(csa_tree_add_110_49_pad_groupi_n_178 ,csa_tree_add_110_49_pad_groupi_n_177);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5789(csa_tree_add_110_49_pad_groupi_n_177 ,csa_tree_add_110_49_pad_groupi_n_511);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5792(csa_tree_add_110_49_pad_groupi_n_176 ,csa_tree_add_110_49_pad_groupi_n_174);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5793(csa_tree_add_110_49_pad_groupi_n_175 ,csa_tree_add_110_49_pad_groupi_n_174);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5794(csa_tree_add_110_49_pad_groupi_n_174 ,csa_tree_add_110_49_pad_groupi_n_301);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5796(csa_tree_add_110_49_pad_groupi_n_173 ,csa_tree_add_110_49_pad_groupi_n_171);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5797(csa_tree_add_110_49_pad_groupi_n_172 ,csa_tree_add_110_49_pad_groupi_n_171);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5798(csa_tree_add_110_49_pad_groupi_n_171 ,csa_tree_add_110_49_pad_groupi_n_277);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5800(csa_tree_add_110_49_pad_groupi_n_170 ,csa_tree_add_110_49_pad_groupi_n_168);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5801(csa_tree_add_110_49_pad_groupi_n_169 ,csa_tree_add_110_49_pad_groupi_n_168);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5802(csa_tree_add_110_49_pad_groupi_n_168 ,csa_tree_add_110_49_pad_groupi_n_277);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5804(csa_tree_add_110_49_pad_groupi_n_167 ,csa_tree_add_110_49_pad_groupi_n_165);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5805(csa_tree_add_110_49_pad_groupi_n_166 ,csa_tree_add_110_49_pad_groupi_n_165);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5806(csa_tree_add_110_49_pad_groupi_n_165 ,csa_tree_add_110_49_pad_groupi_n_301);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5808(csa_tree_add_110_49_pad_groupi_n_164 ,csa_tree_add_110_49_pad_groupi_n_162);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5809(csa_tree_add_110_49_pad_groupi_n_163 ,csa_tree_add_110_49_pad_groupi_n_162);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5810(csa_tree_add_110_49_pad_groupi_n_162 ,csa_tree_add_110_49_pad_groupi_n_391);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5812(csa_tree_add_110_49_pad_groupi_n_161 ,csa_tree_add_110_49_pad_groupi_n_159);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5813(csa_tree_add_110_49_pad_groupi_n_160 ,csa_tree_add_110_49_pad_groupi_n_159);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5814(csa_tree_add_110_49_pad_groupi_n_159 ,csa_tree_add_110_49_pad_groupi_n_390);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5816(csa_tree_add_110_49_pad_groupi_n_158 ,csa_tree_add_110_49_pad_groupi_n_156);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5817(csa_tree_add_110_49_pad_groupi_n_157 ,csa_tree_add_110_49_pad_groupi_n_156);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5818(csa_tree_add_110_49_pad_groupi_n_156 ,csa_tree_add_110_49_pad_groupi_n_390);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5820(csa_tree_add_110_49_pad_groupi_n_155 ,csa_tree_add_110_49_pad_groupi_n_153);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5821(csa_tree_add_110_49_pad_groupi_n_154 ,csa_tree_add_110_49_pad_groupi_n_153);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5822(csa_tree_add_110_49_pad_groupi_n_153 ,csa_tree_add_110_49_pad_groupi_n_514);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5824(csa_tree_add_110_49_pad_groupi_n_152 ,csa_tree_add_110_49_pad_groupi_n_150);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5825(csa_tree_add_110_49_pad_groupi_n_151 ,csa_tree_add_110_49_pad_groupi_n_150);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5826(csa_tree_add_110_49_pad_groupi_n_150 ,csa_tree_add_110_49_pad_groupi_n_514);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5828(csa_tree_add_110_49_pad_groupi_n_149 ,csa_tree_add_110_49_pad_groupi_n_147);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5829(csa_tree_add_110_49_pad_groupi_n_148 ,csa_tree_add_110_49_pad_groupi_n_147);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5830(csa_tree_add_110_49_pad_groupi_n_147 ,csa_tree_add_110_49_pad_groupi_n_391);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5832(csa_tree_add_110_49_pad_groupi_n_146 ,csa_tree_add_110_49_pad_groupi_n_285);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5834(csa_tree_add_110_49_pad_groupi_n_285 ,csa_tree_add_110_49_pad_groupi_n_743);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5836(csa_tree_add_110_49_pad_groupi_n_145 ,csa_tree_add_110_49_pad_groupi_n_283);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5838(csa_tree_add_110_49_pad_groupi_n_283 ,csa_tree_add_110_49_pad_groupi_n_438);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5840(csa_tree_add_110_49_pad_groupi_n_144 ,csa_tree_add_110_49_pad_groupi_n_282);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5842(csa_tree_add_110_49_pad_groupi_n_282 ,csa_tree_add_110_49_pad_groupi_n_438);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5844(csa_tree_add_110_49_pad_groupi_n_143 ,csa_tree_add_110_49_pad_groupi_n_281);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5846(csa_tree_add_110_49_pad_groupi_n_281 ,csa_tree_add_110_49_pad_groupi_n_435);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5848(csa_tree_add_110_49_pad_groupi_n_142 ,csa_tree_add_110_49_pad_groupi_n_280);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5850(csa_tree_add_110_49_pad_groupi_n_280 ,csa_tree_add_110_49_pad_groupi_n_435);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5852(csa_tree_add_110_49_pad_groupi_n_141 ,csa_tree_add_110_49_pad_groupi_n_279);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5854(csa_tree_add_110_49_pad_groupi_n_279 ,csa_tree_add_110_49_pad_groupi_n_386);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5856(csa_tree_add_110_49_pad_groupi_n_140 ,csa_tree_add_110_49_pad_groupi_n_278);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5858(csa_tree_add_110_49_pad_groupi_n_278 ,csa_tree_add_110_49_pad_groupi_n_386);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5861(csa_tree_add_110_49_pad_groupi_n_139 ,csa_tree_add_110_49_pad_groupi_n_138);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5862(csa_tree_add_110_49_pad_groupi_n_138 ,csa_tree_add_110_49_pad_groupi_n_743);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5864(csa_tree_add_110_49_pad_groupi_n_137 ,csa_tree_add_110_49_pad_groupi_n_135);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5865(csa_tree_add_110_49_pad_groupi_n_136 ,csa_tree_add_110_49_pad_groupi_n_135);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5866(csa_tree_add_110_49_pad_groupi_n_135 ,csa_tree_add_110_49_pad_groupi_n_513);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5868(csa_tree_add_110_49_pad_groupi_n_134 ,csa_tree_add_110_49_pad_groupi_n_132);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5869(csa_tree_add_110_49_pad_groupi_n_133 ,csa_tree_add_110_49_pad_groupi_n_132);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5870(csa_tree_add_110_49_pad_groupi_n_132 ,csa_tree_add_110_49_pad_groupi_n_513);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5872(csa_tree_add_110_49_pad_groupi_n_131 ,csa_tree_add_110_49_pad_groupi_n_130);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5874(csa_tree_add_110_49_pad_groupi_n_130 ,csa_tree_add_110_49_pad_groupi_n_274);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5876(csa_tree_add_110_49_pad_groupi_n_129 ,csa_tree_add_110_49_pad_groupi_n_128);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5878(csa_tree_add_110_49_pad_groupi_n_128 ,csa_tree_add_110_49_pad_groupi_n_247);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5880(csa_tree_add_110_49_pad_groupi_n_127 ,csa_tree_add_110_49_pad_groupi_n_126);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5882(csa_tree_add_110_49_pad_groupi_n_126 ,csa_tree_add_110_49_pad_groupi_n_259);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5884(csa_tree_add_110_49_pad_groupi_n_125 ,csa_tree_add_110_49_pad_groupi_n_124);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5886(csa_tree_add_110_49_pad_groupi_n_124 ,csa_tree_add_110_49_pad_groupi_n_260);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5888(csa_tree_add_110_49_pad_groupi_n_123 ,csa_tree_add_110_49_pad_groupi_n_122);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5890(csa_tree_add_110_49_pad_groupi_n_122 ,csa_tree_add_110_49_pad_groupi_n_244);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5892(csa_tree_add_110_49_pad_groupi_n_121 ,csa_tree_add_110_49_pad_groupi_n_120);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5894(csa_tree_add_110_49_pad_groupi_n_120 ,csa_tree_add_110_49_pad_groupi_n_262);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5896(csa_tree_add_110_49_pad_groupi_n_119 ,csa_tree_add_110_49_pad_groupi_n_118);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5898(csa_tree_add_110_49_pad_groupi_n_118 ,csa_tree_add_110_49_pad_groupi_n_236);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5900(csa_tree_add_110_49_pad_groupi_n_117 ,csa_tree_add_110_49_pad_groupi_n_116);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5902(csa_tree_add_110_49_pad_groupi_n_116 ,csa_tree_add_110_49_pad_groupi_n_245);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5904(csa_tree_add_110_49_pad_groupi_n_115 ,csa_tree_add_110_49_pad_groupi_n_114);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5906(csa_tree_add_110_49_pad_groupi_n_114 ,csa_tree_add_110_49_pad_groupi_n_253);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5908(csa_tree_add_110_49_pad_groupi_n_113 ,csa_tree_add_110_49_pad_groupi_n_112);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5910(csa_tree_add_110_49_pad_groupi_n_112 ,csa_tree_add_110_49_pad_groupi_n_241);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5912(csa_tree_add_110_49_pad_groupi_n_111 ,csa_tree_add_110_49_pad_groupi_n_110);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5914(csa_tree_add_110_49_pad_groupi_n_110 ,csa_tree_add_110_49_pad_groupi_n_239);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5916(csa_tree_add_110_49_pad_groupi_n_109 ,csa_tree_add_110_49_pad_groupi_n_108);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5918(csa_tree_add_110_49_pad_groupi_n_108 ,csa_tree_add_110_49_pad_groupi_n_233);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5920(csa_tree_add_110_49_pad_groupi_n_107 ,csa_tree_add_110_49_pad_groupi_n_106);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5922(csa_tree_add_110_49_pad_groupi_n_106 ,csa_tree_add_110_49_pad_groupi_n_242);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5924(csa_tree_add_110_49_pad_groupi_n_105 ,csa_tree_add_110_49_pad_groupi_n_104);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5926(csa_tree_add_110_49_pad_groupi_n_104 ,csa_tree_add_110_49_pad_groupi_n_268);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5928(csa_tree_add_110_49_pad_groupi_n_103 ,csa_tree_add_110_49_pad_groupi_n_102);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5930(csa_tree_add_110_49_pad_groupi_n_102 ,csa_tree_add_110_49_pad_groupi_n_235);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5932(csa_tree_add_110_49_pad_groupi_n_101 ,csa_tree_add_110_49_pad_groupi_n_100);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5934(csa_tree_add_110_49_pad_groupi_n_100 ,csa_tree_add_110_49_pad_groupi_n_256);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5936(csa_tree_add_110_49_pad_groupi_n_99 ,csa_tree_add_110_49_pad_groupi_n_98);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5938(csa_tree_add_110_49_pad_groupi_n_98 ,csa_tree_add_110_49_pad_groupi_n_250);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5940(csa_tree_add_110_49_pad_groupi_n_97 ,csa_tree_add_110_49_pad_groupi_n_96);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5942(csa_tree_add_110_49_pad_groupi_n_96 ,csa_tree_add_110_49_pad_groupi_n_251);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5944(csa_tree_add_110_49_pad_groupi_n_95 ,csa_tree_add_110_49_pad_groupi_n_94);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5946(csa_tree_add_110_49_pad_groupi_n_94 ,csa_tree_add_110_49_pad_groupi_n_266);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5948(csa_tree_add_110_49_pad_groupi_n_93 ,csa_tree_add_110_49_pad_groupi_n_92);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5950(csa_tree_add_110_49_pad_groupi_n_92 ,csa_tree_add_110_49_pad_groupi_n_263);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5952(csa_tree_add_110_49_pad_groupi_n_91 ,csa_tree_add_110_49_pad_groupi_n_90);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5954(csa_tree_add_110_49_pad_groupi_n_90 ,csa_tree_add_110_49_pad_groupi_n_265);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5956(csa_tree_add_110_49_pad_groupi_n_89 ,csa_tree_add_110_49_pad_groupi_n_88);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5958(csa_tree_add_110_49_pad_groupi_n_88 ,csa_tree_add_110_49_pad_groupi_n_257);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5960(csa_tree_add_110_49_pad_groupi_n_87 ,csa_tree_add_110_49_pad_groupi_n_86);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5962(csa_tree_add_110_49_pad_groupi_n_86 ,csa_tree_add_110_49_pad_groupi_n_248);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5964(csa_tree_add_110_49_pad_groupi_n_85 ,csa_tree_add_110_49_pad_groupi_n_84);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5966(csa_tree_add_110_49_pad_groupi_n_84 ,csa_tree_add_110_49_pad_groupi_n_238);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5968(csa_tree_add_110_49_pad_groupi_n_83 ,csa_tree_add_110_49_pad_groupi_n_82);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5970(csa_tree_add_110_49_pad_groupi_n_82 ,csa_tree_add_110_49_pad_groupi_n_254);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5972(csa_tree_add_110_49_pad_groupi_n_81 ,csa_tree_add_110_49_pad_groupi_n_80);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5974(csa_tree_add_110_49_pad_groupi_n_80 ,csa_tree_add_110_49_pad_groupi_n_269);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5976(csa_tree_add_110_49_pad_groupi_n_79 ,csa_tree_add_110_49_pad_groupi_n_78);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5978(csa_tree_add_110_49_pad_groupi_n_78 ,csa_tree_add_110_49_pad_groupi_n_271);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5980(csa_tree_add_110_49_pad_groupi_n_77 ,csa_tree_add_110_49_pad_groupi_n_76);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5982(csa_tree_add_110_49_pad_groupi_n_76 ,csa_tree_add_110_49_pad_groupi_n_272);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5984(csa_tree_add_110_49_pad_groupi_n_75 ,csa_tree_add_110_49_pad_groupi_n_74);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5986(csa_tree_add_110_49_pad_groupi_n_74 ,csa_tree_add_110_49_pad_groupi_n_275);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5988(csa_tree_add_110_49_pad_groupi_n_73 ,csa_tree_add_110_49_pad_groupi_n_71);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5989(csa_tree_add_110_49_pad_groupi_n_72 ,csa_tree_add_110_49_pad_groupi_n_71);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5990(csa_tree_add_110_49_pad_groupi_n_71 ,csa_tree_add_110_49_pad_groupi_n_293);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5992(csa_tree_add_110_49_pad_groupi_n_70 ,csa_tree_add_110_49_pad_groupi_n_68);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5993(csa_tree_add_110_49_pad_groupi_n_69 ,csa_tree_add_110_49_pad_groupi_n_68);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5994(csa_tree_add_110_49_pad_groupi_n_68 ,csa_tree_add_110_49_pad_groupi_n_511);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5996(csa_tree_add_110_49_pad_groupi_n_67 ,csa_tree_add_110_49_pad_groupi_n_65);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5997(csa_tree_add_110_49_pad_groupi_n_66 ,csa_tree_add_110_49_pad_groupi_n_65);
  not csa_tree_add_110_49_pad_groupi_drc_bufs5998(csa_tree_add_110_49_pad_groupi_n_65 ,csa_tree_add_110_49_pad_groupi_n_570);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6000(csa_tree_add_110_49_pad_groupi_n_64 ,csa_tree_add_110_49_pad_groupi_n_62);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6001(csa_tree_add_110_49_pad_groupi_n_63 ,csa_tree_add_110_49_pad_groupi_n_62);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6002(csa_tree_add_110_49_pad_groupi_n_62 ,csa_tree_add_110_49_pad_groupi_n_510);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6004(csa_tree_add_110_49_pad_groupi_n_61 ,csa_tree_add_110_49_pad_groupi_n_59);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6005(csa_tree_add_110_49_pad_groupi_n_60 ,csa_tree_add_110_49_pad_groupi_n_59);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6006(csa_tree_add_110_49_pad_groupi_n_59 ,csa_tree_add_110_49_pad_groupi_n_186);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6008(csa_tree_add_110_49_pad_groupi_n_58 ,csa_tree_add_110_49_pad_groupi_n_56);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6009(csa_tree_add_110_49_pad_groupi_n_57 ,csa_tree_add_110_49_pad_groupi_n_56);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6010(csa_tree_add_110_49_pad_groupi_n_56 ,csa_tree_add_110_49_pad_groupi_n_180);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6012(csa_tree_add_110_49_pad_groupi_n_55 ,csa_tree_add_110_49_pad_groupi_n_53);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6013(csa_tree_add_110_49_pad_groupi_n_54 ,csa_tree_add_110_49_pad_groupi_n_53);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6014(csa_tree_add_110_49_pad_groupi_n_53 ,csa_tree_add_110_49_pad_groupi_n_178);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6016(csa_tree_add_110_49_pad_groupi_n_52 ,csa_tree_add_110_49_pad_groupi_n_50);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6017(csa_tree_add_110_49_pad_groupi_n_51 ,csa_tree_add_110_49_pad_groupi_n_50);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6018(csa_tree_add_110_49_pad_groupi_n_50 ,csa_tree_add_110_49_pad_groupi_n_293);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6020(csa_tree_add_110_49_pad_groupi_n_49 ,csa_tree_add_110_49_pad_groupi_n_47);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6021(csa_tree_add_110_49_pad_groupi_n_48 ,csa_tree_add_110_49_pad_groupi_n_47);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6022(csa_tree_add_110_49_pad_groupi_n_47 ,csa_tree_add_110_49_pad_groupi_n_186);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6024(csa_tree_add_110_49_pad_groupi_n_46 ,csa_tree_add_110_49_pad_groupi_n_44);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6025(csa_tree_add_110_49_pad_groupi_n_45 ,csa_tree_add_110_49_pad_groupi_n_44);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6026(csa_tree_add_110_49_pad_groupi_n_44 ,csa_tree_add_110_49_pad_groupi_n_184);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6028(csa_tree_add_110_49_pad_groupi_n_43 ,csa_tree_add_110_49_pad_groupi_n_41);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6029(csa_tree_add_110_49_pad_groupi_n_42 ,csa_tree_add_110_49_pad_groupi_n_41);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6030(csa_tree_add_110_49_pad_groupi_n_41 ,csa_tree_add_110_49_pad_groupi_n_182);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6032(csa_tree_add_110_49_pad_groupi_n_40 ,csa_tree_add_110_49_pad_groupi_n_38);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6033(csa_tree_add_110_49_pad_groupi_n_39 ,csa_tree_add_110_49_pad_groupi_n_38);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6034(csa_tree_add_110_49_pad_groupi_n_38 ,csa_tree_add_110_49_pad_groupi_n_571);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6036(csa_tree_add_110_49_pad_groupi_n_37 ,csa_tree_add_110_49_pad_groupi_n_35);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6037(csa_tree_add_110_49_pad_groupi_n_36 ,csa_tree_add_110_49_pad_groupi_n_35);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6038(csa_tree_add_110_49_pad_groupi_n_35 ,csa_tree_add_110_49_pad_groupi_n_511);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6040(csa_tree_add_110_49_pad_groupi_n_34 ,csa_tree_add_110_49_pad_groupi_n_32);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6041(csa_tree_add_110_49_pad_groupi_n_33 ,csa_tree_add_110_49_pad_groupi_n_32);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6042(csa_tree_add_110_49_pad_groupi_n_32 ,csa_tree_add_110_49_pad_groupi_n_180);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6044(csa_tree_add_110_49_pad_groupi_n_31 ,csa_tree_add_110_49_pad_groupi_n_29);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6045(csa_tree_add_110_49_pad_groupi_n_30 ,csa_tree_add_110_49_pad_groupi_n_29);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6046(csa_tree_add_110_49_pad_groupi_n_29 ,csa_tree_add_110_49_pad_groupi_n_510);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6048(csa_tree_add_110_49_pad_groupi_n_28 ,csa_tree_add_110_49_pad_groupi_n_26);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6049(csa_tree_add_110_49_pad_groupi_n_27 ,csa_tree_add_110_49_pad_groupi_n_26);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6050(csa_tree_add_110_49_pad_groupi_n_26 ,csa_tree_add_110_49_pad_groupi_n_184);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6052(csa_tree_add_110_49_pad_groupi_n_25 ,csa_tree_add_110_49_pad_groupi_n_23);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6053(csa_tree_add_110_49_pad_groupi_n_24 ,csa_tree_add_110_49_pad_groupi_n_23);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6054(csa_tree_add_110_49_pad_groupi_n_23 ,csa_tree_add_110_49_pad_groupi_n_570);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6056(csa_tree_add_110_49_pad_groupi_n_22 ,csa_tree_add_110_49_pad_groupi_n_20);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6057(csa_tree_add_110_49_pad_groupi_n_21 ,csa_tree_add_110_49_pad_groupi_n_20);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6058(csa_tree_add_110_49_pad_groupi_n_20 ,csa_tree_add_110_49_pad_groupi_n_182);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6060(csa_tree_add_110_49_pad_groupi_n_19 ,csa_tree_add_110_49_pad_groupi_n_17);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6061(csa_tree_add_110_49_pad_groupi_n_18 ,csa_tree_add_110_49_pad_groupi_n_17);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6062(csa_tree_add_110_49_pad_groupi_n_17 ,csa_tree_add_110_49_pad_groupi_n_571);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6064(csa_tree_add_110_49_pad_groupi_n_16 ,csa_tree_add_110_49_pad_groupi_n_14);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6065(csa_tree_add_110_49_pad_groupi_n_15 ,csa_tree_add_110_49_pad_groupi_n_14);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6066(csa_tree_add_110_49_pad_groupi_n_14 ,csa_tree_add_110_49_pad_groupi_n_178);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6068(csa_tree_add_110_49_pad_groupi_n_13 ,csa_tree_add_110_49_pad_groupi_n_12);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6070(csa_tree_add_110_49_pad_groupi_n_12 ,csa_tree_add_110_49_pad_groupi_n_175);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6072(csa_tree_add_110_49_pad_groupi_n_11 ,csa_tree_add_110_49_pad_groupi_n_10);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6074(csa_tree_add_110_49_pad_groupi_n_10 ,csa_tree_add_110_49_pad_groupi_n_73);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6076(csa_tree_add_110_49_pad_groupi_n_9 ,csa_tree_add_110_49_pad_groupi_n_8);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6078(csa_tree_add_110_49_pad_groupi_n_8 ,csa_tree_add_110_49_pad_groupi_n_64);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6080(csa_tree_add_110_49_pad_groupi_n_7 ,csa_tree_add_110_49_pad_groupi_n_6);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6082(csa_tree_add_110_49_pad_groupi_n_6 ,csa_tree_add_110_49_pad_groupi_n_67);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6084(csa_tree_add_110_49_pad_groupi_n_5 ,csa_tree_add_110_49_pad_groupi_n_4);
  not csa_tree_add_110_49_pad_groupi_drc_bufs6086(csa_tree_add_110_49_pad_groupi_n_4 ,csa_tree_add_110_49_pad_groupi_n_70);
  xor csa_tree_add_110_49_pad_groupi_g2(n_140 ,csa_tree_add_110_49_pad_groupi_n_1550 ,csa_tree_add_110_49_pad_groupi_n_1501);
  xor csa_tree_add_110_49_pad_groupi_g6088(n_139 ,csa_tree_add_110_49_pad_groupi_n_1548 ,csa_tree_add_110_49_pad_groupi_n_1518);
  xor csa_tree_add_110_49_pad_groupi_g6089(csa_tree_add_110_49_pad_groupi_n_1 ,csa_tree_add_110_49_pad_groupi_n_1237 ,csa_tree_add_110_49_pad_groupi_n_1418);
  xor csa_tree_add_110_49_pad_groupi_g6090(csa_tree_add_110_49_pad_groupi_n_0 ,csa_tree_add_110_49_pad_groupi_n_904 ,csa_tree_add_110_49_pad_groupi_n_284);
  xnor csa_tree_add_117_21_pad_groupi_g3221(out1[15] ,csa_tree_add_117_21_pad_groupi_n_1045 ,csa_tree_add_117_21_pad_groupi_n_1181);
  nor csa_tree_add_117_21_pad_groupi_g3222(csa_tree_add_117_21_pad_groupi_n_1181 ,csa_tree_add_117_21_pad_groupi_n_1052 ,csa_tree_add_117_21_pad_groupi_n_1179);
  xnor csa_tree_add_117_21_pad_groupi_g3223(out1[14] ,csa_tree_add_117_21_pad_groupi_n_1178 ,csa_tree_add_117_21_pad_groupi_n_1070);
  and csa_tree_add_117_21_pad_groupi_g3224(csa_tree_add_117_21_pad_groupi_n_1179 ,csa_tree_add_117_21_pad_groupi_n_1178 ,csa_tree_add_117_21_pad_groupi_n_1053);
  or csa_tree_add_117_21_pad_groupi_g3225(csa_tree_add_117_21_pad_groupi_n_1178 ,csa_tree_add_117_21_pad_groupi_n_1082 ,csa_tree_add_117_21_pad_groupi_n_1176);
  xnor csa_tree_add_117_21_pad_groupi_g3226(out1[13] ,csa_tree_add_117_21_pad_groupi_n_1175 ,csa_tree_add_117_21_pad_groupi_n_1088);
  nor csa_tree_add_117_21_pad_groupi_g3227(csa_tree_add_117_21_pad_groupi_n_1176 ,csa_tree_add_117_21_pad_groupi_n_1175 ,csa_tree_add_117_21_pad_groupi_n_1080);
  and csa_tree_add_117_21_pad_groupi_g3228(csa_tree_add_117_21_pad_groupi_n_1175 ,csa_tree_add_117_21_pad_groupi_n_1173 ,csa_tree_add_117_21_pad_groupi_n_1101);
  xnor csa_tree_add_117_21_pad_groupi_g3229(out1[12] ,csa_tree_add_117_21_pad_groupi_n_1171 ,csa_tree_add_117_21_pad_groupi_n_1110);
  or csa_tree_add_117_21_pad_groupi_g3230(csa_tree_add_117_21_pad_groupi_n_1173 ,csa_tree_add_117_21_pad_groupi_n_1172 ,csa_tree_add_117_21_pad_groupi_n_1100);
  not csa_tree_add_117_21_pad_groupi_g3231(csa_tree_add_117_21_pad_groupi_n_1172 ,csa_tree_add_117_21_pad_groupi_n_1171);
  or csa_tree_add_117_21_pad_groupi_g3232(csa_tree_add_117_21_pad_groupi_n_1171 ,csa_tree_add_117_21_pad_groupi_n_1169 ,csa_tree_add_117_21_pad_groupi_n_1099);
  xnor csa_tree_add_117_21_pad_groupi_g3233(out1[11] ,csa_tree_add_117_21_pad_groupi_n_1168 ,csa_tree_add_117_21_pad_groupi_n_1111);
  and csa_tree_add_117_21_pad_groupi_g3234(csa_tree_add_117_21_pad_groupi_n_1169 ,csa_tree_add_117_21_pad_groupi_n_1168 ,csa_tree_add_117_21_pad_groupi_n_1102);
  or csa_tree_add_117_21_pad_groupi_g3235(csa_tree_add_117_21_pad_groupi_n_1168 ,csa_tree_add_117_21_pad_groupi_n_1090 ,csa_tree_add_117_21_pad_groupi_n_1166);
  xnor csa_tree_add_117_21_pad_groupi_g3236(csa_tree_add_117_21_pad_groupi_n_1167 ,csa_tree_add_117_21_pad_groupi_n_1165 ,csa_tree_add_117_21_pad_groupi_n_1112);
  and csa_tree_add_117_21_pad_groupi_g3237(csa_tree_add_117_21_pad_groupi_n_1166 ,csa_tree_add_117_21_pad_groupi_n_1089 ,csa_tree_add_117_21_pad_groupi_n_1165);
  or csa_tree_add_117_21_pad_groupi_g3238(csa_tree_add_117_21_pad_groupi_n_1165 ,csa_tree_add_117_21_pad_groupi_n_1121 ,csa_tree_add_117_21_pad_groupi_n_1163);
  xnor csa_tree_add_117_21_pad_groupi_g3239(out1[9] ,csa_tree_add_117_21_pad_groupi_n_1162 ,csa_tree_add_117_21_pad_groupi_n_1134);
  and csa_tree_add_117_21_pad_groupi_g3240(csa_tree_add_117_21_pad_groupi_n_1163 ,csa_tree_add_117_21_pad_groupi_n_1128 ,csa_tree_add_117_21_pad_groupi_n_1162);
  or csa_tree_add_117_21_pad_groupi_g3241(csa_tree_add_117_21_pad_groupi_n_1162 ,csa_tree_add_117_21_pad_groupi_n_1160 ,csa_tree_add_117_21_pad_groupi_n_1118);
  xnor csa_tree_add_117_21_pad_groupi_g3242(out1[8] ,csa_tree_add_117_21_pad_groupi_n_1159 ,csa_tree_add_117_21_pad_groupi_n_1133);
  and csa_tree_add_117_21_pad_groupi_g3243(csa_tree_add_117_21_pad_groupi_n_1160 ,csa_tree_add_117_21_pad_groupi_n_1119 ,csa_tree_add_117_21_pad_groupi_n_1159);
  or csa_tree_add_117_21_pad_groupi_g3244(csa_tree_add_117_21_pad_groupi_n_1159 ,csa_tree_add_117_21_pad_groupi_n_1117 ,csa_tree_add_117_21_pad_groupi_n_1157);
  xnor csa_tree_add_117_21_pad_groupi_g3245(out1[7] ,csa_tree_add_117_21_pad_groupi_n_1156 ,csa_tree_add_117_21_pad_groupi_n_1132);
  and csa_tree_add_117_21_pad_groupi_g3246(csa_tree_add_117_21_pad_groupi_n_1157 ,csa_tree_add_117_21_pad_groupi_n_1116 ,csa_tree_add_117_21_pad_groupi_n_1156);
  or csa_tree_add_117_21_pad_groupi_g3247(csa_tree_add_117_21_pad_groupi_n_1156 ,csa_tree_add_117_21_pad_groupi_n_1115 ,csa_tree_add_117_21_pad_groupi_n_1154);
  xnor csa_tree_add_117_21_pad_groupi_g3248(out1[6] ,csa_tree_add_117_21_pad_groupi_n_1153 ,csa_tree_add_117_21_pad_groupi_n_1131);
  and csa_tree_add_117_21_pad_groupi_g3249(csa_tree_add_117_21_pad_groupi_n_1154 ,csa_tree_add_117_21_pad_groupi_n_1114 ,csa_tree_add_117_21_pad_groupi_n_1153);
  or csa_tree_add_117_21_pad_groupi_g3250(csa_tree_add_117_21_pad_groupi_n_1153 ,csa_tree_add_117_21_pad_groupi_n_1151 ,csa_tree_add_117_21_pad_groupi_n_1126);
  xnor csa_tree_add_117_21_pad_groupi_g3251(out1[5] ,csa_tree_add_117_21_pad_groupi_n_1150 ,csa_tree_add_117_21_pad_groupi_n_1130);
  and csa_tree_add_117_21_pad_groupi_g3252(csa_tree_add_117_21_pad_groupi_n_1151 ,csa_tree_add_117_21_pad_groupi_n_1125 ,csa_tree_add_117_21_pad_groupi_n_1150);
  or csa_tree_add_117_21_pad_groupi_g3253(csa_tree_add_117_21_pad_groupi_n_1150 ,csa_tree_add_117_21_pad_groupi_n_1124 ,csa_tree_add_117_21_pad_groupi_n_1148);
  xnor csa_tree_add_117_21_pad_groupi_g3254(out1[4] ,csa_tree_add_117_21_pad_groupi_n_1147 ,csa_tree_add_117_21_pad_groupi_n_1135);
  and csa_tree_add_117_21_pad_groupi_g3255(csa_tree_add_117_21_pad_groupi_n_1148 ,csa_tree_add_117_21_pad_groupi_n_1123 ,csa_tree_add_117_21_pad_groupi_n_1147);
  or csa_tree_add_117_21_pad_groupi_g3256(csa_tree_add_117_21_pad_groupi_n_1147 ,csa_tree_add_117_21_pad_groupi_n_1145 ,csa_tree_add_117_21_pad_groupi_n_1127);
  xnor csa_tree_add_117_21_pad_groupi_g3257(out1[3] ,csa_tree_add_117_21_pad_groupi_n_1144 ,csa_tree_add_117_21_pad_groupi_n_1136);
  nor csa_tree_add_117_21_pad_groupi_g3258(csa_tree_add_117_21_pad_groupi_n_1145 ,csa_tree_add_117_21_pad_groupi_n_1144 ,csa_tree_add_117_21_pad_groupi_n_1120);
  and csa_tree_add_117_21_pad_groupi_g3259(csa_tree_add_117_21_pad_groupi_n_1144 ,csa_tree_add_117_21_pad_groupi_n_1142 ,csa_tree_add_117_21_pad_groupi_n_1104);
  xnor csa_tree_add_117_21_pad_groupi_g3260(out1[2] ,csa_tree_add_117_21_pad_groupi_n_1140 ,csa_tree_add_117_21_pad_groupi_n_1113);
  or csa_tree_add_117_21_pad_groupi_g3261(csa_tree_add_117_21_pad_groupi_n_1142 ,csa_tree_add_117_21_pad_groupi_n_1103 ,csa_tree_add_117_21_pad_groupi_n_1141);
  not csa_tree_add_117_21_pad_groupi_g3262(csa_tree_add_117_21_pad_groupi_n_1141 ,csa_tree_add_117_21_pad_groupi_n_1140);
  or csa_tree_add_117_21_pad_groupi_g3263(csa_tree_add_117_21_pad_groupi_n_1140 ,csa_tree_add_117_21_pad_groupi_n_1138 ,csa_tree_add_117_21_pad_groupi_n_1063);
  xnor csa_tree_add_117_21_pad_groupi_g3264(csa_tree_add_117_21_pad_groupi_n_1139 ,csa_tree_add_117_21_pad_groupi_n_1137 ,csa_tree_add_117_21_pad_groupi_n_1071);
  and csa_tree_add_117_21_pad_groupi_g3265(csa_tree_add_117_21_pad_groupi_n_1138 ,csa_tree_add_117_21_pad_groupi_n_1067 ,csa_tree_add_117_21_pad_groupi_n_1137);
  or csa_tree_add_117_21_pad_groupi_g3266(csa_tree_add_117_21_pad_groupi_n_1137 ,csa_tree_add_117_21_pad_groupi_n_1031 ,csa_tree_add_117_21_pad_groupi_n_1122);
  xnor csa_tree_add_117_21_pad_groupi_g3267(csa_tree_add_117_21_pad_groupi_n_1136 ,csa_tree_add_117_21_pad_groupi_n_1084 ,csa_tree_add_117_21_pad_groupi_n_1091);
  xnor csa_tree_add_117_21_pad_groupi_g3268(csa_tree_add_117_21_pad_groupi_n_1135 ,csa_tree_add_117_21_pad_groupi_n_1107 ,csa_tree_add_117_21_pad_groupi_n_1092);
  xnor csa_tree_add_117_21_pad_groupi_g3269(csa_tree_add_117_21_pad_groupi_n_1134 ,csa_tree_add_117_21_pad_groupi_n_1109 ,csa_tree_add_117_21_pad_groupi_n_1097);
  xnor csa_tree_add_117_21_pad_groupi_g3270(csa_tree_add_117_21_pad_groupi_n_1133 ,csa_tree_add_117_21_pad_groupi_n_1108 ,csa_tree_add_117_21_pad_groupi_n_1096);
  xnor csa_tree_add_117_21_pad_groupi_g3271(csa_tree_add_117_21_pad_groupi_n_1132 ,csa_tree_add_117_21_pad_groupi_n_1087 ,csa_tree_add_117_21_pad_groupi_n_1095);
  xnor csa_tree_add_117_21_pad_groupi_g3272(csa_tree_add_117_21_pad_groupi_n_1131 ,csa_tree_add_117_21_pad_groupi_n_1106 ,csa_tree_add_117_21_pad_groupi_n_1094);
  xnor csa_tree_add_117_21_pad_groupi_g3273(csa_tree_add_117_21_pad_groupi_n_1130 ,csa_tree_add_117_21_pad_groupi_n_1105 ,csa_tree_add_117_21_pad_groupi_n_1093);
  xnor csa_tree_add_117_21_pad_groupi_g3274(csa_tree_add_117_21_pad_groupi_n_1129 ,csa_tree_add_117_21_pad_groupi_n_1098 ,csa_tree_add_117_21_pad_groupi_n_1047);
  or csa_tree_add_117_21_pad_groupi_g3275(csa_tree_add_117_21_pad_groupi_n_1128 ,csa_tree_add_117_21_pad_groupi_n_1109 ,csa_tree_add_117_21_pad_groupi_n_1097);
  nor csa_tree_add_117_21_pad_groupi_g3276(csa_tree_add_117_21_pad_groupi_n_1127 ,csa_tree_add_117_21_pad_groupi_n_1085 ,csa_tree_add_117_21_pad_groupi_n_1091);
  and csa_tree_add_117_21_pad_groupi_g3277(csa_tree_add_117_21_pad_groupi_n_1126 ,csa_tree_add_117_21_pad_groupi_n_1105 ,csa_tree_add_117_21_pad_groupi_n_1093);
  or csa_tree_add_117_21_pad_groupi_g3278(csa_tree_add_117_21_pad_groupi_n_1125 ,csa_tree_add_117_21_pad_groupi_n_1105 ,csa_tree_add_117_21_pad_groupi_n_1093);
  and csa_tree_add_117_21_pad_groupi_g3279(csa_tree_add_117_21_pad_groupi_n_1124 ,csa_tree_add_117_21_pad_groupi_n_1107 ,csa_tree_add_117_21_pad_groupi_n_1092);
  or csa_tree_add_117_21_pad_groupi_g3280(csa_tree_add_117_21_pad_groupi_n_1123 ,csa_tree_add_117_21_pad_groupi_n_1107 ,csa_tree_add_117_21_pad_groupi_n_1092);
  nor csa_tree_add_117_21_pad_groupi_g3281(csa_tree_add_117_21_pad_groupi_n_1122 ,csa_tree_add_117_21_pad_groupi_n_1035 ,csa_tree_add_117_21_pad_groupi_n_1098);
  and csa_tree_add_117_21_pad_groupi_g3282(csa_tree_add_117_21_pad_groupi_n_1121 ,csa_tree_add_117_21_pad_groupi_n_1109 ,csa_tree_add_117_21_pad_groupi_n_1097);
  and csa_tree_add_117_21_pad_groupi_g3283(csa_tree_add_117_21_pad_groupi_n_1120 ,csa_tree_add_117_21_pad_groupi_n_1085 ,csa_tree_add_117_21_pad_groupi_n_1091);
  or csa_tree_add_117_21_pad_groupi_g3284(csa_tree_add_117_21_pad_groupi_n_1119 ,csa_tree_add_117_21_pad_groupi_n_1108 ,csa_tree_add_117_21_pad_groupi_n_1096);
  and csa_tree_add_117_21_pad_groupi_g3285(csa_tree_add_117_21_pad_groupi_n_1118 ,csa_tree_add_117_21_pad_groupi_n_1108 ,csa_tree_add_117_21_pad_groupi_n_1096);
  and csa_tree_add_117_21_pad_groupi_g3286(csa_tree_add_117_21_pad_groupi_n_1117 ,csa_tree_add_117_21_pad_groupi_n_1087 ,csa_tree_add_117_21_pad_groupi_n_1095);
  or csa_tree_add_117_21_pad_groupi_g3287(csa_tree_add_117_21_pad_groupi_n_1116 ,csa_tree_add_117_21_pad_groupi_n_1087 ,csa_tree_add_117_21_pad_groupi_n_1095);
  and csa_tree_add_117_21_pad_groupi_g3288(csa_tree_add_117_21_pad_groupi_n_1115 ,csa_tree_add_117_21_pad_groupi_n_1106 ,csa_tree_add_117_21_pad_groupi_n_1094);
  or csa_tree_add_117_21_pad_groupi_g3289(csa_tree_add_117_21_pad_groupi_n_1114 ,csa_tree_add_117_21_pad_groupi_n_1106 ,csa_tree_add_117_21_pad_groupi_n_1094);
  xnor csa_tree_add_117_21_pad_groupi_g3290(csa_tree_add_117_21_pad_groupi_n_1113 ,csa_tree_add_117_21_pad_groupi_n_1077 ,csa_tree_add_117_21_pad_groupi_n_996);
  xnor csa_tree_add_117_21_pad_groupi_g3291(csa_tree_add_117_21_pad_groupi_n_1112 ,csa_tree_add_117_21_pad_groupi_n_1086 ,csa_tree_add_117_21_pad_groupi_n_1078);
  xnor csa_tree_add_117_21_pad_groupi_g3292(csa_tree_add_117_21_pad_groupi_n_1111 ,csa_tree_add_117_21_pad_groupi_n_1054 ,csa_tree_add_117_21_pad_groupi_n_1075);
  xnor csa_tree_add_117_21_pad_groupi_g3293(csa_tree_add_117_21_pad_groupi_n_1110 ,csa_tree_add_117_21_pad_groupi_n_1076 ,csa_tree_add_117_21_pad_groupi_n_1068);
  or csa_tree_add_117_21_pad_groupi_g3294(csa_tree_add_117_21_pad_groupi_n_1104 ,csa_tree_add_117_21_pad_groupi_n_996 ,csa_tree_add_117_21_pad_groupi_n_1077);
  and csa_tree_add_117_21_pad_groupi_g3295(csa_tree_add_117_21_pad_groupi_n_1103 ,csa_tree_add_117_21_pad_groupi_n_996 ,csa_tree_add_117_21_pad_groupi_n_1077);
  or csa_tree_add_117_21_pad_groupi_g3296(csa_tree_add_117_21_pad_groupi_n_1102 ,csa_tree_add_117_21_pad_groupi_n_1054 ,csa_tree_add_117_21_pad_groupi_n_1075);
  or csa_tree_add_117_21_pad_groupi_g3297(csa_tree_add_117_21_pad_groupi_n_1101 ,csa_tree_add_117_21_pad_groupi_n_1068 ,csa_tree_add_117_21_pad_groupi_n_1076);
  and csa_tree_add_117_21_pad_groupi_g3298(csa_tree_add_117_21_pad_groupi_n_1100 ,csa_tree_add_117_21_pad_groupi_n_1068 ,csa_tree_add_117_21_pad_groupi_n_1076);
  and csa_tree_add_117_21_pad_groupi_g3299(csa_tree_add_117_21_pad_groupi_n_1099 ,csa_tree_add_117_21_pad_groupi_n_1054 ,csa_tree_add_117_21_pad_groupi_n_1075);
  or csa_tree_add_117_21_pad_groupi_g3300(csa_tree_add_117_21_pad_groupi_n_1109 ,csa_tree_add_117_21_pad_groupi_n_1066 ,csa_tree_add_117_21_pad_groupi_n_1081);
  or csa_tree_add_117_21_pad_groupi_g3301(csa_tree_add_117_21_pad_groupi_n_1108 ,csa_tree_add_117_21_pad_groupi_n_1064 ,csa_tree_add_117_21_pad_groupi_n_1083);
  or csa_tree_add_117_21_pad_groupi_g3302(csa_tree_add_117_21_pad_groupi_n_1107 ,csa_tree_add_117_21_pad_groupi_n_1049 ,csa_tree_add_117_21_pad_groupi_n_1074);
  or csa_tree_add_117_21_pad_groupi_g3303(csa_tree_add_117_21_pad_groupi_n_1106 ,csa_tree_add_117_21_pad_groupi_n_1059 ,csa_tree_add_117_21_pad_groupi_n_1072);
  or csa_tree_add_117_21_pad_groupi_g3304(csa_tree_add_117_21_pad_groupi_n_1105 ,csa_tree_add_117_21_pad_groupi_n_1057 ,csa_tree_add_117_21_pad_groupi_n_1079);
  and csa_tree_add_117_21_pad_groupi_g3305(csa_tree_add_117_21_pad_groupi_n_1090 ,csa_tree_add_117_21_pad_groupi_n_1086 ,csa_tree_add_117_21_pad_groupi_n_1078);
  or csa_tree_add_117_21_pad_groupi_g3306(csa_tree_add_117_21_pad_groupi_n_1089 ,csa_tree_add_117_21_pad_groupi_n_1086 ,csa_tree_add_117_21_pad_groupi_n_1078);
  xnor csa_tree_add_117_21_pad_groupi_g3307(csa_tree_add_117_21_pad_groupi_n_1088 ,csa_tree_add_117_21_pad_groupi_n_1069 ,csa_tree_add_117_21_pad_groupi_n_1013);
  and csa_tree_add_117_21_pad_groupi_g3308(csa_tree_add_117_21_pad_groupi_n_1098 ,csa_tree_add_117_21_pad_groupi_n_998 ,csa_tree_add_117_21_pad_groupi_n_1073);
  xnor csa_tree_add_117_21_pad_groupi_g3309(csa_tree_add_117_21_pad_groupi_n_1097 ,csa_tree_add_117_21_pad_groupi_n_1026 ,csa_tree_add_117_21_pad_groupi_n_1043);
  xnor csa_tree_add_117_21_pad_groupi_g3310(csa_tree_add_117_21_pad_groupi_n_1096 ,csa_tree_add_117_21_pad_groupi_n_1022 ,csa_tree_add_117_21_pad_groupi_n_1042);
  xnor csa_tree_add_117_21_pad_groupi_g3311(csa_tree_add_117_21_pad_groupi_n_1095 ,csa_tree_add_117_21_pad_groupi_n_1017 ,csa_tree_add_117_21_pad_groupi_n_1041);
  xnor csa_tree_add_117_21_pad_groupi_g3312(csa_tree_add_117_21_pad_groupi_n_1094 ,csa_tree_add_117_21_pad_groupi_n_1025 ,csa_tree_add_117_21_pad_groupi_n_1040);
  xnor csa_tree_add_117_21_pad_groupi_g3313(csa_tree_add_117_21_pad_groupi_n_1093 ,csa_tree_add_117_21_pad_groupi_n_1023 ,csa_tree_add_117_21_pad_groupi_n_1048);
  xnor csa_tree_add_117_21_pad_groupi_g3314(csa_tree_add_117_21_pad_groupi_n_1092 ,csa_tree_add_117_21_pad_groupi_n_1016 ,csa_tree_add_117_21_pad_groupi_n_1044);
  xnor csa_tree_add_117_21_pad_groupi_g3315(csa_tree_add_117_21_pad_groupi_n_1091 ,csa_tree_add_117_21_pad_groupi_n_1015 ,csa_tree_add_117_21_pad_groupi_n_1046);
  not csa_tree_add_117_21_pad_groupi_g3316(csa_tree_add_117_21_pad_groupi_n_1085 ,csa_tree_add_117_21_pad_groupi_n_1084);
  nor csa_tree_add_117_21_pad_groupi_g3317(csa_tree_add_117_21_pad_groupi_n_1083 ,csa_tree_add_117_21_pad_groupi_n_1010 ,csa_tree_add_117_21_pad_groupi_n_1061);
  nor csa_tree_add_117_21_pad_groupi_g3318(csa_tree_add_117_21_pad_groupi_n_1082 ,csa_tree_add_117_21_pad_groupi_n_1069 ,csa_tree_add_117_21_pad_groupi_n_1014);
  nor csa_tree_add_117_21_pad_groupi_g3319(csa_tree_add_117_21_pad_groupi_n_1081 ,csa_tree_add_117_21_pad_groupi_n_1008 ,csa_tree_add_117_21_pad_groupi_n_1065);
  and csa_tree_add_117_21_pad_groupi_g3320(csa_tree_add_117_21_pad_groupi_n_1080 ,csa_tree_add_117_21_pad_groupi_n_1069 ,csa_tree_add_117_21_pad_groupi_n_1014);
  nor csa_tree_add_117_21_pad_groupi_g3321(csa_tree_add_117_21_pad_groupi_n_1079 ,csa_tree_add_117_21_pad_groupi_n_1007 ,csa_tree_add_117_21_pad_groupi_n_1056);
  or csa_tree_add_117_21_pad_groupi_g3322(csa_tree_add_117_21_pad_groupi_n_1087 ,csa_tree_add_117_21_pad_groupi_n_1033 ,csa_tree_add_117_21_pad_groupi_n_1060);
  or csa_tree_add_117_21_pad_groupi_g3323(csa_tree_add_117_21_pad_groupi_n_1086 ,csa_tree_add_117_21_pad_groupi_n_1032 ,csa_tree_add_117_21_pad_groupi_n_1055);
  or csa_tree_add_117_21_pad_groupi_g3324(csa_tree_add_117_21_pad_groupi_n_1084 ,csa_tree_add_117_21_pad_groupi_n_927 ,csa_tree_add_117_21_pad_groupi_n_1062);
  nor csa_tree_add_117_21_pad_groupi_g3325(csa_tree_add_117_21_pad_groupi_n_1074 ,csa_tree_add_117_21_pad_groupi_n_1006 ,csa_tree_add_117_21_pad_groupi_n_1051);
  or csa_tree_add_117_21_pad_groupi_g3326(csa_tree_add_117_21_pad_groupi_n_1073 ,csa_tree_add_117_21_pad_groupi_n_989 ,csa_tree_add_117_21_pad_groupi_n_1050);
  nor csa_tree_add_117_21_pad_groupi_g3327(csa_tree_add_117_21_pad_groupi_n_1072 ,csa_tree_add_117_21_pad_groupi_n_1005 ,csa_tree_add_117_21_pad_groupi_n_1058);
  xnor csa_tree_add_117_21_pad_groupi_g3328(csa_tree_add_117_21_pad_groupi_n_1071 ,csa_tree_add_117_21_pad_groupi_n_1019 ,csa_tree_add_117_21_pad_groupi_n_1000);
  xnor csa_tree_add_117_21_pad_groupi_g3329(csa_tree_add_117_21_pad_groupi_n_1070 ,csa_tree_add_117_21_pad_groupi_n_1039 ,csa_tree_add_117_21_pad_groupi_n_1021);
  xnor csa_tree_add_117_21_pad_groupi_g3330(csa_tree_add_117_21_pad_groupi_n_1078 ,csa_tree_add_117_21_pad_groupi_n_1009 ,csa_tree_add_117_21_pad_groupi_n_1027);
  xnor csa_tree_add_117_21_pad_groupi_g3331(csa_tree_add_117_21_pad_groupi_n_1077 ,csa_tree_add_117_21_pad_groupi_n_1024 ,csa_tree_add_117_21_pad_groupi_n_961);
  xnor csa_tree_add_117_21_pad_groupi_g3332(csa_tree_add_117_21_pad_groupi_n_1076 ,csa_tree_add_117_21_pad_groupi_n_933 ,csa_tree_add_117_21_pad_groupi_n_1011);
  xnor csa_tree_add_117_21_pad_groupi_g3333(csa_tree_add_117_21_pad_groupi_n_1075 ,csa_tree_add_117_21_pad_groupi_n_982 ,csa_tree_add_117_21_pad_groupi_n_1012);
  or csa_tree_add_117_21_pad_groupi_g3334(csa_tree_add_117_21_pad_groupi_n_1067 ,csa_tree_add_117_21_pad_groupi_n_999 ,csa_tree_add_117_21_pad_groupi_n_1018);
  nor csa_tree_add_117_21_pad_groupi_g3335(csa_tree_add_117_21_pad_groupi_n_1066 ,csa_tree_add_117_21_pad_groupi_n_878 ,csa_tree_add_117_21_pad_groupi_n_1022);
  and csa_tree_add_117_21_pad_groupi_g3336(csa_tree_add_117_21_pad_groupi_n_1065 ,csa_tree_add_117_21_pad_groupi_n_878 ,csa_tree_add_117_21_pad_groupi_n_1022);
  nor csa_tree_add_117_21_pad_groupi_g3337(csa_tree_add_117_21_pad_groupi_n_1064 ,csa_tree_add_117_21_pad_groupi_n_877 ,csa_tree_add_117_21_pad_groupi_n_1017);
  nor csa_tree_add_117_21_pad_groupi_g3338(csa_tree_add_117_21_pad_groupi_n_1063 ,csa_tree_add_117_21_pad_groupi_n_1000 ,csa_tree_add_117_21_pad_groupi_n_1019);
  and csa_tree_add_117_21_pad_groupi_g3339(csa_tree_add_117_21_pad_groupi_n_1062 ,csa_tree_add_117_21_pad_groupi_n_926 ,csa_tree_add_117_21_pad_groupi_n_1024);
  and csa_tree_add_117_21_pad_groupi_g3340(csa_tree_add_117_21_pad_groupi_n_1061 ,csa_tree_add_117_21_pad_groupi_n_877 ,csa_tree_add_117_21_pad_groupi_n_1017);
  nor csa_tree_add_117_21_pad_groupi_g3341(csa_tree_add_117_21_pad_groupi_n_1060 ,csa_tree_add_117_21_pad_groupi_n_1037 ,csa_tree_add_117_21_pad_groupi_n_1025);
  nor csa_tree_add_117_21_pad_groupi_g3342(csa_tree_add_117_21_pad_groupi_n_1059 ,csa_tree_add_117_21_pad_groupi_n_874 ,csa_tree_add_117_21_pad_groupi_n_1023);
  and csa_tree_add_117_21_pad_groupi_g3343(csa_tree_add_117_21_pad_groupi_n_1058 ,csa_tree_add_117_21_pad_groupi_n_874 ,csa_tree_add_117_21_pad_groupi_n_1023);
  nor csa_tree_add_117_21_pad_groupi_g3344(csa_tree_add_117_21_pad_groupi_n_1057 ,csa_tree_add_117_21_pad_groupi_n_873 ,csa_tree_add_117_21_pad_groupi_n_1016);
  and csa_tree_add_117_21_pad_groupi_g3345(csa_tree_add_117_21_pad_groupi_n_1056 ,csa_tree_add_117_21_pad_groupi_n_873 ,csa_tree_add_117_21_pad_groupi_n_1016);
  nor csa_tree_add_117_21_pad_groupi_g3346(csa_tree_add_117_21_pad_groupi_n_1055 ,csa_tree_add_117_21_pad_groupi_n_1030 ,csa_tree_add_117_21_pad_groupi_n_1026);
  and csa_tree_add_117_21_pad_groupi_g3347(csa_tree_add_117_21_pad_groupi_n_1069 ,csa_tree_add_117_21_pad_groupi_n_993 ,csa_tree_add_117_21_pad_groupi_n_1036);
  and csa_tree_add_117_21_pad_groupi_g3348(csa_tree_add_117_21_pad_groupi_n_1068 ,csa_tree_add_117_21_pad_groupi_n_991 ,csa_tree_add_117_21_pad_groupi_n_1034);
  or csa_tree_add_117_21_pad_groupi_g3349(csa_tree_add_117_21_pad_groupi_n_1053 ,csa_tree_add_117_21_pad_groupi_n_1020 ,csa_tree_add_117_21_pad_groupi_n_1038);
  nor csa_tree_add_117_21_pad_groupi_g3350(csa_tree_add_117_21_pad_groupi_n_1052 ,csa_tree_add_117_21_pad_groupi_n_1021 ,csa_tree_add_117_21_pad_groupi_n_1039);
  nor csa_tree_add_117_21_pad_groupi_g3351(csa_tree_add_117_21_pad_groupi_n_1051 ,csa_tree_add_117_21_pad_groupi_n_872 ,csa_tree_add_117_21_pad_groupi_n_1015);
  nor csa_tree_add_117_21_pad_groupi_g3352(csa_tree_add_117_21_pad_groupi_n_1050 ,csa_tree_add_117_21_pad_groupi_n_929 ,csa_tree_add_117_21_pad_groupi_n_1028);
  and csa_tree_add_117_21_pad_groupi_g3353(csa_tree_add_117_21_pad_groupi_n_1049 ,csa_tree_add_117_21_pad_groupi_n_872 ,csa_tree_add_117_21_pad_groupi_n_1015);
  xor csa_tree_add_117_21_pad_groupi_g3354(csa_tree_add_117_21_pad_groupi_n_1048 ,csa_tree_add_117_21_pad_groupi_n_1005 ,csa_tree_add_117_21_pad_groupi_n_874);
  xnor csa_tree_add_117_21_pad_groupi_g3355(csa_tree_add_117_21_pad_groupi_n_1047 ,csa_tree_add_117_21_pad_groupi_n_983 ,csa_tree_add_117_21_pad_groupi_n_995);
  xnor csa_tree_add_117_21_pad_groupi_g3356(csa_tree_add_117_21_pad_groupi_n_1046 ,csa_tree_add_117_21_pad_groupi_n_872 ,csa_tree_add_117_21_pad_groupi_n_1006);
  xnor csa_tree_add_117_21_pad_groupi_g3357(csa_tree_add_117_21_pad_groupi_n_1045 ,csa_tree_add_117_21_pad_groupi_n_917 ,csa_tree_add_117_21_pad_groupi_n_986);
  xor csa_tree_add_117_21_pad_groupi_g3358(csa_tree_add_117_21_pad_groupi_n_1044 ,csa_tree_add_117_21_pad_groupi_n_1007 ,csa_tree_add_117_21_pad_groupi_n_873);
  xnor csa_tree_add_117_21_pad_groupi_g3359(csa_tree_add_117_21_pad_groupi_n_1043 ,csa_tree_add_117_21_pad_groupi_n_875 ,csa_tree_add_117_21_pad_groupi_n_1003);
  xor csa_tree_add_117_21_pad_groupi_g3360(csa_tree_add_117_21_pad_groupi_n_1042 ,csa_tree_add_117_21_pad_groupi_n_1008 ,csa_tree_add_117_21_pad_groupi_n_878);
  xor csa_tree_add_117_21_pad_groupi_g3361(csa_tree_add_117_21_pad_groupi_n_1041 ,csa_tree_add_117_21_pad_groupi_n_1010 ,csa_tree_add_117_21_pad_groupi_n_877);
  xnor csa_tree_add_117_21_pad_groupi_g3362(csa_tree_add_117_21_pad_groupi_n_1040 ,csa_tree_add_117_21_pad_groupi_n_876 ,csa_tree_add_117_21_pad_groupi_n_1001);
  or csa_tree_add_117_21_pad_groupi_g3363(csa_tree_add_117_21_pad_groupi_n_1054 ,csa_tree_add_117_21_pad_groupi_n_992 ,csa_tree_add_117_21_pad_groupi_n_1029);
  not csa_tree_add_117_21_pad_groupi_g3364(csa_tree_add_117_21_pad_groupi_n_1038 ,csa_tree_add_117_21_pad_groupi_n_1039);
  and csa_tree_add_117_21_pad_groupi_g3365(csa_tree_add_117_21_pad_groupi_n_1037 ,csa_tree_add_117_21_pad_groupi_n_876 ,csa_tree_add_117_21_pad_groupi_n_1002);
  or csa_tree_add_117_21_pad_groupi_g3366(csa_tree_add_117_21_pad_groupi_n_1036 ,csa_tree_add_117_21_pad_groupi_n_933 ,csa_tree_add_117_21_pad_groupi_n_990);
  and csa_tree_add_117_21_pad_groupi_g3367(csa_tree_add_117_21_pad_groupi_n_1035 ,csa_tree_add_117_21_pad_groupi_n_984 ,csa_tree_add_117_21_pad_groupi_n_995);
  or csa_tree_add_117_21_pad_groupi_g3368(csa_tree_add_117_21_pad_groupi_n_1034 ,csa_tree_add_117_21_pad_groupi_n_967 ,csa_tree_add_117_21_pad_groupi_n_988);
  nor csa_tree_add_117_21_pad_groupi_g3369(csa_tree_add_117_21_pad_groupi_n_1033 ,csa_tree_add_117_21_pad_groupi_n_876 ,csa_tree_add_117_21_pad_groupi_n_1002);
  nor csa_tree_add_117_21_pad_groupi_g3370(csa_tree_add_117_21_pad_groupi_n_1032 ,csa_tree_add_117_21_pad_groupi_n_875 ,csa_tree_add_117_21_pad_groupi_n_1004);
  nor csa_tree_add_117_21_pad_groupi_g3371(csa_tree_add_117_21_pad_groupi_n_1031 ,csa_tree_add_117_21_pad_groupi_n_984 ,csa_tree_add_117_21_pad_groupi_n_995);
  and csa_tree_add_117_21_pad_groupi_g3372(csa_tree_add_117_21_pad_groupi_n_1030 ,csa_tree_add_117_21_pad_groupi_n_875 ,csa_tree_add_117_21_pad_groupi_n_1004);
  nor csa_tree_add_117_21_pad_groupi_g3373(csa_tree_add_117_21_pad_groupi_n_1029 ,csa_tree_add_117_21_pad_groupi_n_1009 ,csa_tree_add_117_21_pad_groupi_n_994);
  nor csa_tree_add_117_21_pad_groupi_g3374(csa_tree_add_117_21_pad_groupi_n_1028 ,csa_tree_add_117_21_pad_groupi_n_928 ,csa_tree_add_117_21_pad_groupi_n_997);
  xnor csa_tree_add_117_21_pad_groupi_g3375(csa_tree_add_117_21_pad_groupi_n_1027 ,csa_tree_add_117_21_pad_groupi_n_883 ,csa_tree_add_117_21_pad_groupi_n_965);
  and csa_tree_add_117_21_pad_groupi_g3376(csa_tree_add_117_21_pad_groupi_n_1039 ,csa_tree_add_117_21_pad_groupi_n_921 ,csa_tree_add_117_21_pad_groupi_n_987);
  not csa_tree_add_117_21_pad_groupi_g3377(csa_tree_add_117_21_pad_groupi_n_1021 ,csa_tree_add_117_21_pad_groupi_n_1020);
  not csa_tree_add_117_21_pad_groupi_g3378(csa_tree_add_117_21_pad_groupi_n_1019 ,csa_tree_add_117_21_pad_groupi_n_1018);
  not csa_tree_add_117_21_pad_groupi_g3379(csa_tree_add_117_21_pad_groupi_n_1014 ,csa_tree_add_117_21_pad_groupi_n_1013);
  xnor csa_tree_add_117_21_pad_groupi_g3380(csa_tree_add_117_21_pad_groupi_n_1012 ,csa_tree_add_117_21_pad_groupi_n_910 ,csa_tree_add_117_21_pad_groupi_n_967);
  xnor csa_tree_add_117_21_pad_groupi_g3381(csa_tree_add_117_21_pad_groupi_n_1011 ,csa_tree_add_117_21_pad_groupi_n_964 ,csa_tree_add_117_21_pad_groupi_n_851);
  xnor csa_tree_add_117_21_pad_groupi_g3382(csa_tree_add_117_21_pad_groupi_n_1026 ,csa_tree_add_117_21_pad_groupi_n_850 ,csa_tree_add_117_21_pad_groupi_n_953);
  xnor csa_tree_add_117_21_pad_groupi_g3383(csa_tree_add_117_21_pad_groupi_n_1025 ,csa_tree_add_117_21_pad_groupi_n_863 ,csa_tree_add_117_21_pad_groupi_n_957);
  xnor csa_tree_add_117_21_pad_groupi_g3384(csa_tree_add_117_21_pad_groupi_n_1024 ,csa_tree_add_117_21_pad_groupi_n_853 ,csa_tree_add_117_21_pad_groupi_n_952);
  xnor csa_tree_add_117_21_pad_groupi_g3385(csa_tree_add_117_21_pad_groupi_n_1023 ,csa_tree_add_117_21_pad_groupi_n_861 ,csa_tree_add_117_21_pad_groupi_n_955);
  xnor csa_tree_add_117_21_pad_groupi_g3386(csa_tree_add_117_21_pad_groupi_n_1022 ,csa_tree_add_117_21_pad_groupi_n_859 ,csa_tree_add_117_21_pad_groupi_n_960);
  xnor csa_tree_add_117_21_pad_groupi_g3387(csa_tree_add_117_21_pad_groupi_n_1020 ,csa_tree_add_117_21_pad_groupi_n_911 ,csa_tree_add_117_21_pad_groupi_n_956);
  xnor csa_tree_add_117_21_pad_groupi_g3388(csa_tree_add_117_21_pad_groupi_n_1018 ,csa_tree_add_117_21_pad_groupi_n_902 ,csa_tree_add_117_21_pad_groupi_n_959);
  xnor csa_tree_add_117_21_pad_groupi_g3389(csa_tree_add_117_21_pad_groupi_n_1017 ,csa_tree_add_117_21_pad_groupi_n_864 ,csa_tree_add_117_21_pad_groupi_n_958);
  xnor csa_tree_add_117_21_pad_groupi_g3390(csa_tree_add_117_21_pad_groupi_n_1016 ,csa_tree_add_117_21_pad_groupi_n_860 ,csa_tree_add_117_21_pad_groupi_n_954);
  xnor csa_tree_add_117_21_pad_groupi_g3391(csa_tree_add_117_21_pad_groupi_n_1015 ,csa_tree_add_117_21_pad_groupi_n_849 ,csa_tree_add_117_21_pad_groupi_n_962);
  xnor csa_tree_add_117_21_pad_groupi_g3392(csa_tree_add_117_21_pad_groupi_n_1013 ,csa_tree_add_117_21_pad_groupi_n_985 ,csa_tree_add_117_21_pad_groupi_n_963);
  not csa_tree_add_117_21_pad_groupi_g3393(csa_tree_add_117_21_pad_groupi_n_1004 ,csa_tree_add_117_21_pad_groupi_n_1003);
  not csa_tree_add_117_21_pad_groupi_g3394(csa_tree_add_117_21_pad_groupi_n_1002 ,csa_tree_add_117_21_pad_groupi_n_1001);
  not csa_tree_add_117_21_pad_groupi_g3395(csa_tree_add_117_21_pad_groupi_n_999 ,csa_tree_add_117_21_pad_groupi_n_1000);
  or csa_tree_add_117_21_pad_groupi_g3396(csa_tree_add_117_21_pad_groupi_n_998 ,csa_tree_add_117_21_pad_groupi_n_870 ,csa_tree_add_117_21_pad_groupi_n_968);
  nor csa_tree_add_117_21_pad_groupi_g3397(csa_tree_add_117_21_pad_groupi_n_997 ,csa_tree_add_117_21_pad_groupi_n_2 ,csa_tree_add_117_21_pad_groupi_n_970);
  and csa_tree_add_117_21_pad_groupi_g3398(csa_tree_add_117_21_pad_groupi_n_1010 ,csa_tree_add_117_21_pad_groupi_n_945 ,csa_tree_add_117_21_pad_groupi_n_975);
  and csa_tree_add_117_21_pad_groupi_g3399(csa_tree_add_117_21_pad_groupi_n_1009 ,csa_tree_add_117_21_pad_groupi_n_949 ,csa_tree_add_117_21_pad_groupi_n_977);
  and csa_tree_add_117_21_pad_groupi_g3400(csa_tree_add_117_21_pad_groupi_n_1008 ,csa_tree_add_117_21_pad_groupi_n_947 ,csa_tree_add_117_21_pad_groupi_n_976);
  and csa_tree_add_117_21_pad_groupi_g3401(csa_tree_add_117_21_pad_groupi_n_1007 ,csa_tree_add_117_21_pad_groupi_n_938 ,csa_tree_add_117_21_pad_groupi_n_973);
  and csa_tree_add_117_21_pad_groupi_g3402(csa_tree_add_117_21_pad_groupi_n_1006 ,csa_tree_add_117_21_pad_groupi_n_935 ,csa_tree_add_117_21_pad_groupi_n_979);
  and csa_tree_add_117_21_pad_groupi_g3403(csa_tree_add_117_21_pad_groupi_n_1005 ,csa_tree_add_117_21_pad_groupi_n_940 ,csa_tree_add_117_21_pad_groupi_n_980);
  or csa_tree_add_117_21_pad_groupi_g3404(csa_tree_add_117_21_pad_groupi_n_1003 ,csa_tree_add_117_21_pad_groupi_n_941 ,csa_tree_add_117_21_pad_groupi_n_972);
  or csa_tree_add_117_21_pad_groupi_g3405(csa_tree_add_117_21_pad_groupi_n_1001 ,csa_tree_add_117_21_pad_groupi_n_943 ,csa_tree_add_117_21_pad_groupi_n_974);
  and csa_tree_add_117_21_pad_groupi_g3406(csa_tree_add_117_21_pad_groupi_n_1000 ,csa_tree_add_117_21_pad_groupi_n_942 ,csa_tree_add_117_21_pad_groupi_n_978);
  and csa_tree_add_117_21_pad_groupi_g3407(csa_tree_add_117_21_pad_groupi_n_994 ,csa_tree_add_117_21_pad_groupi_n_883 ,csa_tree_add_117_21_pad_groupi_n_966);
  or csa_tree_add_117_21_pad_groupi_g3408(csa_tree_add_117_21_pad_groupi_n_993 ,csa_tree_add_117_21_pad_groupi_n_851 ,csa_tree_add_117_21_pad_groupi_n_964);
  nor csa_tree_add_117_21_pad_groupi_g3409(csa_tree_add_117_21_pad_groupi_n_992 ,csa_tree_add_117_21_pad_groupi_n_883 ,csa_tree_add_117_21_pad_groupi_n_966);
  or csa_tree_add_117_21_pad_groupi_g3410(csa_tree_add_117_21_pad_groupi_n_991 ,csa_tree_add_117_21_pad_groupi_n_909 ,csa_tree_add_117_21_pad_groupi_n_982);
  and csa_tree_add_117_21_pad_groupi_g3411(csa_tree_add_117_21_pad_groupi_n_990 ,csa_tree_add_117_21_pad_groupi_n_851 ,csa_tree_add_117_21_pad_groupi_n_964);
  and csa_tree_add_117_21_pad_groupi_g3412(csa_tree_add_117_21_pad_groupi_n_989 ,csa_tree_add_117_21_pad_groupi_n_870 ,csa_tree_add_117_21_pad_groupi_n_968);
  nor csa_tree_add_117_21_pad_groupi_g3413(csa_tree_add_117_21_pad_groupi_n_988 ,csa_tree_add_117_21_pad_groupi_n_910 ,csa_tree_add_117_21_pad_groupi_n_981);
  or csa_tree_add_117_21_pad_groupi_g3414(csa_tree_add_117_21_pad_groupi_n_987 ,csa_tree_add_117_21_pad_groupi_n_985 ,csa_tree_add_117_21_pad_groupi_n_919);
  nor csa_tree_add_117_21_pad_groupi_g3415(csa_tree_add_117_21_pad_groupi_n_986 ,csa_tree_add_117_21_pad_groupi_n_920 ,csa_tree_add_117_21_pad_groupi_n_971);
  and csa_tree_add_117_21_pad_groupi_g3416(csa_tree_add_117_21_pad_groupi_n_996 ,csa_tree_add_117_21_pad_groupi_n_918 ,csa_tree_add_117_21_pad_groupi_n_969);
  xnor csa_tree_add_117_21_pad_groupi_g3417(csa_tree_add_117_21_pad_groupi_n_995 ,csa_tree_add_117_21_pad_groupi_n_879 ,csa_tree_add_117_21_pad_groupi_n_916);
  not csa_tree_add_117_21_pad_groupi_g3418(csa_tree_add_117_21_pad_groupi_n_984 ,csa_tree_add_117_21_pad_groupi_n_983);
  not csa_tree_add_117_21_pad_groupi_g3419(csa_tree_add_117_21_pad_groupi_n_981 ,csa_tree_add_117_21_pad_groupi_n_982);
  or csa_tree_add_117_21_pad_groupi_g3420(csa_tree_add_117_21_pad_groupi_n_980 ,csa_tree_add_117_21_pad_groupi_n_840 ,csa_tree_add_117_21_pad_groupi_n_939);
  or csa_tree_add_117_21_pad_groupi_g3421(csa_tree_add_117_21_pad_groupi_n_979 ,csa_tree_add_117_21_pad_groupi_n_854 ,csa_tree_add_117_21_pad_groupi_n_934);
  or csa_tree_add_117_21_pad_groupi_g3422(csa_tree_add_117_21_pad_groupi_n_978 ,csa_tree_add_117_21_pad_groupi_n_852 ,csa_tree_add_117_21_pad_groupi_n_950);
  or csa_tree_add_117_21_pad_groupi_g3423(csa_tree_add_117_21_pad_groupi_n_977 ,csa_tree_add_117_21_pad_groupi_n_839 ,csa_tree_add_117_21_pad_groupi_n_948);
  or csa_tree_add_117_21_pad_groupi_g3424(csa_tree_add_117_21_pad_groupi_n_976 ,csa_tree_add_117_21_pad_groupi_n_837 ,csa_tree_add_117_21_pad_groupi_n_946);
  or csa_tree_add_117_21_pad_groupi_g3425(csa_tree_add_117_21_pad_groupi_n_975 ,csa_tree_add_117_21_pad_groupi_n_833 ,csa_tree_add_117_21_pad_groupi_n_944);
  nor csa_tree_add_117_21_pad_groupi_g3426(csa_tree_add_117_21_pad_groupi_n_974 ,csa_tree_add_117_21_pad_groupi_n_834 ,csa_tree_add_117_21_pad_groupi_n_951);
  or csa_tree_add_117_21_pad_groupi_g3427(csa_tree_add_117_21_pad_groupi_n_973 ,csa_tree_add_117_21_pad_groupi_n_867 ,csa_tree_add_117_21_pad_groupi_n_937);
  nor csa_tree_add_117_21_pad_groupi_g3428(csa_tree_add_117_21_pad_groupi_n_972 ,csa_tree_add_117_21_pad_groupi_n_836 ,csa_tree_add_117_21_pad_groupi_n_936);
  nor csa_tree_add_117_21_pad_groupi_g3429(csa_tree_add_117_21_pad_groupi_n_971 ,csa_tree_add_117_21_pad_groupi_n_911 ,csa_tree_add_117_21_pad_groupi_n_922);
  nor csa_tree_add_117_21_pad_groupi_g3430(csa_tree_add_117_21_pad_groupi_n_970 ,csa_tree_add_117_21_pad_groupi_n_930 ,csa_tree_add_117_21_pad_groupi_n_931);
  or csa_tree_add_117_21_pad_groupi_g3431(csa_tree_add_117_21_pad_groupi_n_969 ,csa_tree_add_117_21_pad_groupi_n_869 ,csa_tree_add_117_21_pad_groupi_n_932);
  and csa_tree_add_117_21_pad_groupi_g3432(csa_tree_add_117_21_pad_groupi_n_985 ,csa_tree_add_117_21_pad_groupi_n_842 ,csa_tree_add_117_21_pad_groupi_n_925);
  or csa_tree_add_117_21_pad_groupi_g3433(csa_tree_add_117_21_pad_groupi_n_983 ,csa_tree_add_117_21_pad_groupi_n_721 ,csa_tree_add_117_21_pad_groupi_n_924);
  and csa_tree_add_117_21_pad_groupi_g3434(csa_tree_add_117_21_pad_groupi_n_982 ,csa_tree_add_117_21_pad_groupi_n_894 ,csa_tree_add_117_21_pad_groupi_n_923);
  not csa_tree_add_117_21_pad_groupi_g3435(csa_tree_add_117_21_pad_groupi_n_966 ,csa_tree_add_117_21_pad_groupi_n_965);
  xnor csa_tree_add_117_21_pad_groupi_g3436(csa_tree_add_117_21_pad_groupi_n_963 ,csa_tree_add_117_21_pad_groupi_n_866 ,csa_tree_add_117_21_pad_groupi_n_906);
  xnor csa_tree_add_117_21_pad_groupi_g3437(csa_tree_add_117_21_pad_groupi_n_962 ,csa_tree_add_117_21_pad_groupi_n_867 ,csa_tree_add_117_21_pad_groupi_n_887);
  xnor csa_tree_add_117_21_pad_groupi_g3438(csa_tree_add_117_21_pad_groupi_n_961 ,csa_tree_add_117_21_pad_groupi_n_904 ,csa_tree_add_117_21_pad_groupi_n_908);
  xnor csa_tree_add_117_21_pad_groupi_g3439(csa_tree_add_117_21_pad_groupi_n_960 ,csa_tree_add_117_21_pad_groupi_n_889 ,csa_tree_add_117_21_pad_groupi_n_836);
  xnor csa_tree_add_117_21_pad_groupi_g3440(csa_tree_add_117_21_pad_groupi_n_959 ,csa_tree_add_117_21_pad_groupi_n_882 ,csa_tree_add_117_21_pad_groupi_n_869);
  xnor csa_tree_add_117_21_pad_groupi_g3441(csa_tree_add_117_21_pad_groupi_n_958 ,csa_tree_add_117_21_pad_groupi_n_898 ,csa_tree_add_117_21_pad_groupi_n_837);
  xnor csa_tree_add_117_21_pad_groupi_g3442(csa_tree_add_117_21_pad_groupi_n_957 ,csa_tree_add_117_21_pad_groupi_n_897 ,csa_tree_add_117_21_pad_groupi_n_833);
  xnor csa_tree_add_117_21_pad_groupi_g3443(csa_tree_add_117_21_pad_groupi_n_956 ,csa_tree_add_117_21_pad_groupi_n_831 ,csa_tree_add_117_21_pad_groupi_n_900);
  xnor csa_tree_add_117_21_pad_groupi_g3444(csa_tree_add_117_21_pad_groupi_n_955 ,csa_tree_add_117_21_pad_groupi_n_880 ,csa_tree_add_117_21_pad_groupi_n_834);
  xnor csa_tree_add_117_21_pad_groupi_g3445(csa_tree_add_117_21_pad_groupi_n_954 ,csa_tree_add_117_21_pad_groupi_n_888 ,csa_tree_add_117_21_pad_groupi_n_840);
  xnor csa_tree_add_117_21_pad_groupi_g3446(csa_tree_add_117_21_pad_groupi_n_953 ,csa_tree_add_117_21_pad_groupi_n_884 ,csa_tree_add_117_21_pad_groupi_n_839);
  xnor csa_tree_add_117_21_pad_groupi_g3447(csa_tree_add_117_21_pad_groupi_n_968 ,csa_tree_add_117_21_pad_groupi_n_912 ,csa_tree_add_117_21_pad_groupi_n_789);
  xnor csa_tree_add_117_21_pad_groupi_g3448(csa_tree_add_117_21_pad_groupi_n_952 ,csa_tree_add_117_21_pad_groupi_n_885 ,csa_tree_add_117_21_pad_groupi_n_620);
  xnor csa_tree_add_117_21_pad_groupi_g3449(csa_tree_add_117_21_pad_groupi_n_967 ,csa_tree_add_117_21_pad_groupi_n_868 ,csa_tree_add_117_21_pad_groupi_n_871);
  xnor csa_tree_add_117_21_pad_groupi_g3450(csa_tree_add_117_21_pad_groupi_n_965 ,csa_tree_add_117_21_pad_groupi_n_862 ,csa_tree_add_117_21_pad_groupi_n_892);
  xnor csa_tree_add_117_21_pad_groupi_g3451(csa_tree_add_117_21_pad_groupi_n_964 ,csa_tree_add_117_21_pad_groupi_n_890 ,csa_tree_add_117_21_pad_groupi_n_891);
  and csa_tree_add_117_21_pad_groupi_g3452(csa_tree_add_117_21_pad_groupi_n_951 ,csa_tree_add_117_21_pad_groupi_n_880 ,csa_tree_add_117_21_pad_groupi_n_861);
  and csa_tree_add_117_21_pad_groupi_g3453(csa_tree_add_117_21_pad_groupi_n_950 ,csa_tree_add_117_21_pad_groupi_n_847 ,csa_tree_add_117_21_pad_groupi_n_879);
  or csa_tree_add_117_21_pad_groupi_g3454(csa_tree_add_117_21_pad_groupi_n_949 ,csa_tree_add_117_21_pad_groupi_n_884 ,csa_tree_add_117_21_pad_groupi_n_850);
  and csa_tree_add_117_21_pad_groupi_g3455(csa_tree_add_117_21_pad_groupi_n_948 ,csa_tree_add_117_21_pad_groupi_n_884 ,csa_tree_add_117_21_pad_groupi_n_850);
  or csa_tree_add_117_21_pad_groupi_g3456(csa_tree_add_117_21_pad_groupi_n_947 ,csa_tree_add_117_21_pad_groupi_n_898 ,csa_tree_add_117_21_pad_groupi_n_864);
  and csa_tree_add_117_21_pad_groupi_g3457(csa_tree_add_117_21_pad_groupi_n_946 ,csa_tree_add_117_21_pad_groupi_n_898 ,csa_tree_add_117_21_pad_groupi_n_864);
  or csa_tree_add_117_21_pad_groupi_g3458(csa_tree_add_117_21_pad_groupi_n_945 ,csa_tree_add_117_21_pad_groupi_n_897 ,csa_tree_add_117_21_pad_groupi_n_863);
  and csa_tree_add_117_21_pad_groupi_g3459(csa_tree_add_117_21_pad_groupi_n_944 ,csa_tree_add_117_21_pad_groupi_n_897 ,csa_tree_add_117_21_pad_groupi_n_863);
  nor csa_tree_add_117_21_pad_groupi_g3460(csa_tree_add_117_21_pad_groupi_n_943 ,csa_tree_add_117_21_pad_groupi_n_880 ,csa_tree_add_117_21_pad_groupi_n_861);
  or csa_tree_add_117_21_pad_groupi_g3461(csa_tree_add_117_21_pad_groupi_n_942 ,csa_tree_add_117_21_pad_groupi_n_847 ,csa_tree_add_117_21_pad_groupi_n_879);
  nor csa_tree_add_117_21_pad_groupi_g3462(csa_tree_add_117_21_pad_groupi_n_941 ,csa_tree_add_117_21_pad_groupi_n_889 ,csa_tree_add_117_21_pad_groupi_n_859);
  or csa_tree_add_117_21_pad_groupi_g3463(csa_tree_add_117_21_pad_groupi_n_940 ,csa_tree_add_117_21_pad_groupi_n_888 ,csa_tree_add_117_21_pad_groupi_n_860);
  and csa_tree_add_117_21_pad_groupi_g3464(csa_tree_add_117_21_pad_groupi_n_939 ,csa_tree_add_117_21_pad_groupi_n_888 ,csa_tree_add_117_21_pad_groupi_n_860);
  or csa_tree_add_117_21_pad_groupi_g3465(csa_tree_add_117_21_pad_groupi_n_938 ,csa_tree_add_117_21_pad_groupi_n_849 ,csa_tree_add_117_21_pad_groupi_n_886);
  nor csa_tree_add_117_21_pad_groupi_g3466(csa_tree_add_117_21_pad_groupi_n_937 ,csa_tree_add_117_21_pad_groupi_n_848 ,csa_tree_add_117_21_pad_groupi_n_887);
  and csa_tree_add_117_21_pad_groupi_g3467(csa_tree_add_117_21_pad_groupi_n_936 ,csa_tree_add_117_21_pad_groupi_n_889 ,csa_tree_add_117_21_pad_groupi_n_859);
  or csa_tree_add_117_21_pad_groupi_g3468(csa_tree_add_117_21_pad_groupi_n_935 ,csa_tree_add_117_21_pad_groupi_n_620 ,csa_tree_add_117_21_pad_groupi_n_885);
  and csa_tree_add_117_21_pad_groupi_g3469(csa_tree_add_117_21_pad_groupi_n_934 ,csa_tree_add_117_21_pad_groupi_n_620 ,csa_tree_add_117_21_pad_groupi_n_885);
  nor csa_tree_add_117_21_pad_groupi_g3470(csa_tree_add_117_21_pad_groupi_n_932 ,csa_tree_add_117_21_pad_groupi_n_881 ,csa_tree_add_117_21_pad_groupi_n_902);
  nor csa_tree_add_117_21_pad_groupi_g3472(csa_tree_add_117_21_pad_groupi_n_931 ,csa_tree_add_117_21_pad_groupi_n_714 ,csa_tree_add_117_21_pad_groupi_n_913);
  nor csa_tree_add_117_21_pad_groupi_g3473(csa_tree_add_117_21_pad_groupi_n_930 ,csa_tree_add_117_21_pad_groupi_n_821 ,csa_tree_add_117_21_pad_groupi_n_893);
  nor csa_tree_add_117_21_pad_groupi_g3474(csa_tree_add_117_21_pad_groupi_n_929 ,csa_tree_add_117_21_pad_groupi_n_855 ,csa_tree_add_117_21_pad_groupi_n_915);
  nor csa_tree_add_117_21_pad_groupi_g3475(csa_tree_add_117_21_pad_groupi_n_928 ,csa_tree_add_117_21_pad_groupi_n_856 ,csa_tree_add_117_21_pad_groupi_n_914);
  nor csa_tree_add_117_21_pad_groupi_g3476(csa_tree_add_117_21_pad_groupi_n_927 ,csa_tree_add_117_21_pad_groupi_n_904 ,csa_tree_add_117_21_pad_groupi_n_907);
  or csa_tree_add_117_21_pad_groupi_g3477(csa_tree_add_117_21_pad_groupi_n_926 ,csa_tree_add_117_21_pad_groupi_n_903 ,csa_tree_add_117_21_pad_groupi_n_908);
  or csa_tree_add_117_21_pad_groupi_g3478(csa_tree_add_117_21_pad_groupi_n_925 ,csa_tree_add_117_21_pad_groupi_n_841 ,csa_tree_add_117_21_pad_groupi_n_890);
  and csa_tree_add_117_21_pad_groupi_g3479(csa_tree_add_117_21_pad_groupi_n_924 ,csa_tree_add_117_21_pad_groupi_n_720 ,csa_tree_add_117_21_pad_groupi_n_912);
  or csa_tree_add_117_21_pad_groupi_g3480(csa_tree_add_117_21_pad_groupi_n_923 ,csa_tree_add_117_21_pad_groupi_n_838 ,csa_tree_add_117_21_pad_groupi_n_895);
  and csa_tree_add_117_21_pad_groupi_g3481(csa_tree_add_117_21_pad_groupi_n_922 ,csa_tree_add_117_21_pad_groupi_n_830 ,csa_tree_add_117_21_pad_groupi_n_900);
  or csa_tree_add_117_21_pad_groupi_g3482(csa_tree_add_117_21_pad_groupi_n_921 ,csa_tree_add_117_21_pad_groupi_n_866 ,csa_tree_add_117_21_pad_groupi_n_905);
  and csa_tree_add_117_21_pad_groupi_g3483(csa_tree_add_117_21_pad_groupi_n_920 ,csa_tree_add_117_21_pad_groupi_n_831 ,csa_tree_add_117_21_pad_groupi_n_899);
  nor csa_tree_add_117_21_pad_groupi_g3484(csa_tree_add_117_21_pad_groupi_n_919 ,csa_tree_add_117_21_pad_groupi_n_865 ,csa_tree_add_117_21_pad_groupi_n_906);
  or csa_tree_add_117_21_pad_groupi_g3485(csa_tree_add_117_21_pad_groupi_n_918 ,csa_tree_add_117_21_pad_groupi_n_882 ,csa_tree_add_117_21_pad_groupi_n_901);
  xnor csa_tree_add_117_21_pad_groupi_g3486(csa_tree_add_117_21_pad_groupi_n_917 ,csa_tree_add_117_21_pad_groupi_n_794 ,csa_tree_add_117_21_pad_groupi_n_857);
  xnor csa_tree_add_117_21_pad_groupi_g3487(csa_tree_add_117_21_pad_groupi_n_916 ,csa_tree_add_117_21_pad_groupi_n_852 ,csa_tree_add_117_21_pad_groupi_n_847);
  and csa_tree_add_117_21_pad_groupi_g3488(csa_tree_add_117_21_pad_groupi_n_933 ,csa_tree_add_117_21_pad_groupi_n_844 ,csa_tree_add_117_21_pad_groupi_n_896);
  not csa_tree_add_117_21_pad_groupi_g3489(csa_tree_add_117_21_pad_groupi_n_915 ,csa_tree_add_117_21_pad_groupi_n_914);
  not csa_tree_add_117_21_pad_groupi_g3491(csa_tree_add_117_21_pad_groupi_n_909 ,csa_tree_add_117_21_pad_groupi_n_910);
  not csa_tree_add_117_21_pad_groupi_g3492(csa_tree_add_117_21_pad_groupi_n_907 ,csa_tree_add_117_21_pad_groupi_n_908);
  not csa_tree_add_117_21_pad_groupi_g3493(csa_tree_add_117_21_pad_groupi_n_905 ,csa_tree_add_117_21_pad_groupi_n_906);
  not csa_tree_add_117_21_pad_groupi_g3494(csa_tree_add_117_21_pad_groupi_n_904 ,csa_tree_add_117_21_pad_groupi_n_903);
  not csa_tree_add_117_21_pad_groupi_g3495(csa_tree_add_117_21_pad_groupi_n_902 ,csa_tree_add_117_21_pad_groupi_n_901);
  not csa_tree_add_117_21_pad_groupi_g3496(csa_tree_add_117_21_pad_groupi_n_899 ,csa_tree_add_117_21_pad_groupi_n_900);
  or csa_tree_add_117_21_pad_groupi_g3497(csa_tree_add_117_21_pad_groupi_n_896 ,csa_tree_add_117_21_pad_groupi_n_845 ,csa_tree_add_117_21_pad_groupi_n_868);
  and csa_tree_add_117_21_pad_groupi_g3498(csa_tree_add_117_21_pad_groupi_n_895 ,csa_tree_add_117_21_pad_groupi_n_806 ,csa_tree_add_117_21_pad_groupi_n_862);
  or csa_tree_add_117_21_pad_groupi_g3499(csa_tree_add_117_21_pad_groupi_n_894 ,csa_tree_add_117_21_pad_groupi_n_806 ,csa_tree_add_117_21_pad_groupi_n_862);
  nor csa_tree_add_117_21_pad_groupi_g3500(csa_tree_add_117_21_pad_groupi_n_893 ,csa_tree_add_117_21_pad_groupi_n_823 ,csa_tree_add_117_21_pad_groupi_n_846);
  xnor csa_tree_add_117_21_pad_groupi_g3501(csa_tree_add_117_21_pad_groupi_n_892 ,csa_tree_add_117_21_pad_groupi_n_838 ,csa_tree_add_117_21_pad_groupi_n_805);
  xnor csa_tree_add_117_21_pad_groupi_g3502(csa_tree_add_117_21_pad_groupi_n_914 ,csa_tree_add_117_21_pad_groupi_n_742 ,csa_tree_add_117_21_pad_groupi_n_779);
  xnor csa_tree_add_117_21_pad_groupi_g3503(csa_tree_add_117_21_pad_groupi_n_913 ,csa_tree_add_117_21_pad_groupi_n_641 ,csa_tree_add_117_21_pad_groupi_n_801);
  xnor csa_tree_add_117_21_pad_groupi_g3504(csa_tree_add_117_21_pad_groupi_n_891 ,csa_tree_add_117_21_pad_groupi_n_829 ,csa_tree_add_117_21_pad_groupi_n_621);
  xnor csa_tree_add_117_21_pad_groupi_g3505(csa_tree_add_117_21_pad_groupi_n_912 ,csa_tree_add_117_21_pad_groupi_n_690 ,csa_tree_add_117_21_pad_groupi_n_802);
  and csa_tree_add_117_21_pad_groupi_g3506(csa_tree_add_117_21_pad_groupi_n_911 ,csa_tree_add_117_21_pad_groupi_n_722 ,csa_tree_add_117_21_pad_groupi_n_843);
  xnor csa_tree_add_117_21_pad_groupi_g3507(csa_tree_add_117_21_pad_groupi_n_910 ,csa_tree_add_117_21_pad_groupi_n_655 ,csa_tree_add_117_21_pad_groupi_n_800);
  xnor csa_tree_add_117_21_pad_groupi_g3508(csa_tree_add_117_21_pad_groupi_n_908 ,csa_tree_add_117_21_pad_groupi_n_625 ,csa_tree_add_117_21_pad_groupi_n_787);
  xnor csa_tree_add_117_21_pad_groupi_g3509(csa_tree_add_117_21_pad_groupi_n_906 ,csa_tree_add_117_21_pad_groupi_n_807 ,csa_tree_add_117_21_pad_groupi_n_799);
  or csa_tree_add_117_21_pad_groupi_g3510(csa_tree_add_117_21_pad_groupi_n_903 ,csa_tree_add_117_21_pad_groupi_n_756 ,csa_tree_add_117_21_pad_groupi_n_858);
  xnor csa_tree_add_117_21_pad_groupi_g3511(csa_tree_add_117_21_pad_groupi_n_901 ,csa_tree_add_117_21_pad_groupi_n_835 ,csa_tree_add_117_21_pad_groupi_n_782);
  xnor csa_tree_add_117_21_pad_groupi_g3512(csa_tree_add_117_21_pad_groupi_n_900 ,csa_tree_add_117_21_pad_groupi_n_622 ,csa_tree_add_117_21_pad_groupi_n_803);
  xnor csa_tree_add_117_21_pad_groupi_g3513(csa_tree_add_117_21_pad_groupi_n_898 ,csa_tree_add_117_21_pad_groupi_n_591 ,csa_tree_add_117_21_pad_groupi_n_797);
  xnor csa_tree_add_117_21_pad_groupi_g3514(csa_tree_add_117_21_pad_groupi_n_897 ,csa_tree_add_117_21_pad_groupi_n_596 ,csa_tree_add_117_21_pad_groupi_n_796);
  not csa_tree_add_117_21_pad_groupi_g3515(csa_tree_add_117_21_pad_groupi_n_887 ,csa_tree_add_117_21_pad_groupi_n_886);
  not csa_tree_add_117_21_pad_groupi_g3516(csa_tree_add_117_21_pad_groupi_n_881 ,csa_tree_add_117_21_pad_groupi_n_882);
  xnor csa_tree_add_117_21_pad_groupi_g3517(csa_tree_add_117_21_pad_groupi_n_871 ,csa_tree_add_117_21_pad_groupi_n_804 ,csa_tree_add_117_21_pad_groupi_n_832);
  xnor csa_tree_add_117_21_pad_groupi_g3518(csa_tree_add_117_21_pad_groupi_n_890 ,csa_tree_add_117_21_pad_groupi_n_632 ,csa_tree_add_117_21_pad_groupi_n_784);
  xnor csa_tree_add_117_21_pad_groupi_g3519(csa_tree_add_117_21_pad_groupi_n_889 ,csa_tree_add_117_21_pad_groupi_n_0 ,csa_tree_add_117_21_pad_groupi_n_792);
  xnor csa_tree_add_117_21_pad_groupi_g3520(csa_tree_add_117_21_pad_groupi_n_888 ,csa_tree_add_117_21_pad_groupi_n_586 ,csa_tree_add_117_21_pad_groupi_n_793);
  xnor csa_tree_add_117_21_pad_groupi_g3521(csa_tree_add_117_21_pad_groupi_n_886 ,csa_tree_add_117_21_pad_groupi_n_604 ,csa_tree_add_117_21_pad_groupi_n_791);
  xnor csa_tree_add_117_21_pad_groupi_g3522(csa_tree_add_117_21_pad_groupi_n_885 ,csa_tree_add_117_21_pad_groupi_n_710 ,csa_tree_add_117_21_pad_groupi_n_790);
  xnor csa_tree_add_117_21_pad_groupi_g3523(csa_tree_add_117_21_pad_groupi_n_884 ,csa_tree_add_117_21_pad_groupi_n_605 ,csa_tree_add_117_21_pad_groupi_n_788);
  xnor csa_tree_add_117_21_pad_groupi_g3524(csa_tree_add_117_21_pad_groupi_n_883 ,csa_tree_add_117_21_pad_groupi_n_659 ,csa_tree_add_117_21_pad_groupi_n_781);
  xnor csa_tree_add_117_21_pad_groupi_g3525(csa_tree_add_117_21_pad_groupi_n_882 ,csa_tree_add_117_21_pad_groupi_n_618 ,csa_tree_add_117_21_pad_groupi_n_783);
  xnor csa_tree_add_117_21_pad_groupi_g3526(csa_tree_add_117_21_pad_groupi_n_880 ,csa_tree_add_117_21_pad_groupi_n_588 ,csa_tree_add_117_21_pad_groupi_n_795);
  xnor csa_tree_add_117_21_pad_groupi_g3527(csa_tree_add_117_21_pad_groupi_n_879 ,csa_tree_add_117_21_pad_groupi_n_692 ,csa_tree_add_117_21_pad_groupi_n_777);
  xnor csa_tree_add_117_21_pad_groupi_g3528(csa_tree_add_117_21_pad_groupi_n_878 ,csa_tree_add_117_21_pad_groupi_n_619 ,csa_tree_add_117_21_pad_groupi_n_780);
  xnor csa_tree_add_117_21_pad_groupi_g3529(csa_tree_add_117_21_pad_groupi_n_877 ,csa_tree_add_117_21_pad_groupi_n_626 ,csa_tree_add_117_21_pad_groupi_n_778);
  xnor csa_tree_add_117_21_pad_groupi_g3530(csa_tree_add_117_21_pad_groupi_n_876 ,csa_tree_add_117_21_pad_groupi_n_623 ,csa_tree_add_117_21_pad_groupi_n_776);
  xnor csa_tree_add_117_21_pad_groupi_g3531(csa_tree_add_117_21_pad_groupi_n_875 ,csa_tree_add_117_21_pad_groupi_n_639 ,csa_tree_add_117_21_pad_groupi_n_775);
  xnor csa_tree_add_117_21_pad_groupi_g3532(csa_tree_add_117_21_pad_groupi_n_874 ,csa_tree_add_117_21_pad_groupi_n_649 ,csa_tree_add_117_21_pad_groupi_n_785);
  xnor csa_tree_add_117_21_pad_groupi_g3533(csa_tree_add_117_21_pad_groupi_n_873 ,csa_tree_add_117_21_pad_groupi_n_642 ,csa_tree_add_117_21_pad_groupi_n_786);
  xnor csa_tree_add_117_21_pad_groupi_g3534(csa_tree_add_117_21_pad_groupi_n_872 ,csa_tree_add_117_21_pad_groupi_n_631 ,csa_tree_add_117_21_pad_groupi_n_798);
  not csa_tree_add_117_21_pad_groupi_g3535(csa_tree_add_117_21_pad_groupi_n_865 ,csa_tree_add_117_21_pad_groupi_n_866);
  nor csa_tree_add_117_21_pad_groupi_g3536(csa_tree_add_117_21_pad_groupi_n_858 ,csa_tree_add_117_21_pad_groupi_n_835 ,csa_tree_add_117_21_pad_groupi_n_734);
  nor csa_tree_add_117_21_pad_groupi_g3537(csa_tree_add_117_21_pad_groupi_n_857 ,csa_tree_add_117_21_pad_groupi_n_772 ,csa_tree_add_117_21_pad_groupi_n_817);
  and csa_tree_add_117_21_pad_groupi_g3538(csa_tree_add_117_21_pad_groupi_n_870 ,csa_tree_add_117_21_pad_groupi_n_754 ,csa_tree_add_117_21_pad_groupi_n_815);
  and csa_tree_add_117_21_pad_groupi_g3539(csa_tree_add_117_21_pad_groupi_n_869 ,csa_tree_add_117_21_pad_groupi_n_758 ,csa_tree_add_117_21_pad_groupi_n_814);
  and csa_tree_add_117_21_pad_groupi_g3540(csa_tree_add_117_21_pad_groupi_n_868 ,csa_tree_add_117_21_pad_groupi_n_716 ,csa_tree_add_117_21_pad_groupi_n_811);
  and csa_tree_add_117_21_pad_groupi_g3541(csa_tree_add_117_21_pad_groupi_n_867 ,csa_tree_add_117_21_pad_groupi_n_760 ,csa_tree_add_117_21_pad_groupi_n_820);
  and csa_tree_add_117_21_pad_groupi_g3542(csa_tree_add_117_21_pad_groupi_n_866 ,csa_tree_add_117_21_pad_groupi_n_765 ,csa_tree_add_117_21_pad_groupi_n_822);
  and csa_tree_add_117_21_pad_groupi_g3543(csa_tree_add_117_21_pad_groupi_n_864 ,csa_tree_add_117_21_pad_groupi_n_749 ,csa_tree_add_117_21_pad_groupi_n_828);
  and csa_tree_add_117_21_pad_groupi_g3544(csa_tree_add_117_21_pad_groupi_n_863 ,csa_tree_add_117_21_pad_groupi_n_751 ,csa_tree_add_117_21_pad_groupi_n_810);
  and csa_tree_add_117_21_pad_groupi_g3545(csa_tree_add_117_21_pad_groupi_n_862 ,csa_tree_add_117_21_pad_groupi_n_755 ,csa_tree_add_117_21_pad_groupi_n_813);
  and csa_tree_add_117_21_pad_groupi_g3546(csa_tree_add_117_21_pad_groupi_n_861 ,csa_tree_add_117_21_pad_groupi_n_747 ,csa_tree_add_117_21_pad_groupi_n_809);
  and csa_tree_add_117_21_pad_groupi_g3547(csa_tree_add_117_21_pad_groupi_n_860 ,csa_tree_add_117_21_pad_groupi_n_741 ,csa_tree_add_117_21_pad_groupi_n_808);
  and csa_tree_add_117_21_pad_groupi_g3548(csa_tree_add_117_21_pad_groupi_n_859 ,csa_tree_add_117_21_pad_groupi_n_739 ,csa_tree_add_117_21_pad_groupi_n_812);
  not csa_tree_add_117_21_pad_groupi_g3549(csa_tree_add_117_21_pad_groupi_n_856 ,csa_tree_add_117_21_pad_groupi_n_855);
  not csa_tree_add_117_21_pad_groupi_g3550(csa_tree_add_117_21_pad_groupi_n_854 ,csa_tree_add_117_21_pad_groupi_n_853);
  not csa_tree_add_117_21_pad_groupi_g3551(csa_tree_add_117_21_pad_groupi_n_848 ,csa_tree_add_117_21_pad_groupi_n_849);
  nor csa_tree_add_117_21_pad_groupi_g3552(csa_tree_add_117_21_pad_groupi_n_846 ,csa_tree_add_117_21_pad_groupi_n_732 ,csa_tree_add_117_21_pad_groupi_n_827);
  and csa_tree_add_117_21_pad_groupi_g3553(csa_tree_add_117_21_pad_groupi_n_845 ,csa_tree_add_117_21_pad_groupi_n_832 ,csa_tree_add_117_21_pad_groupi_n_804);
  or csa_tree_add_117_21_pad_groupi_g3554(csa_tree_add_117_21_pad_groupi_n_844 ,csa_tree_add_117_21_pad_groupi_n_832 ,csa_tree_add_117_21_pad_groupi_n_804);
  or csa_tree_add_117_21_pad_groupi_g3555(csa_tree_add_117_21_pad_groupi_n_843 ,csa_tree_add_117_21_pad_groupi_n_1 ,csa_tree_add_117_21_pad_groupi_n_807);
  or csa_tree_add_117_21_pad_groupi_g3556(csa_tree_add_117_21_pad_groupi_n_842 ,csa_tree_add_117_21_pad_groupi_n_621 ,csa_tree_add_117_21_pad_groupi_n_829);
  and csa_tree_add_117_21_pad_groupi_g3557(csa_tree_add_117_21_pad_groupi_n_841 ,csa_tree_add_117_21_pad_groupi_n_621 ,csa_tree_add_117_21_pad_groupi_n_829);
  and csa_tree_add_117_21_pad_groupi_g3558(csa_tree_add_117_21_pad_groupi_n_855 ,csa_tree_add_117_21_pad_groupi_n_730 ,csa_tree_add_117_21_pad_groupi_n_819);
  or csa_tree_add_117_21_pad_groupi_g3559(csa_tree_add_117_21_pad_groupi_n_853 ,csa_tree_add_117_21_pad_groupi_n_725 ,csa_tree_add_117_21_pad_groupi_n_826);
  and csa_tree_add_117_21_pad_groupi_g3560(csa_tree_add_117_21_pad_groupi_n_852 ,csa_tree_add_117_21_pad_groupi_n_733 ,csa_tree_add_117_21_pad_groupi_n_818);
  and csa_tree_add_117_21_pad_groupi_g3561(csa_tree_add_117_21_pad_groupi_n_851 ,csa_tree_add_117_21_pad_groupi_n_723 ,csa_tree_add_117_21_pad_groupi_n_825);
  and csa_tree_add_117_21_pad_groupi_g3562(csa_tree_add_117_21_pad_groupi_n_850 ,csa_tree_add_117_21_pad_groupi_n_736 ,csa_tree_add_117_21_pad_groupi_n_816);
  and csa_tree_add_117_21_pad_groupi_g3563(csa_tree_add_117_21_pad_groupi_n_849 ,csa_tree_add_117_21_pad_groupi_n_727 ,csa_tree_add_117_21_pad_groupi_n_824);
  xnor csa_tree_add_117_21_pad_groupi_g3564(csa_tree_add_117_21_pad_groupi_n_847 ,csa_tree_add_117_21_pad_groupi_n_613 ,csa_tree_add_117_21_pad_groupi_n_715);
  not csa_tree_add_117_21_pad_groupi_g3565(csa_tree_add_117_21_pad_groupi_n_831 ,csa_tree_add_117_21_pad_groupi_n_830);
  or csa_tree_add_117_21_pad_groupi_g3566(csa_tree_add_117_21_pad_groupi_n_828 ,csa_tree_add_117_21_pad_groupi_n_652 ,csa_tree_add_117_21_pad_groupi_n_753);
  nor csa_tree_add_117_21_pad_groupi_g3567(csa_tree_add_117_21_pad_groupi_n_827 ,csa_tree_add_117_21_pad_groupi_n_717 ,csa_tree_add_117_21_pad_groupi_n_728);
  nor csa_tree_add_117_21_pad_groupi_g3568(csa_tree_add_117_21_pad_groupi_n_826 ,csa_tree_add_117_21_pad_groupi_n_712 ,csa_tree_add_117_21_pad_groupi_n_724);
  or csa_tree_add_117_21_pad_groupi_g3569(csa_tree_add_117_21_pad_groupi_n_825 ,csa_tree_add_117_21_pad_groupi_n_655 ,csa_tree_add_117_21_pad_groupi_n_719);
  or csa_tree_add_117_21_pad_groupi_g3570(csa_tree_add_117_21_pad_groupi_n_824 ,csa_tree_add_117_21_pad_groupi_n_653 ,csa_tree_add_117_21_pad_groupi_n_726);
  nor csa_tree_add_117_21_pad_groupi_g3571(csa_tree_add_117_21_pad_groupi_n_823 ,csa_tree_add_117_21_pad_groupi_n_664 ,csa_tree_add_117_21_pad_groupi_n_744);
  or csa_tree_add_117_21_pad_groupi_g3572(csa_tree_add_117_21_pad_groupi_n_822 ,csa_tree_add_117_21_pad_groupi_n_703 ,csa_tree_add_117_21_pad_groupi_n_763);
  nor csa_tree_add_117_21_pad_groupi_g3573(csa_tree_add_117_21_pad_groupi_n_821 ,csa_tree_add_117_21_pad_groupi_n_663 ,csa_tree_add_117_21_pad_groupi_n_745);
  or csa_tree_add_117_21_pad_groupi_g3574(csa_tree_add_117_21_pad_groupi_n_820 ,csa_tree_add_117_21_pad_groupi_n_711 ,csa_tree_add_117_21_pad_groupi_n_773);
  or csa_tree_add_117_21_pad_groupi_g3575(csa_tree_add_117_21_pad_groupi_n_819 ,csa_tree_add_117_21_pad_groupi_n_661 ,csa_tree_add_117_21_pad_groupi_n_729);
  or csa_tree_add_117_21_pad_groupi_g3576(csa_tree_add_117_21_pad_groupi_n_818 ,csa_tree_add_117_21_pad_groupi_n_704 ,csa_tree_add_117_21_pad_groupi_n_731);
  nor csa_tree_add_117_21_pad_groupi_g3577(csa_tree_add_117_21_pad_groupi_n_817 ,csa_tree_add_117_21_pad_groupi_n_709 ,csa_tree_add_117_21_pad_groupi_n_766);
  or csa_tree_add_117_21_pad_groupi_g3578(csa_tree_add_117_21_pad_groupi_n_816 ,csa_tree_add_117_21_pad_groupi_n_662 ,csa_tree_add_117_21_pad_groupi_n_735);
  or csa_tree_add_117_21_pad_groupi_g3579(csa_tree_add_117_21_pad_groupi_n_815 ,csa_tree_add_117_21_pad_groupi_n_743 ,csa_tree_add_117_21_pad_groupi_n_737);
  or csa_tree_add_117_21_pad_groupi_g3580(csa_tree_add_117_21_pad_groupi_n_814 ,csa_tree_add_117_21_pad_groupi_n_700 ,csa_tree_add_117_21_pad_groupi_n_757);
  or csa_tree_add_117_21_pad_groupi_g3581(csa_tree_add_117_21_pad_groupi_n_813 ,csa_tree_add_117_21_pad_groupi_n_657 ,csa_tree_add_117_21_pad_groupi_n_752);
  or csa_tree_add_117_21_pad_groupi_g3582(csa_tree_add_117_21_pad_groupi_n_812 ,csa_tree_add_117_21_pad_groupi_n_654 ,csa_tree_add_117_21_pad_groupi_n_738);
  or csa_tree_add_117_21_pad_groupi_g3583(csa_tree_add_117_21_pad_groupi_n_811 ,csa_tree_add_117_21_pad_groupi_n_659 ,csa_tree_add_117_21_pad_groupi_n_748);
  or csa_tree_add_117_21_pad_groupi_g3584(csa_tree_add_117_21_pad_groupi_n_810 ,csa_tree_add_117_21_pad_groupi_n_660 ,csa_tree_add_117_21_pad_groupi_n_750);
  or csa_tree_add_117_21_pad_groupi_g3585(csa_tree_add_117_21_pad_groupi_n_809 ,csa_tree_add_117_21_pad_groupi_n_658 ,csa_tree_add_117_21_pad_groupi_n_746);
  or csa_tree_add_117_21_pad_groupi_g3586(csa_tree_add_117_21_pad_groupi_n_808 ,csa_tree_add_117_21_pad_groupi_n_656 ,csa_tree_add_117_21_pad_groupi_n_740);
  and csa_tree_add_117_21_pad_groupi_g3587(csa_tree_add_117_21_pad_groupi_n_840 ,csa_tree_add_117_21_pad_groupi_n_684 ,csa_tree_add_117_21_pad_groupi_n_764);
  and csa_tree_add_117_21_pad_groupi_g3588(csa_tree_add_117_21_pad_groupi_n_839 ,csa_tree_add_117_21_pad_groupi_n_671 ,csa_tree_add_117_21_pad_groupi_n_759);
  and csa_tree_add_117_21_pad_groupi_g3589(csa_tree_add_117_21_pad_groupi_n_838 ,csa_tree_add_117_21_pad_groupi_n_682 ,csa_tree_add_117_21_pad_groupi_n_770);
  and csa_tree_add_117_21_pad_groupi_g3590(csa_tree_add_117_21_pad_groupi_n_837 ,csa_tree_add_117_21_pad_groupi_n_681 ,csa_tree_add_117_21_pad_groupi_n_769);
  and csa_tree_add_117_21_pad_groupi_g3591(csa_tree_add_117_21_pad_groupi_n_836 ,csa_tree_add_117_21_pad_groupi_n_673 ,csa_tree_add_117_21_pad_groupi_n_762);
  and csa_tree_add_117_21_pad_groupi_g3592(csa_tree_add_117_21_pad_groupi_n_835 ,csa_tree_add_117_21_pad_groupi_n_669 ,csa_tree_add_117_21_pad_groupi_n_771);
  and csa_tree_add_117_21_pad_groupi_g3593(csa_tree_add_117_21_pad_groupi_n_834 ,csa_tree_add_117_21_pad_groupi_n_677 ,csa_tree_add_117_21_pad_groupi_n_767);
  and csa_tree_add_117_21_pad_groupi_g3594(csa_tree_add_117_21_pad_groupi_n_833 ,csa_tree_add_117_21_pad_groupi_n_679 ,csa_tree_add_117_21_pad_groupi_n_768);
  and csa_tree_add_117_21_pad_groupi_g3595(csa_tree_add_117_21_pad_groupi_n_832 ,csa_tree_add_117_21_pad_groupi_n_246 ,csa_tree_add_117_21_pad_groupi_n_718);
  and csa_tree_add_117_21_pad_groupi_g3596(csa_tree_add_117_21_pad_groupi_n_830 ,csa_tree_add_117_21_pad_groupi_n_238 ,csa_tree_add_117_21_pad_groupi_n_774);
  and csa_tree_add_117_21_pad_groupi_g3597(csa_tree_add_117_21_pad_groupi_n_829 ,csa_tree_add_117_21_pad_groupi_n_233 ,csa_tree_add_117_21_pad_groupi_n_761);
  not csa_tree_add_117_21_pad_groupi_g3598(csa_tree_add_117_21_pad_groupi_n_806 ,csa_tree_add_117_21_pad_groupi_n_805);
  xnor csa_tree_add_117_21_pad_groupi_g3599(csa_tree_add_117_21_pad_groupi_n_803 ,csa_tree_add_117_21_pad_groupi_n_709 ,in4[14]);
  xnor csa_tree_add_117_21_pad_groupi_g3600(csa_tree_add_117_21_pad_groupi_n_802 ,csa_tree_add_117_21_pad_groupi_n_609 ,csa_tree_add_117_21_pad_groupi_n_704);
  xnor csa_tree_add_117_21_pad_groupi_g3601(csa_tree_add_117_21_pad_groupi_n_801 ,csa_tree_add_117_21_pad_groupi_n_607 ,csa_tree_add_117_21_pad_groupi_n_661);
  xnor csa_tree_add_117_21_pad_groupi_g3602(csa_tree_add_117_21_pad_groupi_n_800 ,csa_tree_add_117_21_pad_groupi_n_695 ,csa_tree_add_117_21_pad_groupi_n_651);
  xnor csa_tree_add_117_21_pad_groupi_g3603(csa_tree_add_117_21_pad_groupi_n_799 ,csa_tree_add_117_21_pad_groupi_n_637 ,csa_tree_add_117_21_pad_groupi_n_643);
  xnor csa_tree_add_117_21_pad_groupi_g3604(csa_tree_add_117_21_pad_groupi_n_798 ,csa_tree_add_117_21_pad_groupi_n_634 ,csa_tree_add_117_21_pad_groupi_n_656);
  xnor csa_tree_add_117_21_pad_groupi_g3605(csa_tree_add_117_21_pad_groupi_n_797 ,csa_tree_add_117_21_pad_groupi_n_699 ,in4[7]);
  xnor csa_tree_add_117_21_pad_groupi_g3606(csa_tree_add_117_21_pad_groupi_n_796 ,csa_tree_add_117_21_pad_groupi_n_708 ,in4[6]);
  xnor csa_tree_add_117_21_pad_groupi_g3607(csa_tree_add_117_21_pad_groupi_n_795 ,csa_tree_add_117_21_pad_groupi_n_707 ,in4[5]);
  xnor csa_tree_add_117_21_pad_groupi_g3608(csa_tree_add_117_21_pad_groupi_n_794 ,csa_tree_add_117_21_pad_groupi_n_667 ,csa_tree_add_117_21_pad_groupi_n_616);
  xnor csa_tree_add_117_21_pad_groupi_g3609(csa_tree_add_117_21_pad_groupi_n_793 ,csa_tree_add_117_21_pad_groupi_n_705 ,in4[4]);
  xnor csa_tree_add_117_21_pad_groupi_g3610(csa_tree_add_117_21_pad_groupi_n_792 ,csa_tree_add_117_21_pad_groupi_n_702 ,in4[8]);
  xnor csa_tree_add_117_21_pad_groupi_g3611(csa_tree_add_117_21_pad_groupi_n_791 ,csa_tree_add_117_21_pad_groupi_n_701 ,in4[3]);
  xnor csa_tree_add_117_21_pad_groupi_g3612(csa_tree_add_117_21_pad_groupi_n_790 ,csa_tree_add_117_21_pad_groupi_n_688 ,in4[2]);
  xnor csa_tree_add_117_21_pad_groupi_g3613(csa_tree_add_117_21_pad_groupi_n_789 ,csa_tree_add_117_21_pad_groupi_n_686 ,csa_tree_add_117_21_pad_groupi_n_636);
  xnor csa_tree_add_117_21_pad_groupi_g3614(csa_tree_add_117_21_pad_groupi_n_788 ,csa_tree_add_117_21_pad_groupi_n_713 ,in4[9]);
  xnor csa_tree_add_117_21_pad_groupi_g3615(csa_tree_add_117_21_pad_groupi_n_787 ,csa_tree_add_117_21_pad_groupi_n_593 ,csa_tree_add_117_21_pad_groupi_n_653);
  xnor csa_tree_add_117_21_pad_groupi_g3616(csa_tree_add_117_21_pad_groupi_n_786 ,csa_tree_add_117_21_pad_groupi_n_658 ,csa_tree_add_117_21_pad_groupi_n_644);
  xnor csa_tree_add_117_21_pad_groupi_g3617(csa_tree_add_117_21_pad_groupi_n_785 ,csa_tree_add_117_21_pad_groupi_n_660 ,csa_tree_add_117_21_pad_groupi_n_617);
  xnor csa_tree_add_117_21_pad_groupi_g3618(csa_tree_add_117_21_pad_groupi_n_784 ,csa_tree_add_117_21_pad_groupi_n_703 ,in4[12]);
  xnor csa_tree_add_117_21_pad_groupi_g3619(csa_tree_add_117_21_pad_groupi_n_783 ,csa_tree_add_117_21_pad_groupi_n_712 ,csa_tree_add_117_21_pad_groupi_n_589);
  xnor csa_tree_add_117_21_pad_groupi_g3620(csa_tree_add_117_21_pad_groupi_n_782 ,csa_tree_add_117_21_pad_groupi_n_691 ,csa_tree_add_117_21_pad_groupi_n_696);
  xnor csa_tree_add_117_21_pad_groupi_g3621(csa_tree_add_117_21_pad_groupi_n_781 ,csa_tree_add_117_21_pad_groupi_n_647 ,csa_tree_add_117_21_pad_groupi_n_645);
  xnor csa_tree_add_117_21_pad_groupi_g3622(csa_tree_add_117_21_pad_groupi_n_780 ,csa_tree_add_117_21_pad_groupi_n_662 ,csa_tree_add_117_21_pad_groupi_n_628);
  xnor csa_tree_add_117_21_pad_groupi_g3623(csa_tree_add_117_21_pad_groupi_n_779 ,csa_tree_add_117_21_pad_groupi_n_646 ,csa_tree_add_117_21_pad_groupi_n_648);
  xnor csa_tree_add_117_21_pad_groupi_g3624(csa_tree_add_117_21_pad_groupi_n_778 ,csa_tree_add_117_21_pad_groupi_n_654 ,csa_tree_add_117_21_pad_groupi_n_627);
  xnor csa_tree_add_117_21_pad_groupi_g3625(csa_tree_add_117_21_pad_groupi_n_777 ,csa_tree_add_117_21_pad_groupi_n_700 ,csa_tree_add_117_21_pad_groupi_n_693);
  xnor csa_tree_add_117_21_pad_groupi_g3626(csa_tree_add_117_21_pad_groupi_n_776 ,csa_tree_add_117_21_pad_groupi_n_652 ,csa_tree_add_117_21_pad_groupi_n_629);
  xnor csa_tree_add_117_21_pad_groupi_g3627(csa_tree_add_117_21_pad_groupi_n_775 ,csa_tree_add_117_21_pad_groupi_n_657 ,csa_tree_add_117_21_pad_groupi_n_638);
  xnor csa_tree_add_117_21_pad_groupi_g3628(csa_tree_add_117_21_pad_groupi_n_807 ,csa_tree_add_117_21_pad_groupi_n_697 ,csa_tree_add_117_21_pad_groupi_n_266);
  xnor csa_tree_add_117_21_pad_groupi_g3629(csa_tree_add_117_21_pad_groupi_n_805 ,csa_tree_add_117_21_pad_groupi_n_706 ,csa_tree_add_117_21_pad_groupi_n_268);
  xnor csa_tree_add_117_21_pad_groupi_g3630(csa_tree_add_117_21_pad_groupi_n_804 ,csa_tree_add_117_21_pad_groupi_n_698 ,csa_tree_add_117_21_pad_groupi_n_267);
  or csa_tree_add_117_21_pad_groupi_g3631(csa_tree_add_117_21_pad_groupi_n_774 ,csa_tree_add_117_21_pad_groupi_n_234 ,csa_tree_add_117_21_pad_groupi_n_697);
  nor csa_tree_add_117_21_pad_groupi_g3632(csa_tree_add_117_21_pad_groupi_n_773 ,in4[2] ,csa_tree_add_117_21_pad_groupi_n_687);
  nor csa_tree_add_117_21_pad_groupi_g3633(csa_tree_add_117_21_pad_groupi_n_772 ,in4[14] ,csa_tree_add_117_21_pad_groupi_n_622);
  or csa_tree_add_117_21_pad_groupi_g3634(csa_tree_add_117_21_pad_groupi_n_771 ,csa_tree_add_117_21_pad_groupi_n_675 ,csa_tree_add_117_21_pad_groupi_n_613);
  or csa_tree_add_117_21_pad_groupi_g3635(csa_tree_add_117_21_pad_groupi_n_770 ,csa_tree_add_117_21_pad_groupi_n_683 ,csa_tree_add_117_21_pad_groupi_n_713);
  or csa_tree_add_117_21_pad_groupi_g3636(csa_tree_add_117_21_pad_groupi_n_769 ,csa_tree_add_117_21_pad_groupi_n_680 ,csa_tree_add_117_21_pad_groupi_n_708);
  or csa_tree_add_117_21_pad_groupi_g3637(csa_tree_add_117_21_pad_groupi_n_768 ,csa_tree_add_117_21_pad_groupi_n_678 ,csa_tree_add_117_21_pad_groupi_n_707);
  or csa_tree_add_117_21_pad_groupi_g3638(csa_tree_add_117_21_pad_groupi_n_767 ,csa_tree_add_117_21_pad_groupi_n_676 ,csa_tree_add_117_21_pad_groupi_n_705);
  and csa_tree_add_117_21_pad_groupi_g3639(csa_tree_add_117_21_pad_groupi_n_766 ,in4[14] ,csa_tree_add_117_21_pad_groupi_n_622);
  or csa_tree_add_117_21_pad_groupi_g3640(csa_tree_add_117_21_pad_groupi_n_765 ,in4[12] ,csa_tree_add_117_21_pad_groupi_n_632);
  or csa_tree_add_117_21_pad_groupi_g3641(csa_tree_add_117_21_pad_groupi_n_764 ,csa_tree_add_117_21_pad_groupi_n_674 ,csa_tree_add_117_21_pad_groupi_n_701);
  and csa_tree_add_117_21_pad_groupi_g3642(csa_tree_add_117_21_pad_groupi_n_763 ,in4[12] ,csa_tree_add_117_21_pad_groupi_n_632);
  or csa_tree_add_117_21_pad_groupi_g3643(csa_tree_add_117_21_pad_groupi_n_762 ,csa_tree_add_117_21_pad_groupi_n_672 ,csa_tree_add_117_21_pad_groupi_n_699);
  or csa_tree_add_117_21_pad_groupi_g3644(csa_tree_add_117_21_pad_groupi_n_761 ,csa_tree_add_117_21_pad_groupi_n_236 ,csa_tree_add_117_21_pad_groupi_n_698);
  or csa_tree_add_117_21_pad_groupi_g3645(csa_tree_add_117_21_pad_groupi_n_760 ,csa_tree_add_117_21_pad_groupi_n_218 ,csa_tree_add_117_21_pad_groupi_n_688);
  or csa_tree_add_117_21_pad_groupi_g3646(csa_tree_add_117_21_pad_groupi_n_759 ,csa_tree_add_117_21_pad_groupi_n_670 ,csa_tree_add_117_21_pad_groupi_n_702);
  or csa_tree_add_117_21_pad_groupi_g3647(csa_tree_add_117_21_pad_groupi_n_758 ,csa_tree_add_117_21_pad_groupi_n_693 ,csa_tree_add_117_21_pad_groupi_n_692);
  and csa_tree_add_117_21_pad_groupi_g3648(csa_tree_add_117_21_pad_groupi_n_757 ,csa_tree_add_117_21_pad_groupi_n_693 ,csa_tree_add_117_21_pad_groupi_n_692);
  nor csa_tree_add_117_21_pad_groupi_g3649(csa_tree_add_117_21_pad_groupi_n_756 ,csa_tree_add_117_21_pad_groupi_n_696 ,csa_tree_add_117_21_pad_groupi_n_691);
  or csa_tree_add_117_21_pad_groupi_g3650(csa_tree_add_117_21_pad_groupi_n_755 ,csa_tree_add_117_21_pad_groupi_n_638 ,csa_tree_add_117_21_pad_groupi_n_639);
  or csa_tree_add_117_21_pad_groupi_g3651(csa_tree_add_117_21_pad_groupi_n_754 ,csa_tree_add_117_21_pad_groupi_n_648 ,csa_tree_add_117_21_pad_groupi_n_646);
  and csa_tree_add_117_21_pad_groupi_g3652(csa_tree_add_117_21_pad_groupi_n_753 ,csa_tree_add_117_21_pad_groupi_n_629 ,csa_tree_add_117_21_pad_groupi_n_623);
  and csa_tree_add_117_21_pad_groupi_g3653(csa_tree_add_117_21_pad_groupi_n_752 ,csa_tree_add_117_21_pad_groupi_n_638 ,csa_tree_add_117_21_pad_groupi_n_639);
  or csa_tree_add_117_21_pad_groupi_g3654(csa_tree_add_117_21_pad_groupi_n_751 ,csa_tree_add_117_21_pad_groupi_n_617 ,csa_tree_add_117_21_pad_groupi_n_649);
  and csa_tree_add_117_21_pad_groupi_g3655(csa_tree_add_117_21_pad_groupi_n_750 ,csa_tree_add_117_21_pad_groupi_n_617 ,csa_tree_add_117_21_pad_groupi_n_649);
  or csa_tree_add_117_21_pad_groupi_g3656(csa_tree_add_117_21_pad_groupi_n_749 ,csa_tree_add_117_21_pad_groupi_n_629 ,csa_tree_add_117_21_pad_groupi_n_623);
  and csa_tree_add_117_21_pad_groupi_g3657(csa_tree_add_117_21_pad_groupi_n_748 ,csa_tree_add_117_21_pad_groupi_n_645 ,csa_tree_add_117_21_pad_groupi_n_647);
  or csa_tree_add_117_21_pad_groupi_g3658(csa_tree_add_117_21_pad_groupi_n_747 ,csa_tree_add_117_21_pad_groupi_n_644 ,csa_tree_add_117_21_pad_groupi_n_642);
  and csa_tree_add_117_21_pad_groupi_g3659(csa_tree_add_117_21_pad_groupi_n_746 ,csa_tree_add_117_21_pad_groupi_n_644 ,csa_tree_add_117_21_pad_groupi_n_642);
  not csa_tree_add_117_21_pad_groupi_g3660(csa_tree_add_117_21_pad_groupi_n_745 ,csa_tree_add_117_21_pad_groupi_n_744);
  not csa_tree_add_117_21_pad_groupi_g3661(csa_tree_add_117_21_pad_groupi_n_743 ,csa_tree_add_117_21_pad_groupi_n_742);
  or csa_tree_add_117_21_pad_groupi_g3662(csa_tree_add_117_21_pad_groupi_n_741 ,csa_tree_add_117_21_pad_groupi_n_633 ,csa_tree_add_117_21_pad_groupi_n_631);
  nor csa_tree_add_117_21_pad_groupi_g3663(csa_tree_add_117_21_pad_groupi_n_740 ,csa_tree_add_117_21_pad_groupi_n_634 ,csa_tree_add_117_21_pad_groupi_n_630);
  or csa_tree_add_117_21_pad_groupi_g3664(csa_tree_add_117_21_pad_groupi_n_739 ,csa_tree_add_117_21_pad_groupi_n_627 ,csa_tree_add_117_21_pad_groupi_n_626);
  and csa_tree_add_117_21_pad_groupi_g3665(csa_tree_add_117_21_pad_groupi_n_738 ,csa_tree_add_117_21_pad_groupi_n_627 ,csa_tree_add_117_21_pad_groupi_n_626);
  and csa_tree_add_117_21_pad_groupi_g3666(csa_tree_add_117_21_pad_groupi_n_737 ,csa_tree_add_117_21_pad_groupi_n_648 ,csa_tree_add_117_21_pad_groupi_n_646);
  or csa_tree_add_117_21_pad_groupi_g3667(csa_tree_add_117_21_pad_groupi_n_736 ,csa_tree_add_117_21_pad_groupi_n_628 ,csa_tree_add_117_21_pad_groupi_n_619);
  and csa_tree_add_117_21_pad_groupi_g3668(csa_tree_add_117_21_pad_groupi_n_735 ,csa_tree_add_117_21_pad_groupi_n_628 ,csa_tree_add_117_21_pad_groupi_n_619);
  and csa_tree_add_117_21_pad_groupi_g3669(csa_tree_add_117_21_pad_groupi_n_734 ,csa_tree_add_117_21_pad_groupi_n_696 ,csa_tree_add_117_21_pad_groupi_n_691);
  or csa_tree_add_117_21_pad_groupi_g3670(csa_tree_add_117_21_pad_groupi_n_733 ,csa_tree_add_117_21_pad_groupi_n_608 ,csa_tree_add_117_21_pad_groupi_n_690);
  nor csa_tree_add_117_21_pad_groupi_g3671(csa_tree_add_117_21_pad_groupi_n_732 ,csa_tree_add_117_21_pad_groupi_n_615 ,csa_tree_add_117_21_pad_groupi_n_665);
  nor csa_tree_add_117_21_pad_groupi_g3672(csa_tree_add_117_21_pad_groupi_n_731 ,csa_tree_add_117_21_pad_groupi_n_609 ,csa_tree_add_117_21_pad_groupi_n_689);
  or csa_tree_add_117_21_pad_groupi_g3673(csa_tree_add_117_21_pad_groupi_n_730 ,csa_tree_add_117_21_pad_groupi_n_606 ,csa_tree_add_117_21_pad_groupi_n_641);
  nor csa_tree_add_117_21_pad_groupi_g3674(csa_tree_add_117_21_pad_groupi_n_729 ,csa_tree_add_117_21_pad_groupi_n_607 ,csa_tree_add_117_21_pad_groupi_n_640);
  nor csa_tree_add_117_21_pad_groupi_g3675(csa_tree_add_117_21_pad_groupi_n_728 ,csa_tree_add_117_21_pad_groupi_n_614 ,csa_tree_add_117_21_pad_groupi_n_666);
  or csa_tree_add_117_21_pad_groupi_g3676(csa_tree_add_117_21_pad_groupi_n_727 ,csa_tree_add_117_21_pad_groupi_n_592 ,csa_tree_add_117_21_pad_groupi_n_625);
  nor csa_tree_add_117_21_pad_groupi_g3677(csa_tree_add_117_21_pad_groupi_n_726 ,csa_tree_add_117_21_pad_groupi_n_593 ,csa_tree_add_117_21_pad_groupi_n_624);
  nor csa_tree_add_117_21_pad_groupi_g3678(csa_tree_add_117_21_pad_groupi_n_725 ,csa_tree_add_117_21_pad_groupi_n_589 ,csa_tree_add_117_21_pad_groupi_n_618);
  and csa_tree_add_117_21_pad_groupi_g3679(csa_tree_add_117_21_pad_groupi_n_724 ,csa_tree_add_117_21_pad_groupi_n_589 ,csa_tree_add_117_21_pad_groupi_n_618);
  or csa_tree_add_117_21_pad_groupi_g3680(csa_tree_add_117_21_pad_groupi_n_723 ,csa_tree_add_117_21_pad_groupi_n_694 ,csa_tree_add_117_21_pad_groupi_n_651);
  or csa_tree_add_117_21_pad_groupi_g3681(csa_tree_add_117_21_pad_groupi_n_722 ,csa_tree_add_117_21_pad_groupi_n_637 ,csa_tree_add_117_21_pad_groupi_n_211);
  nor csa_tree_add_117_21_pad_groupi_g3682(csa_tree_add_117_21_pad_groupi_n_721 ,csa_tree_add_117_21_pad_groupi_n_685 ,csa_tree_add_117_21_pad_groupi_n_636);
  or csa_tree_add_117_21_pad_groupi_g3683(csa_tree_add_117_21_pad_groupi_n_720 ,csa_tree_add_117_21_pad_groupi_n_686 ,csa_tree_add_117_21_pad_groupi_n_635);
  nor csa_tree_add_117_21_pad_groupi_g3684(csa_tree_add_117_21_pad_groupi_n_719 ,csa_tree_add_117_21_pad_groupi_n_695 ,csa_tree_add_117_21_pad_groupi_n_650);
  or csa_tree_add_117_21_pad_groupi_g3686(csa_tree_add_117_21_pad_groupi_n_718 ,csa_tree_add_117_21_pad_groupi_n_241 ,csa_tree_add_117_21_pad_groupi_n_706);
  or csa_tree_add_117_21_pad_groupi_g3687(csa_tree_add_117_21_pad_groupi_n_717 ,csa_tree_add_117_21_pad_groupi_n_4 ,csa_tree_add_117_21_pad_groupi_n_668);
  or csa_tree_add_117_21_pad_groupi_g3688(csa_tree_add_117_21_pad_groupi_n_716 ,csa_tree_add_117_21_pad_groupi_n_645 ,csa_tree_add_117_21_pad_groupi_n_647);
  xnor csa_tree_add_117_21_pad_groupi_g3689(csa_tree_add_117_21_pad_groupi_n_715 ,csa_tree_add_117_21_pad_groupi_n_602 ,in4[0]);
  xnor csa_tree_add_117_21_pad_groupi_g3690(csa_tree_add_117_21_pad_groupi_n_744 ,csa_tree_add_117_21_pad_groupi_n_599 ,csa_tree_add_117_21_pad_groupi_n_611);
  xnor csa_tree_add_117_21_pad_groupi_g3691(csa_tree_add_117_21_pad_groupi_n_742 ,csa_tree_add_117_21_pad_groupi_n_597 ,csa_tree_add_117_21_pad_groupi_n_610);
  not csa_tree_add_117_21_pad_groupi_g3693(csa_tree_add_117_21_pad_groupi_n_711 ,csa_tree_add_117_21_pad_groupi_n_710);
  not csa_tree_add_117_21_pad_groupi_g3694(csa_tree_add_117_21_pad_groupi_n_694 ,csa_tree_add_117_21_pad_groupi_n_695);
  not csa_tree_add_117_21_pad_groupi_g3695(csa_tree_add_117_21_pad_groupi_n_689 ,csa_tree_add_117_21_pad_groupi_n_690);
  not csa_tree_add_117_21_pad_groupi_g3696(csa_tree_add_117_21_pad_groupi_n_687 ,csa_tree_add_117_21_pad_groupi_n_688);
  not csa_tree_add_117_21_pad_groupi_g3697(csa_tree_add_117_21_pad_groupi_n_686 ,csa_tree_add_117_21_pad_groupi_n_685);
  or csa_tree_add_117_21_pad_groupi_g3698(csa_tree_add_117_21_pad_groupi_n_684 ,csa_tree_add_117_21_pad_groupi_n_215 ,csa_tree_add_117_21_pad_groupi_n_603);
  and csa_tree_add_117_21_pad_groupi_g3699(csa_tree_add_117_21_pad_groupi_n_683 ,in4[9] ,csa_tree_add_117_21_pad_groupi_n_605);
  or csa_tree_add_117_21_pad_groupi_g3700(csa_tree_add_117_21_pad_groupi_n_682 ,in4[9] ,csa_tree_add_117_21_pad_groupi_n_605);
  or csa_tree_add_117_21_pad_groupi_g3701(csa_tree_add_117_21_pad_groupi_n_681 ,csa_tree_add_117_21_pad_groupi_n_227 ,csa_tree_add_117_21_pad_groupi_n_595);
  nor csa_tree_add_117_21_pad_groupi_g3702(csa_tree_add_117_21_pad_groupi_n_680 ,in4[6] ,csa_tree_add_117_21_pad_groupi_n_596);
  or csa_tree_add_117_21_pad_groupi_g3703(csa_tree_add_117_21_pad_groupi_n_679 ,csa_tree_add_117_21_pad_groupi_n_226 ,csa_tree_add_117_21_pad_groupi_n_587);
  nor csa_tree_add_117_21_pad_groupi_g3704(csa_tree_add_117_21_pad_groupi_n_678 ,in4[5] ,csa_tree_add_117_21_pad_groupi_n_588);
  or csa_tree_add_117_21_pad_groupi_g3705(csa_tree_add_117_21_pad_groupi_n_677 ,csa_tree_add_117_21_pad_groupi_n_216 ,csa_tree_add_117_21_pad_groupi_n_585);
  nor csa_tree_add_117_21_pad_groupi_g3706(csa_tree_add_117_21_pad_groupi_n_676 ,in4[4] ,csa_tree_add_117_21_pad_groupi_n_586);
  nor csa_tree_add_117_21_pad_groupi_g3707(csa_tree_add_117_21_pad_groupi_n_675 ,in4[0] ,csa_tree_add_117_21_pad_groupi_n_602);
  nor csa_tree_add_117_21_pad_groupi_g3708(csa_tree_add_117_21_pad_groupi_n_674 ,in4[3] ,csa_tree_add_117_21_pad_groupi_n_604);
  or csa_tree_add_117_21_pad_groupi_g3709(csa_tree_add_117_21_pad_groupi_n_673 ,csa_tree_add_117_21_pad_groupi_n_217 ,csa_tree_add_117_21_pad_groupi_n_590);
  nor csa_tree_add_117_21_pad_groupi_g3710(csa_tree_add_117_21_pad_groupi_n_672 ,in4[7] ,csa_tree_add_117_21_pad_groupi_n_591);
  or csa_tree_add_117_21_pad_groupi_g3711(csa_tree_add_117_21_pad_groupi_n_671 ,csa_tree_add_117_21_pad_groupi_n_223 ,csa_tree_add_117_21_pad_groupi_n_594);
  nor csa_tree_add_117_21_pad_groupi_g3712(csa_tree_add_117_21_pad_groupi_n_670 ,in4[8] ,csa_tree_add_117_21_pad_groupi_n_0);
  or csa_tree_add_117_21_pad_groupi_g3713(csa_tree_add_117_21_pad_groupi_n_669 ,csa_tree_add_117_21_pad_groupi_n_224 ,csa_tree_add_117_21_pad_groupi_n_601);
  or csa_tree_add_117_21_pad_groupi_g3714(csa_tree_add_117_21_pad_groupi_n_668 ,csa_tree_add_117_21_pad_groupi_n_344 ,csa_tree_add_117_21_pad_groupi_n_584);
  and csa_tree_add_117_21_pad_groupi_g3716(csa_tree_add_117_21_pad_groupi_n_714 ,csa_tree_add_117_21_pad_groupi_n_599 ,csa_tree_add_117_21_pad_groupi_n_612);
  xnor csa_tree_add_117_21_pad_groupi_g3718(csa_tree_add_117_21_pad_groupi_n_712 ,csa_tree_add_117_21_pad_groupi_n_550 ,csa_tree_add_117_21_pad_groupi_n_354);
  xnor csa_tree_add_117_21_pad_groupi_g3725(csa_tree_add_117_21_pad_groupi_n_704 ,csa_tree_add_117_21_pad_groupi_n_544 ,csa_tree_add_117_21_pad_groupi_n_191);
  xnor csa_tree_add_117_21_pad_groupi_g3729(csa_tree_add_117_21_pad_groupi_n_700 ,csa_tree_add_117_21_pad_groupi_n_578 ,csa_tree_add_117_21_pad_groupi_n_167);
  xnor csa_tree_add_117_21_pad_groupi_g3733(csa_tree_add_117_21_pad_groupi_n_696 ,csa_tree_add_117_21_pad_groupi_n_527 ,csa_tree_add_117_21_pad_groupi_n_173);
  xnor csa_tree_add_117_21_pad_groupi_g3734(csa_tree_add_117_21_pad_groupi_n_695 ,csa_tree_add_117_21_pad_groupi_n_163 ,csa_tree_add_117_21_pad_groupi_n_560);
  xnor csa_tree_add_117_21_pad_groupi_g3735(csa_tree_add_117_21_pad_groupi_n_693 ,csa_tree_add_117_21_pad_groupi_n_580 ,csa_tree_add_117_21_pad_groupi_n_184);
  xnor csa_tree_add_117_21_pad_groupi_g3736(csa_tree_add_117_21_pad_groupi_n_692 ,csa_tree_add_117_21_pad_groupi_n_557 ,csa_tree_add_117_21_pad_groupi_n_176);
  xnor csa_tree_add_117_21_pad_groupi_g3737(csa_tree_add_117_21_pad_groupi_n_691 ,csa_tree_add_117_21_pad_groupi_n_582 ,csa_tree_add_117_21_pad_groupi_n_196);
  xnor csa_tree_add_117_21_pad_groupi_g3738(csa_tree_add_117_21_pad_groupi_n_690 ,csa_tree_add_117_21_pad_groupi_n_573 ,csa_tree_add_117_21_pad_groupi_n_170);
  or csa_tree_add_117_21_pad_groupi_g3740(csa_tree_add_117_21_pad_groupi_n_685 ,csa_tree_add_117_21_pad_groupi_n_598 ,csa_tree_add_117_21_pad_groupi_n_610);
  not csa_tree_add_117_21_pad_groupi_g3741(csa_tree_add_117_21_pad_groupi_n_666 ,csa_tree_add_117_21_pad_groupi_n_665);
  not csa_tree_add_117_21_pad_groupi_g3742(csa_tree_add_117_21_pad_groupi_n_664 ,csa_tree_add_117_21_pad_groupi_n_663);
  not csa_tree_add_117_21_pad_groupi_g3743(csa_tree_add_117_21_pad_groupi_n_650 ,csa_tree_add_117_21_pad_groupi_n_651);
  not csa_tree_add_117_21_pad_groupi_g3745(csa_tree_add_117_21_pad_groupi_n_640 ,csa_tree_add_117_21_pad_groupi_n_641);
  not csa_tree_add_117_21_pad_groupi_g3747(csa_tree_add_117_21_pad_groupi_n_635 ,csa_tree_add_117_21_pad_groupi_n_636);
  not csa_tree_add_117_21_pad_groupi_g3748(csa_tree_add_117_21_pad_groupi_n_634 ,csa_tree_add_117_21_pad_groupi_n_633);
  not csa_tree_add_117_21_pad_groupi_g3749(csa_tree_add_117_21_pad_groupi_n_630 ,csa_tree_add_117_21_pad_groupi_n_631);
  not csa_tree_add_117_21_pad_groupi_g3750(csa_tree_add_117_21_pad_groupi_n_624 ,csa_tree_add_117_21_pad_groupi_n_625);
  xnor csa_tree_add_117_21_pad_groupi_g3751(csa_tree_add_117_21_pad_groupi_n_665 ,csa_tree_add_117_21_pad_groupi_n_546 ,csa_tree_add_117_21_pad_groupi_n_184);
  xnor csa_tree_add_117_21_pad_groupi_g3752(csa_tree_add_117_21_pad_groupi_n_663 ,csa_tree_add_117_21_pad_groupi_n_559 ,csa_tree_add_117_21_pad_groupi_n_188);
  xnor csa_tree_add_117_21_pad_groupi_g3753(csa_tree_add_117_21_pad_groupi_n_616 ,csa_tree_add_117_21_pad_groupi_n_520 ,csa_tree_add_117_21_pad_groupi_n_196);
  xnor csa_tree_add_117_21_pad_groupi_g3754(csa_tree_add_117_21_pad_groupi_n_662 ,csa_tree_add_117_21_pad_groupi_n_532 ,csa_tree_add_117_21_pad_groupi_n_194);
  xnor csa_tree_add_117_21_pad_groupi_g3755(csa_tree_add_117_21_pad_groupi_n_661 ,csa_tree_add_117_21_pad_groupi_n_548 ,csa_tree_add_117_21_pad_groupi_n_181);
  xnor csa_tree_add_117_21_pad_groupi_g3756(csa_tree_add_117_21_pad_groupi_n_660 ,csa_tree_add_117_21_pad_groupi_n_553 ,csa_tree_add_117_21_pad_groupi_n_334);
  xnor csa_tree_add_117_21_pad_groupi_g3757(csa_tree_add_117_21_pad_groupi_n_659 ,csa_tree_add_117_21_pad_groupi_n_540 ,csa_tree_add_117_21_pad_groupi_n_190);
  xnor csa_tree_add_117_21_pad_groupi_g3758(csa_tree_add_117_21_pad_groupi_n_658 ,csa_tree_add_117_21_pad_groupi_n_539 ,csa_tree_add_117_21_pad_groupi_n_334);
  xnor csa_tree_add_117_21_pad_groupi_g3759(csa_tree_add_117_21_pad_groupi_n_657 ,csa_tree_add_117_21_pad_groupi_n_533 ,csa_tree_add_117_21_pad_groupi_n_193);
  xnor csa_tree_add_117_21_pad_groupi_g3760(csa_tree_add_117_21_pad_groupi_n_656 ,csa_tree_add_117_21_pad_groupi_n_528 ,csa_tree_add_117_21_pad_groupi_n_190);
  xnor csa_tree_add_117_21_pad_groupi_g3761(csa_tree_add_117_21_pad_groupi_n_655 ,csa_tree_add_117_21_pad_groupi_n_536 ,csa_tree_add_117_21_pad_groupi_n_197);
  xnor csa_tree_add_117_21_pad_groupi_g3762(csa_tree_add_117_21_pad_groupi_n_654 ,csa_tree_add_117_21_pad_groupi_n_518 ,csa_tree_add_117_21_pad_groupi_n_194);
  xnor csa_tree_add_117_21_pad_groupi_g3763(csa_tree_add_117_21_pad_groupi_n_653 ,csa_tree_add_117_21_pad_groupi_n_519 ,csa_tree_add_117_21_pad_groupi_n_193);
  xnor csa_tree_add_117_21_pad_groupi_g3764(csa_tree_add_117_21_pad_groupi_n_652 ,csa_tree_add_117_21_pad_groupi_n_571 ,csa_tree_add_117_21_pad_groupi_n_197);
  xnor csa_tree_add_117_21_pad_groupi_g3765(csa_tree_add_117_21_pad_groupi_n_651 ,csa_tree_add_117_21_pad_groupi_n_583 ,csa_tree_add_117_21_pad_groupi_n_181);
  xnor csa_tree_add_117_21_pad_groupi_g3766(csa_tree_add_117_21_pad_groupi_n_649 ,csa_tree_add_117_21_pad_groupi_n_566 ,csa_tree_add_117_21_pad_groupi_n_179);
  xnor csa_tree_add_117_21_pad_groupi_g3767(csa_tree_add_117_21_pad_groupi_n_648 ,csa_tree_add_117_21_pad_groupi_n_568 ,csa_tree_add_117_21_pad_groupi_n_331);
  xnor csa_tree_add_117_21_pad_groupi_g3768(csa_tree_add_117_21_pad_groupi_n_647 ,csa_tree_add_117_21_pad_groupi_n_552 ,csa_tree_add_117_21_pad_groupi_n_328);
  xnor csa_tree_add_117_21_pad_groupi_g3769(csa_tree_add_117_21_pad_groupi_n_646 ,csa_tree_add_117_21_pad_groupi_n_581 ,csa_tree_add_117_21_pad_groupi_n_175);
  xnor csa_tree_add_117_21_pad_groupi_g3770(csa_tree_add_117_21_pad_groupi_n_645 ,csa_tree_add_117_21_pad_groupi_n_172 ,csa_tree_add_117_21_pad_groupi_n_572);
  xnor csa_tree_add_117_21_pad_groupi_g3771(csa_tree_add_117_21_pad_groupi_n_644 ,csa_tree_add_117_21_pad_groupi_n_541 ,csa_tree_add_117_21_pad_groupi_n_331);
  xnor csa_tree_add_117_21_pad_groupi_g3772(csa_tree_add_117_21_pad_groupi_n_643 ,csa_tree_add_117_21_pad_groupi_n_576 ,csa_tree_add_117_21_pad_groupi_n_328);
  xnor csa_tree_add_117_21_pad_groupi_g3773(csa_tree_add_117_21_pad_groupi_n_642 ,csa_tree_add_117_21_pad_groupi_n_562 ,csa_tree_add_117_21_pad_groupi_n_178);
  xnor csa_tree_add_117_21_pad_groupi_g3774(csa_tree_add_117_21_pad_groupi_n_641 ,csa_tree_add_117_21_pad_groupi_n_534 ,csa_tree_add_117_21_pad_groupi_n_187);
  xnor csa_tree_add_117_21_pad_groupi_g3775(csa_tree_add_117_21_pad_groupi_n_639 ,csa_tree_add_117_21_pad_groupi_n_538 ,csa_tree_add_117_21_pad_groupi_n_175);
  xnor csa_tree_add_117_21_pad_groupi_g3776(csa_tree_add_117_21_pad_groupi_n_638 ,csa_tree_add_117_21_pad_groupi_n_521 ,csa_tree_add_117_21_pad_groupi_n_172);
  xnor csa_tree_add_117_21_pad_groupi_g3777(csa_tree_add_117_21_pad_groupi_n_637 ,csa_tree_add_117_21_pad_groupi_n_574 ,csa_tree_add_117_21_pad_groupi_n_166);
  xnor csa_tree_add_117_21_pad_groupi_g3778(csa_tree_add_117_21_pad_groupi_n_636 ,csa_tree_add_117_21_pad_groupi_n_570 ,csa_tree_add_117_21_pad_groupi_n_185);
  xnor csa_tree_add_117_21_pad_groupi_g3779(csa_tree_add_117_21_pad_groupi_n_633 ,csa_tree_add_117_21_pad_groupi_n_531 ,csa_tree_add_117_21_pad_groupi_n_188);
  xnor csa_tree_add_117_21_pad_groupi_g3780(csa_tree_add_117_21_pad_groupi_n_632 ,csa_tree_add_117_21_pad_groupi_n_529 ,csa_tree_add_117_21_pad_groupi_n_182);
  xnor csa_tree_add_117_21_pad_groupi_g3781(csa_tree_add_117_21_pad_groupi_n_631 ,csa_tree_add_117_21_pad_groupi_n_530 ,csa_tree_add_117_21_pad_groupi_n_179);
  xnor csa_tree_add_117_21_pad_groupi_g3782(csa_tree_add_117_21_pad_groupi_n_629 ,csa_tree_add_117_21_pad_groupi_n_535 ,csa_tree_add_117_21_pad_groupi_n_187);
  xnor csa_tree_add_117_21_pad_groupi_g3783(csa_tree_add_117_21_pad_groupi_n_628 ,csa_tree_add_117_21_pad_groupi_n_516 ,csa_tree_add_117_21_pad_groupi_n_185);
  xnor csa_tree_add_117_21_pad_groupi_g3784(csa_tree_add_117_21_pad_groupi_n_627 ,csa_tree_add_117_21_pad_groupi_n_523 ,csa_tree_add_117_21_pad_groupi_n_163);
  xnor csa_tree_add_117_21_pad_groupi_g3785(csa_tree_add_117_21_pad_groupi_n_626 ,csa_tree_add_117_21_pad_groupi_n_577 ,csa_tree_add_117_21_pad_groupi_n_178);
  xnor csa_tree_add_117_21_pad_groupi_g3786(csa_tree_add_117_21_pad_groupi_n_625 ,csa_tree_add_117_21_pad_groupi_n_524 ,csa_tree_add_117_21_pad_groupi_n_182);
  xnor csa_tree_add_117_21_pad_groupi_g3787(csa_tree_add_117_21_pad_groupi_n_623 ,csa_tree_add_117_21_pad_groupi_n_555 ,csa_tree_add_117_21_pad_groupi_n_169);
  xnor csa_tree_add_117_21_pad_groupi_g3788(csa_tree_add_117_21_pad_groupi_n_622 ,csa_tree_add_117_21_pad_groupi_n_543 ,csa_tree_add_117_21_pad_groupi_n_191);
  xnor csa_tree_add_117_21_pad_groupi_g3789(csa_tree_add_117_21_pad_groupi_n_621 ,csa_tree_add_117_21_pad_groupi_n_517 ,csa_tree_add_117_21_pad_groupi_n_167);
  xnor csa_tree_add_117_21_pad_groupi_g3790(csa_tree_add_117_21_pad_groupi_n_620 ,csa_tree_add_117_21_pad_groupi_n_575 ,csa_tree_add_117_21_pad_groupi_n_173);
  xnor csa_tree_add_117_21_pad_groupi_g3791(csa_tree_add_117_21_pad_groupi_n_619 ,csa_tree_add_117_21_pad_groupi_n_551 ,csa_tree_add_117_21_pad_groupi_n_176);
  xnor csa_tree_add_117_21_pad_groupi_g3792(csa_tree_add_117_21_pad_groupi_n_618 ,csa_tree_add_117_21_pad_groupi_n_569 ,csa_tree_add_117_21_pad_groupi_n_170);
  xnor csa_tree_add_117_21_pad_groupi_g3793(csa_tree_add_117_21_pad_groupi_n_617 ,csa_tree_add_117_21_pad_groupi_n_563 ,csa_tree_add_117_21_pad_groupi_n_164);
  not csa_tree_add_117_21_pad_groupi_g3794(csa_tree_add_117_21_pad_groupi_n_615 ,csa_tree_add_117_21_pad_groupi_n_614);
  not csa_tree_add_117_21_pad_groupi_g3795(csa_tree_add_117_21_pad_groupi_n_612 ,csa_tree_add_117_21_pad_groupi_n_611);
  not csa_tree_add_117_21_pad_groupi_g3796(csa_tree_add_117_21_pad_groupi_n_608 ,csa_tree_add_117_21_pad_groupi_n_609);
  not csa_tree_add_117_21_pad_groupi_g3797(csa_tree_add_117_21_pad_groupi_n_606 ,csa_tree_add_117_21_pad_groupi_n_607);
  not csa_tree_add_117_21_pad_groupi_g3798(csa_tree_add_117_21_pad_groupi_n_603 ,csa_tree_add_117_21_pad_groupi_n_604);
  not csa_tree_add_117_21_pad_groupi_g3799(csa_tree_add_117_21_pad_groupi_n_601 ,csa_tree_add_117_21_pad_groupi_n_602);
  nor csa_tree_add_117_21_pad_groupi_g3800(csa_tree_add_117_21_pad_groupi_n_600 ,csa_tree_add_117_21_pad_groupi_n_352 ,csa_tree_add_117_21_pad_groupi_n_550);
  xnor csa_tree_add_117_21_pad_groupi_g3801(csa_tree_add_117_21_pad_groupi_n_614 ,csa_tree_add_117_21_pad_groupi_n_446 ,csa_tree_add_117_21_pad_groupi_n_53);
  or csa_tree_add_117_21_pad_groupi_g3802(csa_tree_add_117_21_pad_groupi_n_613 ,csa_tree_add_117_21_pad_groupi_n_74 ,csa_tree_add_117_21_pad_groupi_n_545);
  or csa_tree_add_117_21_pad_groupi_g3803(csa_tree_add_117_21_pad_groupi_n_611 ,csa_tree_add_117_21_pad_groupi_n_75 ,csa_tree_add_117_21_pad_groupi_n_547);
  or csa_tree_add_117_21_pad_groupi_g3804(csa_tree_add_117_21_pad_groupi_n_610 ,csa_tree_add_117_21_pad_groupi_n_76 ,csa_tree_add_117_21_pad_groupi_n_549);
  xnor csa_tree_add_117_21_pad_groupi_g3805(csa_tree_add_117_21_pad_groupi_n_609 ,csa_tree_add_117_21_pad_groupi_n_451 ,csa_tree_add_117_21_pad_groupi_n_44);
  xnor csa_tree_add_117_21_pad_groupi_g3806(csa_tree_add_117_21_pad_groupi_n_607 ,csa_tree_add_117_21_pad_groupi_n_442 ,csa_tree_add_117_21_pad_groupi_n_44);
  xnor csa_tree_add_117_21_pad_groupi_g3807(csa_tree_add_117_21_pad_groupi_n_605 ,csa_tree_add_117_21_pad_groupi_n_448 ,csa_tree_add_117_21_pad_groupi_n_47);
  xnor csa_tree_add_117_21_pad_groupi_g3808(csa_tree_add_117_21_pad_groupi_n_604 ,csa_tree_add_117_21_pad_groupi_n_439 ,csa_tree_add_117_21_pad_groupi_n_52);
  xnor csa_tree_add_117_21_pad_groupi_g3809(csa_tree_add_117_21_pad_groupi_n_602 ,csa_tree_add_117_21_pad_groupi_n_449 ,csa_tree_add_117_21_pad_groupi_n_50);
  not csa_tree_add_117_21_pad_groupi_g3810(csa_tree_add_117_21_pad_groupi_n_598 ,csa_tree_add_117_21_pad_groupi_n_597);
  not csa_tree_add_117_21_pad_groupi_g3811(csa_tree_add_117_21_pad_groupi_n_595 ,csa_tree_add_117_21_pad_groupi_n_596);
  not csa_tree_add_117_21_pad_groupi_g3812(csa_tree_add_117_21_pad_groupi_n_594 ,csa_tree_add_117_21_pad_groupi_n_0);
  not csa_tree_add_117_21_pad_groupi_g3813(csa_tree_add_117_21_pad_groupi_n_592 ,csa_tree_add_117_21_pad_groupi_n_593);
  not csa_tree_add_117_21_pad_groupi_g3814(csa_tree_add_117_21_pad_groupi_n_590 ,csa_tree_add_117_21_pad_groupi_n_591);
  not csa_tree_add_117_21_pad_groupi_g3815(csa_tree_add_117_21_pad_groupi_n_587 ,csa_tree_add_117_21_pad_groupi_n_588);
  not csa_tree_add_117_21_pad_groupi_g3816(csa_tree_add_117_21_pad_groupi_n_585 ,csa_tree_add_117_21_pad_groupi_n_586);
  xor csa_tree_add_117_21_pad_groupi_g3817(csa_tree_add_117_21_pad_groupi_n_584 ,csa_tree_add_117_21_pad_groupi_n_445 ,csa_tree_add_117_21_pad_groupi_n_6);
  xnor csa_tree_add_117_21_pad_groupi_g3818(csa_tree_add_117_21_pad_groupi_n_599 ,csa_tree_add_117_21_pad_groupi_n_447 ,csa_tree_add_117_21_pad_groupi_n_47);
  xnor csa_tree_add_117_21_pad_groupi_g3819(csa_tree_add_117_21_pad_groupi_n_597 ,csa_tree_add_117_21_pad_groupi_n_450 ,csa_tree_add_117_21_pad_groupi_n_50);
  xnor csa_tree_add_117_21_pad_groupi_g3820(csa_tree_add_117_21_pad_groupi_n_596 ,csa_tree_add_117_21_pad_groupi_n_443 ,csa_tree_add_117_21_pad_groupi_n_48);
  xnor csa_tree_add_117_21_pad_groupi_g3822(csa_tree_add_117_21_pad_groupi_n_593 ,csa_tree_add_117_21_pad_groupi_n_444 ,csa_tree_add_117_21_pad_groupi_n_48);
  xnor csa_tree_add_117_21_pad_groupi_g3823(csa_tree_add_117_21_pad_groupi_n_591 ,csa_tree_add_117_21_pad_groupi_n_438 ,csa_tree_add_117_21_pad_groupi_n_45);
  xor csa_tree_add_117_21_pad_groupi_g3824(csa_tree_add_117_21_pad_groupi_n_589 ,csa_tree_add_117_21_pad_groupi_n_441 ,csa_tree_add_117_21_pad_groupi_n_4);
  xnor csa_tree_add_117_21_pad_groupi_g3825(csa_tree_add_117_21_pad_groupi_n_588 ,csa_tree_add_117_21_pad_groupi_n_437 ,csa_tree_add_117_21_pad_groupi_n_6);
  xnor csa_tree_add_117_21_pad_groupi_g3826(csa_tree_add_117_21_pad_groupi_n_586 ,csa_tree_add_117_21_pad_groupi_n_452 ,csa_tree_add_117_21_pad_groupi_n_52);
  or csa_tree_add_117_21_pad_groupi_g3827(csa_tree_add_117_21_pad_groupi_n_583 ,csa_tree_add_117_21_pad_groupi_n_408 ,csa_tree_add_117_21_pad_groupi_n_480);
  or csa_tree_add_117_21_pad_groupi_g3828(csa_tree_add_117_21_pad_groupi_n_582 ,csa_tree_add_117_21_pad_groupi_n_413 ,csa_tree_add_117_21_pad_groupi_n_482);
  or csa_tree_add_117_21_pad_groupi_g3829(csa_tree_add_117_21_pad_groupi_n_581 ,csa_tree_add_117_21_pad_groupi_n_410 ,csa_tree_add_117_21_pad_groupi_n_505);
  or csa_tree_add_117_21_pad_groupi_g3830(csa_tree_add_117_21_pad_groupi_n_580 ,csa_tree_add_117_21_pad_groupi_n_363 ,csa_tree_add_117_21_pad_groupi_n_510);
  or csa_tree_add_117_21_pad_groupi_g3832(csa_tree_add_117_21_pad_groupi_n_578 ,csa_tree_add_117_21_pad_groupi_n_430 ,csa_tree_add_117_21_pad_groupi_n_471);
  or csa_tree_add_117_21_pad_groupi_g3833(csa_tree_add_117_21_pad_groupi_n_577 ,csa_tree_add_117_21_pad_groupi_n_411 ,csa_tree_add_117_21_pad_groupi_n_508);
  or csa_tree_add_117_21_pad_groupi_g3834(csa_tree_add_117_21_pad_groupi_n_576 ,csa_tree_add_117_21_pad_groupi_n_435 ,csa_tree_add_117_21_pad_groupi_n_493);
  or csa_tree_add_117_21_pad_groupi_g3835(csa_tree_add_117_21_pad_groupi_n_575 ,csa_tree_add_117_21_pad_groupi_n_368 ,csa_tree_add_117_21_pad_groupi_n_503);
  or csa_tree_add_117_21_pad_groupi_g3836(csa_tree_add_117_21_pad_groupi_n_574 ,csa_tree_add_117_21_pad_groupi_n_414 ,csa_tree_add_117_21_pad_groupi_n_513);
  or csa_tree_add_117_21_pad_groupi_g3837(csa_tree_add_117_21_pad_groupi_n_573 ,csa_tree_add_117_21_pad_groupi_n_421 ,csa_tree_add_117_21_pad_groupi_n_489);
  or csa_tree_add_117_21_pad_groupi_g3838(csa_tree_add_117_21_pad_groupi_n_572 ,csa_tree_add_117_21_pad_groupi_n_394 ,csa_tree_add_117_21_pad_groupi_n_511);
  or csa_tree_add_117_21_pad_groupi_g3839(csa_tree_add_117_21_pad_groupi_n_571 ,csa_tree_add_117_21_pad_groupi_n_424 ,csa_tree_add_117_21_pad_groupi_n_498);
  or csa_tree_add_117_21_pad_groupi_g3840(csa_tree_add_117_21_pad_groupi_n_570 ,csa_tree_add_117_21_pad_groupi_n_365 ,csa_tree_add_117_21_pad_groupi_n_476);
  or csa_tree_add_117_21_pad_groupi_g3841(csa_tree_add_117_21_pad_groupi_n_569 ,csa_tree_add_117_21_pad_groupi_n_416 ,csa_tree_add_117_21_pad_groupi_n_507);
  or csa_tree_add_117_21_pad_groupi_g3842(csa_tree_add_117_21_pad_groupi_n_568 ,csa_tree_add_117_21_pad_groupi_n_370 ,csa_tree_add_117_21_pad_groupi_n_512);
  or csa_tree_add_117_21_pad_groupi_g3844(csa_tree_add_117_21_pad_groupi_n_566 ,csa_tree_add_117_21_pad_groupi_n_406 ,csa_tree_add_117_21_pad_groupi_n_472);
  or csa_tree_add_117_21_pad_groupi_g3847(csa_tree_add_117_21_pad_groupi_n_563 ,csa_tree_add_117_21_pad_groupi_n_360 ,csa_tree_add_117_21_pad_groupi_n_492);
  or csa_tree_add_117_21_pad_groupi_g3848(csa_tree_add_117_21_pad_groupi_n_562 ,csa_tree_add_117_21_pad_groupi_n_427 ,csa_tree_add_117_21_pad_groupi_n_486);
  or csa_tree_add_117_21_pad_groupi_g3850(csa_tree_add_117_21_pad_groupi_n_560 ,csa_tree_add_117_21_pad_groupi_n_394 ,csa_tree_add_117_21_pad_groupi_n_490);
  or csa_tree_add_117_21_pad_groupi_g3851(csa_tree_add_117_21_pad_groupi_n_559 ,csa_tree_add_117_21_pad_groupi_n_372 ,csa_tree_add_117_21_pad_groupi_n_499);
  or csa_tree_add_117_21_pad_groupi_g3853(csa_tree_add_117_21_pad_groupi_n_557 ,csa_tree_add_117_21_pad_groupi_n_429 ,csa_tree_add_117_21_pad_groupi_n_509);
  or csa_tree_add_117_21_pad_groupi_g3855(csa_tree_add_117_21_pad_groupi_n_555 ,csa_tree_add_117_21_pad_groupi_n_428 ,csa_tree_add_117_21_pad_groupi_n_473);
  or csa_tree_add_117_21_pad_groupi_g3857(csa_tree_add_117_21_pad_groupi_n_553 ,csa_tree_add_117_21_pad_groupi_n_425 ,csa_tree_add_117_21_pad_groupi_n_500);
  or csa_tree_add_117_21_pad_groupi_g3858(csa_tree_add_117_21_pad_groupi_n_552 ,csa_tree_add_117_21_pad_groupi_n_412 ,csa_tree_add_117_21_pad_groupi_n_514);
  or csa_tree_add_117_21_pad_groupi_g3859(csa_tree_add_117_21_pad_groupi_n_551 ,csa_tree_add_117_21_pad_groupi_n_426 ,csa_tree_add_117_21_pad_groupi_n_468);
  not csa_tree_add_117_21_pad_groupi_g3860(csa_tree_add_117_21_pad_groupi_n_549 ,csa_tree_add_117_21_pad_groupi_n_548);
  not csa_tree_add_117_21_pad_groupi_g3861(csa_tree_add_117_21_pad_groupi_n_547 ,csa_tree_add_117_21_pad_groupi_n_546);
  not csa_tree_add_117_21_pad_groupi_g3862(csa_tree_add_117_21_pad_groupi_n_545 ,csa_tree_add_117_21_pad_groupi_n_544);
  or csa_tree_add_117_21_pad_groupi_g3863(csa_tree_add_117_21_pad_groupi_n_543 ,csa_tree_add_117_21_pad_groupi_n_436 ,csa_tree_add_117_21_pad_groupi_n_477);
  or csa_tree_add_117_21_pad_groupi_g3865(csa_tree_add_117_21_pad_groupi_n_541 ,csa_tree_add_117_21_pad_groupi_n_373 ,csa_tree_add_117_21_pad_groupi_n_487);
  or csa_tree_add_117_21_pad_groupi_g3866(csa_tree_add_117_21_pad_groupi_n_540 ,csa_tree_add_117_21_pad_groupi_n_433 ,csa_tree_add_117_21_pad_groupi_n_504);
  or csa_tree_add_117_21_pad_groupi_g3867(csa_tree_add_117_21_pad_groupi_n_539 ,csa_tree_add_117_21_pad_groupi_n_418 ,csa_tree_add_117_21_pad_groupi_n_484);
  or csa_tree_add_117_21_pad_groupi_g3868(csa_tree_add_117_21_pad_groupi_n_538 ,csa_tree_add_117_21_pad_groupi_n_432 ,csa_tree_add_117_21_pad_groupi_n_495);
  or csa_tree_add_117_21_pad_groupi_g3870(csa_tree_add_117_21_pad_groupi_n_536 ,csa_tree_add_117_21_pad_groupi_n_422 ,csa_tree_add_117_21_pad_groupi_n_488);
  or csa_tree_add_117_21_pad_groupi_g3871(csa_tree_add_117_21_pad_groupi_n_535 ,csa_tree_add_117_21_pad_groupi_n_389 ,csa_tree_add_117_21_pad_groupi_n_497);
  or csa_tree_add_117_21_pad_groupi_g3872(csa_tree_add_117_21_pad_groupi_n_534 ,csa_tree_add_117_21_pad_groupi_n_374 ,csa_tree_add_117_21_pad_groupi_n_502);
  or csa_tree_add_117_21_pad_groupi_g3873(csa_tree_add_117_21_pad_groupi_n_533 ,csa_tree_add_117_21_pad_groupi_n_415 ,csa_tree_add_117_21_pad_groupi_n_481);
  or csa_tree_add_117_21_pad_groupi_g3874(csa_tree_add_117_21_pad_groupi_n_532 ,csa_tree_add_117_21_pad_groupi_n_405 ,csa_tree_add_117_21_pad_groupi_n_474);
  or csa_tree_add_117_21_pad_groupi_g3875(csa_tree_add_117_21_pad_groupi_n_531 ,csa_tree_add_117_21_pad_groupi_n_369 ,csa_tree_add_117_21_pad_groupi_n_483);
  or csa_tree_add_117_21_pad_groupi_g3876(csa_tree_add_117_21_pad_groupi_n_530 ,csa_tree_add_117_21_pad_groupi_n_420 ,csa_tree_add_117_21_pad_groupi_n_496);
  or csa_tree_add_117_21_pad_groupi_g3877(csa_tree_add_117_21_pad_groupi_n_529 ,csa_tree_add_117_21_pad_groupi_n_435 ,csa_tree_add_117_21_pad_groupi_n_470);
  or csa_tree_add_117_21_pad_groupi_g3878(csa_tree_add_117_21_pad_groupi_n_528 ,csa_tree_add_117_21_pad_groupi_n_419 ,csa_tree_add_117_21_pad_groupi_n_478);
  or csa_tree_add_117_21_pad_groupi_g3879(csa_tree_add_117_21_pad_groupi_n_527 ,csa_tree_add_117_21_pad_groupi_n_356 ,csa_tree_add_117_21_pad_groupi_n_456);
  or csa_tree_add_117_21_pad_groupi_g3882(csa_tree_add_117_21_pad_groupi_n_524 ,csa_tree_add_117_21_pad_groupi_n_407 ,csa_tree_add_117_21_pad_groupi_n_467);
  or csa_tree_add_117_21_pad_groupi_g3883(csa_tree_add_117_21_pad_groupi_n_523 ,csa_tree_add_117_21_pad_groupi_n_375 ,csa_tree_add_117_21_pad_groupi_n_506);
  or csa_tree_add_117_21_pad_groupi_g3885(csa_tree_add_117_21_pad_groupi_n_521 ,csa_tree_add_117_21_pad_groupi_n_358 ,csa_tree_add_117_21_pad_groupi_n_501);
  or csa_tree_add_117_21_pad_groupi_g3886(csa_tree_add_117_21_pad_groupi_n_520 ,csa_tree_add_117_21_pad_groupi_n_436 ,csa_tree_add_117_21_pad_groupi_n_485);
  or csa_tree_add_117_21_pad_groupi_g3887(csa_tree_add_117_21_pad_groupi_n_519 ,csa_tree_add_117_21_pad_groupi_n_417 ,csa_tree_add_117_21_pad_groupi_n_494);
  or csa_tree_add_117_21_pad_groupi_g3888(csa_tree_add_117_21_pad_groupi_n_518 ,csa_tree_add_117_21_pad_groupi_n_409 ,csa_tree_add_117_21_pad_groupi_n_491);
  or csa_tree_add_117_21_pad_groupi_g3889(csa_tree_add_117_21_pad_groupi_n_517 ,csa_tree_add_117_21_pad_groupi_n_431 ,csa_tree_add_117_21_pad_groupi_n_479);
  or csa_tree_add_117_21_pad_groupi_g3890(csa_tree_add_117_21_pad_groupi_n_516 ,csa_tree_add_117_21_pad_groupi_n_361 ,csa_tree_add_117_21_pad_groupi_n_469);
  xnor csa_tree_add_117_21_pad_groupi_g3893(csa_tree_add_117_21_pad_groupi_n_548 ,csa_tree_add_117_21_pad_groupi_n_169 ,csa_tree_add_117_21_pad_groupi_n_395);
  xnor csa_tree_add_117_21_pad_groupi_g3894(csa_tree_add_117_21_pad_groupi_n_546 ,csa_tree_add_117_21_pad_groupi_n_164 ,csa_tree_add_117_21_pad_groupi_n_353);
  xnor csa_tree_add_117_21_pad_groupi_g3895(csa_tree_add_117_21_pad_groupi_n_544 ,csa_tree_add_117_21_pad_groupi_n_166 ,csa_tree_add_117_21_pad_groupi_n_397);
  and csa_tree_add_117_21_pad_groupi_g3896(csa_tree_add_117_21_pad_groupi_n_514 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_30);
  and csa_tree_add_117_21_pad_groupi_g3897(csa_tree_add_117_21_pad_groupi_n_513 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_15);
  and csa_tree_add_117_21_pad_groupi_g3898(csa_tree_add_117_21_pad_groupi_n_512 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_36);
  and csa_tree_add_117_21_pad_groupi_g3899(csa_tree_add_117_21_pad_groupi_n_511 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_18);
  and csa_tree_add_117_21_pad_groupi_g3900(csa_tree_add_117_21_pad_groupi_n_510 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_35);
  and csa_tree_add_117_21_pad_groupi_g3901(csa_tree_add_117_21_pad_groupi_n_509 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_42);
  and csa_tree_add_117_21_pad_groupi_g3902(csa_tree_add_117_21_pad_groupi_n_508 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_29);
  and csa_tree_add_117_21_pad_groupi_g3903(csa_tree_add_117_21_pad_groupi_n_507 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_9);
  and csa_tree_add_117_21_pad_groupi_g3904(csa_tree_add_117_21_pad_groupi_n_506 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_21);
  and csa_tree_add_117_21_pad_groupi_g3905(csa_tree_add_117_21_pad_groupi_n_505 ,in3[0] ,csa_tree_add_117_21_pad_groupi_n_8);
  and csa_tree_add_117_21_pad_groupi_g3906(csa_tree_add_117_21_pad_groupi_n_504 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_24);
  and csa_tree_add_117_21_pad_groupi_g3907(csa_tree_add_117_21_pad_groupi_n_503 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_20);
  and csa_tree_add_117_21_pad_groupi_g3908(csa_tree_add_117_21_pad_groupi_n_502 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_36);
  and csa_tree_add_117_21_pad_groupi_g3909(csa_tree_add_117_21_pad_groupi_n_501 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_35);
  and csa_tree_add_117_21_pad_groupi_g3910(csa_tree_add_117_21_pad_groupi_n_500 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_14);
  and csa_tree_add_117_21_pad_groupi_g3911(csa_tree_add_117_21_pad_groupi_n_499 ,in3[0] ,csa_tree_add_117_21_pad_groupi_n_38);
  and csa_tree_add_117_21_pad_groupi_g3912(csa_tree_add_117_21_pad_groupi_n_498 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_27);
  and csa_tree_add_117_21_pad_groupi_g3913(csa_tree_add_117_21_pad_groupi_n_497 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_39);
  and csa_tree_add_117_21_pad_groupi_g3914(csa_tree_add_117_21_pad_groupi_n_496 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_30);
  and csa_tree_add_117_21_pad_groupi_g3915(csa_tree_add_117_21_pad_groupi_n_495 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_29);
  and csa_tree_add_117_21_pad_groupi_g3916(csa_tree_add_117_21_pad_groupi_n_494 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_26);
  and csa_tree_add_117_21_pad_groupi_g3917(csa_tree_add_117_21_pad_groupi_n_493 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_32);
  and csa_tree_add_117_21_pad_groupi_g3918(csa_tree_add_117_21_pad_groupi_n_492 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_39);
  and csa_tree_add_117_21_pad_groupi_g3919(csa_tree_add_117_21_pad_groupi_n_491 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_15);
  and csa_tree_add_117_21_pad_groupi_g3920(csa_tree_add_117_21_pad_groupi_n_490 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_21);
  and csa_tree_add_117_21_pad_groupi_g3921(csa_tree_add_117_21_pad_groupi_n_489 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_33);
  and csa_tree_add_117_21_pad_groupi_g3922(csa_tree_add_117_21_pad_groupi_n_488 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_14);
  and csa_tree_add_117_21_pad_groupi_g3923(csa_tree_add_117_21_pad_groupi_n_487 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_38);
  and csa_tree_add_117_21_pad_groupi_g3924(csa_tree_add_117_21_pad_groupi_n_486 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_33);
  and csa_tree_add_117_21_pad_groupi_g3925(csa_tree_add_117_21_pad_groupi_n_485 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_11);
  and csa_tree_add_117_21_pad_groupi_g3926(csa_tree_add_117_21_pad_groupi_n_484 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_12);
  and csa_tree_add_117_21_pad_groupi_g3927(csa_tree_add_117_21_pad_groupi_n_483 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_17);
  and csa_tree_add_117_21_pad_groupi_g3928(csa_tree_add_117_21_pad_groupi_n_482 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_12);
  and csa_tree_add_117_21_pad_groupi_g3929(csa_tree_add_117_21_pad_groupi_n_481 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_27);
  and csa_tree_add_117_21_pad_groupi_g3930(csa_tree_add_117_21_pad_groupi_n_480 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_9);
  and csa_tree_add_117_21_pad_groupi_g3931(csa_tree_add_117_21_pad_groupi_n_479 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_11);
  and csa_tree_add_117_21_pad_groupi_g3932(csa_tree_add_117_21_pad_groupi_n_478 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_23);
  and csa_tree_add_117_21_pad_groupi_g3933(csa_tree_add_117_21_pad_groupi_n_477 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_23);
  and csa_tree_add_117_21_pad_groupi_g3934(csa_tree_add_117_21_pad_groupi_n_476 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_17);
  and csa_tree_add_117_21_pad_groupi_g3936(csa_tree_add_117_21_pad_groupi_n_474 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_24);
  and csa_tree_add_117_21_pad_groupi_g3937(csa_tree_add_117_21_pad_groupi_n_473 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_32);
  and csa_tree_add_117_21_pad_groupi_g3938(csa_tree_add_117_21_pad_groupi_n_472 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_41);
  and csa_tree_add_117_21_pad_groupi_g3939(csa_tree_add_117_21_pad_groupi_n_471 ,in3[0] ,csa_tree_add_117_21_pad_groupi_n_26);
  and csa_tree_add_117_21_pad_groupi_g3940(csa_tree_add_117_21_pad_groupi_n_470 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_41);
  and csa_tree_add_117_21_pad_groupi_g3941(csa_tree_add_117_21_pad_groupi_n_469 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_18);
  and csa_tree_add_117_21_pad_groupi_g3942(csa_tree_add_117_21_pad_groupi_n_468 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_42);
  and csa_tree_add_117_21_pad_groupi_g3943(csa_tree_add_117_21_pad_groupi_n_467 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_8);
  and csa_tree_add_117_21_pad_groupi_g3954(csa_tree_add_117_21_pad_groupi_n_456 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_20);
  or csa_tree_add_117_21_pad_groupi_g3958(csa_tree_add_117_21_pad_groupi_n_452 ,csa_tree_add_117_21_pad_groupi_n_305 ,csa_tree_add_117_21_pad_groupi_n_379);
  or csa_tree_add_117_21_pad_groupi_g3959(csa_tree_add_117_21_pad_groupi_n_451 ,csa_tree_add_117_21_pad_groupi_n_301 ,csa_tree_add_117_21_pad_groupi_n_377);
  or csa_tree_add_117_21_pad_groupi_g3960(csa_tree_add_117_21_pad_groupi_n_450 ,csa_tree_add_117_21_pad_groupi_n_306 ,csa_tree_add_117_21_pad_groupi_n_367);
  or csa_tree_add_117_21_pad_groupi_g3961(csa_tree_add_117_21_pad_groupi_n_449 ,csa_tree_add_117_21_pad_groupi_n_288 ,csa_tree_add_117_21_pad_groupi_n_382);
  or csa_tree_add_117_21_pad_groupi_g3962(csa_tree_add_117_21_pad_groupi_n_448 ,csa_tree_add_117_21_pad_groupi_n_308 ,csa_tree_add_117_21_pad_groupi_n_364);
  or csa_tree_add_117_21_pad_groupi_g3963(csa_tree_add_117_21_pad_groupi_n_447 ,csa_tree_add_117_21_pad_groupi_n_287 ,csa_tree_add_117_21_pad_groupi_n_371);
  or csa_tree_add_117_21_pad_groupi_g3964(csa_tree_add_117_21_pad_groupi_n_446 ,csa_tree_add_117_21_pad_groupi_n_286 ,csa_tree_add_117_21_pad_groupi_n_359);
  or csa_tree_add_117_21_pad_groupi_g3965(csa_tree_add_117_21_pad_groupi_n_445 ,csa_tree_add_117_21_pad_groupi_n_302 ,csa_tree_add_117_21_pad_groupi_n_384);
  or csa_tree_add_117_21_pad_groupi_g3966(csa_tree_add_117_21_pad_groupi_n_444 ,csa_tree_add_117_21_pad_groupi_n_299 ,csa_tree_add_117_21_pad_groupi_n_380);
  or csa_tree_add_117_21_pad_groupi_g3967(csa_tree_add_117_21_pad_groupi_n_443 ,csa_tree_add_117_21_pad_groupi_n_285 ,csa_tree_add_117_21_pad_groupi_n_383);
  or csa_tree_add_117_21_pad_groupi_g3968(csa_tree_add_117_21_pad_groupi_n_442 ,csa_tree_add_117_21_pad_groupi_n_298 ,csa_tree_add_117_21_pad_groupi_n_376);
  or csa_tree_add_117_21_pad_groupi_g3969(csa_tree_add_117_21_pad_groupi_n_441 ,csa_tree_add_117_21_pad_groupi_n_303 ,csa_tree_add_117_21_pad_groupi_n_366);
  or csa_tree_add_117_21_pad_groupi_g3970(csa_tree_add_117_21_pad_groupi_n_440 ,csa_tree_add_117_21_pad_groupi_n_308 ,csa_tree_add_117_21_pad_groupi_n_381);
  or csa_tree_add_117_21_pad_groupi_g3971(csa_tree_add_117_21_pad_groupi_n_439 ,csa_tree_add_117_21_pad_groupi_n_307 ,csa_tree_add_117_21_pad_groupi_n_385);
  or csa_tree_add_117_21_pad_groupi_g3972(csa_tree_add_117_21_pad_groupi_n_438 ,csa_tree_add_117_21_pad_groupi_n_300 ,csa_tree_add_117_21_pad_groupi_n_357);
  or csa_tree_add_117_21_pad_groupi_g3973(csa_tree_add_117_21_pad_groupi_n_437 ,csa_tree_add_117_21_pad_groupi_n_304 ,csa_tree_add_117_21_pad_groupi_n_362);
  and csa_tree_add_117_21_pad_groupi_g3974(csa_tree_add_117_21_pad_groupi_n_434 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_96);
  and csa_tree_add_117_21_pad_groupi_g3975(csa_tree_add_117_21_pad_groupi_n_433 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_155);
  and csa_tree_add_117_21_pad_groupi_g3976(csa_tree_add_117_21_pad_groupi_n_432 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_161);
  and csa_tree_add_117_21_pad_groupi_g3977(csa_tree_add_117_21_pad_groupi_n_431 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_148);
  and csa_tree_add_117_21_pad_groupi_g3978(csa_tree_add_117_21_pad_groupi_n_430 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_139);
  and csa_tree_add_117_21_pad_groupi_g3979(csa_tree_add_117_21_pad_groupi_n_429 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_151);
  and csa_tree_add_117_21_pad_groupi_g3980(csa_tree_add_117_21_pad_groupi_n_428 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_145);
  and csa_tree_add_117_21_pad_groupi_g3981(csa_tree_add_117_21_pad_groupi_n_427 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_152);
  and csa_tree_add_117_21_pad_groupi_g3982(csa_tree_add_117_21_pad_groupi_n_426 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_145);
  and csa_tree_add_117_21_pad_groupi_g3983(csa_tree_add_117_21_pad_groupi_n_425 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_149);
  and csa_tree_add_117_21_pad_groupi_g3984(csa_tree_add_117_21_pad_groupi_n_424 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_139);
  and csa_tree_add_117_21_pad_groupi_g3985(csa_tree_add_117_21_pad_groupi_n_423 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_96);
  and csa_tree_add_117_21_pad_groupi_g3986(csa_tree_add_117_21_pad_groupi_n_422 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_140);
  and csa_tree_add_117_21_pad_groupi_g3987(csa_tree_add_117_21_pad_groupi_n_421 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_146);
  and csa_tree_add_117_21_pad_groupi_g3988(csa_tree_add_117_21_pad_groupi_n_420 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_146);
  and csa_tree_add_117_21_pad_groupi_g3989(csa_tree_add_117_21_pad_groupi_n_419 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_140);
  and csa_tree_add_117_21_pad_groupi_g3990(csa_tree_add_117_21_pad_groupi_n_418 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_149);
  and csa_tree_add_117_21_pad_groupi_g3991(csa_tree_add_117_21_pad_groupi_n_417 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_121);
  and csa_tree_add_117_21_pad_groupi_g3992(csa_tree_add_117_21_pad_groupi_n_416 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_152);
  and csa_tree_add_117_21_pad_groupi_g3993(csa_tree_add_117_21_pad_groupi_n_415 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_120);
  and csa_tree_add_117_21_pad_groupi_g3994(csa_tree_add_117_21_pad_groupi_n_414 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_148);
  and csa_tree_add_117_21_pad_groupi_g3995(csa_tree_add_117_21_pad_groupi_n_413 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_155);
  and csa_tree_add_117_21_pad_groupi_g3996(csa_tree_add_117_21_pad_groupi_n_412 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_124);
  and csa_tree_add_117_21_pad_groupi_g3997(csa_tree_add_117_21_pad_groupi_n_411 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_123);
  and csa_tree_add_117_21_pad_groupi_g3998(csa_tree_add_117_21_pad_groupi_n_410 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_151);
  and csa_tree_add_117_21_pad_groupi_g3999(csa_tree_add_117_21_pad_groupi_n_409 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_121);
  and csa_tree_add_117_21_pad_groupi_g4000(csa_tree_add_117_21_pad_groupi_n_408 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_161);
  and csa_tree_add_117_21_pad_groupi_g4001(csa_tree_add_117_21_pad_groupi_n_407 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_124);
  and csa_tree_add_117_21_pad_groupi_g4002(csa_tree_add_117_21_pad_groupi_n_406 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_160);
  and csa_tree_add_117_21_pad_groupi_g4003(csa_tree_add_117_21_pad_groupi_n_405 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_154);
  and csa_tree_add_117_21_pad_groupi_g4004(csa_tree_add_117_21_pad_groupi_n_404 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_67);
  and csa_tree_add_117_21_pad_groupi_g4005(csa_tree_add_117_21_pad_groupi_n_403 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_102);
  and csa_tree_add_117_21_pad_groupi_g4006(csa_tree_add_117_21_pad_groupi_n_402 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_68);
  and csa_tree_add_117_21_pad_groupi_g4007(csa_tree_add_117_21_pad_groupi_n_401 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_100);
  and csa_tree_add_117_21_pad_groupi_g4008(csa_tree_add_117_21_pad_groupi_n_400 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_100);
  and csa_tree_add_117_21_pad_groupi_g4009(csa_tree_add_117_21_pad_groupi_n_399 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_102);
  and csa_tree_add_117_21_pad_groupi_g4010(csa_tree_add_117_21_pad_groupi_n_398 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_99);
  and csa_tree_add_117_21_pad_groupi_g4011(csa_tree_add_117_21_pad_groupi_n_436 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_154);
  or csa_tree_add_117_21_pad_groupi_g4012(csa_tree_add_117_21_pad_groupi_n_397 ,csa_tree_add_117_21_pad_groupi_n_56 ,csa_tree_add_117_21_pad_groupi_n_77);
  or csa_tree_add_117_21_pad_groupi_g4013(csa_tree_add_117_21_pad_groupi_n_396 ,csa_tree_add_117_21_pad_groupi_n_73 ,csa_tree_add_117_21_pad_groupi_n_341);
  or csa_tree_add_117_21_pad_groupi_g4014(csa_tree_add_117_21_pad_groupi_n_395 ,csa_tree_add_117_21_pad_groupi_n_73 ,csa_tree_add_117_21_pad_groupi_n_81);
  and csa_tree_add_117_21_pad_groupi_g4015(csa_tree_add_117_21_pad_groupi_n_435 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_160);
  and csa_tree_add_117_21_pad_groupi_g4016(csa_tree_add_117_21_pad_groupi_n_389 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_137);
  and csa_tree_add_117_21_pad_groupi_g4017(csa_tree_add_117_21_pad_groupi_n_388 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_68);
  and csa_tree_add_117_21_pad_groupi_g4018(csa_tree_add_117_21_pad_groupi_n_387 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_97);
  and csa_tree_add_117_21_pad_groupi_g4019(csa_tree_add_117_21_pad_groupi_n_386 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_103);
  and csa_tree_add_117_21_pad_groupi_g4020(csa_tree_add_117_21_pad_groupi_n_385 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_90);
  nor csa_tree_add_117_21_pad_groupi_g4021(csa_tree_add_117_21_pad_groupi_n_384 ,csa_tree_add_117_21_pad_groupi_n_221 ,csa_tree_add_117_21_pad_groupi_n_348);
  and csa_tree_add_117_21_pad_groupi_g4022(csa_tree_add_117_21_pad_groupi_n_383 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_93);
  and csa_tree_add_117_21_pad_groupi_g4023(csa_tree_add_117_21_pad_groupi_n_382 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_90);
  and csa_tree_add_117_21_pad_groupi_g4024(csa_tree_add_117_21_pad_groupi_n_381 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_64);
  and csa_tree_add_117_21_pad_groupi_g4025(csa_tree_add_117_21_pad_groupi_n_380 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_94);
  and csa_tree_add_117_21_pad_groupi_g4026(csa_tree_add_117_21_pad_groupi_n_379 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_65);
  and csa_tree_add_117_21_pad_groupi_g4027(csa_tree_add_117_21_pad_groupi_n_378 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_99);
  and csa_tree_add_117_21_pad_groupi_g4028(csa_tree_add_117_21_pad_groupi_n_377 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_88);
  and csa_tree_add_117_21_pad_groupi_g4029(csa_tree_add_117_21_pad_groupi_n_376 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_88);
  and csa_tree_add_117_21_pad_groupi_g4030(csa_tree_add_117_21_pad_groupi_n_375 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_142);
  and csa_tree_add_117_21_pad_groupi_g4031(csa_tree_add_117_21_pad_groupi_n_374 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_157);
  and csa_tree_add_117_21_pad_groupi_g4032(csa_tree_add_117_21_pad_groupi_n_373 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_143);
  and csa_tree_add_117_21_pad_groupi_g4033(csa_tree_add_117_21_pad_groupi_n_372 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_157);
  and csa_tree_add_117_21_pad_groupi_g4034(csa_tree_add_117_21_pad_groupi_n_371 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_93);
  and csa_tree_add_117_21_pad_groupi_g4035(csa_tree_add_117_21_pad_groupi_n_370 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_158);
  and csa_tree_add_117_21_pad_groupi_g4036(csa_tree_add_117_21_pad_groupi_n_369 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_158);
  and csa_tree_add_117_21_pad_groupi_g4037(csa_tree_add_117_21_pad_groupi_n_368 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_143);
  and csa_tree_add_117_21_pad_groupi_g4038(csa_tree_add_117_21_pad_groupi_n_367 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_87);
  and csa_tree_add_117_21_pad_groupi_g4039(csa_tree_add_117_21_pad_groupi_n_366 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_65);
  and csa_tree_add_117_21_pad_groupi_g4040(csa_tree_add_117_21_pad_groupi_n_365 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_118);
  and csa_tree_add_117_21_pad_groupi_g4041(csa_tree_add_117_21_pad_groupi_n_364 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_91);
  and csa_tree_add_117_21_pad_groupi_g4042(csa_tree_add_117_21_pad_groupi_n_363 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_117);
  and csa_tree_add_117_21_pad_groupi_g4043(csa_tree_add_117_21_pad_groupi_n_362 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_91);
  and csa_tree_add_117_21_pad_groupi_g4044(csa_tree_add_117_21_pad_groupi_n_361 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_142);
  and csa_tree_add_117_21_pad_groupi_g4045(csa_tree_add_117_21_pad_groupi_n_360 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_137);
  and csa_tree_add_117_21_pad_groupi_g4046(csa_tree_add_117_21_pad_groupi_n_359 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_87);
  and csa_tree_add_117_21_pad_groupi_g4047(csa_tree_add_117_21_pad_groupi_n_358 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_118);
  and csa_tree_add_117_21_pad_groupi_g4048(csa_tree_add_117_21_pad_groupi_n_357 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_94);
  and csa_tree_add_117_21_pad_groupi_g4049(csa_tree_add_117_21_pad_groupi_n_356 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_136);
  and csa_tree_add_117_21_pad_groupi_g4050(csa_tree_add_117_21_pad_groupi_n_355 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_97);
  and csa_tree_add_117_21_pad_groupi_g4051(csa_tree_add_117_21_pad_groupi_n_394 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_136);
  or csa_tree_add_117_21_pad_groupi_g4053(csa_tree_add_117_21_pad_groupi_n_353 ,csa_tree_add_117_21_pad_groupi_n_56 ,csa_tree_add_117_21_pad_groupi_n_82);
  and csa_tree_add_117_21_pad_groupi_g4055(csa_tree_add_117_21_pad_groupi_n_392 ,csa_tree_add_117_21_pad_groupi_n_324 ,csa_tree_add_117_21_pad_groupi_n_78);
  and csa_tree_add_117_21_pad_groupi_g4056(csa_tree_add_117_21_pad_groupi_n_391 ,csa_tree_add_117_21_pad_groupi_n_323 ,csa_tree_add_117_21_pad_groupi_n_80);
  and csa_tree_add_117_21_pad_groupi_g4057(csa_tree_add_117_21_pad_groupi_n_390 ,csa_tree_add_117_21_pad_groupi_n_325 ,csa_tree_add_117_21_pad_groupi_n_79);
  not csa_tree_add_117_21_pad_groupi_g4060(csa_tree_add_117_21_pad_groupi_n_350 ,csa_tree_add_117_21_pad_groupi_n_348);
  not csa_tree_add_117_21_pad_groupi_g4061(csa_tree_add_117_21_pad_groupi_n_349 ,csa_tree_add_117_21_pad_groupi_n_348);
  or csa_tree_add_117_21_pad_groupi_g4062(csa_tree_add_117_21_pad_groupi_n_348 ,csa_tree_add_117_21_pad_groupi_n_70 ,csa_tree_add_117_21_pad_groupi_n_320);
  not csa_tree_add_117_21_pad_groupi_g4063(csa_tree_add_117_21_pad_groupi_n_347 ,csa_tree_add_117_21_pad_groupi_n_82);
  not csa_tree_add_117_21_pad_groupi_g4064(csa_tree_add_117_21_pad_groupi_n_346 ,csa_tree_add_117_21_pad_groupi_n_78);
  xnor csa_tree_add_117_21_pad_groupi_g4067(csa_tree_add_117_21_pad_groupi_n_345 ,csa_tree_add_117_21_pad_groupi_n_289 ,csa_tree_add_117_21_pad_groupi_n_309);
  xnor csa_tree_add_117_21_pad_groupi_g4068(csa_tree_add_117_21_pad_groupi_n_344 ,csa_tree_add_117_21_pad_groupi_n_296 ,csa_tree_add_117_21_pad_groupi_n_45);
  not csa_tree_add_117_21_pad_groupi_g4069(csa_tree_add_117_21_pad_groupi_n_343 ,csa_tree_add_117_21_pad_groupi_n_341);
  not csa_tree_add_117_21_pad_groupi_g4070(csa_tree_add_117_21_pad_groupi_n_342 ,csa_tree_add_117_21_pad_groupi_n_341);
  not csa_tree_add_117_21_pad_groupi_g4072(csa_tree_add_117_21_pad_groupi_n_340 ,csa_tree_add_117_21_pad_groupi_n_81);
  not csa_tree_add_117_21_pad_groupi_g4073(csa_tree_add_117_21_pad_groupi_n_339 ,csa_tree_add_117_21_pad_groupi_n_80);
  xnor csa_tree_add_117_21_pad_groupi_g4076(csa_tree_add_117_21_pad_groupi_n_338 ,csa_tree_add_117_21_pad_groupi_n_319 ,csa_tree_add_117_21_pad_groupi_n_312);
  not csa_tree_add_117_21_pad_groupi_g4077(csa_tree_add_117_21_pad_groupi_n_337 ,csa_tree_add_117_21_pad_groupi_n_77);
  not csa_tree_add_117_21_pad_groupi_g4078(csa_tree_add_117_21_pad_groupi_n_336 ,csa_tree_add_117_21_pad_groupi_n_79);
  xnor csa_tree_add_117_21_pad_groupi_g4081(csa_tree_add_117_21_pad_groupi_n_335 ,csa_tree_add_117_21_pad_groupi_n_318 ,csa_tree_add_117_21_pad_groupi_n_310);
  not csa_tree_add_117_21_pad_groupi_g4082(csa_tree_add_117_21_pad_groupi_n_334 ,csa_tree_add_117_21_pad_groupi_n_333);
  not csa_tree_add_117_21_pad_groupi_g4085(csa_tree_add_117_21_pad_groupi_n_332 ,csa_tree_add_117_21_pad_groupi_n_74);
  and csa_tree_add_117_21_pad_groupi_g4087(csa_tree_add_117_21_pad_groupi_n_333 ,csa_tree_add_117_21_pad_groupi_n_314 ,csa_tree_add_117_21_pad_groupi_n_315);
  not csa_tree_add_117_21_pad_groupi_g4088(csa_tree_add_117_21_pad_groupi_n_331 ,csa_tree_add_117_21_pad_groupi_n_330);
  not csa_tree_add_117_21_pad_groupi_g4091(csa_tree_add_117_21_pad_groupi_n_329 ,csa_tree_add_117_21_pad_groupi_n_75);
  and csa_tree_add_117_21_pad_groupi_g4093(csa_tree_add_117_21_pad_groupi_n_330 ,csa_tree_add_117_21_pad_groupi_n_319 ,csa_tree_add_117_21_pad_groupi_n_317);
  not csa_tree_add_117_21_pad_groupi_g4094(csa_tree_add_117_21_pad_groupi_n_328 ,csa_tree_add_117_21_pad_groupi_n_327);
  not csa_tree_add_117_21_pad_groupi_g4097(csa_tree_add_117_21_pad_groupi_n_326 ,csa_tree_add_117_21_pad_groupi_n_76);
  and csa_tree_add_117_21_pad_groupi_g4099(csa_tree_add_117_21_pad_groupi_n_327 ,csa_tree_add_117_21_pad_groupi_n_318 ,csa_tree_add_117_21_pad_groupi_n_316);
  xnor csa_tree_add_117_21_pad_groupi_g4100(csa_tree_add_117_21_pad_groupi_n_325 ,csa_tree_add_117_21_pad_groupi_n_257 ,csa_tree_add_117_21_pad_groupi_n_283);
  xnor csa_tree_add_117_21_pad_groupi_g4101(csa_tree_add_117_21_pad_groupi_n_324 ,csa_tree_add_117_21_pad_groupi_n_259 ,csa_tree_add_117_21_pad_groupi_n_279);
  xnor csa_tree_add_117_21_pad_groupi_g4102(csa_tree_add_117_21_pad_groupi_n_323 ,csa_tree_add_117_21_pad_groupi_n_261 ,csa_tree_add_117_21_pad_groupi_n_281);
  xnor csa_tree_add_117_21_pad_groupi_g4105(csa_tree_add_117_21_pad_groupi_n_320 ,csa_tree_add_117_21_pad_groupi_n_297 ,csa_tree_add_117_21_pad_groupi_n_255);
  or csa_tree_add_117_21_pad_groupi_g4106(csa_tree_add_117_21_pad_groupi_n_317 ,csa_tree_add_117_21_pad_groupi_n_259 ,csa_tree_add_117_21_pad_groupi_n_292);
  or csa_tree_add_117_21_pad_groupi_g4107(csa_tree_add_117_21_pad_groupi_n_316 ,csa_tree_add_117_21_pad_groupi_n_261 ,csa_tree_add_117_21_pad_groupi_n_290);
  or csa_tree_add_117_21_pad_groupi_g4108(csa_tree_add_117_21_pad_groupi_n_315 ,csa_tree_add_117_21_pad_groupi_n_257 ,csa_tree_add_117_21_pad_groupi_n_294);
  or csa_tree_add_117_21_pad_groupi_g4109(csa_tree_add_117_21_pad_groupi_n_319 ,csa_tree_add_117_21_pad_groupi_n_258 ,csa_tree_add_117_21_pad_groupi_n_293);
  or csa_tree_add_117_21_pad_groupi_g4110(csa_tree_add_117_21_pad_groupi_n_318 ,csa_tree_add_117_21_pad_groupi_n_260 ,csa_tree_add_117_21_pad_groupi_n_291);
  xnor csa_tree_add_117_21_pad_groupi_g4111(csa_tree_add_117_21_pad_groupi_n_312 ,csa_tree_add_117_21_pad_groupi_n_277 ,csa_tree_add_117_21_pad_groupi_n_239);
  xnor csa_tree_add_117_21_pad_groupi_g4113(csa_tree_add_117_21_pad_groupi_n_310 ,csa_tree_add_117_21_pad_groupi_n_262 ,csa_tree_add_117_21_pad_groupi_n_229);
  xnor csa_tree_add_117_21_pad_groupi_g4114(csa_tree_add_117_21_pad_groupi_n_309 ,csa_tree_add_117_21_pad_groupi_n_264 ,csa_tree_add_117_21_pad_groupi_n_240);
  or csa_tree_add_117_21_pad_groupi_g4115(csa_tree_add_117_21_pad_groupi_n_314 ,csa_tree_add_117_21_pad_groupi_n_256 ,csa_tree_add_117_21_pad_groupi_n_295);
  and csa_tree_add_117_21_pad_groupi_g4116(csa_tree_add_117_21_pad_groupi_n_313 ,csa_tree_add_117_21_pad_groupi_n_284 ,csa_tree_add_117_21_pad_groupi_n_289);
  and csa_tree_add_117_21_pad_groupi_g4117(csa_tree_add_117_21_pad_groupi_n_307 ,in3[10] ,csa_tree_add_117_21_pad_groupi_n_133);
  and csa_tree_add_117_21_pad_groupi_g4118(csa_tree_add_117_21_pad_groupi_n_306 ,in3[5] ,csa_tree_add_117_21_pad_groupi_n_58);
  and csa_tree_add_117_21_pad_groupi_g4119(csa_tree_add_117_21_pad_groupi_n_305 ,in3[11] ,csa_tree_add_117_21_pad_groupi_n_62);
  and csa_tree_add_117_21_pad_groupi_g4120(csa_tree_add_117_21_pad_groupi_n_304 ,in3[12] ,csa_tree_add_117_21_pad_groupi_n_133);
  and csa_tree_add_117_21_pad_groupi_g4121(csa_tree_add_117_21_pad_groupi_n_303 ,in3[8] ,csa_tree_add_117_21_pad_groupi_n_84);
  and csa_tree_add_117_21_pad_groupi_g4122(csa_tree_add_117_21_pad_groupi_n_302 ,in3[1] ,csa_tree_add_117_21_pad_groupi_n_59);
  and csa_tree_add_117_21_pad_groupi_g4123(csa_tree_add_117_21_pad_groupi_n_301 ,in3[6] ,csa_tree_add_117_21_pad_groupi_n_62);
  and csa_tree_add_117_21_pad_groupi_g4124(csa_tree_add_117_21_pad_groupi_n_300 ,in3[14] ,csa_tree_add_117_21_pad_groupi_n_85);
  and csa_tree_add_117_21_pad_groupi_g4125(csa_tree_add_117_21_pad_groupi_n_299 ,in3[9] ,csa_tree_add_117_21_pad_groupi_n_59);
  and csa_tree_add_117_21_pad_groupi_g4126(csa_tree_add_117_21_pad_groupi_n_298 ,in3[4] ,csa_tree_add_117_21_pad_groupi_n_61);
  nor csa_tree_add_117_21_pad_groupi_g4127(csa_tree_add_117_21_pad_groupi_n_297 ,n_471 ,csa_tree_add_117_21_pad_groupi_n_71);
  and csa_tree_add_117_21_pad_groupi_g4128(csa_tree_add_117_21_pad_groupi_n_308 ,in3[15] ,csa_tree_add_117_21_pad_groupi_n_70);
  or csa_tree_add_117_21_pad_groupi_g4129(csa_tree_add_117_21_pad_groupi_n_296 ,csa_tree_add_117_21_pad_groupi_n_55 ,csa_tree_add_117_21_pad_groupi_n_131);
  not csa_tree_add_117_21_pad_groupi_g4130(csa_tree_add_117_21_pad_groupi_n_295 ,csa_tree_add_117_21_pad_groupi_n_294);
  not csa_tree_add_117_21_pad_groupi_g4131(csa_tree_add_117_21_pad_groupi_n_293 ,csa_tree_add_117_21_pad_groupi_n_292);
  not csa_tree_add_117_21_pad_groupi_g4132(csa_tree_add_117_21_pad_groupi_n_291 ,csa_tree_add_117_21_pad_groupi_n_290);
  and csa_tree_add_117_21_pad_groupi_g4133(csa_tree_add_117_21_pad_groupi_n_288 ,in3[7] ,csa_tree_add_117_21_pad_groupi_n_134);
  and csa_tree_add_117_21_pad_groupi_g4134(csa_tree_add_117_21_pad_groupi_n_287 ,in3[3] ,csa_tree_add_117_21_pad_groupi_n_84);
  and csa_tree_add_117_21_pad_groupi_g4135(csa_tree_add_117_21_pad_groupi_n_286 ,in3[2] ,csa_tree_add_117_21_pad_groupi_n_85);
  and csa_tree_add_117_21_pad_groupi_g4136(csa_tree_add_117_21_pad_groupi_n_285 ,in3[13] ,csa_tree_add_117_21_pad_groupi_n_134);
  or csa_tree_add_117_21_pad_groupi_g4137(csa_tree_add_117_21_pad_groupi_n_284 ,csa_tree_add_117_21_pad_groupi_n_248 ,csa_tree_add_117_21_pad_groupi_n_255);
  or csa_tree_add_117_21_pad_groupi_g4138(csa_tree_add_117_21_pad_groupi_n_283 ,csa_tree_add_117_21_pad_groupi_n_263 ,csa_tree_add_117_21_pad_groupi_n_250);
  or csa_tree_add_117_21_pad_groupi_g4140(csa_tree_add_117_21_pad_groupi_n_281 ,csa_tree_add_117_21_pad_groupi_n_278 ,csa_tree_add_117_21_pad_groupi_n_249);
  or csa_tree_add_117_21_pad_groupi_g4141(csa_tree_add_117_21_pad_groupi_n_294 ,csa_tree_add_117_21_pad_groupi_n_231 ,csa_tree_add_117_21_pad_groupi_n_271);
  or csa_tree_add_117_21_pad_groupi_g4143(csa_tree_add_117_21_pad_groupi_n_292 ,csa_tree_add_117_21_pad_groupi_n_232 ,csa_tree_add_117_21_pad_groupi_n_272);
  or csa_tree_add_117_21_pad_groupi_g4144(csa_tree_add_117_21_pad_groupi_n_290 ,csa_tree_add_117_21_pad_groupi_n_235 ,csa_tree_add_117_21_pad_groupi_n_273);
  or csa_tree_add_117_21_pad_groupi_g4145(csa_tree_add_117_21_pad_groupi_n_279 ,csa_tree_add_117_21_pad_groupi_n_265 ,csa_tree_add_117_21_pad_groupi_n_269);
  or csa_tree_add_117_21_pad_groupi_g4146(csa_tree_add_117_21_pad_groupi_n_289 ,csa_tree_add_117_21_pad_groupi_n_247 ,csa_tree_add_117_21_pad_groupi_n_254);
  not csa_tree_add_117_21_pad_groupi_g4147(csa_tree_add_117_21_pad_groupi_n_278 ,csa_tree_add_117_21_pad_groupi_n_277);
  not csa_tree_add_117_21_pad_groupi_g4148(csa_tree_add_117_21_pad_groupi_n_276 ,csa_tree_add_117_21_pad_groupi_n_274);
  not csa_tree_add_117_21_pad_groupi_g4149(csa_tree_add_117_21_pad_groupi_n_275 ,csa_tree_add_117_21_pad_groupi_n_131);
  and csa_tree_add_117_21_pad_groupi_g4151(csa_tree_add_117_21_pad_groupi_n_273 ,n_467 ,csa_tree_add_117_21_pad_groupi_n_243);
  and csa_tree_add_117_21_pad_groupi_g4152(csa_tree_add_117_21_pad_groupi_n_272 ,n_469 ,csa_tree_add_117_21_pad_groupi_n_245);
  and csa_tree_add_117_21_pad_groupi_g4153(csa_tree_add_117_21_pad_groupi_n_271 ,n_465 ,csa_tree_add_117_21_pad_groupi_n_237);
  xnor csa_tree_add_117_21_pad_groupi_g4156(csa_tree_add_117_21_pad_groupi_n_268 ,in4[10] ,in4[9]);
  xnor csa_tree_add_117_21_pad_groupi_g4157(csa_tree_add_117_21_pad_groupi_n_267 ,in4[11] ,in4[10]);
  xnor csa_tree_add_117_21_pad_groupi_g4158(csa_tree_add_117_21_pad_groupi_n_266 ,in4[13] ,in4[12]);
  xnor csa_tree_add_117_21_pad_groupi_g4159(csa_tree_add_117_21_pad_groupi_n_277 ,n_467 ,n_458);
  xnor csa_tree_add_117_21_pad_groupi_g4160(csa_tree_add_117_21_pad_groupi_n_274 ,n_471 ,n_462);
  not csa_tree_add_117_21_pad_groupi_g4161(csa_tree_add_117_21_pad_groupi_n_265 ,csa_tree_add_117_21_pad_groupi_n_264);
  not csa_tree_add_117_21_pad_groupi_g4162(csa_tree_add_117_21_pad_groupi_n_263 ,csa_tree_add_117_21_pad_groupi_n_262);
  not csa_tree_add_117_21_pad_groupi_g4163(csa_tree_add_117_21_pad_groupi_n_260 ,csa_tree_add_117_21_pad_groupi_n_261);
  not csa_tree_add_117_21_pad_groupi_g4164(csa_tree_add_117_21_pad_groupi_n_258 ,csa_tree_add_117_21_pad_groupi_n_259);
  not csa_tree_add_117_21_pad_groupi_g4165(csa_tree_add_117_21_pad_groupi_n_256 ,csa_tree_add_117_21_pad_groupi_n_257);
  not csa_tree_add_117_21_pad_groupi_g4166(csa_tree_add_117_21_pad_groupi_n_254 ,csa_tree_add_117_21_pad_groupi_n_255);
  xor csa_tree_add_117_21_pad_groupi_g4169(csa_tree_add_117_21_pad_groupi_n_250 ,n_465 ,n_466);
  xor csa_tree_add_117_21_pad_groupi_g4170(csa_tree_add_117_21_pad_groupi_n_249 ,n_467 ,n_468);
  xnor csa_tree_add_117_21_pad_groupi_g4171(csa_tree_add_117_21_pad_groupi_n_264 ,n_469 ,n_460);
  xnor csa_tree_add_117_21_pad_groupi_g4172(csa_tree_add_117_21_pad_groupi_n_262 ,n_465 ,n_456);
  xnor csa_tree_add_117_21_pad_groupi_g4173(csa_tree_add_117_21_pad_groupi_n_261 ,csa_tree_add_117_21_pad_groupi_n_129 ,n_466);
  xnor csa_tree_add_117_21_pad_groupi_g4174(csa_tree_add_117_21_pad_groupi_n_259 ,csa_tree_add_117_21_pad_groupi_n_126 ,n_468);
  xnor csa_tree_add_117_21_pad_groupi_g4176(csa_tree_add_117_21_pad_groupi_n_255 ,n_470 ,in1[0]);
  not csa_tree_add_117_21_pad_groupi_g4178(csa_tree_add_117_21_pad_groupi_n_248 ,csa_tree_add_117_21_pad_groupi_n_247);
  or csa_tree_add_117_21_pad_groupi_g4179(csa_tree_add_117_21_pad_groupi_n_246 ,csa_tree_add_117_21_pad_groupi_n_213 ,in4[10]);
  or csa_tree_add_117_21_pad_groupi_g4180(csa_tree_add_117_21_pad_groupi_n_245 ,n_460 ,in1[0]);
  or csa_tree_add_117_21_pad_groupi_g4182(csa_tree_add_117_21_pad_groupi_n_243 ,n_458 ,csa_tree_add_117_21_pad_groupi_n_126);
  nor csa_tree_add_117_21_pad_groupi_g4184(csa_tree_add_117_21_pad_groupi_n_241 ,csa_tree_add_117_21_pad_groupi_n_222 ,in4[9]);
  nor csa_tree_add_117_21_pad_groupi_g4185(csa_tree_add_117_21_pad_groupi_n_240 ,in1[0] ,n_470);
  nor csa_tree_add_117_21_pad_groupi_g4186(csa_tree_add_117_21_pad_groupi_n_239 ,csa_tree_add_117_21_pad_groupi_n_127 ,n_468);
  or csa_tree_add_117_21_pad_groupi_g4187(csa_tree_add_117_21_pad_groupi_n_247 ,csa_tree_add_117_21_pad_groupi_n_220 ,csa_tree_add_117_21_pad_groupi_n_219);
  or csa_tree_add_117_21_pad_groupi_g4188(csa_tree_add_117_21_pad_groupi_n_238 ,csa_tree_add_117_21_pad_groupi_n_225 ,csa_tree_add_117_21_pad_groupi_n_214);
  or csa_tree_add_117_21_pad_groupi_g4189(csa_tree_add_117_21_pad_groupi_n_237 ,n_456 ,csa_tree_add_117_21_pad_groupi_n_129);
  nor csa_tree_add_117_21_pad_groupi_g4190(csa_tree_add_117_21_pad_groupi_n_236 ,in4[11] ,in4[10]);
  and csa_tree_add_117_21_pad_groupi_g4191(csa_tree_add_117_21_pad_groupi_n_235 ,n_458 ,csa_tree_add_117_21_pad_groupi_n_127);
  nor csa_tree_add_117_21_pad_groupi_g4192(csa_tree_add_117_21_pad_groupi_n_234 ,in4[13] ,in4[12]);
  or csa_tree_add_117_21_pad_groupi_g4193(csa_tree_add_117_21_pad_groupi_n_233 ,csa_tree_add_117_21_pad_groupi_n_228 ,csa_tree_add_117_21_pad_groupi_n_222);
  and csa_tree_add_117_21_pad_groupi_g4194(csa_tree_add_117_21_pad_groupi_n_232 ,n_460 ,in1[0]);
  and csa_tree_add_117_21_pad_groupi_g4195(csa_tree_add_117_21_pad_groupi_n_231 ,n_456 ,csa_tree_add_117_21_pad_groupi_n_130);
  nor csa_tree_add_117_21_pad_groupi_g4197(csa_tree_add_117_21_pad_groupi_n_229 ,csa_tree_add_117_21_pad_groupi_n_130 ,n_466);
  not csa_tree_add_117_21_pad_groupi_g4198(csa_tree_add_117_21_pad_groupi_n_228 ,in4[11]);
  not csa_tree_add_117_21_pad_groupi_g4199(csa_tree_add_117_21_pad_groupi_n_227 ,in4[6]);
  not csa_tree_add_117_21_pad_groupi_g4200(csa_tree_add_117_21_pad_groupi_n_226 ,in4[5]);
  not csa_tree_add_117_21_pad_groupi_g4201(csa_tree_add_117_21_pad_groupi_n_225 ,in4[13]);
  not csa_tree_add_117_21_pad_groupi_g4202(csa_tree_add_117_21_pad_groupi_n_224 ,in4[0]);
  not csa_tree_add_117_21_pad_groupi_g4203(csa_tree_add_117_21_pad_groupi_n_223 ,in4[8]);
  not csa_tree_add_117_21_pad_groupi_g4204(csa_tree_add_117_21_pad_groupi_n_222 ,in4[10]);
  not csa_tree_add_117_21_pad_groupi_g4205(csa_tree_add_117_21_pad_groupi_n_221 ,in3[0]);
  not csa_tree_add_117_21_pad_groupi_g4206(csa_tree_add_117_21_pad_groupi_n_220 ,n_462);
  not csa_tree_add_117_21_pad_groupi_g4207(csa_tree_add_117_21_pad_groupi_n_219 ,n_471);
  not csa_tree_add_117_21_pad_groupi_g4208(csa_tree_add_117_21_pad_groupi_n_218 ,in4[2]);
  not csa_tree_add_117_21_pad_groupi_g4209(csa_tree_add_117_21_pad_groupi_n_217 ,in4[7]);
  not csa_tree_add_117_21_pad_groupi_g4210(csa_tree_add_117_21_pad_groupi_n_216 ,in4[4]);
  not csa_tree_add_117_21_pad_groupi_g4211(csa_tree_add_117_21_pad_groupi_n_215 ,in4[3]);
  not csa_tree_add_117_21_pad_groupi_g4212(csa_tree_add_117_21_pad_groupi_n_214 ,in4[12]);
  not csa_tree_add_117_21_pad_groupi_g4213(csa_tree_add_117_21_pad_groupi_n_213 ,in4[9]);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4295(csa_tree_add_117_21_pad_groupi_n_197 ,csa_tree_add_117_21_pad_groupi_n_195);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4296(csa_tree_add_117_21_pad_groupi_n_196 ,csa_tree_add_117_21_pad_groupi_n_195);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4297(csa_tree_add_117_21_pad_groupi_n_195 ,csa_tree_add_117_21_pad_groupi_n_332);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4299(csa_tree_add_117_21_pad_groupi_n_194 ,csa_tree_add_117_21_pad_groupi_n_192);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4300(csa_tree_add_117_21_pad_groupi_n_193 ,csa_tree_add_117_21_pad_groupi_n_192);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4301(csa_tree_add_117_21_pad_groupi_n_192 ,csa_tree_add_117_21_pad_groupi_n_203);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4303(csa_tree_add_117_21_pad_groupi_n_191 ,csa_tree_add_117_21_pad_groupi_n_189);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4304(csa_tree_add_117_21_pad_groupi_n_190 ,csa_tree_add_117_21_pad_groupi_n_189);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4305(csa_tree_add_117_21_pad_groupi_n_189 ,csa_tree_add_117_21_pad_groupi_n_204);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4307(csa_tree_add_117_21_pad_groupi_n_188 ,csa_tree_add_117_21_pad_groupi_n_186);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4308(csa_tree_add_117_21_pad_groupi_n_187 ,csa_tree_add_117_21_pad_groupi_n_186);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4309(csa_tree_add_117_21_pad_groupi_n_186 ,csa_tree_add_117_21_pad_groupi_n_329);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4311(csa_tree_add_117_21_pad_groupi_n_185 ,csa_tree_add_117_21_pad_groupi_n_183);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4312(csa_tree_add_117_21_pad_groupi_n_184 ,csa_tree_add_117_21_pad_groupi_n_183);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4313(csa_tree_add_117_21_pad_groupi_n_183 ,csa_tree_add_117_21_pad_groupi_n_202);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4315(csa_tree_add_117_21_pad_groupi_n_182 ,csa_tree_add_117_21_pad_groupi_n_180);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4316(csa_tree_add_117_21_pad_groupi_n_181 ,csa_tree_add_117_21_pad_groupi_n_180);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4317(csa_tree_add_117_21_pad_groupi_n_180 ,csa_tree_add_117_21_pad_groupi_n_326);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4319(csa_tree_add_117_21_pad_groupi_n_179 ,csa_tree_add_117_21_pad_groupi_n_177);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4320(csa_tree_add_117_21_pad_groupi_n_178 ,csa_tree_add_117_21_pad_groupi_n_177);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4321(csa_tree_add_117_21_pad_groupi_n_177 ,csa_tree_add_117_21_pad_groupi_n_199);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4323(csa_tree_add_117_21_pad_groupi_n_176 ,csa_tree_add_117_21_pad_groupi_n_174);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4324(csa_tree_add_117_21_pad_groupi_n_175 ,csa_tree_add_117_21_pad_groupi_n_174);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4325(csa_tree_add_117_21_pad_groupi_n_174 ,csa_tree_add_117_21_pad_groupi_n_200);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4327(csa_tree_add_117_21_pad_groupi_n_173 ,csa_tree_add_117_21_pad_groupi_n_171);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4328(csa_tree_add_117_21_pad_groupi_n_172 ,csa_tree_add_117_21_pad_groupi_n_171);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4329(csa_tree_add_117_21_pad_groupi_n_171 ,csa_tree_add_117_21_pad_groupi_n_201);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4331(csa_tree_add_117_21_pad_groupi_n_170 ,csa_tree_add_117_21_pad_groupi_n_168);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4332(csa_tree_add_117_21_pad_groupi_n_169 ,csa_tree_add_117_21_pad_groupi_n_168);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4333(csa_tree_add_117_21_pad_groupi_n_168 ,csa_tree_add_117_21_pad_groupi_n_200);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4335(csa_tree_add_117_21_pad_groupi_n_167 ,csa_tree_add_117_21_pad_groupi_n_165);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4336(csa_tree_add_117_21_pad_groupi_n_166 ,csa_tree_add_117_21_pad_groupi_n_165);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4337(csa_tree_add_117_21_pad_groupi_n_165 ,csa_tree_add_117_21_pad_groupi_n_204);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4339(csa_tree_add_117_21_pad_groupi_n_164 ,csa_tree_add_117_21_pad_groupi_n_162);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4340(csa_tree_add_117_21_pad_groupi_n_163 ,csa_tree_add_117_21_pad_groupi_n_162);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4341(csa_tree_add_117_21_pad_groupi_n_162 ,csa_tree_add_117_21_pad_groupi_n_202);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4343(csa_tree_add_117_21_pad_groupi_n_161 ,csa_tree_add_117_21_pad_groupi_n_159);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4344(csa_tree_add_117_21_pad_groupi_n_160 ,csa_tree_add_117_21_pad_groupi_n_159);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4345(csa_tree_add_117_21_pad_groupi_n_159 ,csa_tree_add_117_21_pad_groupi_n_339);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4347(csa_tree_add_117_21_pad_groupi_n_158 ,csa_tree_add_117_21_pad_groupi_n_156);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4348(csa_tree_add_117_21_pad_groupi_n_157 ,csa_tree_add_117_21_pad_groupi_n_156);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4349(csa_tree_add_117_21_pad_groupi_n_156 ,csa_tree_add_117_21_pad_groupi_n_209);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4351(csa_tree_add_117_21_pad_groupi_n_155 ,csa_tree_add_117_21_pad_groupi_n_153);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4352(csa_tree_add_117_21_pad_groupi_n_154 ,csa_tree_add_117_21_pad_groupi_n_153);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4353(csa_tree_add_117_21_pad_groupi_n_153 ,csa_tree_add_117_21_pad_groupi_n_336);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4355(csa_tree_add_117_21_pad_groupi_n_152 ,csa_tree_add_117_21_pad_groupi_n_150);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4356(csa_tree_add_117_21_pad_groupi_n_151 ,csa_tree_add_117_21_pad_groupi_n_150);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4357(csa_tree_add_117_21_pad_groupi_n_150 ,csa_tree_add_117_21_pad_groupi_n_340);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4359(csa_tree_add_117_21_pad_groupi_n_149 ,csa_tree_add_117_21_pad_groupi_n_147);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4360(csa_tree_add_117_21_pad_groupi_n_148 ,csa_tree_add_117_21_pad_groupi_n_147);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4361(csa_tree_add_117_21_pad_groupi_n_147 ,csa_tree_add_117_21_pad_groupi_n_337);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4363(csa_tree_add_117_21_pad_groupi_n_146 ,csa_tree_add_117_21_pad_groupi_n_144);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4364(csa_tree_add_117_21_pad_groupi_n_145 ,csa_tree_add_117_21_pad_groupi_n_144);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4365(csa_tree_add_117_21_pad_groupi_n_144 ,csa_tree_add_117_21_pad_groupi_n_207);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4367(csa_tree_add_117_21_pad_groupi_n_143 ,csa_tree_add_117_21_pad_groupi_n_141);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4368(csa_tree_add_117_21_pad_groupi_n_142 ,csa_tree_add_117_21_pad_groupi_n_141);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4369(csa_tree_add_117_21_pad_groupi_n_141 ,csa_tree_add_117_21_pad_groupi_n_347);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4371(csa_tree_add_117_21_pad_groupi_n_140 ,csa_tree_add_117_21_pad_groupi_n_138);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4372(csa_tree_add_117_21_pad_groupi_n_139 ,csa_tree_add_117_21_pad_groupi_n_138);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4373(csa_tree_add_117_21_pad_groupi_n_138 ,csa_tree_add_117_21_pad_groupi_n_205);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4375(csa_tree_add_117_21_pad_groupi_n_137 ,csa_tree_add_117_21_pad_groupi_n_135);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4376(csa_tree_add_117_21_pad_groupi_n_136 ,csa_tree_add_117_21_pad_groupi_n_135);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4377(csa_tree_add_117_21_pad_groupi_n_135 ,csa_tree_add_117_21_pad_groupi_n_346);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4379(csa_tree_add_117_21_pad_groupi_n_134 ,csa_tree_add_117_21_pad_groupi_n_132);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4380(csa_tree_add_117_21_pad_groupi_n_133 ,csa_tree_add_117_21_pad_groupi_n_132);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4381(csa_tree_add_117_21_pad_groupi_n_132 ,csa_tree_add_117_21_pad_groupi_n_198);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4384(csa_tree_add_117_21_pad_groupi_n_131 ,csa_tree_add_117_21_pad_groupi_n_198);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4385(csa_tree_add_117_21_pad_groupi_n_198 ,csa_tree_add_117_21_pad_groupi_n_274);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4387(csa_tree_add_117_21_pad_groupi_n_130 ,csa_tree_add_117_21_pad_groupi_n_128);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4388(csa_tree_add_117_21_pad_groupi_n_129 ,csa_tree_add_117_21_pad_groupi_n_128);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4389(csa_tree_add_117_21_pad_groupi_n_128 ,n_457);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4391(csa_tree_add_117_21_pad_groupi_n_127 ,csa_tree_add_117_21_pad_groupi_n_125);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4392(csa_tree_add_117_21_pad_groupi_n_126 ,csa_tree_add_117_21_pad_groupi_n_125);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4393(csa_tree_add_117_21_pad_groupi_n_125 ,n_459);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4395(csa_tree_add_117_21_pad_groupi_n_124 ,csa_tree_add_117_21_pad_groupi_n_122);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4396(csa_tree_add_117_21_pad_groupi_n_123 ,csa_tree_add_117_21_pad_groupi_n_122);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4397(csa_tree_add_117_21_pad_groupi_n_122 ,csa_tree_add_117_21_pad_groupi_n_208);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4399(csa_tree_add_117_21_pad_groupi_n_121 ,csa_tree_add_117_21_pad_groupi_n_119);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4400(csa_tree_add_117_21_pad_groupi_n_120 ,csa_tree_add_117_21_pad_groupi_n_119);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4401(csa_tree_add_117_21_pad_groupi_n_119 ,csa_tree_add_117_21_pad_groupi_n_206);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4403(csa_tree_add_117_21_pad_groupi_n_118 ,csa_tree_add_117_21_pad_groupi_n_116);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4404(csa_tree_add_117_21_pad_groupi_n_117 ,csa_tree_add_117_21_pad_groupi_n_116);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4405(csa_tree_add_117_21_pad_groupi_n_116 ,csa_tree_add_117_21_pad_groupi_n_210);
  buf csa_tree_add_117_21_pad_groupi_drc_bufs4408(out1[1] ,csa_tree_add_117_21_pad_groupi_n_1139);
  buf csa_tree_add_117_21_pad_groupi_drc_bufs4409(out1[10] ,csa_tree_add_117_21_pad_groupi_n_1167);
  buf csa_tree_add_117_21_pad_groupi_drc_bufs4410(out1[0] ,csa_tree_add_117_21_pad_groupi_n_1129);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4413(csa_tree_add_117_21_pad_groupi_n_211 ,csa_tree_add_117_21_pad_groupi_n_643);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4420(csa_tree_add_117_21_pad_groupi_n_112 ,csa_tree_add_117_21_pad_groupi_n_110);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4421(csa_tree_add_117_21_pad_groupi_n_111 ,csa_tree_add_117_21_pad_groupi_n_110);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4422(csa_tree_add_117_21_pad_groupi_n_110 ,csa_tree_add_117_21_pad_groupi_n_313);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4440(csa_tree_add_117_21_pad_groupi_n_109 ,csa_tree_add_117_21_pad_groupi_n_108);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4442(csa_tree_add_117_21_pad_groupi_n_108 ,csa_tree_add_117_21_pad_groupi_n_392);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4445(csa_tree_add_117_21_pad_groupi_n_107 ,csa_tree_add_117_21_pad_groupi_n_106);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4447(csa_tree_add_117_21_pad_groupi_n_106 ,csa_tree_add_117_21_pad_groupi_n_391);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4450(csa_tree_add_117_21_pad_groupi_n_105 ,csa_tree_add_117_21_pad_groupi_n_104);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4452(csa_tree_add_117_21_pad_groupi_n_104 ,csa_tree_add_117_21_pad_groupi_n_390);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4455(csa_tree_add_117_21_pad_groupi_n_103 ,csa_tree_add_117_21_pad_groupi_n_101);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4456(csa_tree_add_117_21_pad_groupi_n_102 ,csa_tree_add_117_21_pad_groupi_n_101);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4457(csa_tree_add_117_21_pad_groupi_n_101 ,csa_tree_add_117_21_pad_groupi_n_343);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4459(csa_tree_add_117_21_pad_groupi_n_100 ,csa_tree_add_117_21_pad_groupi_n_98);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4460(csa_tree_add_117_21_pad_groupi_n_99 ,csa_tree_add_117_21_pad_groupi_n_98);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4461(csa_tree_add_117_21_pad_groupi_n_98 ,csa_tree_add_117_21_pad_groupi_n_342);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4463(csa_tree_add_117_21_pad_groupi_n_97 ,csa_tree_add_117_21_pad_groupi_n_95);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4464(csa_tree_add_117_21_pad_groupi_n_96 ,csa_tree_add_117_21_pad_groupi_n_95);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4465(csa_tree_add_117_21_pad_groupi_n_95 ,csa_tree_add_117_21_pad_groupi_n_343);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4467(csa_tree_add_117_21_pad_groupi_n_94 ,csa_tree_add_117_21_pad_groupi_n_92);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4468(csa_tree_add_117_21_pad_groupi_n_93 ,csa_tree_add_117_21_pad_groupi_n_92);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4469(csa_tree_add_117_21_pad_groupi_n_92 ,csa_tree_add_117_21_pad_groupi_n_350);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4471(csa_tree_add_117_21_pad_groupi_n_91 ,csa_tree_add_117_21_pad_groupi_n_89);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4472(csa_tree_add_117_21_pad_groupi_n_90 ,csa_tree_add_117_21_pad_groupi_n_89);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4473(csa_tree_add_117_21_pad_groupi_n_89 ,csa_tree_add_117_21_pad_groupi_n_350);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4475(csa_tree_add_117_21_pad_groupi_n_88 ,csa_tree_add_117_21_pad_groupi_n_86);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4476(csa_tree_add_117_21_pad_groupi_n_87 ,csa_tree_add_117_21_pad_groupi_n_86);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4477(csa_tree_add_117_21_pad_groupi_n_86 ,csa_tree_add_117_21_pad_groupi_n_349);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4479(csa_tree_add_117_21_pad_groupi_n_85 ,csa_tree_add_117_21_pad_groupi_n_83);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4480(csa_tree_add_117_21_pad_groupi_n_84 ,csa_tree_add_117_21_pad_groupi_n_83);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4481(csa_tree_add_117_21_pad_groupi_n_83 ,csa_tree_add_117_21_pad_groupi_n_275);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4485(csa_tree_add_117_21_pad_groupi_n_204 ,csa_tree_add_117_21_pad_groupi_n_333);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4489(csa_tree_add_117_21_pad_groupi_n_202 ,csa_tree_add_117_21_pad_groupi_n_330);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4493(csa_tree_add_117_21_pad_groupi_n_200 ,csa_tree_add_117_21_pad_groupi_n_327);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4495(csa_tree_add_117_21_pad_groupi_n_82 ,csa_tree_add_117_21_pad_groupi_n_210);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4497(csa_tree_add_117_21_pad_groupi_n_210 ,csa_tree_add_117_21_pad_groupi_n_345);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4499(csa_tree_add_117_21_pad_groupi_n_81 ,csa_tree_add_117_21_pad_groupi_n_208);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4501(csa_tree_add_117_21_pad_groupi_n_208 ,csa_tree_add_117_21_pad_groupi_n_338);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4503(csa_tree_add_117_21_pad_groupi_n_80 ,csa_tree_add_117_21_pad_groupi_n_207);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4505(csa_tree_add_117_21_pad_groupi_n_207 ,csa_tree_add_117_21_pad_groupi_n_338);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4507(csa_tree_add_117_21_pad_groupi_n_79 ,csa_tree_add_117_21_pad_groupi_n_205);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4509(csa_tree_add_117_21_pad_groupi_n_205 ,csa_tree_add_117_21_pad_groupi_n_335);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4511(csa_tree_add_117_21_pad_groupi_n_78 ,csa_tree_add_117_21_pad_groupi_n_209);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4513(csa_tree_add_117_21_pad_groupi_n_209 ,csa_tree_add_117_21_pad_groupi_n_345);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4515(csa_tree_add_117_21_pad_groupi_n_77 ,csa_tree_add_117_21_pad_groupi_n_206);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4517(csa_tree_add_117_21_pad_groupi_n_206 ,csa_tree_add_117_21_pad_groupi_n_335);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4519(csa_tree_add_117_21_pad_groupi_n_76 ,csa_tree_add_117_21_pad_groupi_n_199);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4521(csa_tree_add_117_21_pad_groupi_n_199 ,csa_tree_add_117_21_pad_groupi_n_327);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4523(csa_tree_add_117_21_pad_groupi_n_75 ,csa_tree_add_117_21_pad_groupi_n_201);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4525(csa_tree_add_117_21_pad_groupi_n_201 ,csa_tree_add_117_21_pad_groupi_n_330);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4527(csa_tree_add_117_21_pad_groupi_n_74 ,csa_tree_add_117_21_pad_groupi_n_203);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4529(csa_tree_add_117_21_pad_groupi_n_203 ,csa_tree_add_117_21_pad_groupi_n_333);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4532(csa_tree_add_117_21_pad_groupi_n_73 ,csa_tree_add_117_21_pad_groupi_n_72);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4533(csa_tree_add_117_21_pad_groupi_n_72 ,csa_tree_add_117_21_pad_groupi_n_221);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4535(csa_tree_add_117_21_pad_groupi_n_71 ,csa_tree_add_117_21_pad_groupi_n_69);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4536(csa_tree_add_117_21_pad_groupi_n_70 ,csa_tree_add_117_21_pad_groupi_n_69);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4537(csa_tree_add_117_21_pad_groupi_n_69 ,csa_tree_add_117_21_pad_groupi_n_275);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4539(csa_tree_add_117_21_pad_groupi_n_68 ,csa_tree_add_117_21_pad_groupi_n_66);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4540(csa_tree_add_117_21_pad_groupi_n_67 ,csa_tree_add_117_21_pad_groupi_n_66);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4541(csa_tree_add_117_21_pad_groupi_n_66 ,csa_tree_add_117_21_pad_groupi_n_342);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4543(csa_tree_add_117_21_pad_groupi_n_65 ,csa_tree_add_117_21_pad_groupi_n_63);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4544(csa_tree_add_117_21_pad_groupi_n_64 ,csa_tree_add_117_21_pad_groupi_n_63);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4545(csa_tree_add_117_21_pad_groupi_n_63 ,csa_tree_add_117_21_pad_groupi_n_349);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4547(csa_tree_add_117_21_pad_groupi_n_62 ,csa_tree_add_117_21_pad_groupi_n_60);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4548(csa_tree_add_117_21_pad_groupi_n_61 ,csa_tree_add_117_21_pad_groupi_n_60);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4549(csa_tree_add_117_21_pad_groupi_n_60 ,csa_tree_add_117_21_pad_groupi_n_276);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4551(csa_tree_add_117_21_pad_groupi_n_59 ,csa_tree_add_117_21_pad_groupi_n_57);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4552(csa_tree_add_117_21_pad_groupi_n_58 ,csa_tree_add_117_21_pad_groupi_n_57);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4553(csa_tree_add_117_21_pad_groupi_n_57 ,csa_tree_add_117_21_pad_groupi_n_276);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4555(csa_tree_add_117_21_pad_groupi_n_56 ,csa_tree_add_117_21_pad_groupi_n_54);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4556(csa_tree_add_117_21_pad_groupi_n_55 ,csa_tree_add_117_21_pad_groupi_n_54);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4557(csa_tree_add_117_21_pad_groupi_n_54 ,csa_tree_add_117_21_pad_groupi_n_221);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4559(csa_tree_add_117_21_pad_groupi_n_53 ,csa_tree_add_117_21_pad_groupi_n_51);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4560(csa_tree_add_117_21_pad_groupi_n_52 ,csa_tree_add_117_21_pad_groupi_n_51);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4561(csa_tree_add_117_21_pad_groupi_n_51 ,csa_tree_add_117_21_pad_groupi_n_313);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4564(csa_tree_add_117_21_pad_groupi_n_50 ,csa_tree_add_117_21_pad_groupi_n_49);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4565(csa_tree_add_117_21_pad_groupi_n_49 ,csa_tree_add_117_21_pad_groupi_n_112);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4567(csa_tree_add_117_21_pad_groupi_n_48 ,csa_tree_add_117_21_pad_groupi_n_46);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4568(csa_tree_add_117_21_pad_groupi_n_47 ,csa_tree_add_117_21_pad_groupi_n_46);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4569(csa_tree_add_117_21_pad_groupi_n_46 ,csa_tree_add_117_21_pad_groupi_n_313);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4571(csa_tree_add_117_21_pad_groupi_n_45 ,csa_tree_add_117_21_pad_groupi_n_43);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4572(csa_tree_add_117_21_pad_groupi_n_44 ,csa_tree_add_117_21_pad_groupi_n_43);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4573(csa_tree_add_117_21_pad_groupi_n_43 ,csa_tree_add_117_21_pad_groupi_n_111);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4575(csa_tree_add_117_21_pad_groupi_n_42 ,csa_tree_add_117_21_pad_groupi_n_40);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4576(csa_tree_add_117_21_pad_groupi_n_41 ,csa_tree_add_117_21_pad_groupi_n_40);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4577(csa_tree_add_117_21_pad_groupi_n_40 ,csa_tree_add_117_21_pad_groupi_n_107);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4579(csa_tree_add_117_21_pad_groupi_n_39 ,csa_tree_add_117_21_pad_groupi_n_37);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4580(csa_tree_add_117_21_pad_groupi_n_38 ,csa_tree_add_117_21_pad_groupi_n_37);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4581(csa_tree_add_117_21_pad_groupi_n_37 ,csa_tree_add_117_21_pad_groupi_n_109);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4583(csa_tree_add_117_21_pad_groupi_n_36 ,csa_tree_add_117_21_pad_groupi_n_34);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4584(csa_tree_add_117_21_pad_groupi_n_35 ,csa_tree_add_117_21_pad_groupi_n_34);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4585(csa_tree_add_117_21_pad_groupi_n_34 ,csa_tree_add_117_21_pad_groupi_n_109);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4587(csa_tree_add_117_21_pad_groupi_n_33 ,csa_tree_add_117_21_pad_groupi_n_31);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4588(csa_tree_add_117_21_pad_groupi_n_32 ,csa_tree_add_117_21_pad_groupi_n_31);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4589(csa_tree_add_117_21_pad_groupi_n_31 ,csa_tree_add_117_21_pad_groupi_n_391);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4591(csa_tree_add_117_21_pad_groupi_n_30 ,csa_tree_add_117_21_pad_groupi_n_28);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4592(csa_tree_add_117_21_pad_groupi_n_29 ,csa_tree_add_117_21_pad_groupi_n_28);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4593(csa_tree_add_117_21_pad_groupi_n_28 ,csa_tree_add_117_21_pad_groupi_n_391);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4595(csa_tree_add_117_21_pad_groupi_n_27 ,csa_tree_add_117_21_pad_groupi_n_25);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4596(csa_tree_add_117_21_pad_groupi_n_26 ,csa_tree_add_117_21_pad_groupi_n_25);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4597(csa_tree_add_117_21_pad_groupi_n_25 ,csa_tree_add_117_21_pad_groupi_n_390);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4599(csa_tree_add_117_21_pad_groupi_n_24 ,csa_tree_add_117_21_pad_groupi_n_22);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4600(csa_tree_add_117_21_pad_groupi_n_23 ,csa_tree_add_117_21_pad_groupi_n_22);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4601(csa_tree_add_117_21_pad_groupi_n_22 ,csa_tree_add_117_21_pad_groupi_n_390);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4603(csa_tree_add_117_21_pad_groupi_n_21 ,csa_tree_add_117_21_pad_groupi_n_19);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4604(csa_tree_add_117_21_pad_groupi_n_20 ,csa_tree_add_117_21_pad_groupi_n_19);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4605(csa_tree_add_117_21_pad_groupi_n_19 ,csa_tree_add_117_21_pad_groupi_n_392);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4607(csa_tree_add_117_21_pad_groupi_n_18 ,csa_tree_add_117_21_pad_groupi_n_16);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4608(csa_tree_add_117_21_pad_groupi_n_17 ,csa_tree_add_117_21_pad_groupi_n_16);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4609(csa_tree_add_117_21_pad_groupi_n_16 ,csa_tree_add_117_21_pad_groupi_n_392);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4611(csa_tree_add_117_21_pad_groupi_n_15 ,csa_tree_add_117_21_pad_groupi_n_13);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4612(csa_tree_add_117_21_pad_groupi_n_14 ,csa_tree_add_117_21_pad_groupi_n_13);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4613(csa_tree_add_117_21_pad_groupi_n_13 ,csa_tree_add_117_21_pad_groupi_n_105);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4615(csa_tree_add_117_21_pad_groupi_n_12 ,csa_tree_add_117_21_pad_groupi_n_10);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4616(csa_tree_add_117_21_pad_groupi_n_11 ,csa_tree_add_117_21_pad_groupi_n_10);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4617(csa_tree_add_117_21_pad_groupi_n_10 ,csa_tree_add_117_21_pad_groupi_n_105);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4619(csa_tree_add_117_21_pad_groupi_n_9 ,csa_tree_add_117_21_pad_groupi_n_7);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4620(csa_tree_add_117_21_pad_groupi_n_8 ,csa_tree_add_117_21_pad_groupi_n_7);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4621(csa_tree_add_117_21_pad_groupi_n_7 ,csa_tree_add_117_21_pad_groupi_n_107);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4623(csa_tree_add_117_21_pad_groupi_n_6 ,csa_tree_add_117_21_pad_groupi_n_5);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4625(csa_tree_add_117_21_pad_groupi_n_5 ,csa_tree_add_117_21_pad_groupi_n_53);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4627(csa_tree_add_117_21_pad_groupi_n_4 ,csa_tree_add_117_21_pad_groupi_n_3);
  not csa_tree_add_117_21_pad_groupi_drc_bufs4629(csa_tree_add_117_21_pad_groupi_n_3 ,csa_tree_add_117_21_pad_groupi_n_112);
  and csa_tree_add_117_21_pad_groupi_g2(csa_tree_add_117_21_pad_groupi_n_2 ,csa_tree_add_117_21_pad_groupi_n_714 ,csa_tree_add_117_21_pad_groupi_n_913);
  and csa_tree_add_117_21_pad_groupi_g4631(csa_tree_add_117_21_pad_groupi_n_1 ,csa_tree_add_117_21_pad_groupi_n_211 ,csa_tree_add_117_21_pad_groupi_n_637);
  xor csa_tree_add_117_21_pad_groupi_g4632(csa_tree_add_117_21_pad_groupi_n_0 ,csa_tree_add_117_21_pad_groupi_n_440 ,csa_tree_add_117_21_pad_groupi_n_3);
  xnor csa_tree_add_118_30_groupi_g641(out2[15] ,csa_tree_add_118_30_groupi_n_211 ,csa_tree_add_118_30_groupi_n_144);
  or csa_tree_add_118_30_groupi_g642(csa_tree_add_118_30_groupi_n_211 ,csa_tree_add_118_30_groupi_n_126 ,csa_tree_add_118_30_groupi_n_209);
  xnor csa_tree_add_118_30_groupi_g643(out2[14] ,csa_tree_add_118_30_groupi_n_208 ,csa_tree_add_118_30_groupi_n_153);
  and csa_tree_add_118_30_groupi_g644(csa_tree_add_118_30_groupi_n_209 ,csa_tree_add_118_30_groupi_n_130 ,csa_tree_add_118_30_groupi_n_208);
  or csa_tree_add_118_30_groupi_g645(csa_tree_add_118_30_groupi_n_208 ,csa_tree_add_118_30_groupi_n_136 ,csa_tree_add_118_30_groupi_n_206);
  xnor csa_tree_add_118_30_groupi_g646(out2[13] ,csa_tree_add_118_30_groupi_n_205 ,csa_tree_add_118_30_groupi_n_152);
  and csa_tree_add_118_30_groupi_g647(csa_tree_add_118_30_groupi_n_206 ,csa_tree_add_118_30_groupi_n_128 ,csa_tree_add_118_30_groupi_n_205);
  or csa_tree_add_118_30_groupi_g648(csa_tree_add_118_30_groupi_n_205 ,csa_tree_add_118_30_groupi_n_131 ,csa_tree_add_118_30_groupi_n_203);
  xnor csa_tree_add_118_30_groupi_g649(out2[12] ,csa_tree_add_118_30_groupi_n_202 ,csa_tree_add_118_30_groupi_n_147);
  and csa_tree_add_118_30_groupi_g650(csa_tree_add_118_30_groupi_n_203 ,csa_tree_add_118_30_groupi_n_138 ,csa_tree_add_118_30_groupi_n_202);
  or csa_tree_add_118_30_groupi_g651(csa_tree_add_118_30_groupi_n_202 ,csa_tree_add_118_30_groupi_n_137 ,csa_tree_add_118_30_groupi_n_200);
  xnor csa_tree_add_118_30_groupi_g652(out2[11] ,csa_tree_add_118_30_groupi_n_199 ,csa_tree_add_118_30_groupi_n_150);
  and csa_tree_add_118_30_groupi_g653(csa_tree_add_118_30_groupi_n_200 ,csa_tree_add_118_30_groupi_n_135 ,csa_tree_add_118_30_groupi_n_199);
  or csa_tree_add_118_30_groupi_g654(csa_tree_add_118_30_groupi_n_199 ,csa_tree_add_118_30_groupi_n_134 ,csa_tree_add_118_30_groupi_n_197);
  xnor csa_tree_add_118_30_groupi_g655(out2[10] ,csa_tree_add_118_30_groupi_n_196 ,csa_tree_add_118_30_groupi_n_149);
  and csa_tree_add_118_30_groupi_g656(csa_tree_add_118_30_groupi_n_197 ,csa_tree_add_118_30_groupi_n_129 ,csa_tree_add_118_30_groupi_n_196);
  or csa_tree_add_118_30_groupi_g657(csa_tree_add_118_30_groupi_n_196 ,csa_tree_add_118_30_groupi_n_127 ,csa_tree_add_118_30_groupi_n_194);
  xnor csa_tree_add_118_30_groupi_g658(out2[9] ,csa_tree_add_118_30_groupi_n_193 ,csa_tree_add_118_30_groupi_n_148);
  and csa_tree_add_118_30_groupi_g659(csa_tree_add_118_30_groupi_n_194 ,csa_tree_add_118_30_groupi_n_123 ,csa_tree_add_118_30_groupi_n_193);
  or csa_tree_add_118_30_groupi_g660(csa_tree_add_118_30_groupi_n_193 ,csa_tree_add_118_30_groupi_n_124 ,csa_tree_add_118_30_groupi_n_191);
  xnor csa_tree_add_118_30_groupi_g661(out2[8] ,csa_tree_add_118_30_groupi_n_190 ,csa_tree_add_118_30_groupi_n_145);
  and csa_tree_add_118_30_groupi_g662(csa_tree_add_118_30_groupi_n_191 ,csa_tree_add_118_30_groupi_n_140 ,csa_tree_add_118_30_groupi_n_190);
  or csa_tree_add_118_30_groupi_g663(csa_tree_add_118_30_groupi_n_190 ,csa_tree_add_118_30_groupi_n_139 ,csa_tree_add_118_30_groupi_n_188);
  xnor csa_tree_add_118_30_groupi_g664(out2[7] ,csa_tree_add_118_30_groupi_n_187 ,csa_tree_add_118_30_groupi_n_146);
  and csa_tree_add_118_30_groupi_g665(csa_tree_add_118_30_groupi_n_188 ,csa_tree_add_118_30_groupi_n_125 ,csa_tree_add_118_30_groupi_n_187);
  or csa_tree_add_118_30_groupi_g666(csa_tree_add_118_30_groupi_n_187 ,csa_tree_add_118_30_groupi_n_177 ,csa_tree_add_118_30_groupi_n_185);
  xnor csa_tree_add_118_30_groupi_g667(out2[6] ,csa_tree_add_118_30_groupi_n_184 ,csa_tree_add_118_30_groupi_n_179);
  and csa_tree_add_118_30_groupi_g668(csa_tree_add_118_30_groupi_n_185 ,csa_tree_add_118_30_groupi_n_176 ,csa_tree_add_118_30_groupi_n_184);
  or csa_tree_add_118_30_groupi_g669(csa_tree_add_118_30_groupi_n_184 ,csa_tree_add_118_30_groupi_n_175 ,csa_tree_add_118_30_groupi_n_182);
  xnor csa_tree_add_118_30_groupi_g670(out2[5] ,csa_tree_add_118_30_groupi_n_181 ,csa_tree_add_118_30_groupi_n_180);
  and csa_tree_add_118_30_groupi_g671(csa_tree_add_118_30_groupi_n_182 ,csa_tree_add_118_30_groupi_n_174 ,csa_tree_add_118_30_groupi_n_181);
  or csa_tree_add_118_30_groupi_g672(csa_tree_add_118_30_groupi_n_181 ,csa_tree_add_118_30_groupi_n_166 ,csa_tree_add_118_30_groupi_n_173);
  xnor csa_tree_add_118_30_groupi_g673(csa_tree_add_118_30_groupi_n_180 ,csa_tree_add_118_30_groupi_n_168 ,n_116);
  xnor csa_tree_add_118_30_groupi_g674(csa_tree_add_118_30_groupi_n_179 ,csa_tree_add_118_30_groupi_n_122 ,csa_tree_add_118_30_groupi_n_172);
  xnor csa_tree_add_118_30_groupi_g675(out2[4] ,csa_tree_add_118_30_groupi_n_171 ,csa_tree_add_118_30_groupi_n_170);
  and csa_tree_add_118_30_groupi_g676(csa_tree_add_118_30_groupi_n_177 ,csa_tree_add_118_30_groupi_n_122 ,csa_tree_add_118_30_groupi_n_172);
  or csa_tree_add_118_30_groupi_g677(csa_tree_add_118_30_groupi_n_176 ,csa_tree_add_118_30_groupi_n_122 ,csa_tree_add_118_30_groupi_n_172);
  and csa_tree_add_118_30_groupi_g678(csa_tree_add_118_30_groupi_n_175 ,n_116 ,csa_tree_add_118_30_groupi_n_168);
  or csa_tree_add_118_30_groupi_g679(csa_tree_add_118_30_groupi_n_174 ,n_116 ,csa_tree_add_118_30_groupi_n_168);
  and csa_tree_add_118_30_groupi_g680(csa_tree_add_118_30_groupi_n_173 ,csa_tree_add_118_30_groupi_n_165 ,csa_tree_add_118_30_groupi_n_171);
  or csa_tree_add_118_30_groupi_g681(csa_tree_add_118_30_groupi_n_172 ,csa_tree_add_118_30_groupi_n_43 ,csa_tree_add_118_30_groupi_n_167);
  or csa_tree_add_118_30_groupi_g682(csa_tree_add_118_30_groupi_n_171 ,csa_tree_add_118_30_groupi_n_156 ,csa_tree_add_118_30_groupi_n_164);
  xnor csa_tree_add_118_30_groupi_g683(csa_tree_add_118_30_groupi_n_170 ,csa_tree_add_118_30_groupi_n_159 ,n_115);
  xnor csa_tree_add_118_30_groupi_g684(out2[3] ,csa_tree_add_118_30_groupi_n_161 ,csa_tree_add_118_30_groupi_n_160);
  xnor csa_tree_add_118_30_groupi_g685(csa_tree_add_118_30_groupi_n_168 ,csa_tree_add_118_30_groupi_n_162 ,csa_tree_add_118_30_groupi_n_0);
  and csa_tree_add_118_30_groupi_g686(csa_tree_add_118_30_groupi_n_167 ,csa_tree_add_118_30_groupi_n_63 ,csa_tree_add_118_30_groupi_n_162);
  and csa_tree_add_118_30_groupi_g687(csa_tree_add_118_30_groupi_n_166 ,n_115 ,csa_tree_add_118_30_groupi_n_159);
  or csa_tree_add_118_30_groupi_g688(csa_tree_add_118_30_groupi_n_165 ,n_115 ,csa_tree_add_118_30_groupi_n_159);
  and csa_tree_add_118_30_groupi_g689(csa_tree_add_118_30_groupi_n_164 ,csa_tree_add_118_30_groupi_n_157 ,csa_tree_add_118_30_groupi_n_161);
  xor csa_tree_add_118_30_groupi_g690(out2[2] ,csa_tree_add_118_30_groupi_n_133 ,csa_tree_add_118_30_groupi_n_154);
  or csa_tree_add_118_30_groupi_g691(csa_tree_add_118_30_groupi_n_162 ,csa_tree_add_118_30_groupi_n_65 ,csa_tree_add_118_30_groupi_n_155);
  or csa_tree_add_118_30_groupi_g692(csa_tree_add_118_30_groupi_n_161 ,csa_tree_add_118_30_groupi_n_142 ,csa_tree_add_118_30_groupi_n_158);
  xnor csa_tree_add_118_30_groupi_g693(csa_tree_add_118_30_groupi_n_160 ,csa_tree_add_118_30_groupi_n_132 ,n_114);
  xnor csa_tree_add_118_30_groupi_g694(csa_tree_add_118_30_groupi_n_159 ,csa_tree_add_118_30_groupi_n_143 ,csa_tree_add_118_30_groupi_n_2);
  and csa_tree_add_118_30_groupi_g695(csa_tree_add_118_30_groupi_n_158 ,csa_tree_add_118_30_groupi_n_141 ,csa_tree_add_118_30_groupi_n_133);
  or csa_tree_add_118_30_groupi_g696(csa_tree_add_118_30_groupi_n_157 ,n_114 ,csa_tree_add_118_30_groupi_n_132);
  and csa_tree_add_118_30_groupi_g697(csa_tree_add_118_30_groupi_n_156 ,n_114 ,csa_tree_add_118_30_groupi_n_132);
  and csa_tree_add_118_30_groupi_g698(csa_tree_add_118_30_groupi_n_155 ,csa_tree_add_118_30_groupi_n_56 ,csa_tree_add_118_30_groupi_n_143);
  xnor csa_tree_add_118_30_groupi_g699(csa_tree_add_118_30_groupi_n_154 ,csa_tree_add_118_30_groupi_n_111 ,n_113);
  xnor csa_tree_add_118_30_groupi_g700(csa_tree_add_118_30_groupi_n_153 ,csa_tree_add_118_30_groupi_n_96 ,csa_tree_add_118_30_groupi_n_113);
  xnor csa_tree_add_118_30_groupi_g701(csa_tree_add_118_30_groupi_n_152 ,csa_tree_add_118_30_groupi_n_103 ,csa_tree_add_118_30_groupi_n_109);
  xor csa_tree_add_118_30_groupi_g702(out2[1] ,csa_tree_add_118_30_groupi_n_99 ,csa_tree_add_118_30_groupi_n_116);
  xnor csa_tree_add_118_30_groupi_g703(csa_tree_add_118_30_groupi_n_150 ,csa_tree_add_118_30_groupi_n_105 ,csa_tree_add_118_30_groupi_n_114);
  xnor csa_tree_add_118_30_groupi_g704(csa_tree_add_118_30_groupi_n_149 ,csa_tree_add_118_30_groupi_n_106 ,csa_tree_add_118_30_groupi_n_115);
  xnor csa_tree_add_118_30_groupi_g705(csa_tree_add_118_30_groupi_n_148 ,csa_tree_add_118_30_groupi_n_98 ,csa_tree_add_118_30_groupi_n_112);
  xnor csa_tree_add_118_30_groupi_g706(csa_tree_add_118_30_groupi_n_147 ,csa_tree_add_118_30_groupi_n_97 ,csa_tree_add_118_30_groupi_n_121);
  xnor csa_tree_add_118_30_groupi_g707(csa_tree_add_118_30_groupi_n_146 ,csa_tree_add_118_30_groupi_n_104 ,csa_tree_add_118_30_groupi_n_120);
  xnor csa_tree_add_118_30_groupi_g708(csa_tree_add_118_30_groupi_n_145 ,csa_tree_add_118_30_groupi_n_95 ,csa_tree_add_118_30_groupi_n_119);
  xnor csa_tree_add_118_30_groupi_g709(csa_tree_add_118_30_groupi_n_144 ,csa_tree_add_118_30_groupi_n_94 ,csa_tree_add_118_30_groupi_n_107);
  nor csa_tree_add_118_30_groupi_g710(csa_tree_add_118_30_groupi_n_142 ,csa_tree_add_118_30_groupi_n_36 ,csa_tree_add_118_30_groupi_n_111);
  or csa_tree_add_118_30_groupi_g711(csa_tree_add_118_30_groupi_n_141 ,n_113 ,csa_tree_add_118_30_groupi_n_110);
  or csa_tree_add_118_30_groupi_g712(csa_tree_add_118_30_groupi_n_140 ,csa_tree_add_118_30_groupi_n_95 ,csa_tree_add_118_30_groupi_n_119);
  and csa_tree_add_118_30_groupi_g713(csa_tree_add_118_30_groupi_n_139 ,csa_tree_add_118_30_groupi_n_104 ,csa_tree_add_118_30_groupi_n_120);
  or csa_tree_add_118_30_groupi_g714(csa_tree_add_118_30_groupi_n_138 ,csa_tree_add_118_30_groupi_n_97 ,csa_tree_add_118_30_groupi_n_121);
  and csa_tree_add_118_30_groupi_g715(csa_tree_add_118_30_groupi_n_137 ,csa_tree_add_118_30_groupi_n_105 ,csa_tree_add_118_30_groupi_n_114);
  and csa_tree_add_118_30_groupi_g716(csa_tree_add_118_30_groupi_n_136 ,csa_tree_add_118_30_groupi_n_103 ,csa_tree_add_118_30_groupi_n_109);
  or csa_tree_add_118_30_groupi_g717(csa_tree_add_118_30_groupi_n_135 ,csa_tree_add_118_30_groupi_n_105 ,csa_tree_add_118_30_groupi_n_114);
  and csa_tree_add_118_30_groupi_g718(csa_tree_add_118_30_groupi_n_134 ,csa_tree_add_118_30_groupi_n_106 ,csa_tree_add_118_30_groupi_n_115);
  or csa_tree_add_118_30_groupi_g719(csa_tree_add_118_30_groupi_n_143 ,csa_tree_add_118_30_groupi_n_55 ,csa_tree_add_118_30_groupi_n_117);
  and csa_tree_add_118_30_groupi_g720(csa_tree_add_118_30_groupi_n_131 ,csa_tree_add_118_30_groupi_n_97 ,csa_tree_add_118_30_groupi_n_121);
  or csa_tree_add_118_30_groupi_g721(csa_tree_add_118_30_groupi_n_130 ,csa_tree_add_118_30_groupi_n_96 ,csa_tree_add_118_30_groupi_n_113);
  or csa_tree_add_118_30_groupi_g722(csa_tree_add_118_30_groupi_n_129 ,csa_tree_add_118_30_groupi_n_106 ,csa_tree_add_118_30_groupi_n_115);
  or csa_tree_add_118_30_groupi_g723(csa_tree_add_118_30_groupi_n_128 ,csa_tree_add_118_30_groupi_n_103 ,csa_tree_add_118_30_groupi_n_109);
  and csa_tree_add_118_30_groupi_g724(csa_tree_add_118_30_groupi_n_127 ,csa_tree_add_118_30_groupi_n_98 ,csa_tree_add_118_30_groupi_n_112);
  and csa_tree_add_118_30_groupi_g725(csa_tree_add_118_30_groupi_n_126 ,csa_tree_add_118_30_groupi_n_96 ,csa_tree_add_118_30_groupi_n_113);
  or csa_tree_add_118_30_groupi_g726(csa_tree_add_118_30_groupi_n_125 ,csa_tree_add_118_30_groupi_n_104 ,csa_tree_add_118_30_groupi_n_120);
  and csa_tree_add_118_30_groupi_g727(csa_tree_add_118_30_groupi_n_124 ,csa_tree_add_118_30_groupi_n_95 ,csa_tree_add_118_30_groupi_n_119);
  or csa_tree_add_118_30_groupi_g728(csa_tree_add_118_30_groupi_n_123 ,csa_tree_add_118_30_groupi_n_98 ,csa_tree_add_118_30_groupi_n_112);
  or csa_tree_add_118_30_groupi_g729(csa_tree_add_118_30_groupi_n_133 ,csa_tree_add_118_30_groupi_n_102 ,csa_tree_add_118_30_groupi_n_118);
  xnor csa_tree_add_118_30_groupi_g730(csa_tree_add_118_30_groupi_n_132 ,csa_tree_add_118_30_groupi_n_100 ,csa_tree_add_118_30_groupi_n_1);
  and csa_tree_add_118_30_groupi_g731(csa_tree_add_118_30_groupi_n_118 ,csa_tree_add_118_30_groupi_n_99 ,csa_tree_add_118_30_groupi_n_101);
  and csa_tree_add_118_30_groupi_g732(csa_tree_add_118_30_groupi_n_117 ,csa_tree_add_118_30_groupi_n_64 ,csa_tree_add_118_30_groupi_n_100);
  xnor csa_tree_add_118_30_groupi_g733(csa_tree_add_118_30_groupi_n_116 ,csa_tree_add_118_30_groupi_n_80 ,n_112);
  xnor csa_tree_add_118_30_groupi_g734(csa_tree_add_118_30_groupi_n_122 ,csa_tree_add_118_30_groupi_n_74 ,n_117);
  xnor csa_tree_add_118_30_groupi_g735(csa_tree_add_118_30_groupi_n_121 ,csa_tree_add_118_30_groupi_n_73 ,n_123);
  xnor csa_tree_add_118_30_groupi_g736(csa_tree_add_118_30_groupi_n_120 ,csa_tree_add_118_30_groupi_n_78 ,n_118);
  xnor csa_tree_add_118_30_groupi_g737(csa_tree_add_118_30_groupi_n_119 ,csa_tree_add_118_30_groupi_n_77 ,n_119);
  not csa_tree_add_118_30_groupi_g738(csa_tree_add_118_30_groupi_n_110 ,csa_tree_add_118_30_groupi_n_111);
  xnor csa_tree_add_118_30_groupi_g739(out2[0] ,csa_tree_add_118_30_groupi_n_82 ,out1[0]);
  xnor csa_tree_add_118_30_groupi_g740(csa_tree_add_118_30_groupi_n_107 ,csa_tree_add_118_30_groupi_n_69 ,n_126);
  xnor csa_tree_add_118_30_groupi_g741(csa_tree_add_118_30_groupi_n_115 ,csa_tree_add_118_30_groupi_n_71 ,n_121);
  xnor csa_tree_add_118_30_groupi_g742(csa_tree_add_118_30_groupi_n_114 ,csa_tree_add_118_30_groupi_n_75 ,n_122);
  xnor csa_tree_add_118_30_groupi_g743(csa_tree_add_118_30_groupi_n_113 ,csa_tree_add_118_30_groupi_n_76 ,n_125);
  xnor csa_tree_add_118_30_groupi_g744(csa_tree_add_118_30_groupi_n_112 ,csa_tree_add_118_30_groupi_n_70 ,n_120);
  xnor csa_tree_add_118_30_groupi_g745(csa_tree_add_118_30_groupi_n_111 ,csa_tree_add_118_30_groupi_n_68 ,csa_tree_add_118_30_groupi_n_81);
  xnor csa_tree_add_118_30_groupi_g746(csa_tree_add_118_30_groupi_n_109 ,csa_tree_add_118_30_groupi_n_72 ,n_124);
  nor csa_tree_add_118_30_groupi_g747(csa_tree_add_118_30_groupi_n_102 ,csa_tree_add_118_30_groupi_n_38 ,csa_tree_add_118_30_groupi_n_80);
  or csa_tree_add_118_30_groupi_g748(csa_tree_add_118_30_groupi_n_101 ,n_112 ,csa_tree_add_118_30_groupi_n_79);
  or csa_tree_add_118_30_groupi_g749(csa_tree_add_118_30_groupi_n_106 ,csa_tree_add_118_30_groupi_n_61 ,csa_tree_add_118_30_groupi_n_88);
  or csa_tree_add_118_30_groupi_g750(csa_tree_add_118_30_groupi_n_105 ,csa_tree_add_118_30_groupi_n_54 ,csa_tree_add_118_30_groupi_n_90);
  or csa_tree_add_118_30_groupi_g751(csa_tree_add_118_30_groupi_n_104 ,csa_tree_add_118_30_groupi_n_62 ,csa_tree_add_118_30_groupi_n_86);
  or csa_tree_add_118_30_groupi_g752(csa_tree_add_118_30_groupi_n_103 ,csa_tree_add_118_30_groupi_n_57 ,csa_tree_add_118_30_groupi_n_89);
  or csa_tree_add_118_30_groupi_g753(csa_tree_add_118_30_groupi_n_94 ,csa_tree_add_118_30_groupi_n_59 ,csa_tree_add_118_30_groupi_n_91);
  or csa_tree_add_118_30_groupi_g754(csa_tree_add_118_30_groupi_n_100 ,csa_tree_add_118_30_groupi_n_53 ,csa_tree_add_118_30_groupi_n_83);
  or csa_tree_add_118_30_groupi_g755(csa_tree_add_118_30_groupi_n_99 ,csa_tree_add_118_30_groupi_n_51 ,csa_tree_add_118_30_groupi_n_84);
  or csa_tree_add_118_30_groupi_g756(csa_tree_add_118_30_groupi_n_98 ,csa_tree_add_118_30_groupi_n_46 ,csa_tree_add_118_30_groupi_n_87);
  or csa_tree_add_118_30_groupi_g757(csa_tree_add_118_30_groupi_n_97 ,csa_tree_add_118_30_groupi_n_49 ,csa_tree_add_118_30_groupi_n_85);
  or csa_tree_add_118_30_groupi_g758(csa_tree_add_118_30_groupi_n_96 ,csa_tree_add_118_30_groupi_n_41 ,csa_tree_add_118_30_groupi_n_92);
  or csa_tree_add_118_30_groupi_g759(csa_tree_add_118_30_groupi_n_95 ,csa_tree_add_118_30_groupi_n_47 ,csa_tree_add_118_30_groupi_n_93);
  and csa_tree_add_118_30_groupi_g760(csa_tree_add_118_30_groupi_n_93 ,n_118 ,csa_tree_add_118_30_groupi_n_48);
  and csa_tree_add_118_30_groupi_g761(csa_tree_add_118_30_groupi_n_92 ,n_300 ,csa_tree_add_118_30_groupi_n_40);
  and csa_tree_add_118_30_groupi_g762(csa_tree_add_118_30_groupi_n_91 ,n_301 ,csa_tree_add_118_30_groupi_n_67);
  and csa_tree_add_118_30_groupi_g763(csa_tree_add_118_30_groupi_n_90 ,out1[10] ,csa_tree_add_118_30_groupi_n_60);
  and csa_tree_add_118_30_groupi_g764(csa_tree_add_118_30_groupi_n_89 ,n_299 ,csa_tree_add_118_30_groupi_n_50);
  and csa_tree_add_118_30_groupi_g765(csa_tree_add_118_30_groupi_n_88 ,n_296 ,csa_tree_add_118_30_groupi_n_45);
  and csa_tree_add_118_30_groupi_g766(csa_tree_add_118_30_groupi_n_87 ,n_295 ,csa_tree_add_118_30_groupi_n_66);
  and csa_tree_add_118_30_groupi_g767(csa_tree_add_118_30_groupi_n_86 ,n_117 ,csa_tree_add_118_30_groupi_n_52);
  and csa_tree_add_118_30_groupi_g768(csa_tree_add_118_30_groupi_n_85 ,n_298 ,csa_tree_add_118_30_groupi_n_58);
  and csa_tree_add_118_30_groupi_g769(csa_tree_add_118_30_groupi_n_84 ,out1[0] ,csa_tree_add_118_30_groupi_n_44);
  nor csa_tree_add_118_30_groupi_g770(csa_tree_add_118_30_groupi_n_83 ,csa_tree_add_118_30_groupi_n_68 ,csa_tree_add_118_30_groupi_n_42);
  xnor csa_tree_add_118_30_groupi_g771(csa_tree_add_118_30_groupi_n_82 ,n_287 ,n_111);
  xnor csa_tree_add_118_30_groupi_g772(csa_tree_add_118_30_groupi_n_81 ,n_289 ,csa_tree_add_118_30_groupi_n_35);
  not csa_tree_add_118_30_groupi_g773(csa_tree_add_118_30_groupi_n_79 ,csa_tree_add_118_30_groupi_n_80);
  xnor csa_tree_add_118_30_groupi_g774(csa_tree_add_118_30_groupi_n_78 ,csa_tree_add_118_30_groupi_n_17 ,n_294);
  xnor csa_tree_add_118_30_groupi_g775(csa_tree_add_118_30_groupi_n_77 ,csa_tree_add_118_30_groupi_n_26 ,n_295);
  xnor csa_tree_add_118_30_groupi_g776(csa_tree_add_118_30_groupi_n_76 ,csa_tree_add_118_30_groupi_n_5 ,n_301);
  xnor csa_tree_add_118_30_groupi_g777(csa_tree_add_118_30_groupi_n_75 ,csa_tree_add_118_30_groupi_n_23 ,n_298);
  xnor csa_tree_add_118_30_groupi_g778(csa_tree_add_118_30_groupi_n_74 ,csa_tree_add_118_30_groupi_n_8 ,n_293);
  xnor csa_tree_add_118_30_groupi_g780(csa_tree_add_118_30_groupi_n_73 ,csa_tree_add_118_30_groupi_n_14 ,n_299);
  xnor csa_tree_add_118_30_groupi_g782(csa_tree_add_118_30_groupi_n_72 ,csa_tree_add_118_30_groupi_n_20 ,n_300);
  xnor csa_tree_add_118_30_groupi_g783(csa_tree_add_118_30_groupi_n_71 ,n_297 ,out1[10]);
  xnor csa_tree_add_118_30_groupi_g785(csa_tree_add_118_30_groupi_n_70 ,csa_tree_add_118_30_groupi_n_11 ,n_296);
  xnor csa_tree_add_118_30_groupi_g786(csa_tree_add_118_30_groupi_n_69 ,n_302 ,out1[15]);
  xnor csa_tree_add_118_30_groupi_g787(csa_tree_add_118_30_groupi_n_80 ,n_288 ,out1[1]);
  or csa_tree_add_118_30_groupi_g788(csa_tree_add_118_30_groupi_n_67 ,csa_tree_add_118_30_groupi_n_4 ,n_125);
  or csa_tree_add_118_30_groupi_g789(csa_tree_add_118_30_groupi_n_66 ,csa_tree_add_118_30_groupi_n_25 ,n_119);
  and csa_tree_add_118_30_groupi_g790(csa_tree_add_118_30_groupi_n_65 ,n_291 ,csa_tree_add_118_30_groupi_n_32);
  or csa_tree_add_118_30_groupi_g791(csa_tree_add_118_30_groupi_n_64 ,n_290 ,csa_tree_add_118_30_groupi_n_30);
  or csa_tree_add_118_30_groupi_g792(csa_tree_add_118_30_groupi_n_63 ,n_292 ,csa_tree_add_118_30_groupi_n_28);
  and csa_tree_add_118_30_groupi_g793(csa_tree_add_118_30_groupi_n_62 ,n_293 ,csa_tree_add_118_30_groupi_n_7);
  and csa_tree_add_118_30_groupi_g794(csa_tree_add_118_30_groupi_n_61 ,csa_tree_add_118_30_groupi_n_10 ,n_120);
  or csa_tree_add_118_30_groupi_g795(csa_tree_add_118_30_groupi_n_60 ,n_297 ,n_121);
  and csa_tree_add_118_30_groupi_g796(csa_tree_add_118_30_groupi_n_59 ,csa_tree_add_118_30_groupi_n_5 ,n_125);
  or csa_tree_add_118_30_groupi_g797(csa_tree_add_118_30_groupi_n_58 ,csa_tree_add_118_30_groupi_n_22 ,n_122);
  and csa_tree_add_118_30_groupi_g798(csa_tree_add_118_30_groupi_n_57 ,csa_tree_add_118_30_groupi_n_13 ,n_123);
  or csa_tree_add_118_30_groupi_g799(csa_tree_add_118_30_groupi_n_56 ,n_291 ,csa_tree_add_118_30_groupi_n_32);
  and csa_tree_add_118_30_groupi_g800(csa_tree_add_118_30_groupi_n_55 ,n_290 ,csa_tree_add_118_30_groupi_n_30);
  or csa_tree_add_118_30_groupi_g801(csa_tree_add_118_30_groupi_n_68 ,csa_tree_add_118_30_groupi_n_37 ,csa_tree_add_118_30_groupi_n_39);
  and csa_tree_add_118_30_groupi_g802(csa_tree_add_118_30_groupi_n_54 ,n_297 ,n_121);
  and csa_tree_add_118_30_groupi_g803(csa_tree_add_118_30_groupi_n_53 ,n_289 ,csa_tree_add_118_30_groupi_n_35);
  or csa_tree_add_118_30_groupi_g804(csa_tree_add_118_30_groupi_n_52 ,n_293 ,csa_tree_add_118_30_groupi_n_8);
  and csa_tree_add_118_30_groupi_g805(csa_tree_add_118_30_groupi_n_51 ,n_287 ,n_111);
  or csa_tree_add_118_30_groupi_g806(csa_tree_add_118_30_groupi_n_50 ,csa_tree_add_118_30_groupi_n_14 ,n_123);
  and csa_tree_add_118_30_groupi_g807(csa_tree_add_118_30_groupi_n_49 ,csa_tree_add_118_30_groupi_n_23 ,n_122);
  or csa_tree_add_118_30_groupi_g808(csa_tree_add_118_30_groupi_n_48 ,n_294 ,csa_tree_add_118_30_groupi_n_16);
  and csa_tree_add_118_30_groupi_g809(csa_tree_add_118_30_groupi_n_47 ,n_294 ,csa_tree_add_118_30_groupi_n_17);
  and csa_tree_add_118_30_groupi_g810(csa_tree_add_118_30_groupi_n_46 ,csa_tree_add_118_30_groupi_n_26 ,n_119);
  or csa_tree_add_118_30_groupi_g811(csa_tree_add_118_30_groupi_n_45 ,csa_tree_add_118_30_groupi_n_11 ,n_120);
  or csa_tree_add_118_30_groupi_g812(csa_tree_add_118_30_groupi_n_44 ,n_287 ,n_111);
  and csa_tree_add_118_30_groupi_g813(csa_tree_add_118_30_groupi_n_43 ,n_292 ,csa_tree_add_118_30_groupi_n_28);
  nor csa_tree_add_118_30_groupi_g814(csa_tree_add_118_30_groupi_n_42 ,n_289 ,csa_tree_add_118_30_groupi_n_34);
  and csa_tree_add_118_30_groupi_g815(csa_tree_add_118_30_groupi_n_41 ,csa_tree_add_118_30_groupi_n_19 ,n_124);
  or csa_tree_add_118_30_groupi_g816(csa_tree_add_118_30_groupi_n_40 ,csa_tree_add_118_30_groupi_n_20 ,n_124);
  not csa_tree_add_118_30_groupi_g817(csa_tree_add_118_30_groupi_n_39 ,out1[1]);
  not csa_tree_add_118_30_groupi_g818(csa_tree_add_118_30_groupi_n_38 ,n_112);
  not csa_tree_add_118_30_groupi_g819(csa_tree_add_118_30_groupi_n_37 ,n_288);
  not csa_tree_add_118_30_groupi_g820(csa_tree_add_118_30_groupi_n_36 ,n_113);
  not csa_tree_add_118_30_groupi_drc_bufs(csa_tree_add_118_30_groupi_n_35 ,csa_tree_add_118_30_groupi_n_33);
  not csa_tree_add_118_30_groupi_drc_bufs821(csa_tree_add_118_30_groupi_n_34 ,csa_tree_add_118_30_groupi_n_33);
  not csa_tree_add_118_30_groupi_drc_bufs822(csa_tree_add_118_30_groupi_n_33 ,out1[2]);
  not csa_tree_add_118_30_groupi_drc_bufs825(csa_tree_add_118_30_groupi_n_32 ,csa_tree_add_118_30_groupi_n_31);
  not csa_tree_add_118_30_groupi_drc_bufs826(csa_tree_add_118_30_groupi_n_31 ,out1[4]);
  not csa_tree_add_118_30_groupi_drc_bufs829(csa_tree_add_118_30_groupi_n_30 ,csa_tree_add_118_30_groupi_n_29);
  not csa_tree_add_118_30_groupi_drc_bufs830(csa_tree_add_118_30_groupi_n_29 ,out1[3]);
  not csa_tree_add_118_30_groupi_drc_bufs833(csa_tree_add_118_30_groupi_n_28 ,csa_tree_add_118_30_groupi_n_27);
  not csa_tree_add_118_30_groupi_drc_bufs834(csa_tree_add_118_30_groupi_n_27 ,out1[5]);
  not csa_tree_add_118_30_groupi_drc_bufs836(csa_tree_add_118_30_groupi_n_26 ,csa_tree_add_118_30_groupi_n_24);
  not csa_tree_add_118_30_groupi_drc_bufs837(csa_tree_add_118_30_groupi_n_25 ,csa_tree_add_118_30_groupi_n_24);
  not csa_tree_add_118_30_groupi_drc_bufs838(csa_tree_add_118_30_groupi_n_24 ,out1[8]);
  not csa_tree_add_118_30_groupi_drc_bufs840(csa_tree_add_118_30_groupi_n_23 ,csa_tree_add_118_30_groupi_n_21);
  not csa_tree_add_118_30_groupi_drc_bufs841(csa_tree_add_118_30_groupi_n_22 ,csa_tree_add_118_30_groupi_n_21);
  not csa_tree_add_118_30_groupi_drc_bufs842(csa_tree_add_118_30_groupi_n_21 ,out1[11]);
  not csa_tree_add_118_30_groupi_drc_bufs844(csa_tree_add_118_30_groupi_n_20 ,csa_tree_add_118_30_groupi_n_18);
  not csa_tree_add_118_30_groupi_drc_bufs845(csa_tree_add_118_30_groupi_n_19 ,csa_tree_add_118_30_groupi_n_18);
  not csa_tree_add_118_30_groupi_drc_bufs846(csa_tree_add_118_30_groupi_n_18 ,out1[13]);
  not csa_tree_add_118_30_groupi_drc_bufs848(csa_tree_add_118_30_groupi_n_17 ,csa_tree_add_118_30_groupi_n_15);
  not csa_tree_add_118_30_groupi_drc_bufs849(csa_tree_add_118_30_groupi_n_16 ,csa_tree_add_118_30_groupi_n_15);
  not csa_tree_add_118_30_groupi_drc_bufs850(csa_tree_add_118_30_groupi_n_15 ,out1[7]);
  not csa_tree_add_118_30_groupi_drc_bufs852(csa_tree_add_118_30_groupi_n_14 ,csa_tree_add_118_30_groupi_n_12);
  not csa_tree_add_118_30_groupi_drc_bufs853(csa_tree_add_118_30_groupi_n_13 ,csa_tree_add_118_30_groupi_n_12);
  not csa_tree_add_118_30_groupi_drc_bufs854(csa_tree_add_118_30_groupi_n_12 ,out1[12]);
  not csa_tree_add_118_30_groupi_drc_bufs856(csa_tree_add_118_30_groupi_n_11 ,csa_tree_add_118_30_groupi_n_9);
  not csa_tree_add_118_30_groupi_drc_bufs857(csa_tree_add_118_30_groupi_n_10 ,csa_tree_add_118_30_groupi_n_9);
  not csa_tree_add_118_30_groupi_drc_bufs858(csa_tree_add_118_30_groupi_n_9 ,out1[9]);
  not csa_tree_add_118_30_groupi_drc_bufs860(csa_tree_add_118_30_groupi_n_8 ,csa_tree_add_118_30_groupi_n_6);
  not csa_tree_add_118_30_groupi_drc_bufs861(csa_tree_add_118_30_groupi_n_7 ,csa_tree_add_118_30_groupi_n_6);
  not csa_tree_add_118_30_groupi_drc_bufs862(csa_tree_add_118_30_groupi_n_6 ,out1[6]);
  not csa_tree_add_118_30_groupi_drc_bufs864(csa_tree_add_118_30_groupi_n_5 ,csa_tree_add_118_30_groupi_n_3);
  not csa_tree_add_118_30_groupi_drc_bufs865(csa_tree_add_118_30_groupi_n_4 ,csa_tree_add_118_30_groupi_n_3);
  not csa_tree_add_118_30_groupi_drc_bufs866(csa_tree_add_118_30_groupi_n_3 ,out1[14]);
  xor csa_tree_add_118_30_groupi_g2(csa_tree_add_118_30_groupi_n_2 ,n_291 ,csa_tree_add_118_30_groupi_n_31);
  xor csa_tree_add_118_30_groupi_g868(csa_tree_add_118_30_groupi_n_1 ,n_290 ,csa_tree_add_118_30_groupi_n_29);
  xor csa_tree_add_118_30_groupi_g869(csa_tree_add_118_30_groupi_n_0 ,n_292 ,csa_tree_add_118_30_groupi_n_27);
  xnor csa_tree_sub_77_21_g192(csa_tree_sub_77_21_n_32 ,in1[6] ,in2[6]);
  xnor csa_tree_sub_77_21_g193(csa_tree_sub_77_21_n_31 ,in1[1] ,in2[1]);
  xnor csa_tree_sub_77_21_g194(csa_tree_sub_77_21_n_30 ,in1[5] ,in2[5]);
  xnor csa_tree_sub_77_21_g195(csa_tree_sub_77_21_n_29 ,in1[4] ,in2[4]);
  xnor csa_tree_sub_77_21_g196(csa_tree_sub_77_21_n_28 ,in1[3] ,in2[3]);
  xnor csa_tree_sub_77_21_g197(csa_tree_sub_77_21_n_27 ,in1[2] ,in2[2]);
  and csa_tree_sub_77_21_g198(csa_tree_sub_77_21_n_26 ,in1[5] ,csa_tree_sub_77_21_n_17);
  and csa_tree_sub_77_21_g199(csa_tree_sub_77_21_n_25 ,in1[3] ,csa_tree_sub_77_21_n_20);
  and csa_tree_sub_77_21_g200(csa_tree_sub_77_21_n_24 ,in2[6] ,csa_tree_sub_77_21_n_19);
  and csa_tree_sub_77_21_g201(n_457 ,in1[4] ,csa_tree_sub_77_21_n_15);
  and csa_tree_sub_77_21_g202(n_459 ,in1[2] ,csa_tree_sub_77_21_n_13);
  and csa_tree_sub_77_21_g203(csa_tree_sub_77_21_n_21 ,in1[1] ,csa_tree_sub_77_21_n_18);
  not csa_tree_sub_77_21_g204(csa_tree_sub_77_21_n_20 ,in2[3]);
  not csa_tree_sub_77_21_g205(csa_tree_sub_77_21_n_19 ,in1[6]);
  not csa_tree_sub_77_21_g206(csa_tree_sub_77_21_n_18 ,in2[1]);
  not csa_tree_sub_77_21_g207(csa_tree_sub_77_21_n_17 ,in2[5]);
  not csa_tree_sub_77_21_g208(n_462 ,in2[0]);
  not csa_tree_sub_77_21_g209(csa_tree_sub_77_21_n_15 ,in2[4]);
  not csa_tree_sub_77_21_g210(csa_tree_sub_77_21_n_14 ,in1[0]);
  not csa_tree_sub_77_21_g211(csa_tree_sub_77_21_n_13 ,in2[2]);
  buf csa_tree_sub_77_21_drc_bufs(n_466 ,csa_tree_sub_77_21_n_30);
  buf csa_tree_sub_77_21_drc_bufs212(n_468 ,csa_tree_sub_77_21_n_28);
  buf csa_tree_sub_77_21_drc_bufs213(n_470 ,csa_tree_sub_77_21_n_31);
  buf csa_tree_sub_77_21_drc_bufs214(n_458 ,csa_tree_sub_77_21_n_25);
  buf csa_tree_sub_77_21_drc_bufs215(n_460 ,csa_tree_sub_77_21_n_21);
  buf csa_tree_sub_77_21_drc_bufs216(n_456 ,csa_tree_sub_77_21_n_26);
  buf csa_tree_sub_77_21_drc_bufs217(n_469 ,csa_tree_sub_77_21_n_27);
  buf csa_tree_sub_77_21_drc_bufs218(n_467 ,csa_tree_sub_77_21_n_29);
  buf csa_tree_sub_77_21_drc_bufs219(n_465 ,csa_tree_sub_77_21_n_32);
  buf csa_tree_sub_77_21_drc_bufs220(n_464 ,csa_tree_sub_77_21_n_24);
  buf csa_tree_sub_77_21_drc_bufs221(n_471 ,csa_tree_sub_77_21_n_14);
  xnor csa_tree_sub_80_22_g130(n_679 ,in10[4] ,in11[4]);
  xnor csa_tree_sub_80_22_g131(n_680 ,in10[3] ,in11[3]);
  xnor csa_tree_sub_80_22_g132(n_681 ,in10[2] ,in11[2]);
  xnor csa_tree_sub_80_22_g133(n_682 ,in10[1] ,in11[1]);
  and csa_tree_sub_80_22_g134(n_672 ,in10[3] ,csa_tree_sub_80_22_n_6);
  and csa_tree_sub_80_22_g135(n_674 ,in10[1] ,csa_tree_sub_80_22_n_4);
  and csa_tree_sub_80_22_g136(n_673 ,in10[2] ,csa_tree_sub_80_22_n_3);
  and csa_tree_sub_80_22_g137(n_678 ,in11[4] ,csa_tree_sub_80_22_n_2);
  not csa_tree_sub_80_22_g138(n_676 ,in11[0]);
  not csa_tree_sub_80_22_g139(csa_tree_sub_80_22_n_6 ,in11[3]);
  not csa_tree_sub_80_22_g140(n_683 ,in10[0]);
  not csa_tree_sub_80_22_g141(csa_tree_sub_80_22_n_4 ,in11[1]);
  not csa_tree_sub_80_22_g142(csa_tree_sub_80_22_n_3 ,in11[2]);
  not csa_tree_sub_80_22_g143(csa_tree_sub_80_22_n_2 ,in10[4]);
  xnor csa_tree_sub_86_22_g130(n_725 ,in14[4] ,in15[4]);
  xnor csa_tree_sub_86_22_g131(n_726 ,in14[3] ,in15[3]);
  xnor csa_tree_sub_86_22_g132(n_727 ,in14[2] ,in15[2]);
  xnor csa_tree_sub_86_22_g133(n_728 ,in14[1] ,in15[1]);
  and csa_tree_sub_86_22_g134(n_718 ,in14[3] ,csa_tree_sub_86_22_n_6);
  and csa_tree_sub_86_22_g135(n_720 ,in14[1] ,csa_tree_sub_86_22_n_4);
  and csa_tree_sub_86_22_g136(n_719 ,in14[2] ,csa_tree_sub_86_22_n_3);
  and csa_tree_sub_86_22_g137(n_724 ,in15[4] ,csa_tree_sub_86_22_n_2);
  not csa_tree_sub_86_22_g138(n_722 ,in15[0]);
  not csa_tree_sub_86_22_g139(csa_tree_sub_86_22_n_6 ,in15[3]);
  not csa_tree_sub_86_22_g140(n_729 ,in14[0]);
  not csa_tree_sub_86_22_g141(csa_tree_sub_86_22_n_4 ,in15[1]);
  not csa_tree_sub_86_22_g142(csa_tree_sub_86_22_n_3 ,in15[2]);
  not csa_tree_sub_86_22_g143(csa_tree_sub_86_22_n_2 ,in14[4]);
  xnor csa_tree_sub_92_22_g130(n_557 ,in18[4] ,in19[4]);
  xnor csa_tree_sub_92_22_g131(n_558 ,in18[3] ,in19[3]);
  xnor csa_tree_sub_92_22_g132(n_559 ,in18[2] ,in19[2]);
  xnor csa_tree_sub_92_22_g133(n_560 ,in18[1] ,in19[1]);
  and csa_tree_sub_92_22_g134(n_550 ,in18[3] ,csa_tree_sub_92_22_n_6);
  and csa_tree_sub_92_22_g135(n_552 ,in18[1] ,csa_tree_sub_92_22_n_4);
  and csa_tree_sub_92_22_g136(n_551 ,in18[2] ,csa_tree_sub_92_22_n_3);
  and csa_tree_sub_92_22_g137(n_556 ,in19[4] ,csa_tree_sub_92_22_n_2);
  not csa_tree_sub_92_22_g138(n_554 ,in19[0]);
  not csa_tree_sub_92_22_g139(csa_tree_sub_92_22_n_6 ,in19[3]);
  not csa_tree_sub_92_22_g140(n_561 ,in18[0]);
  not csa_tree_sub_92_22_g141(csa_tree_sub_92_22_n_4 ,in19[1]);
  not csa_tree_sub_92_22_g142(csa_tree_sub_92_22_n_3 ,in19[2]);
  not csa_tree_sub_92_22_g143(csa_tree_sub_92_22_n_2 ,in18[4]);
  xnor csa_tree_sub_98_22_g130(n_633 ,in22[4] ,in23[4]);
  xnor csa_tree_sub_98_22_g131(n_634 ,in22[3] ,in23[3]);
  xnor csa_tree_sub_98_22_g132(n_635 ,in22[2] ,in23[2]);
  xnor csa_tree_sub_98_22_g133(n_636 ,in22[1] ,in23[1]);
  and csa_tree_sub_98_22_g134(n_626 ,in22[3] ,csa_tree_sub_98_22_n_6);
  and csa_tree_sub_98_22_g135(n_628 ,in22[1] ,csa_tree_sub_98_22_n_4);
  and csa_tree_sub_98_22_g136(n_627 ,in22[2] ,csa_tree_sub_98_22_n_3);
  and csa_tree_sub_98_22_g137(n_632 ,in23[4] ,csa_tree_sub_98_22_n_2);
  not csa_tree_sub_98_22_g138(n_630 ,in23[0]);
  not csa_tree_sub_98_22_g139(csa_tree_sub_98_22_n_6 ,in23[3]);
  not csa_tree_sub_98_22_g140(n_637 ,in22[0]);
  not csa_tree_sub_98_22_g141(csa_tree_sub_98_22_n_4 ,in23[1]);
  not csa_tree_sub_98_22_g142(csa_tree_sub_98_22_n_3 ,in23[2]);
  not csa_tree_sub_98_22_g143(csa_tree_sub_98_22_n_2 ,in22[4]);
  xnor csa_tree_sub_104_22_g130(n_587 ,in26[4] ,in27[4]);
  xnor csa_tree_sub_104_22_g131(n_588 ,in26[3] ,in27[3]);
  xnor csa_tree_sub_104_22_g132(n_589 ,in26[2] ,in27[2]);
  xnor csa_tree_sub_104_22_g133(n_590 ,in26[1] ,in27[1]);
  and csa_tree_sub_104_22_g134(n_580 ,in26[3] ,csa_tree_sub_104_22_n_6);
  and csa_tree_sub_104_22_g135(n_582 ,in26[1] ,csa_tree_sub_104_22_n_4);
  and csa_tree_sub_104_22_g136(n_581 ,in26[2] ,csa_tree_sub_104_22_n_3);
  and csa_tree_sub_104_22_g137(n_586 ,in27[4] ,csa_tree_sub_104_22_n_2);
  not csa_tree_sub_104_22_g138(n_584 ,in27[0]);
  not csa_tree_sub_104_22_g139(csa_tree_sub_104_22_n_6 ,in27[3]);
  not csa_tree_sub_104_22_g140(n_591 ,in26[0]);
  not csa_tree_sub_104_22_g141(csa_tree_sub_104_22_n_4 ,in27[1]);
  not csa_tree_sub_104_22_g142(csa_tree_sub_104_22_n_3 ,in27[2]);
  not csa_tree_sub_104_22_g143(csa_tree_sub_104_22_n_2 ,in26[4]);
  xnor mul_84_22_g2868(n_190 ,mul_84_22_n_984 ,mul_84_22_n_1157);
  nor mul_84_22_g2869(mul_84_22_n_1157 ,mul_84_22_n_1026 ,mul_84_22_n_1155);
  xnor mul_84_22_g2870(mul_84_22_n_1156 ,mul_84_22_n_1154 ,mul_84_22_n_1040);
  and mul_84_22_g2871(mul_84_22_n_1155 ,mul_84_22_n_1027 ,mul_84_22_n_1154);
  or mul_84_22_g2872(mul_84_22_n_1154 ,mul_84_22_n_1050 ,mul_84_22_n_1152);
  xnor mul_84_22_g2873(mul_84_22_n_1153 ,mul_84_22_n_1151 ,mul_84_22_n_1061);
  and mul_84_22_g2874(mul_84_22_n_1152 ,mul_84_22_n_1051 ,mul_84_22_n_1151);
  or mul_84_22_g2875(mul_84_22_n_1151 ,mul_84_22_n_1079 ,mul_84_22_n_1149);
  xnor mul_84_22_g2876(mul_84_22_n_1150 ,mul_84_22_n_1148 ,mul_84_22_n_1081);
  nor mul_84_22_g2877(mul_84_22_n_1149 ,mul_84_22_n_1072 ,mul_84_22_n_1148);
  and mul_84_22_g2878(mul_84_22_n_1148 ,mul_84_22_n_1094 ,mul_84_22_n_1146);
  xnor mul_84_22_g2879(mul_84_22_n_1147 ,mul_84_22_n_1144 ,mul_84_22_n_1106);
  or mul_84_22_g2880(mul_84_22_n_1146 ,mul_84_22_n_1093 ,mul_84_22_n_1145);
  not mul_84_22_g2881(mul_84_22_n_1145 ,mul_84_22_n_1144);
  or mul_84_22_g2882(mul_84_22_n_1144 ,mul_84_22_n_1073 ,mul_84_22_n_1142);
  xnor mul_84_22_g2883(mul_84_22_n_1143 ,mul_84_22_n_1141 ,mul_84_22_n_1082);
  and mul_84_22_g2884(mul_84_22_n_1142 ,mul_84_22_n_1080 ,mul_84_22_n_1141);
  or mul_84_22_g2885(mul_84_22_n_1141 ,mul_84_22_n_1087 ,mul_84_22_n_1139);
  xnor mul_84_22_g2886(mul_84_22_n_1140 ,mul_84_22_n_1138 ,mul_84_22_n_1105);
  and mul_84_22_g2887(mul_84_22_n_1139 ,mul_84_22_n_1086 ,mul_84_22_n_1138);
  or mul_84_22_g2888(mul_84_22_n_1138 ,mul_84_22_n_1085 ,mul_84_22_n_1136);
  xnor mul_84_22_g2889(mul_84_22_n_1137 ,mul_84_22_n_1135 ,mul_84_22_n_1104);
  nor mul_84_22_g2890(mul_84_22_n_1136 ,mul_84_22_n_1135 ,mul_84_22_n_1099);
  and mul_84_22_g2891(mul_84_22_n_1135 ,mul_84_22_n_1092 ,mul_84_22_n_1133);
  xnor mul_84_22_g2892(mul_84_22_n_1134 ,mul_84_22_n_1131 ,mul_84_22_n_1103);
  or mul_84_22_g2893(mul_84_22_n_1133 ,mul_84_22_n_1090 ,mul_84_22_n_1132);
  not mul_84_22_g2894(mul_84_22_n_1132 ,mul_84_22_n_1131);
  or mul_84_22_g2895(mul_84_22_n_1131 ,mul_84_22_n_1089 ,mul_84_22_n_1129);
  xnor mul_84_22_g2896(mul_84_22_n_1130 ,mul_84_22_n_1128 ,mul_84_22_n_1102);
  and mul_84_22_g2897(mul_84_22_n_1129 ,mul_84_22_n_1088 ,mul_84_22_n_1128);
  or mul_84_22_g2898(mul_84_22_n_1128 ,mul_84_22_n_1075 ,mul_84_22_n_1126);
  xnor mul_84_22_g2899(mul_84_22_n_1127 ,mul_84_22_n_1125 ,mul_84_22_n_1084);
  and mul_84_22_g2900(mul_84_22_n_1126 ,mul_84_22_n_1074 ,mul_84_22_n_1125);
  or mul_84_22_g2901(mul_84_22_n_1125 ,mul_84_22_n_1098 ,mul_84_22_n_1123);
  xnor mul_84_22_g2902(mul_84_22_n_1124 ,mul_84_22_n_1122 ,mul_84_22_n_1101);
  and mul_84_22_g2903(mul_84_22_n_1123 ,mul_84_22_n_1097 ,mul_84_22_n_1122);
  or mul_84_22_g2904(mul_84_22_n_1122 ,mul_84_22_n_1078 ,mul_84_22_n_1120);
  xnor mul_84_22_g2905(mul_84_22_n_1121 ,mul_84_22_n_1119 ,mul_84_22_n_1083);
  and mul_84_22_g2906(mul_84_22_n_1120 ,mul_84_22_n_1077 ,mul_84_22_n_1119);
  or mul_84_22_g2907(mul_84_22_n_1119 ,mul_84_22_n_1096 ,mul_84_22_n_1117);
  xnor mul_84_22_g2908(mul_84_22_n_1118 ,mul_84_22_n_1116 ,mul_84_22_n_1100);
  and mul_84_22_g2909(mul_84_22_n_1117 ,mul_84_22_n_1095 ,mul_84_22_n_1116);
  or mul_84_22_g2910(mul_84_22_n_1116 ,mul_84_22_n_1041 ,mul_84_22_n_1114);
  xnor mul_84_22_g2911(mul_84_22_n_1115 ,mul_84_22_n_1113 ,mul_84_22_n_1060);
  and mul_84_22_g2912(mul_84_22_n_1114 ,mul_84_22_n_1042 ,mul_84_22_n_1113);
  or mul_84_22_g2913(mul_84_22_n_1113 ,mul_84_22_n_1043 ,mul_84_22_n_1111);
  xnor mul_84_22_g2914(mul_84_22_n_1112 ,mul_84_22_n_1110 ,mul_84_22_n_1059);
  and mul_84_22_g2915(mul_84_22_n_1111 ,mul_84_22_n_1044 ,mul_84_22_n_1110);
  or mul_84_22_g2916(mul_84_22_n_1110 ,mul_84_22_n_6 ,mul_84_22_n_1109);
  nor mul_84_22_g2917(mul_84_22_n_1109 ,mul_84_22_n_1016 ,mul_84_22_n_1108);
  nor mul_84_22_g2918(mul_84_22_n_1108 ,mul_84_22_n_5 ,mul_84_22_n_1107);
  nor mul_84_22_g2919(mul_84_22_n_1107 ,mul_84_22_n_1003 ,mul_84_22_n_1091);
  xnor mul_84_22_g2920(mul_84_22_n_1106 ,mul_84_22_n_1062 ,mul_84_22_n_1039);
  xnor mul_84_22_g2921(mul_84_22_n_1105 ,mul_84_22_n_1019 ,mul_84_22_n_1063);
  xnor mul_84_22_g2922(mul_84_22_n_1104 ,mul_84_22_n_1038 ,mul_84_22_n_1070);
  xnor mul_84_22_g2923(mul_84_22_n_1103 ,mul_84_22_n_1037 ,mul_84_22_n_1069);
  xnor mul_84_22_g2924(mul_84_22_n_1102 ,mul_84_22_n_1055 ,mul_84_22_n_1066);
  xnor mul_84_22_g2925(mul_84_22_n_1101 ,mul_84_22_n_1065 ,mul_84_22_n_1058);
  xnor mul_84_22_g2926(mul_84_22_n_1100 ,mul_84_22_n_1035 ,mul_84_22_n_1067);
  and mul_84_22_g2927(mul_84_22_n_1099 ,mul_84_22_n_1038 ,mul_84_22_n_1071);
  nor mul_84_22_g2928(mul_84_22_n_1098 ,mul_84_22_n_1058 ,mul_84_22_n_1065);
  or mul_84_22_g2929(mul_84_22_n_1097 ,mul_84_22_n_1057 ,mul_84_22_n_1064);
  and mul_84_22_g2930(mul_84_22_n_1096 ,mul_84_22_n_1035 ,mul_84_22_n_1067);
  or mul_84_22_g2931(mul_84_22_n_1095 ,mul_84_22_n_1035 ,mul_84_22_n_1067);
  or mul_84_22_g2932(mul_84_22_n_1094 ,mul_84_22_n_1039 ,mul_84_22_n_1062);
  and mul_84_22_g2933(mul_84_22_n_1093 ,mul_84_22_n_1039 ,mul_84_22_n_1062);
  or mul_84_22_g2934(mul_84_22_n_1092 ,mul_84_22_n_1036 ,mul_84_22_n_1068);
  nor mul_84_22_g2935(mul_84_22_n_1091 ,mul_84_22_n_1000 ,mul_84_22_n_1076);
  nor mul_84_22_g2936(mul_84_22_n_1090 ,mul_84_22_n_1037 ,mul_84_22_n_1069);
  and mul_84_22_g2937(mul_84_22_n_1089 ,mul_84_22_n_1055 ,mul_84_22_n_1066);
  or mul_84_22_g2938(mul_84_22_n_1088 ,mul_84_22_n_1055 ,mul_84_22_n_1066);
  and mul_84_22_g2939(mul_84_22_n_1087 ,mul_84_22_n_1019 ,mul_84_22_n_1063);
  or mul_84_22_g2940(mul_84_22_n_1086 ,mul_84_22_n_1019 ,mul_84_22_n_1063);
  nor mul_84_22_g2941(mul_84_22_n_1085 ,mul_84_22_n_1038 ,mul_84_22_n_1071);
  xnor mul_84_22_g2942(mul_84_22_n_1084 ,mul_84_22_n_1056 ,mul_84_22_n_1045);
  xnor mul_84_22_g2943(mul_84_22_n_1083 ,mul_84_22_n_1047 ,mul_84_22_n_1053);
  xnor mul_84_22_g2944(mul_84_22_n_1082 ,mul_84_22_n_1034 ,mul_84_22_n_1048);
  xnor mul_84_22_g2945(mul_84_22_n_1081 ,mul_84_22_n_1054 ,mul_84_22_n_1017);
  or mul_84_22_g2946(mul_84_22_n_1080 ,mul_84_22_n_1034 ,mul_84_22_n_1048);
  nor mul_84_22_g2947(mul_84_22_n_1079 ,mul_84_22_n_1054 ,mul_84_22_n_1018);
  nor mul_84_22_g2948(mul_84_22_n_1078 ,mul_84_22_n_1053 ,mul_84_22_n_1047);
  or mul_84_22_g2949(mul_84_22_n_1077 ,mul_84_22_n_1052 ,mul_84_22_n_1046);
  nor mul_84_22_g2950(mul_84_22_n_1076 ,mul_84_22_n_999 ,mul_84_22_n_1049);
  and mul_84_22_g2951(mul_84_22_n_1075 ,mul_84_22_n_1056 ,mul_84_22_n_1045);
  or mul_84_22_g2952(mul_84_22_n_1074 ,mul_84_22_n_1056 ,mul_84_22_n_1045);
  and mul_84_22_g2953(mul_84_22_n_1073 ,mul_84_22_n_1034 ,mul_84_22_n_1048);
  and mul_84_22_g2954(mul_84_22_n_1072 ,mul_84_22_n_1054 ,mul_84_22_n_1018);
  not mul_84_22_g2955(mul_84_22_n_1071 ,mul_84_22_n_1070);
  not mul_84_22_g2956(mul_84_22_n_1069 ,mul_84_22_n_1068);
  not mul_84_22_g2957(mul_84_22_n_1065 ,mul_84_22_n_1064);
  xnor mul_84_22_g2958(mul_84_22_n_1061 ,mul_84_22_n_1023 ,mul_84_22_n_1033);
  xnor mul_84_22_g2959(mul_84_22_n_1060 ,mul_84_22_n_1009 ,mul_84_22_n_1021);
  xnor mul_84_22_g2960(mul_84_22_n_1059 ,mul_84_22_n_1010 ,mul_84_22_n_1020);
  xnor mul_84_22_g2961(mul_84_22_n_1070 ,mul_84_22_n_941 ,mul_84_22_n_1011);
  xnor mul_84_22_g2962(mul_84_22_n_1068 ,mul_84_22_n_925 ,mul_84_22_n_4);
  xnor mul_84_22_g2963(mul_84_22_n_1067 ,mul_84_22_n_945 ,mul_84_22_n_1014);
  xnor mul_84_22_g2964(mul_84_22_n_1066 ,mul_84_22_n_942 ,mul_84_22_n_3);
  xnor mul_84_22_g2965(mul_84_22_n_1064 ,mul_84_22_n_912 ,mul_84_22_n_1012);
  xnor mul_84_22_g2966(mul_84_22_n_1063 ,mul_84_22_n_939 ,mul_84_22_n_1013);
  xnor mul_84_22_g2967(mul_84_22_n_1062 ,mul_84_22_n_944 ,mul_84_22_n_1015);
  not mul_84_22_g2968(mul_84_22_n_1057 ,mul_84_22_n_1058);
  not mul_84_22_g2969(mul_84_22_n_1052 ,mul_84_22_n_1053);
  or mul_84_22_g2970(mul_84_22_n_1051 ,mul_84_22_n_1032 ,mul_84_22_n_1022);
  nor mul_84_22_g2971(mul_84_22_n_1050 ,mul_84_22_n_1033 ,mul_84_22_n_1023);
  nor mul_84_22_g2972(mul_84_22_n_1049 ,mul_84_22_n_921 ,mul_84_22_n_1031);
  and mul_84_22_g2973(mul_84_22_n_1058 ,mul_84_22_n_993 ,mul_84_22_n_1024);
  or mul_84_22_g2974(mul_84_22_n_1056 ,mul_84_22_n_1005 ,mul_84_22_n_1030);
  or mul_84_22_g2975(mul_84_22_n_1055 ,mul_84_22_n_997 ,mul_84_22_n_1025);
  and mul_84_22_g2976(mul_84_22_n_1054 ,mul_84_22_n_1007 ,mul_84_22_n_1029);
  and mul_84_22_g2977(mul_84_22_n_1053 ,mul_84_22_n_991 ,mul_84_22_n_1028);
  not mul_84_22_g2978(mul_84_22_n_1047 ,mul_84_22_n_1046);
  or mul_84_22_g2979(mul_84_22_n_1044 ,mul_84_22_n_1010 ,mul_84_22_n_1020);
  and mul_84_22_g2980(mul_84_22_n_1043 ,mul_84_22_n_1010 ,mul_84_22_n_1020);
  or mul_84_22_g2981(mul_84_22_n_1042 ,mul_84_22_n_1009 ,mul_84_22_n_1021);
  and mul_84_22_g2982(mul_84_22_n_1041 ,mul_84_22_n_1009 ,mul_84_22_n_1021);
  xnor mul_84_22_g2983(mul_84_22_n_1040 ,mul_84_22_n_927 ,mul_84_22_n_995);
  xnor mul_84_22_g2984(mul_84_22_n_1048 ,mul_84_22_n_940 ,mul_84_22_n_2);
  xnor mul_84_22_g2985(mul_84_22_n_1046 ,mul_84_22_n_956 ,mul_84_22_n_983);
  xnor mul_84_22_g2986(mul_84_22_n_1045 ,mul_84_22_n_952 ,mul_84_22_n_985);
  not mul_84_22_g2987(mul_84_22_n_1037 ,mul_84_22_n_1036);
  not mul_84_22_g2988(mul_84_22_n_1033 ,mul_84_22_n_1032);
  nor mul_84_22_g2989(mul_84_22_n_1031 ,mul_84_22_n_920 ,mul_84_22_n_1002);
  and mul_84_22_g2990(mul_84_22_n_1030 ,mul_84_22_n_912 ,mul_84_22_n_987);
  or mul_84_22_g2991(mul_84_22_n_1029 ,mul_84_22_n_944 ,mul_84_22_n_1004);
  or mul_84_22_g2992(mul_84_22_n_1028 ,mul_84_22_n_945 ,mul_84_22_n_990);
  or mul_84_22_g2993(mul_84_22_n_1027 ,mul_84_22_n_927 ,mul_84_22_n_995);
  and mul_84_22_g2994(mul_84_22_n_1026 ,mul_84_22_n_927 ,mul_84_22_n_995);
  nor mul_84_22_g2995(mul_84_22_n_1025 ,mul_84_22_n_943 ,mul_84_22_n_1001);
  or mul_84_22_g2996(mul_84_22_n_1024 ,mul_84_22_n_929 ,mul_84_22_n_992);
  and mul_84_22_g2997(mul_84_22_n_1039 ,mul_84_22_n_973 ,mul_84_22_n_994);
  and mul_84_22_g2998(mul_84_22_n_1038 ,mul_84_22_n_969 ,mul_84_22_n_989);
  and mul_84_22_g2999(mul_84_22_n_1036 ,mul_84_22_n_971 ,mul_84_22_n_998);
  or mul_84_22_g3000(mul_84_22_n_1035 ,mul_84_22_n_976 ,mul_84_22_n_986);
  or mul_84_22_g3001(mul_84_22_n_1034 ,mul_84_22_n_978 ,mul_84_22_n_1006);
  or mul_84_22_g3002(mul_84_22_n_1032 ,mul_84_22_n_937 ,mul_84_22_n_1008);
  not mul_84_22_g3003(mul_84_22_n_1022 ,mul_84_22_n_1023);
  not mul_84_22_g3004(mul_84_22_n_1018 ,mul_84_22_n_1017);
  nor mul_84_22_g3006(mul_84_22_n_1016 ,mul_84_22_n_982 ,mul_84_22_n_996);
  xnor mul_84_22_g3007(mul_84_22_n_1015 ,mul_84_22_n_959 ,mul_84_22_n_862);
  xnor mul_84_22_g3008(mul_84_22_n_1014 ,mul_84_22_n_794 ,mul_84_22_n_954);
  xnor mul_84_22_g3009(mul_84_22_n_1013 ,mul_84_22_n_878 ,mul_84_22_n_962);
  xnor mul_84_22_g3010(mul_84_22_n_1012 ,mul_84_22_n_958 ,mul_84_22_n_885);
  xnor mul_84_22_g3011(mul_84_22_n_1011 ,mul_84_22_n_906 ,mul_84_22_n_961);
  xnor mul_84_22_g3014(mul_84_22_n_1023 ,mul_84_22_n_842 ,mul_84_22_n_947);
  xnor mul_84_22_g3015(mul_84_22_n_1021 ,mul_84_22_n_926 ,mul_84_22_n_946);
  xnor mul_84_22_g3016(mul_84_22_n_1020 ,mul_84_22_n_928 ,mul_84_22_n_948);
  or mul_84_22_g3017(mul_84_22_n_1019 ,mul_84_22_n_951 ,mul_84_22_n_988);
  xnor mul_84_22_g3018(mul_84_22_n_1017 ,mul_84_22_n_981 ,mul_84_22_n_949);
  and mul_84_22_g3020(mul_84_22_n_1008 ,mul_84_22_n_981 ,mul_84_22_n_931);
  or mul_84_22_g3021(mul_84_22_n_1007 ,mul_84_22_n_862 ,mul_84_22_n_959);
  and mul_84_22_g3022(mul_84_22_n_1006 ,mul_84_22_n_962 ,mul_84_22_n_977);
  nor mul_84_22_g3023(mul_84_22_n_1005 ,mul_84_22_n_182 ,mul_84_22_n_958);
  and mul_84_22_g3024(mul_84_22_n_1004 ,mul_84_22_n_862 ,mul_84_22_n_959);
  nor mul_84_22_g3025(mul_84_22_n_1003 ,mul_84_22_n_913 ,mul_84_22_n_966);
  nor mul_84_22_g3026(mul_84_22_n_1002 ,mul_84_22_n_935 ,mul_84_22_n_979);
  and mul_84_22_g3027(mul_84_22_n_1001 ,mul_84_22_n_886 ,mul_84_22_n_952);
  nor mul_84_22_g3028(mul_84_22_n_1000 ,mul_84_22_n_848 ,mul_84_22_n_965);
  nor mul_84_22_g3029(mul_84_22_n_999 ,mul_84_22_n_849 ,mul_84_22_n_964);
  or mul_84_22_g3030(mul_84_22_n_998 ,mul_84_22_n_970 ,mul_84_22_n_960);
  nor mul_84_22_g3031(mul_84_22_n_997 ,mul_84_22_n_886 ,mul_84_22_n_952);
  or mul_84_22_g3032(mul_84_22_n_1010 ,mul_84_22_n_923 ,mul_84_22_n_972);
  or mul_84_22_g3033(mul_84_22_n_1009 ,mul_84_22_n_918 ,mul_84_22_n_974);
  or mul_84_22_g3035(mul_84_22_n_994 ,mul_84_22_n_930 ,mul_84_22_n_980);
  or mul_84_22_g3036(mul_84_22_n_993 ,mul_84_22_n_884 ,mul_84_22_n_955);
  nor mul_84_22_g3037(mul_84_22_n_992 ,mul_84_22_n_883 ,mul_84_22_n_956);
  or mul_84_22_g3038(mul_84_22_n_991 ,mul_84_22_n_794 ,mul_84_22_n_953);
  nor mul_84_22_g3039(mul_84_22_n_990 ,mul_84_22_n_793 ,mul_84_22_n_954);
  or mul_84_22_g3040(mul_84_22_n_989 ,mul_84_22_n_968 ,mul_84_22_n_963);
  nor mul_84_22_g3041(mul_84_22_n_988 ,mul_84_22_n_950 ,mul_84_22_n_961);
  or mul_84_22_g3042(mul_84_22_n_987 ,mul_84_22_n_308 ,mul_84_22_n_957);
  nor mul_84_22_g3043(mul_84_22_n_986 ,mul_84_22_n_840 ,mul_84_22_n_975);
  xor mul_84_22_g3044(mul_84_22_n_985 ,mul_84_22_n_943 ,mul_84_22_n_886);
  xnor mul_84_22_g3046(mul_84_22_n_984 ,mul_84_22_n_0 ,mul_84_22_n_916);
  xnor mul_84_22_g3047(mul_84_22_n_996 ,mul_84_22_n_876 ,mul_84_22_n_1);
  xnor mul_84_22_g3048(mul_84_22_n_983 ,mul_84_22_n_929 ,mul_84_22_n_884);
  or mul_84_22_g3049(mul_84_22_n_995 ,mul_84_22_n_933 ,mul_84_22_n_967);
  and mul_84_22_g3051(mul_84_22_n_980 ,mul_84_22_n_890 ,mul_84_22_n_940);
  and mul_84_22_g3052(mul_84_22_n_979 ,mul_84_22_n_802 ,mul_84_22_n_934);
  nor mul_84_22_g3053(mul_84_22_n_978 ,mul_84_22_n_878 ,mul_84_22_n_939);
  or mul_84_22_g3054(mul_84_22_n_977 ,mul_84_22_n_877 ,mul_84_22_n_938);
  nor mul_84_22_g3055(mul_84_22_n_976 ,mul_84_22_n_905 ,mul_84_22_n_926);
  and mul_84_22_g3056(mul_84_22_n_975 ,mul_84_22_n_905 ,mul_84_22_n_926);
  and mul_84_22_g3057(mul_84_22_n_974 ,mul_84_22_n_928 ,mul_84_22_n_917);
  or mul_84_22_g3058(mul_84_22_n_973 ,mul_84_22_n_890 ,mul_84_22_n_940);
  nor mul_84_22_g3059(mul_84_22_n_972 ,mul_84_22_n_847 ,mul_84_22_n_919);
  or mul_84_22_g3060(mul_84_22_n_971 ,mul_84_22_n_889 ,mul_84_22_n_942);
  and mul_84_22_g3061(mul_84_22_n_970 ,mul_84_22_n_889 ,mul_84_22_n_942);
  or mul_84_22_g3062(mul_84_22_n_969 ,mul_84_22_n_882 ,mul_84_22_n_924);
  nor mul_84_22_g3063(mul_84_22_n_968 ,mul_84_22_n_881 ,mul_84_22_n_925);
  and mul_84_22_g3064(mul_84_22_n_967 ,mul_84_22_n_842 ,mul_84_22_n_936);
  or mul_84_22_g3065(mul_84_22_n_982 ,mul_84_22_n_705 ,mul_84_22_n_922);
  or mul_84_22_g3066(mul_84_22_n_981 ,mul_84_22_n_746 ,mul_84_22_n_932);
  not mul_84_22_g3068(mul_84_22_n_965 ,mul_84_22_n_964);
  not mul_84_22_g3071(mul_84_22_n_958 ,mul_84_22_n_957);
  not mul_84_22_g3072(mul_84_22_n_956 ,mul_84_22_n_955);
  not mul_84_22_g3073(mul_84_22_n_953 ,mul_84_22_n_954);
  nor mul_84_22_g3074(mul_84_22_n_951 ,mul_84_22_n_907 ,mul_84_22_n_941);
  and mul_84_22_g3075(mul_84_22_n_950 ,mul_84_22_n_907 ,mul_84_22_n_941);
  xnor mul_84_22_g3076(mul_84_22_n_966 ,mul_84_22_n_910 ,mul_84_22_n_780);
  xnor mul_84_22_g3077(mul_84_22_n_964 ,mul_84_22_n_602 ,mul_84_22_n_875);
  xnor mul_84_22_g3078(mul_84_22_n_949 ,mul_84_22_n_888 ,mul_84_22_n_839);
  xnor mul_84_22_g3079(mul_84_22_n_948 ,mul_84_22_n_880 ,mul_84_22_n_909);
  xnor mul_84_22_g3080(mul_84_22_n_947 ,mul_84_22_n_904 ,mul_84_22_n_649);
  xor mul_84_22_g3081(mul_84_22_n_946 ,mul_84_22_n_905 ,mul_84_22_n_840);
  xnor mul_84_22_g3082(mul_84_22_n_963 ,mul_84_22_n_841 ,mul_84_22_n_868);
  xnor mul_84_22_g3083(mul_84_22_n_962 ,mul_84_22_n_867 ,mul_84_22_n_870);
  xnor mul_84_22_g3084(mul_84_22_n_961 ,mul_84_22_n_866 ,mul_84_22_n_869);
  xnor mul_84_22_g3085(mul_84_22_n_960 ,mul_84_22_n_845 ,mul_84_22_n_874);
  xnor mul_84_22_g3086(mul_84_22_n_959 ,mul_84_22_n_911 ,mul_84_22_n_787);
  xnor mul_84_22_g3087(mul_84_22_n_957 ,mul_84_22_n_865 ,mul_84_22_n_872);
  xnor mul_84_22_g3088(mul_84_22_n_955 ,mul_84_22_n_762 ,mul_84_22_n_871);
  xnor mul_84_22_g3089(mul_84_22_n_954 ,mul_84_22_n_843 ,mul_84_22_n_893);
  xnor mul_84_22_g3090(mul_84_22_n_952 ,mul_84_22_n_864 ,mul_84_22_n_873);
  not mul_84_22_g3091(mul_84_22_n_939 ,mul_84_22_n_938);
  nor mul_84_22_g3092(mul_84_22_n_937 ,mul_84_22_n_839 ,mul_84_22_n_888);
  or mul_84_22_g3093(mul_84_22_n_936 ,mul_84_22_n_204 ,mul_84_22_n_904);
  nor mul_84_22_g3094(mul_84_22_n_935 ,mul_84_22_n_643 ,mul_84_22_n_914);
  or mul_84_22_g3095(mul_84_22_n_934 ,mul_84_22_n_644 ,mul_84_22_n_915);
  and mul_84_22_g3096(mul_84_22_n_933 ,mul_84_22_n_203 ,mul_84_22_n_904);
  and mul_84_22_g3097(mul_84_22_n_932 ,mul_84_22_n_755 ,mul_84_22_n_911);
  or mul_84_22_g3098(mul_84_22_n_931 ,mul_84_22_n_838 ,mul_84_22_n_887);
  and mul_84_22_g3099(mul_84_22_n_945 ,mul_84_22_n_754 ,mul_84_22_n_899);
  and mul_84_22_g3100(mul_84_22_n_944 ,mul_84_22_n_804 ,mul_84_22_n_897);
  and mul_84_22_g3101(mul_84_22_n_943 ,mul_84_22_n_857 ,mul_84_22_n_901);
  and mul_84_22_g3102(mul_84_22_n_942 ,mul_84_22_n_861 ,mul_84_22_n_902);
  and mul_84_22_g3103(mul_84_22_n_941 ,mul_84_22_n_832 ,mul_84_22_n_898);
  and mul_84_22_g3104(mul_84_22_n_940 ,mul_84_22_n_855 ,mul_84_22_n_903);
  or mul_84_22_g3105(mul_84_22_n_938 ,mul_84_22_n_854 ,mul_84_22_n_900);
  not mul_84_22_g3107(mul_84_22_n_924 ,mul_84_22_n_925);
  nor mul_84_22_g3108(mul_84_22_n_923 ,mul_84_22_n_599 ,mul_84_22_n_876);
  and mul_84_22_g3109(mul_84_22_n_922 ,mul_84_22_n_704 ,mul_84_22_n_910);
  nor mul_84_22_g3110(mul_84_22_n_921 ,mul_84_22_n_769 ,mul_84_22_n_891);
  nor mul_84_22_g3111(mul_84_22_n_920 ,mul_84_22_n_768 ,mul_84_22_n_892);
  and mul_84_22_g3112(mul_84_22_n_919 ,mul_84_22_n_599 ,mul_84_22_n_876);
  nor mul_84_22_g3113(mul_84_22_n_918 ,mul_84_22_n_909 ,mul_84_22_n_880);
  or mul_84_22_g3114(mul_84_22_n_917 ,mul_84_22_n_908 ,mul_84_22_n_879);
  or mul_84_22_g3116(mul_84_22_n_916 ,mul_84_22_n_719 ,mul_84_22_n_894);
  xnor mul_84_22_g3117(mul_84_22_n_930 ,mul_84_22_n_844 ,mul_84_22_n_830);
  and mul_84_22_g3118(mul_84_22_n_929 ,mul_84_22_n_851 ,mul_84_22_n_895);
  xnor mul_84_22_g3119(mul_84_22_n_928 ,mul_84_22_n_606 ,mul_84_22_n_831);
  xnor mul_84_22_g3120(mul_84_22_n_927 ,mul_84_22_n_863 ,mul_84_22_n_782);
  xnor mul_84_22_g3121(mul_84_22_n_926 ,mul_84_22_n_846 ,mul_84_22_n_783);
  or mul_84_22_g3122(mul_84_22_n_925 ,mul_84_22_n_835 ,mul_84_22_n_896);
  not mul_84_22_g3123(mul_84_22_n_915 ,mul_84_22_n_914);
  not mul_84_22_g3125(mul_84_22_n_908 ,mul_84_22_n_909);
  not mul_84_22_g3126(mul_84_22_n_907 ,mul_84_22_n_906);
  or mul_84_22_g3127(mul_84_22_n_903 ,mul_84_22_n_858 ,mul_84_22_n_867);
  or mul_84_22_g3128(mul_84_22_n_902 ,mul_84_22_n_860 ,mul_84_22_n_864);
  or mul_84_22_g3129(mul_84_22_n_901 ,mul_84_22_n_856 ,mul_84_22_n_865);
  nor mul_84_22_g3130(mul_84_22_n_900 ,mul_84_22_n_852 ,mul_84_22_n_866);
  or mul_84_22_g3131(mul_84_22_n_899 ,mul_84_22_n_726 ,mul_84_22_n_846);
  or mul_84_22_g3132(mul_84_22_n_898 ,mul_84_22_n_837 ,mul_84_22_n_841);
  or mul_84_22_g3133(mul_84_22_n_897 ,mul_84_22_n_803 ,mul_84_22_n_844);
  nor mul_84_22_g3134(mul_84_22_n_896 ,mul_84_22_n_834 ,mul_84_22_n_845);
  or mul_84_22_g3135(mul_84_22_n_895 ,mul_84_22_n_843 ,mul_84_22_n_850);
  and mul_84_22_g3136(mul_84_22_n_894 ,mul_84_22_n_720 ,mul_84_22_n_863);
  and mul_84_22_g3137(mul_84_22_n_914 ,mul_84_22_n_753 ,mul_84_22_n_859);
  xnor mul_84_22_g3138(mul_84_22_n_893 ,mul_84_22_n_663 ,mul_84_22_n_792);
  xnor mul_84_22_g3139(mul_84_22_n_913 ,mul_84_22_n_731 ,mul_84_22_n_774);
  or mul_84_22_g3140(mul_84_22_n_912 ,mul_84_22_n_816 ,mul_84_22_n_853);
  xnor mul_84_22_g3141(mul_84_22_n_911 ,mul_84_22_n_692 ,mul_84_22_n_800);
  or mul_84_22_g3142(mul_84_22_n_910 ,mul_84_22_n_703 ,mul_84_22_n_833);
  and mul_84_22_g3143(mul_84_22_n_909 ,mul_84_22_n_713 ,mul_84_22_n_836);
  xnor mul_84_22_g3144(mul_84_22_n_906 ,mul_84_22_n_672 ,mul_84_22_n_785);
  xnor mul_84_22_g3145(mul_84_22_n_905 ,mul_84_22_n_661 ,mul_84_22_n_779);
  xnor mul_84_22_g3146(mul_84_22_n_904 ,mul_84_22_n_687 ,mul_84_22_n_777);
  not mul_84_22_g3147(mul_84_22_n_892 ,mul_84_22_n_891);
  not mul_84_22_g3148(mul_84_22_n_888 ,mul_84_22_n_887);
  not mul_84_22_g3150(mul_84_22_n_883 ,mul_84_22_n_884);
  not mul_84_22_g3151(mul_84_22_n_881 ,mul_84_22_n_882);
  not mul_84_22_g3152(mul_84_22_n_879 ,mul_84_22_n_880);
  not mul_84_22_g3153(mul_84_22_n_877 ,mul_84_22_n_878);
  xnor mul_84_22_g3154(mul_84_22_n_875 ,mul_84_22_n_618 ,mul_84_22_n_797);
  xnor mul_84_22_g3155(mul_84_22_n_874 ,mul_84_22_n_758 ,mul_84_22_n_796);
  xnor mul_84_22_g3156(mul_84_22_n_873 ,mul_84_22_n_764 ,mul_84_22_n_829);
  xnor mul_84_22_g3157(mul_84_22_n_872 ,mul_84_22_n_760 ,mul_84_22_n_827);
  xnor mul_84_22_g3158(mul_84_22_n_871 ,mul_84_22_n_767 ,mul_84_22_n_799);
  xnor mul_84_22_g3159(mul_84_22_n_870 ,mul_84_22_n_757 ,mul_84_22_n_825);
  xnor mul_84_22_g3160(mul_84_22_n_869 ,mul_84_22_n_765 ,mul_84_22_n_795);
  xnor mul_84_22_g3161(mul_84_22_n_868 ,mul_84_22_n_730 ,mul_84_22_n_790);
  xnor mul_84_22_g3162(mul_84_22_n_891 ,mul_84_22_n_641 ,mul_84_22_n_775);
  xnor mul_84_22_g3164(mul_84_22_n_890 ,mul_84_22_n_697 ,mul_84_22_n_781);
  xnor mul_84_22_g3165(mul_84_22_n_889 ,mul_84_22_n_608 ,mul_84_22_n_778);
  xnor mul_84_22_g3166(mul_84_22_n_887 ,mul_84_22_n_786 ,mul_84_22_n_204);
  xnor mul_84_22_g3167(mul_84_22_n_886 ,mul_84_22_n_621 ,mul_84_22_n_773);
  xnor mul_84_22_g3168(mul_84_22_n_885 ,mul_84_22_n_632 ,mul_84_22_n_771);
  xnor mul_84_22_g3169(mul_84_22_n_884 ,mul_84_22_n_627 ,mul_84_22_n_770);
  xnor mul_84_22_g3170(mul_84_22_n_882 ,mul_84_22_n_664 ,mul_84_22_n_788);
  xnor mul_84_22_g3171(mul_84_22_n_880 ,mul_84_22_n_631 ,mul_84_22_n_776);
  xnor mul_84_22_g3172(mul_84_22_n_878 ,mul_84_22_n_633 ,mul_84_22_n_772);
  xnor mul_84_22_g3173(mul_84_22_n_876 ,mul_84_22_n_798 ,mul_84_22_n_784);
  or mul_84_22_g3174(mul_84_22_n_861 ,mul_84_22_n_763 ,mul_84_22_n_828);
  nor mul_84_22_g3175(mul_84_22_n_860 ,mul_84_22_n_764 ,mul_84_22_n_829);
  or mul_84_22_g3176(mul_84_22_n_859 ,mul_84_22_n_821 ,mul_84_22_n_751);
  nor mul_84_22_g3177(mul_84_22_n_858 ,mul_84_22_n_757 ,mul_84_22_n_824);
  or mul_84_22_g3178(mul_84_22_n_857 ,mul_84_22_n_760 ,mul_84_22_n_826);
  nor mul_84_22_g3179(mul_84_22_n_856 ,mul_84_22_n_759 ,mul_84_22_n_827);
  or mul_84_22_g3180(mul_84_22_n_855 ,mul_84_22_n_756 ,mul_84_22_n_825);
  and mul_84_22_g3181(mul_84_22_n_854 ,mul_84_22_n_765 ,mul_84_22_n_795);
  and mul_84_22_g3182(mul_84_22_n_853 ,mul_84_22_n_799 ,mul_84_22_n_815);
  nor mul_84_22_g3183(mul_84_22_n_852 ,mul_84_22_n_765 ,mul_84_22_n_795);
  or mul_84_22_g3184(mul_84_22_n_851 ,mul_84_22_n_663 ,mul_84_22_n_791);
  nor mul_84_22_g3185(mul_84_22_n_850 ,mul_84_22_n_662 ,mul_84_22_n_792);
  and mul_84_22_g3186(mul_84_22_n_867 ,mul_84_22_n_715 ,mul_84_22_n_820);
  and mul_84_22_g3187(mul_84_22_n_866 ,mul_84_22_n_736 ,mul_84_22_n_814);
  and mul_84_22_g3188(mul_84_22_n_865 ,mul_84_22_n_743 ,mul_84_22_n_817);
  and mul_84_22_g3189(mul_84_22_n_864 ,mul_84_22_n_752 ,mul_84_22_n_819);
  or mul_84_22_g3190(mul_84_22_n_863 ,mul_84_22_n_741 ,mul_84_22_n_818);
  and mul_84_22_g3191(mul_84_22_n_862 ,mul_84_22_n_737 ,mul_84_22_n_813);
  not mul_84_22_g3192(mul_84_22_n_849 ,mul_84_22_n_848);
  not mul_84_22_g3193(mul_84_22_n_838 ,mul_84_22_n_839);
  nor mul_84_22_g3194(mul_84_22_n_837 ,mul_84_22_n_730 ,mul_84_22_n_790);
  or mul_84_22_g3195(mul_84_22_n_836 ,mul_84_22_n_711 ,mul_84_22_n_798);
  and mul_84_22_g3196(mul_84_22_n_835 ,mul_84_22_n_758 ,mul_84_22_n_796);
  nor mul_84_22_g3197(mul_84_22_n_834 ,mul_84_22_n_758 ,mul_84_22_n_796);
  and mul_84_22_g3198(mul_84_22_n_833 ,mul_84_22_n_750 ,mul_84_22_n_797);
  or mul_84_22_g3199(mul_84_22_n_832 ,mul_84_22_n_729 ,mul_84_22_n_789);
  and mul_84_22_g3200(mul_84_22_n_848 ,mul_84_22_n_747 ,mul_84_22_n_822);
  xnor mul_84_22_g3201(mul_84_22_n_831 ,mul_84_22_n_598 ,mul_84_22_n_733);
  xnor mul_84_22_g3202(mul_84_22_n_830 ,mul_84_22_n_728 ,mul_84_22_n_648);
  and mul_84_22_g3203(mul_84_22_n_847 ,mul_84_22_n_709 ,mul_84_22_n_809);
  and mul_84_22_g3204(mul_84_22_n_846 ,mul_84_22_n_735 ,mul_84_22_n_812);
  and mul_84_22_g3205(mul_84_22_n_845 ,mul_84_22_n_710 ,mul_84_22_n_808);
  and mul_84_22_g3206(mul_84_22_n_844 ,mul_84_22_n_745 ,mul_84_22_n_807);
  and mul_84_22_g3207(mul_84_22_n_843 ,mul_84_22_n_738 ,mul_84_22_n_806);
  or mul_84_22_g3208(mul_84_22_n_842 ,mul_84_22_n_725 ,mul_84_22_n_805);
  and mul_84_22_g3209(mul_84_22_n_841 ,mul_84_22_n_722 ,mul_84_22_n_811);
  and mul_84_22_g3210(mul_84_22_n_840 ,mul_84_22_n_721 ,mul_84_22_n_810);
  and mul_84_22_g3211(mul_84_22_n_839 ,mul_84_22_n_706 ,mul_84_22_n_823);
  not mul_84_22_g3212(mul_84_22_n_828 ,mul_84_22_n_829);
  not mul_84_22_g3213(mul_84_22_n_826 ,mul_84_22_n_827);
  not mul_84_22_g3214(mul_84_22_n_824 ,mul_84_22_n_825);
  or mul_84_22_g3215(mul_84_22_n_823 ,mul_84_22_n_692 ,mul_84_22_n_749);
  or mul_84_22_g3216(mul_84_22_n_822 ,mul_84_22_n_641 ,mul_84_22_n_716);
  or mul_84_22_g3217(mul_84_22_n_821 ,mul_84_22_n_327 ,mul_84_22_n_727);
  or mul_84_22_g3218(mul_84_22_n_820 ,mul_84_22_n_630 ,mul_84_22_n_744);
  or mul_84_22_g3219(mul_84_22_n_819 ,mul_84_22_n_632 ,mul_84_22_n_718);
  and mul_84_22_g3220(mul_84_22_n_818 ,mul_84_22_n_687 ,mul_84_22_n_748);
  or mul_84_22_g3221(mul_84_22_n_817 ,mul_84_22_n_627 ,mul_84_22_n_742);
  nor mul_84_22_g3222(mul_84_22_n_816 ,mul_84_22_n_767 ,mul_84_22_n_761);
  or mul_84_22_g3223(mul_84_22_n_815 ,mul_84_22_n_766 ,mul_84_22_n_762);
  or mul_84_22_g3224(mul_84_22_n_814 ,mul_84_22_n_624 ,mul_84_22_n_739);
  or mul_84_22_g3225(mul_84_22_n_813 ,mul_84_22_n_697 ,mul_84_22_n_723);
  or mul_84_22_g3226(mul_84_22_n_812 ,mul_84_22_n_631 ,mul_84_22_n_724);
  or mul_84_22_g3227(mul_84_22_n_811 ,mul_84_22_n_622 ,mul_84_22_n_714);
  or mul_84_22_g3228(mul_84_22_n_810 ,mul_84_22_n_734 ,mul_84_22_n_717);
  or mul_84_22_g3229(mul_84_22_n_809 ,mul_84_22_n_708 ,mul_84_22_n_732);
  or mul_84_22_g3230(mul_84_22_n_808 ,mul_84_22_n_621 ,mul_84_22_n_707);
  or mul_84_22_g3231(mul_84_22_n_807 ,mul_84_22_n_633 ,mul_84_22_n_702);
  or mul_84_22_g3232(mul_84_22_n_806 ,mul_84_22_n_623 ,mul_84_22_n_740);
  nor mul_84_22_g3233(mul_84_22_n_805 ,mul_84_22_n_203 ,mul_84_22_n_712);
  or mul_84_22_g3234(mul_84_22_n_804 ,mul_84_22_n_156 ,mul_84_22_n_728);
  and mul_84_22_g3235(mul_84_22_n_803 ,mul_84_22_n_157 ,mul_84_22_n_728);
  xnor mul_84_22_g3236(mul_84_22_n_802 ,mul_84_22_n_698 ,mul_84_22_n_547);
  xnor mul_84_22_g3237(mul_84_22_n_801 ,mul_84_22_n_647 ,mul_84_22_n_646);
  xnor mul_84_22_g3238(mul_84_22_n_800 ,mul_84_22_n_604 ,mul_84_22_n_656);
  xnor mul_84_22_g3239(mul_84_22_n_829 ,mul_84_22_n_628 ,mul_84_22_n_636);
  xnor mul_84_22_g3240(mul_84_22_n_827 ,mul_84_22_n_679 ,mul_84_22_n_696);
  xnor mul_84_22_g3241(mul_84_22_n_825 ,mul_84_22_n_645 ,mul_84_22_n_700);
  not mul_84_22_g3242(mul_84_22_n_793 ,mul_84_22_n_794);
  not mul_84_22_g3243(mul_84_22_n_791 ,mul_84_22_n_792);
  not mul_84_22_g3244(mul_84_22_n_789 ,mul_84_22_n_790);
  xnor mul_84_22_g3245(mul_84_22_n_788 ,mul_84_22_n_667 ,mul_84_22_n_624);
  xnor mul_84_22_g3246(mul_84_22_n_787 ,mul_84_22_n_677 ,mul_84_22_n_157);
  xnor mul_84_22_g3247(mul_84_22_n_786 ,mul_84_22_n_670 ,mul_84_22_n_611);
  xor mul_84_22_g3248(mul_84_22_n_785 ,mul_84_22_n_666 ,mul_84_22_n_630);
  xnor mul_84_22_g3249(mul_84_22_n_784 ,mul_84_22_n_609 ,mul_84_22_n_669);
  xnor mul_84_22_g3250(mul_84_22_n_783 ,mul_84_22_n_674 ,mul_84_22_n_654);
  xnor mul_84_22_g3251(mul_84_22_n_782 ,mul_84_22_n_614 ,mul_84_22_n_650);
  xnor mul_84_22_g3252(mul_84_22_n_781 ,mul_84_22_n_657 ,mul_84_22_n_612);
  xnor mul_84_22_g3253(mul_84_22_n_780 ,mul_84_22_n_594 ,mul_84_22_n_596);
  xor mul_84_22_g3254(mul_84_22_n_779 ,mul_84_22_n_659 ,mul_84_22_n_623);
  xnor mul_84_22_g3255(mul_84_22_n_778 ,mul_84_22_n_600 ,mul_84_22_n_622);
  xnor mul_84_22_g3256(mul_84_22_n_777 ,mul_84_22_n_616 ,mul_84_22_n_653);
  xnor mul_84_22_g3257(mul_84_22_n_776 ,mul_84_22_n_449 ,mul_84_22_n_673);
  xnor mul_84_22_g3258(mul_84_22_n_775 ,mul_84_22_n_451 ,mul_84_22_n_651);
  xnor mul_84_22_g3259(mul_84_22_n_774 ,mul_84_22_n_450 ,mul_84_22_n_605);
  xnor mul_84_22_g3260(mul_84_22_n_773 ,mul_84_22_n_592 ,mul_84_22_n_597);
  xnor mul_84_22_g3261(mul_84_22_n_772 ,mul_84_22_n_607 ,mul_84_22_n_665);
  xnor mul_84_22_g3262(mul_84_22_n_771 ,mul_84_22_n_610 ,mul_84_22_n_668);
  xnor mul_84_22_g3263(mul_84_22_n_770 ,mul_84_22_n_678 ,mul_84_22_n_675);
  xnor mul_84_22_g3264(mul_84_22_n_799 ,mul_84_22_n_684 ,mul_84_22_n_682);
  xnor mul_84_22_g3265(mul_84_22_n_798 ,mul_84_22_n_639 ,mul_84_22_n_544);
  xnor mul_84_22_g3266(mul_84_22_n_797 ,mul_84_22_n_546 ,mul_84_22_n_634);
  xnor mul_84_22_g3267(mul_84_22_n_796 ,mul_84_22_n_619 ,mul_84_22_n_629);
  xnor mul_84_22_g3268(mul_84_22_n_795 ,mul_84_22_n_694 ,mul_84_22_n_693);
  xnor mul_84_22_g3269(mul_84_22_n_794 ,mul_84_22_n_690 ,mul_84_22_n_625);
  xnor mul_84_22_g3270(mul_84_22_n_792 ,mul_84_22_n_681 ,mul_84_22_n_685);
  xnor mul_84_22_g3271(mul_84_22_n_790 ,mul_84_22_n_638 ,mul_84_22_n_688);
  not mul_84_22_g3272(mul_84_22_n_769 ,mul_84_22_n_768);
  not mul_84_22_g3273(mul_84_22_n_767 ,mul_84_22_n_766);
  not mul_84_22_g3274(mul_84_22_n_764 ,mul_84_22_n_763);
  not mul_84_22_g3275(mul_84_22_n_761 ,mul_84_22_n_762);
  not mul_84_22_g3276(mul_84_22_n_760 ,mul_84_22_n_759);
  not mul_84_22_g3277(mul_84_22_n_757 ,mul_84_22_n_756);
  or mul_84_22_g3278(mul_84_22_n_755 ,mul_84_22_n_156 ,mul_84_22_n_676);
  or mul_84_22_g3279(mul_84_22_n_754 ,mul_84_22_n_654 ,mul_84_22_n_674);
  or mul_84_22_g3280(mul_84_22_n_753 ,mul_84_22_n_456 ,mul_84_22_n_642);
  or mul_84_22_g3281(mul_84_22_n_752 ,mul_84_22_n_668 ,mul_84_22_n_610);
  and mul_84_22_g3282(mul_84_22_n_751 ,mul_84_22_n_456 ,mul_84_22_n_642);
  or mul_84_22_g3283(mul_84_22_n_750 ,mul_84_22_n_601 ,mul_84_22_n_617);
  nor mul_84_22_g3284(mul_84_22_n_749 ,mul_84_22_n_604 ,mul_84_22_n_655);
  or mul_84_22_g3285(mul_84_22_n_748 ,mul_84_22_n_652 ,mul_84_22_n_615);
  or mul_84_22_g3286(mul_84_22_n_747 ,mul_84_22_n_451 ,mul_84_22_n_651);
  nor mul_84_22_g3287(mul_84_22_n_746 ,mul_84_22_n_306 ,mul_84_22_n_677);
  or mul_84_22_g3288(mul_84_22_n_745 ,mul_84_22_n_665 ,mul_84_22_n_607);
  and mul_84_22_g3289(mul_84_22_n_744 ,mul_84_22_n_672 ,mul_84_22_n_666);
  or mul_84_22_g3290(mul_84_22_n_743 ,mul_84_22_n_675 ,mul_84_22_n_678);
  and mul_84_22_g3291(mul_84_22_n_742 ,mul_84_22_n_675 ,mul_84_22_n_678);
  nor mul_84_22_g3292(mul_84_22_n_741 ,mul_84_22_n_653 ,mul_84_22_n_616);
  nor mul_84_22_g3293(mul_84_22_n_740 ,mul_84_22_n_661 ,mul_84_22_n_658);
  and mul_84_22_g3294(mul_84_22_n_739 ,mul_84_22_n_667 ,mul_84_22_n_664);
  or mul_84_22_g3295(mul_84_22_n_738 ,mul_84_22_n_660 ,mul_84_22_n_659);
  or mul_84_22_g3296(mul_84_22_n_737 ,mul_84_22_n_612 ,mul_84_22_n_657);
  or mul_84_22_g3297(mul_84_22_n_736 ,mul_84_22_n_667 ,mul_84_22_n_664);
  or mul_84_22_g3298(mul_84_22_n_735 ,mul_84_22_n_449 ,mul_84_22_n_673);
  and mul_84_22_g3299(mul_84_22_n_768 ,mul_84_22_n_547 ,mul_84_22_n_699);
  and mul_84_22_g3300(mul_84_22_n_766 ,mul_84_22_n_681 ,mul_84_22_n_686);
  and mul_84_22_g3301(mul_84_22_n_765 ,mul_84_22_n_638 ,mul_84_22_n_689);
  or mul_84_22_g3302(mul_84_22_n_763 ,mul_84_22_n_680 ,mul_84_22_n_696);
  and mul_84_22_g3303(mul_84_22_n_762 ,mul_84_22_n_626 ,mul_84_22_n_691);
  and mul_84_22_g3304(mul_84_22_n_759 ,mul_84_22_n_684 ,mul_84_22_n_683);
  and mul_84_22_g3305(mul_84_22_n_758 ,mul_84_22_n_628 ,mul_84_22_n_637);
  or mul_84_22_g3306(mul_84_22_n_756 ,mul_84_22_n_695 ,mul_84_22_n_693);
  not mul_84_22_g3307(mul_84_22_n_734 ,mul_84_22_n_733);
  not mul_84_22_g3308(mul_84_22_n_732 ,mul_84_22_n_731);
  not mul_84_22_g3309(mul_84_22_n_730 ,mul_84_22_n_729);
  or mul_84_22_g3310(mul_84_22_n_727 ,mul_84_22_n_311 ,mul_84_22_n_591);
  and mul_84_22_g3311(mul_84_22_n_726 ,mul_84_22_n_654 ,mul_84_22_n_674);
  nor mul_84_22_g3312(mul_84_22_n_725 ,mul_84_22_n_671 ,mul_84_22_n_611);
  and mul_84_22_g3313(mul_84_22_n_724 ,mul_84_22_n_449 ,mul_84_22_n_673);
  and mul_84_22_g3314(mul_84_22_n_723 ,mul_84_22_n_612 ,mul_84_22_n_657);
  or mul_84_22_g3315(mul_84_22_n_722 ,mul_84_22_n_600 ,mul_84_22_n_608);
  or mul_84_22_g3316(mul_84_22_n_721 ,mul_84_22_n_598 ,mul_84_22_n_606);
  or mul_84_22_g3317(mul_84_22_n_720 ,mul_84_22_n_307 ,mul_84_22_n_613);
  nor mul_84_22_g3318(mul_84_22_n_719 ,mul_84_22_n_650 ,mul_84_22_n_614);
  and mul_84_22_g3319(mul_84_22_n_718 ,mul_84_22_n_668 ,mul_84_22_n_610);
  and mul_84_22_g3320(mul_84_22_n_717 ,mul_84_22_n_598 ,mul_84_22_n_606);
  and mul_84_22_g3321(mul_84_22_n_716 ,mul_84_22_n_451 ,mul_84_22_n_651);
  or mul_84_22_g3322(mul_84_22_n_715 ,mul_84_22_n_672 ,mul_84_22_n_666);
  and mul_84_22_g3323(mul_84_22_n_714 ,mul_84_22_n_600 ,mul_84_22_n_608);
  or mul_84_22_g3324(mul_84_22_n_713 ,mul_84_22_n_669 ,mul_84_22_n_609);
  and mul_84_22_g3325(mul_84_22_n_712 ,mul_84_22_n_671 ,mul_84_22_n_611);
  and mul_84_22_g3326(mul_84_22_n_711 ,mul_84_22_n_669 ,mul_84_22_n_609);
  or mul_84_22_g3327(mul_84_22_n_710 ,mul_84_22_n_597 ,mul_84_22_n_592);
  or mul_84_22_g3328(mul_84_22_n_709 ,mul_84_22_n_450 ,mul_84_22_n_605);
  and mul_84_22_g3329(mul_84_22_n_708 ,mul_84_22_n_450 ,mul_84_22_n_605);
  and mul_84_22_g3330(mul_84_22_n_707 ,mul_84_22_n_597 ,mul_84_22_n_592);
  or mul_84_22_g3331(mul_84_22_n_706 ,mul_84_22_n_603 ,mul_84_22_n_656);
  nor mul_84_22_g3332(mul_84_22_n_705 ,mul_84_22_n_596 ,mul_84_22_n_594);
  or mul_84_22_g3333(mul_84_22_n_704 ,mul_84_22_n_595 ,mul_84_22_n_593);
  nor mul_84_22_g3334(mul_84_22_n_703 ,mul_84_22_n_602 ,mul_84_22_n_618);
  and mul_84_22_g3335(mul_84_22_n_702 ,mul_84_22_n_665 ,mul_84_22_n_607);
  and mul_84_22_g3336(mul_84_22_n_733 ,mul_84_22_n_545 ,mul_84_22_n_640);
  and mul_84_22_g3337(mul_84_22_n_731 ,mul_84_22_n_546 ,mul_84_22_n_635);
  or mul_84_22_g3338(mul_84_22_n_729 ,mul_84_22_n_620 ,mul_84_22_n_629);
  and mul_84_22_g3339(mul_84_22_n_728 ,mul_84_22_n_645 ,mul_84_22_n_701);
  not mul_84_22_g3340(mul_84_22_n_701 ,mul_84_22_n_700);
  not mul_84_22_g3341(mul_84_22_n_699 ,mul_84_22_n_698);
  not mul_84_22_g3342(mul_84_22_n_695 ,mul_84_22_n_694);
  not mul_84_22_g3343(mul_84_22_n_691 ,mul_84_22_n_690);
  not mul_84_22_g3344(mul_84_22_n_689 ,mul_84_22_n_688);
  not mul_84_22_g3345(mul_84_22_n_686 ,mul_84_22_n_685);
  not mul_84_22_g3346(mul_84_22_n_683 ,mul_84_22_n_682);
  not mul_84_22_g3347(mul_84_22_n_680 ,mul_84_22_n_679);
  not mul_84_22_g3348(mul_84_22_n_676 ,mul_84_22_n_677);
  not mul_84_22_g3349(mul_84_22_n_671 ,mul_84_22_n_670);
  not mul_84_22_g3350(mul_84_22_n_662 ,mul_84_22_n_663);
  not mul_84_22_g3351(mul_84_22_n_660 ,mul_84_22_n_661);
  not mul_84_22_g3352(mul_84_22_n_658 ,mul_84_22_n_659);
  not mul_84_22_g3353(mul_84_22_n_655 ,mul_84_22_n_656);
  not mul_84_22_g3354(mul_84_22_n_652 ,mul_84_22_n_653);
  or mul_84_22_g3358(mul_84_22_n_700 ,mul_84_22_n_502 ,mul_84_22_n_578);
  and mul_84_22_g3359(mul_84_22_n_698 ,mul_84_22_n_422 ,mul_84_22_n_536);
  or mul_84_22_g3360(mul_84_22_n_647 ,mul_84_22_n_457 ,mul_84_22_n_506);
  or mul_84_22_g3361(mul_84_22_n_646 ,mul_84_22_n_497 ,mul_84_22_n_580);
  and mul_84_22_g3362(mul_84_22_n_697 ,mul_84_22_n_429 ,mul_84_22_n_565);
  and mul_84_22_g3363(mul_84_22_n_696 ,mul_84_22_n_460 ,mul_84_22_n_561);
  or mul_84_22_g3364(mul_84_22_n_694 ,mul_84_22_n_500 ,mul_84_22_n_588);
  and mul_84_22_g3365(mul_84_22_n_693 ,mul_84_22_n_466 ,mul_84_22_n_573);
  and mul_84_22_g3366(mul_84_22_n_692 ,mul_84_22_n_461 ,mul_84_22_n_517);
  and mul_84_22_g3367(mul_84_22_n_690 ,mul_84_22_n_470 ,mul_84_22_n_526);
  and mul_84_22_g3368(mul_84_22_n_688 ,mul_84_22_n_472 ,mul_84_22_n_562);
  or mul_84_22_g3369(mul_84_22_n_687 ,mul_84_22_n_495 ,mul_84_22_n_587);
  and mul_84_22_g3370(mul_84_22_n_685 ,mul_84_22_n_412 ,mul_84_22_n_563);
  or mul_84_22_g3371(mul_84_22_n_684 ,mul_84_22_n_499 ,mul_84_22_n_585);
  and mul_84_22_g3372(mul_84_22_n_682 ,mul_84_22_n_441 ,mul_84_22_n_568);
  or mul_84_22_g3373(mul_84_22_n_681 ,mul_84_22_n_491 ,mul_84_22_n_582);
  or mul_84_22_g3374(mul_84_22_n_679 ,mul_84_22_n_501 ,mul_84_22_n_589);
  and mul_84_22_g3375(mul_84_22_n_678 ,mul_84_22_n_471 ,mul_84_22_n_528);
  and mul_84_22_g3376(mul_84_22_n_677 ,mul_84_22_n_440 ,mul_84_22_n_567);
  and mul_84_22_g3377(mul_84_22_n_675 ,mul_84_22_n_464 ,mul_84_22_n_529);
  and mul_84_22_g3378(mul_84_22_n_674 ,mul_84_22_n_467 ,mul_84_22_n_538);
  and mul_84_22_g3379(mul_84_22_n_673 ,mul_84_22_n_443 ,mul_84_22_n_555);
  and mul_84_22_g3380(mul_84_22_n_672 ,mul_84_22_n_459 ,mul_84_22_n_521);
  or mul_84_22_g3381(mul_84_22_n_670 ,mul_84_22_n_492 ,mul_84_22_n_579);
  and mul_84_22_g3382(mul_84_22_n_669 ,mul_84_22_n_434 ,mul_84_22_n_514);
  and mul_84_22_g3383(mul_84_22_n_668 ,mul_84_22_n_462 ,mul_84_22_n_535);
  and mul_84_22_g3384(mul_84_22_n_667 ,mul_84_22_n_473 ,mul_84_22_n_524);
  and mul_84_22_g3385(mul_84_22_n_666 ,mul_84_22_n_436 ,mul_84_22_n_533);
  and mul_84_22_g3386(mul_84_22_n_665 ,mul_84_22_n_432 ,mul_84_22_n_552);
  and mul_84_22_g3387(mul_84_22_n_664 ,mul_84_22_n_423 ,mul_84_22_n_523);
  and mul_84_22_g3388(mul_84_22_n_663 ,mul_84_22_n_426 ,mul_84_22_n_518);
  or mul_84_22_g3389(mul_84_22_n_661 ,mul_84_22_n_494 ,mul_84_22_n_540);
  and mul_84_22_g3390(mul_84_22_n_659 ,mul_84_22_n_433 ,mul_84_22_n_558);
  and mul_84_22_g3391(mul_84_22_n_657 ,mul_84_22_n_431 ,mul_84_22_n_531);
  or mul_84_22_g3392(mul_84_22_n_656 ,mul_84_22_n_454 ,mul_84_22_n_504);
  and mul_84_22_g3393(mul_84_22_n_654 ,mul_84_22_n_418 ,mul_84_22_n_527);
  or mul_84_22_g3394(mul_84_22_n_653 ,mul_84_22_n_452 ,mul_84_22_n_505);
  and mul_84_22_g3395(mul_84_22_n_651 ,mul_84_22_n_413 ,mul_84_22_n_532);
  or mul_84_22_g3396(mul_84_22_n_650 ,mul_84_22_n_493 ,mul_84_22_n_577);
  and mul_84_22_g3397(mul_84_22_n_649 ,mul_84_22_n_425 ,mul_84_22_n_559);
  or mul_84_22_g3398(mul_84_22_n_648 ,mul_84_22_n_498 ,mul_84_22_n_584);
  not mul_84_22_g3399(mul_84_22_n_644 ,mul_84_22_n_643);
  not mul_84_22_g3400(mul_84_22_n_640 ,mul_84_22_n_639);
  not mul_84_22_g3401(mul_84_22_n_637 ,mul_84_22_n_636);
  not mul_84_22_g3402(mul_84_22_n_635 ,mul_84_22_n_634);
  not mul_84_22_g3403(mul_84_22_n_626 ,mul_84_22_n_625);
  not mul_84_22_g3404(mul_84_22_n_620 ,mul_84_22_n_619);
  not mul_84_22_g3405(mul_84_22_n_617 ,mul_84_22_n_618);
  not mul_84_22_g3406(mul_84_22_n_615 ,mul_84_22_n_616);
  not mul_84_22_g3407(mul_84_22_n_613 ,mul_84_22_n_614);
  not mul_84_22_g3408(mul_84_22_n_603 ,mul_84_22_n_604);
  not mul_84_22_g3409(mul_84_22_n_601 ,mul_84_22_n_602);
  not mul_84_22_g3411(mul_84_22_n_595 ,mul_84_22_n_596);
  not mul_84_22_g3412(mul_84_22_n_593 ,mul_84_22_n_594);
  nor mul_84_22_g3413(mul_84_22_n_591 ,mul_84_22_n_486 ,mul_84_22_n_574);
  or mul_84_22_g3414(mul_84_22_n_645 ,mul_84_22_n_324 ,mul_84_22_n_507);
  and mul_84_22_g3415(mul_84_22_n_643 ,mul_84_22_n_488 ,mul_84_22_n_571);
  and mul_84_22_g3416(mul_84_22_n_642 ,mul_84_22_n_478 ,mul_84_22_n_570);
  and mul_84_22_g3417(mul_84_22_n_641 ,mul_84_22_n_481 ,mul_84_22_n_572);
  and mul_84_22_g3418(mul_84_22_n_639 ,mul_84_22_n_421 ,mul_84_22_n_575);
  or mul_84_22_g3419(mul_84_22_n_638 ,mul_84_22_n_490 ,mul_84_22_n_581);
  and mul_84_22_g3420(mul_84_22_n_636 ,mul_84_22_n_428 ,mul_84_22_n_512);
  and mul_84_22_g3421(mul_84_22_n_634 ,mul_84_22_n_468 ,mul_84_22_n_539);
  and mul_84_22_g3422(mul_84_22_n_633 ,mul_84_22_n_430 ,mul_84_22_n_509);
  and mul_84_22_g3423(mul_84_22_n_632 ,mul_84_22_n_484 ,mul_84_22_n_590);
  and mul_84_22_g3424(mul_84_22_n_631 ,mul_84_22_n_437 ,mul_84_22_n_520);
  and mul_84_22_g3425(mul_84_22_n_630 ,mul_84_22_n_325 ,mul_84_22_n_556);
  and mul_84_22_g3426(mul_84_22_n_629 ,mul_84_22_n_427 ,mul_84_22_n_519);
  or mul_84_22_g3427(mul_84_22_n_628 ,mul_84_22_n_496 ,mul_84_22_n_569);
  and mul_84_22_g3428(mul_84_22_n_627 ,mul_84_22_n_482 ,mul_84_22_n_566);
  and mul_84_22_g3429(mul_84_22_n_625 ,mul_84_22_n_479 ,mul_84_22_n_560);
  and mul_84_22_g3430(mul_84_22_n_624 ,mul_84_22_n_477 ,mul_84_22_n_576);
  and mul_84_22_g3431(mul_84_22_n_623 ,mul_84_22_n_475 ,mul_84_22_n_557);
  and mul_84_22_g3432(mul_84_22_n_622 ,mul_84_22_n_474 ,mul_84_22_n_553);
  and mul_84_22_g3433(mul_84_22_n_621 ,mul_84_22_n_487 ,mul_84_22_n_541);
  or mul_84_22_g3434(mul_84_22_n_619 ,mul_84_22_n_503 ,mul_84_22_n_583);
  and mul_84_22_g3435(mul_84_22_n_618 ,mul_84_22_n_416 ,mul_84_22_n_530);
  and mul_84_22_g3436(mul_84_22_n_616 ,mul_84_22_n_420 ,mul_84_22_n_542);
  and mul_84_22_g3437(mul_84_22_n_614 ,mul_84_22_n_458 ,mul_84_22_n_564);
  and mul_84_22_g3438(mul_84_22_n_612 ,mul_84_22_n_455 ,mul_84_22_n_543);
  and mul_84_22_g3439(mul_84_22_n_611 ,mul_84_22_n_453 ,mul_84_22_n_515);
  and mul_84_22_g3440(mul_84_22_n_610 ,mul_84_22_n_438 ,mul_84_22_n_534);
  and mul_84_22_g3441(mul_84_22_n_609 ,mul_84_22_n_469 ,mul_84_22_n_513);
  and mul_84_22_g3442(mul_84_22_n_608 ,mul_84_22_n_442 ,mul_84_22_n_537);
  and mul_84_22_g3443(mul_84_22_n_607 ,mul_84_22_n_419 ,mul_84_22_n_510);
  and mul_84_22_g3444(mul_84_22_n_606 ,mul_84_22_n_463 ,mul_84_22_n_516);
  and mul_84_22_g3445(mul_84_22_n_605 ,mul_84_22_n_465 ,mul_84_22_n_511);
  or mul_84_22_g3446(mul_84_22_n_604 ,mul_84_22_n_489 ,mul_84_22_n_586);
  and mul_84_22_g3447(mul_84_22_n_602 ,mul_84_22_n_485 ,mul_84_22_n_522);
  and mul_84_22_g3448(mul_84_22_n_600 ,mul_84_22_n_435 ,mul_84_22_n_548);
  and mul_84_22_g3449(mul_84_22_n_599 ,mul_84_22_n_483 ,mul_84_22_n_551);
  and mul_84_22_g3450(mul_84_22_n_598 ,mul_84_22_n_476 ,mul_84_22_n_554);
  and mul_84_22_g3451(mul_84_22_n_597 ,mul_84_22_n_417 ,mul_84_22_n_550);
  and mul_84_22_g3452(mul_84_22_n_596 ,mul_84_22_n_480 ,mul_84_22_n_549);
  and mul_84_22_g3453(mul_84_22_n_594 ,mul_84_22_n_411 ,mul_84_22_n_525);
  and mul_84_22_g3454(mul_84_22_n_592 ,mul_84_22_n_414 ,mul_84_22_n_508);
  or mul_84_22_g3455(mul_84_22_n_590 ,mul_84_22_n_353 ,mul_84_22_n_66);
  and mul_84_22_g3456(mul_84_22_n_589 ,mul_84_22_n_140 ,mul_84_22_n_33);
  and mul_84_22_g3457(mul_84_22_n_588 ,mul_84_22_n_90 ,mul_84_22_n_45);
  and mul_84_22_g3458(mul_84_22_n_587 ,mul_84_22_n_132 ,mul_84_22_n_16);
  and mul_84_22_g3459(mul_84_22_n_586 ,mul_84_22_n_128 ,mul_84_22_n_33);
  and mul_84_22_g3460(mul_84_22_n_585 ,mul_84_22_n_110 ,mul_84_22_n_34);
  and mul_84_22_g3461(mul_84_22_n_584 ,mul_84_22_n_92 ,mul_84_22_n_46);
  and mul_84_22_g3462(mul_84_22_n_583 ,mul_84_22_n_142 ,mul_84_22_n_22);
  and mul_84_22_g3463(mul_84_22_n_582 ,mul_84_22_n_144 ,mul_84_22_n_21);
  and mul_84_22_g3464(mul_84_22_n_581 ,mul_84_22_n_134 ,mul_84_22_n_34);
  and mul_84_22_g3465(mul_84_22_n_580 ,mul_84_22_n_138 ,mul_84_22_n_21);
  and mul_84_22_g3466(mul_84_22_n_579 ,mul_84_22_n_120 ,mul_84_22_n_46);
  and mul_84_22_g3467(mul_84_22_n_578 ,mul_84_22_n_94 ,mul_84_22_n_45);
  and mul_84_22_g3468(mul_84_22_n_577 ,mul_84_22_n_126 ,mul_84_22_n_170);
  or mul_84_22_g3469(mul_84_22_n_576 ,mul_84_22_n_351 ,mul_84_22_n_76);
  or mul_84_22_g3470(mul_84_22_n_575 ,mul_84_22_n_328 ,mul_84_22_n_25);
  nor mul_84_22_g3471(mul_84_22_n_574 ,mul_84_22_n_76 ,mul_84_22_n_330);
  or mul_84_22_g3472(mul_84_22_n_573 ,mul_84_22_n_344 ,mul_84_22_n_58);
  or mul_84_22_g3473(mul_84_22_n_572 ,mul_84_22_n_338 ,mul_84_22_n_75);
  or mul_84_22_g3474(mul_84_22_n_571 ,mul_84_22_n_347 ,mul_84_22_n_40);
  or mul_84_22_g3475(mul_84_22_n_570 ,mul_84_22_n_365 ,mul_84_22_n_39);
  and mul_84_22_g3476(mul_84_22_n_569 ,mul_84_22_n_136 ,mul_84_22_n_22);
  or mul_84_22_g3477(mul_84_22_n_568 ,mul_84_22_n_362 ,mul_84_22_n_37);
  or mul_84_22_g3478(mul_84_22_n_567 ,mul_84_22_n_349 ,mul_84_22_n_57);
  or mul_84_22_g3479(mul_84_22_n_566 ,mul_84_22_n_360 ,mul_84_22_n_40);
  or mul_84_22_g3480(mul_84_22_n_565 ,mul_84_22_n_341 ,mul_84_22_n_81);
  or mul_84_22_g3481(mul_84_22_n_564 ,mul_84_22_n_346 ,mul_84_22_n_36);
  or mul_84_22_g3482(mul_84_22_n_563 ,mul_84_22_n_366 ,mul_84_22_n_25);
  or mul_84_22_g3483(mul_84_22_n_562 ,mul_84_22_n_354 ,mul_84_22_n_24);
  or mul_84_22_g3484(mul_84_22_n_561 ,mul_84_22_n_369 ,mul_84_22_n_24);
  or mul_84_22_g3485(mul_84_22_n_560 ,mul_84_22_n_350 ,mul_84_22_n_14);
  or mul_84_22_g3486(mul_84_22_n_559 ,mul_84_22_n_368 ,mul_84_22_n_37);
  or mul_84_22_g3487(mul_84_22_n_558 ,mul_84_22_n_345 ,mul_84_22_n_57);
  or mul_84_22_g3488(mul_84_22_n_557 ,mul_84_22_n_355 ,mul_84_22_n_88);
  or mul_84_22_g3489(mul_84_22_n_556 ,mul_84_22_n_364 ,mul_84_22_n_39);
  or mul_84_22_g3490(mul_84_22_n_555 ,mul_84_22_n_358 ,mul_84_22_n_81);
  or mul_84_22_g3491(mul_84_22_n_554 ,mul_84_22_n_352 ,mul_84_22_n_66);
  or mul_84_22_g3492(mul_84_22_n_553 ,mul_84_22_n_337 ,mul_84_22_n_75);
  or mul_84_22_g3493(mul_84_22_n_552 ,mul_84_22_n_343 ,mul_84_22_n_36);
  or mul_84_22_g3494(mul_84_22_n_551 ,mul_84_22_n_361 ,mul_84_22_n_67);
  or mul_84_22_g3495(mul_84_22_n_550 ,mul_84_22_n_359 ,mul_84_22_n_10);
  or mul_84_22_g3496(mul_84_22_n_549 ,mul_84_22_n_357 ,mul_84_22_n_87);
  or mul_84_22_g3497(mul_84_22_n_548 ,mul_84_22_n_342 ,mul_84_22_n_10);
  not mul_84_22_g3498(mul_84_22_n_545 ,mul_84_22_n_544);
  or mul_84_22_g3499(mul_84_22_n_543 ,mul_84_22_n_392 ,mul_84_22_n_49);
  or mul_84_22_g3500(mul_84_22_n_542 ,mul_84_22_n_356 ,mul_84_22_n_82);
  or mul_84_22_g3501(mul_84_22_n_541 ,mul_84_22_n_340 ,mul_84_22_n_87);
  and mul_84_22_g3502(mul_84_22_n_540 ,mul_84_22_n_165 ,mul_84_22_n_16);
  or mul_84_22_g3503(mul_84_22_n_539 ,mul_84_22_n_377 ,mul_84_22_n_31);
  or mul_84_22_g3504(mul_84_22_n_538 ,mul_84_22_n_388 ,mul_84_22_n_64);
  or mul_84_22_g3505(mul_84_22_n_537 ,mul_84_22_n_407 ,mul_84_22_n_28);
  or mul_84_22_g3506(mul_84_22_n_536 ,mul_84_22_n_370 ,mul_84_22_n_63);
  or mul_84_22_g3507(mul_84_22_n_535 ,mul_84_22_n_405 ,mul_84_22_n_61);
  or mul_84_22_g3508(mul_84_22_n_534 ,mul_84_22_n_404 ,mul_84_22_n_84);
  or mul_84_22_g3509(mul_84_22_n_533 ,mul_84_22_n_386 ,mul_84_22_n_27);
  or mul_84_22_g3510(mul_84_22_n_532 ,mul_84_22_n_399 ,mul_84_22_n_49);
  or mul_84_22_g3511(mul_84_22_n_531 ,mul_84_22_n_390 ,mul_84_22_n_52);
  or mul_84_22_g3512(mul_84_22_n_530 ,mul_84_22_n_339 ,mul_84_22_n_48);
  or mul_84_22_g3513(mul_84_22_n_529 ,mul_84_22_n_410 ,mul_84_22_n_60);
  or mul_84_22_g3514(mul_84_22_n_528 ,mul_84_22_n_385 ,mul_84_22_n_48);
  or mul_84_22_g3515(mul_84_22_n_527 ,mul_84_22_n_389 ,mul_84_22_n_78);
  or mul_84_22_g3516(mul_84_22_n_526 ,mul_84_22_n_408 ,mul_84_22_n_28);
  or mul_84_22_g3517(mul_84_22_n_525 ,mul_84_22_n_397 ,mul_84_22_n_63);
  or mul_84_22_g3518(mul_84_22_n_524 ,mul_84_22_n_395 ,mul_84_22_n_51);
  or mul_84_22_g3519(mul_84_22_n_523 ,mul_84_22_n_403 ,mul_84_22_n_84);
  or mul_84_22_g3520(mul_84_22_n_522 ,mul_84_22_n_348 ,mul_84_22_n_14);
  or mul_84_22_g3521(mul_84_22_n_521 ,mul_84_22_n_406 ,mul_84_22_n_31);
  or mul_84_22_g3522(mul_84_22_n_520 ,mul_84_22_n_396 ,mul_84_22_n_30);
  or mul_84_22_g3523(mul_84_22_n_519 ,mul_84_22_n_363 ,mul_84_22_n_30);
  or mul_84_22_g3524(mul_84_22_n_518 ,mul_84_22_n_391 ,mul_84_22_n_52);
  or mul_84_22_g3525(mul_84_22_n_517 ,mul_84_22_n_394 ,mul_84_22_n_60);
  or mul_84_22_g3526(mul_84_22_n_516 ,mul_84_22_n_400 ,mul_84_22_n_27);
  or mul_84_22_g3527(mul_84_22_n_515 ,mul_84_22_n_387 ,mul_84_22_n_78);
  or mul_84_22_g3528(mul_84_22_n_514 ,mul_84_22_n_384 ,mul_84_22_n_51);
  or mul_84_22_g3529(mul_84_22_n_513 ,mul_84_22_n_409 ,mul_84_22_n_8);
  or mul_84_22_g3530(mul_84_22_n_512 ,mul_84_22_n_393 ,mul_84_22_n_12);
  or mul_84_22_g3531(mul_84_22_n_511 ,mul_84_22_n_401 ,mul_84_22_n_12);
  or mul_84_22_g3532(mul_84_22_n_510 ,mul_84_22_n_367 ,mul_84_22_n_79);
  or mul_84_22_g3533(mul_84_22_n_509 ,mul_84_22_n_402 ,mul_84_22_n_8);
  or mul_84_22_g3534(mul_84_22_n_508 ,mul_84_22_n_398 ,mul_84_22_n_85);
  nor mul_84_22_g3535(mul_84_22_n_507 ,mul_84_22_n_67 ,mul_84_22_n_311);
  nor mul_84_22_g3536(mul_84_22_n_506 ,mul_84_22_n_58 ,mul_84_22_n_310);
  nor mul_84_22_g3537(mul_84_22_n_505 ,mul_84_22_n_61 ,mul_84_22_n_315);
  nor mul_84_22_g3538(mul_84_22_n_504 ,mul_84_22_n_64 ,mul_84_22_n_316);
  and mul_84_22_g3539(mul_84_22_n_547 ,in7[3] ,mul_84_22_n_439);
  and mul_84_22_g3540(mul_84_22_n_546 ,in7[5] ,mul_84_22_n_415);
  or mul_84_22_g3541(mul_84_22_n_544 ,mul_84_22_n_310 ,mul_84_22_n_424);
  and mul_84_22_g3542(mul_84_22_n_503 ,mul_84_22_n_134 ,mul_84_22_n_246);
  and mul_84_22_g3543(mul_84_22_n_502 ,mul_84_22_n_92 ,mul_84_22_n_236);
  and mul_84_22_g3544(mul_84_22_n_501 ,mul_84_22_n_136 ,mul_84_22_n_209);
  and mul_84_22_g3545(mul_84_22_n_500 ,mul_84_22_n_94 ,mul_84_22_n_237);
  and mul_84_22_g3546(mul_84_22_n_499 ,mul_84_22_n_140 ,mul_84_22_n_209);
  and mul_84_22_g3547(mul_84_22_n_498 ,mul_84_22_n_128 ,mul_84_22_n_210);
  and mul_84_22_g3548(mul_84_22_n_497 ,mul_84_22_n_252 ,mul_84_22_n_210);
  and mul_84_22_g3549(mul_84_22_n_496 ,mul_84_22_n_142 ,mul_84_22_n_237);
  and mul_84_22_g3550(mul_84_22_n_495 ,mul_84_22_n_126 ,mul_84_22_n_200);
  and mul_84_22_g3551(mul_84_22_n_494 ,mul_84_22_n_144 ,mul_84_22_n_199);
  and mul_84_22_g3552(mul_84_22_n_493 ,mul_84_22_n_138 ,mul_84_22_n_236);
  and mul_84_22_g3553(mul_84_22_n_492 ,mul_84_22_n_132 ,mul_84_22_n_246);
  and mul_84_22_g3554(mul_84_22_n_491 ,mul_84_22_n_110 ,mul_84_22_n_200);
  and mul_84_22_g3555(mul_84_22_n_490 ,mul_84_22_n_90 ,mul_84_22_n_245);
  and mul_84_22_g3556(mul_84_22_n_489 ,mul_84_22_n_120 ,mul_84_22_n_245);
  or mul_84_22_g3557(mul_84_22_n_488 ,mul_84_22_n_70 ,mul_84_22_n_338);
  or mul_84_22_g3558(mul_84_22_n_487 ,mul_84_22_n_42 ,mul_84_22_n_337);
  nor mul_84_22_g3559(mul_84_22_n_486 ,mul_84_22_n_73 ,mul_84_22_n_365);
  or mul_84_22_g3560(mul_84_22_n_485 ,mul_84_22_n_54 ,mul_84_22_n_357);
  or mul_84_22_g3561(mul_84_22_n_484 ,mul_84_22_n_72 ,mul_84_22_n_340);
  or mul_84_22_g3562(mul_84_22_n_483 ,mul_84_22_n_69 ,mul_84_22_n_352);
  or mul_84_22_g3563(mul_84_22_n_482 ,mul_84_22_n_43 ,mul_84_22_n_353);
  or mul_84_22_g3564(mul_84_22_n_481 ,mul_84_22_n_55 ,mul_84_22_n_348);
  or mul_84_22_g3565(mul_84_22_n_480 ,mul_84_22_n_72 ,mul_84_22_n_361);
  or mul_84_22_g3566(mul_84_22_n_479 ,mul_84_22_n_69 ,mul_84_22_n_360);
  or mul_84_22_g3567(mul_84_22_n_478 ,mul_84_22_n_42 ,mul_84_22_n_347);
  or mul_84_22_g3568(mul_84_22_n_477 ,mul_84_22_n_54 ,mul_84_22_n_364);
  or mul_84_22_g3569(mul_84_22_n_476 ,mul_84_22_n_55 ,mul_84_22_n_355);
  or mul_84_22_g3570(mul_84_22_n_475 ,mul_84_22_n_43 ,mul_84_22_n_350);
  or mul_84_22_g3571(mul_84_22_n_474 ,mul_84_22_n_73 ,mul_84_22_n_351);
  or mul_84_22_g3572(mul_84_22_n_473 ,mul_84_22_n_406 ,mul_84_22_n_224);
  or mul_84_22_g3573(mul_84_22_n_472 ,mul_84_22_n_344 ,mul_84_22_n_215);
  or mul_84_22_g3574(mul_84_22_n_471 ,mul_84_22_n_404 ,mul_84_22_n_239);
  or mul_84_22_g3575(mul_84_22_n_470 ,mul_84_22_n_385 ,mul_84_22_n_206);
  or mul_84_22_g3576(mul_84_22_n_469 ,mul_84_22_n_400 ,mul_84_22_n_206);
  or mul_84_22_g3577(mul_84_22_n_468 ,mul_84_22_n_401 ,mul_84_22_n_233);
  or mul_84_22_g3578(mul_84_22_n_467 ,mul_84_22_n_408 ,mul_84_22_n_240);
  or mul_84_22_g3579(mul_84_22_n_466 ,mul_84_22_n_343 ,mul_84_22_n_218);
  or mul_84_22_g3580(mul_84_22_n_465 ,mul_84_22_n_384 ,mul_84_22_n_233);
  or mul_84_22_g3581(mul_84_22_n_464 ,mul_84_22_n_405 ,mul_84_22_n_225);
  or mul_84_22_g3582(mul_84_22_n_463 ,mul_84_22_n_388 ,mul_84_22_n_243);
  or mul_84_22_g3583(mul_84_22_n_462 ,mul_84_22_n_393 ,mul_84_22_n_228);
  or mul_84_22_g3584(mul_84_22_n_461 ,mul_84_22_n_387 ,mul_84_22_n_224);
  or mul_84_22_g3585(mul_84_22_n_460 ,mul_84_22_n_359 ,mul_84_22_n_218);
  or mul_84_22_g3586(mul_84_22_n_459 ,mul_84_22_n_367 ,mul_84_22_n_227);
  not mul_84_22_g3587(mul_84_22_n_458 ,mul_84_22_n_457);
  not mul_84_22_g3588(mul_84_22_n_455 ,mul_84_22_n_454);
  not mul_84_22_g3589(mul_84_22_n_453 ,mul_84_22_n_452);
  or mul_84_22_g3590(mul_84_22_n_443 ,mul_84_22_n_345 ,mul_84_22_n_216);
  or mul_84_22_g3591(mul_84_22_n_442 ,mul_84_22_n_403 ,mul_84_22_n_239);
  or mul_84_22_g3592(mul_84_22_n_441 ,mul_84_22_n_369 ,mul_84_22_n_249);
  or mul_84_22_g3593(mul_84_22_n_440 ,mul_84_22_n_368 ,mul_84_22_n_215);
  or mul_84_22_g3594(mul_84_22_n_439 ,mul_84_22_n_321 ,mul_84_22_n_376);
  or mul_84_22_g3595(mul_84_22_n_438 ,mul_84_22_n_398 ,mul_84_22_n_242);
  or mul_84_22_g3596(mul_84_22_n_437 ,mul_84_22_n_389 ,mul_84_22_n_230);
  or mul_84_22_g3597(mul_84_22_n_436 ,mul_84_22_n_402 ,mul_84_22_n_212);
  or mul_84_22_g3598(mul_84_22_n_435 ,mul_84_22_n_354 ,mul_84_22_n_248);
  or mul_84_22_g3599(mul_84_22_n_434 ,mul_84_22_n_396 ,mul_84_22_n_230);
  or mul_84_22_g3600(mul_84_22_n_433 ,mul_84_22_n_366 ,mul_84_22_n_221);
  or mul_84_22_g3601(mul_84_22_n_432 ,mul_84_22_n_341 ,mul_84_22_n_221);
  or mul_84_22_g3602(mul_84_22_n_431 ,mul_84_22_n_394 ,mul_84_22_n_227);
  or mul_84_22_g3603(mul_84_22_n_430 ,mul_84_22_n_392 ,mul_84_22_n_212);
  or mul_84_22_g3604(mul_84_22_n_429 ,mul_84_22_n_349 ,mul_84_22_n_248);
  or mul_84_22_g3605(mul_84_22_n_428 ,mul_84_22_n_363 ,mul_84_22_n_234);
  or mul_84_22_g3606(mul_84_22_n_427 ,mul_84_22_n_395 ,mul_84_22_n_228);
  or mul_84_22_g3607(mul_84_22_n_426 ,mul_84_22_n_410 ,mul_84_22_n_231);
  or mul_84_22_g3608(mul_84_22_n_425 ,mul_84_22_n_356 ,mul_84_22_n_219);
  nor mul_84_22_g3609(mul_84_22_n_424 ,mul_84_22_n_320 ,mul_84_22_n_374);
  or mul_84_22_g3610(mul_84_22_n_423 ,mul_84_22_n_386 ,mul_84_22_n_242);
  or mul_84_22_g3611(mul_84_22_n_422 ,mul_84_22_n_399 ,mul_84_22_n_207);
  or mul_84_22_g3612(mul_84_22_n_421 ,mul_84_22_n_358 ,mul_84_22_n_249);
  or mul_84_22_g3613(mul_84_22_n_420 ,mul_84_22_n_346 ,mul_84_22_n_222);
  or mul_84_22_g3614(mul_84_22_n_419 ,mul_84_22_n_390 ,mul_84_22_n_225);
  or mul_84_22_g3615(mul_84_22_n_418 ,mul_84_22_n_391 ,mul_84_22_n_234);
  or mul_84_22_g3616(mul_84_22_n_417 ,mul_84_22_n_342 ,mul_84_22_n_216);
  or mul_84_22_g3617(mul_84_22_n_416 ,mul_84_22_n_397 ,mul_84_22_n_243);
  or mul_84_22_g3618(mul_84_22_n_415 ,mul_84_22_n_326 ,mul_84_22_n_373);
  or mul_84_22_g3619(mul_84_22_n_414 ,mul_84_22_n_407 ,mul_84_22_n_213);
  or mul_84_22_g3620(mul_84_22_n_413 ,mul_84_22_n_339 ,mul_84_22_n_240);
  or mul_84_22_g3621(mul_84_22_n_412 ,mul_84_22_n_362 ,mul_84_22_n_219);
  or mul_84_22_g3622(mul_84_22_n_411 ,mul_84_22_n_409 ,mul_84_22_n_207);
  and mul_84_22_g3623(mul_84_22_n_457 ,in7[7] ,mul_84_22_n_150);
  or mul_84_22_g3624(mul_84_22_n_456 ,mul_84_22_n_159 ,mul_84_22_n_213);
  and mul_84_22_g3625(mul_84_22_n_454 ,in7[3] ,mul_84_22_n_154);
  and mul_84_22_g3626(mul_84_22_n_452 ,in7[5] ,mul_84_22_n_152);
  or mul_84_22_g3627(mul_84_22_n_451 ,mul_84_22_n_163 ,mul_84_22_n_231);
  or mul_84_22_g3628(mul_84_22_n_450 ,mul_84_22_n_162 ,mul_84_22_n_222);
  or mul_84_22_g3629(mul_84_22_n_449 ,mul_84_22_n_162 ,mul_84_22_n_148);
  and mul_84_22_g3630(mul_84_22_n_448 ,in7[8] ,mul_84_22_n_147);
  or mul_84_22_g3631(mul_84_22_n_447 ,mul_84_22_n_371 ,mul_84_22_n_151);
  or mul_84_22_g3632(mul_84_22_n_446 ,in7[0] ,mul_84_22_n_375);
  or mul_84_22_g3633(mul_84_22_n_445 ,mul_84_22_n_329 ,mul_84_22_n_149);
  or mul_84_22_g3634(mul_84_22_n_444 ,mul_84_22_n_372 ,mul_84_22_n_153);
  not mul_84_22_g3635(mul_84_22_n_383 ,mul_84_22_n_152);
  not mul_84_22_g3636(mul_84_22_n_382 ,mul_84_22_n_151);
  not mul_84_22_g3639(mul_84_22_n_380 ,mul_84_22_n_150);
  not mul_84_22_g3640(mul_84_22_n_379 ,mul_84_22_n_149);
  xnor mul_84_22_g3643(mul_84_22_n_377 ,mul_84_22_n_18 ,in7[5]);
  and mul_84_22_g3644(mul_84_22_n_376 ,mul_84_22_n_202 ,mul_84_22_n_322);
  and mul_84_22_g3646(mul_84_22_n_374 ,mul_84_22_n_315 ,mul_84_22_n_319);
  and mul_84_22_g3647(mul_84_22_n_373 ,mul_84_22_n_316 ,mul_84_22_n_323);
  xnor mul_84_22_g3648(mul_84_22_n_372 ,in7[3] ,in7[2]);
  xnor mul_84_22_g3649(mul_84_22_n_371 ,in7[5] ,in7[4]);
  xnor mul_84_22_g3650(mul_84_22_n_370 ,mul_84_22_n_18 ,in7[3]);
  xnor mul_84_22_g3651(mul_84_22_n_410 ,mul_84_22_n_260 ,in7[5]);
  xnor mul_84_22_g3652(mul_84_22_n_409 ,mul_84_22_n_281 ,in7[3]);
  xnor mul_84_22_g3653(mul_84_22_n_408 ,mul_84_22_n_287 ,in7[3]);
  xnor mul_84_22_g3654(mul_84_22_n_407 ,mul_84_22_n_269 ,in7[3]);
  xnor mul_84_22_g3655(mul_84_22_n_406 ,mul_84_22_n_270 ,in7[5]);
  xnor mul_84_22_g3656(mul_84_22_n_405 ,mul_84_22_n_288 ,in7[5]);
  xnor mul_84_22_g3657(mul_84_22_n_404 ,mul_84_22_n_278 ,in7[3]);
  xnor mul_84_22_g3658(mul_84_22_n_403 ,mul_84_22_n_263 ,in7[3]);
  xnor mul_84_22_g3659(mul_84_22_n_402 ,mul_84_22_n_254 ,in7[3]);
  xnor mul_84_22_g3660(mul_84_22_n_401 ,mul_84_22_n_290 ,in7[5]);
  xnor mul_84_22_g3661(mul_84_22_n_400 ,mul_84_22_n_272 ,in7[3]);
  xnor mul_84_22_g3662(mul_84_22_n_399 ,mul_84_22_n_291 ,in7[3]);
  xnor mul_84_22_g3663(mul_84_22_n_398 ,mul_84_22_n_275 ,in7[3]);
  xnor mul_84_22_g3664(mul_84_22_n_397 ,mul_84_22_n_293 ,in7[3]);
  xnor mul_84_22_g3665(mul_84_22_n_396 ,mul_84_22_n_294 ,in7[5]);
  xnor mul_84_22_g3666(mul_84_22_n_395 ,mul_84_22_n_276 ,in7[5]);
  xnor mul_84_22_g3667(mul_84_22_n_394 ,mul_84_22_n_255 ,in7[5]);
  xnor mul_84_22_g3668(mul_84_22_n_393 ,mul_84_22_n_284 ,in7[5]);
  xnor mul_84_22_g3669(mul_84_22_n_392 ,mul_84_22_n_251 ,in7[3]);
  xnor mul_84_22_g3670(mul_84_22_n_391 ,mul_84_22_n_273 ,in7[5]);
  xnor mul_84_22_g3671(mul_84_22_n_390 ,mul_84_22_n_257 ,in7[5]);
  xnor mul_84_22_g3672(mul_84_22_n_389 ,mul_84_22_n_282 ,in7[5]);
  xnor mul_84_22_g3673(mul_84_22_n_388 ,mul_84_22_n_261 ,in7[3]);
  xnor mul_84_22_g3674(mul_84_22_n_387 ,mul_84_22_n_122 ,in7[5]);
  xnor mul_84_22_g3675(mul_84_22_n_386 ,mul_84_22_n_258 ,in7[3]);
  xnor mul_84_22_g3676(mul_84_22_n_385 ,mul_84_22_n_285 ,in7[3]);
  xnor mul_84_22_g3677(mul_84_22_n_384 ,mul_84_22_n_266 ,in7[5]);
  xnor mul_84_22_g3678(mul_84_22_n_381 ,mul_84_22_n_316 ,in7[4]);
  xnor mul_84_22_g3679(mul_84_22_n_378 ,mul_84_22_n_315 ,in7[6]);
  not mul_84_22_g3680(mul_84_22_n_336 ,mul_84_22_n_148);
  not mul_84_22_g3681(mul_84_22_n_335 ,mul_84_22_n_147);
  not mul_84_22_g3684(mul_84_22_n_333 ,mul_84_22_n_154);
  not mul_84_22_g3685(mul_84_22_n_332 ,mul_84_22_n_153);
  xnor mul_84_22_g3689(mul_84_22_n_329 ,in7[7] ,in7[6]);
  xnor mul_84_22_g3690(mul_84_22_n_328 ,mul_84_22_n_168 ,in7[7]);
  xnor mul_84_22_g3691(mul_84_22_n_369 ,mul_84_22_n_98 ,in7[7]);
  xnor mul_84_22_g3692(mul_84_22_n_368 ,mul_84_22_n_100 ,in7[7]);
  xnor mul_84_22_g3693(mul_84_22_n_367 ,mul_84_22_n_264 ,in7[5]);
  xnor mul_84_22_g3694(mul_84_22_n_366 ,mul_84_22_n_112 ,in7[7]);
  xnor mul_84_22_g3695(mul_84_22_n_365 ,mul_84_22_n_114 ,in7[1]);
  xnor mul_84_22_g3696(mul_84_22_n_364 ,mul_84_22_n_251 ,in7[1]);
  xnor mul_84_22_g3697(mul_84_22_n_363 ,mul_84_22_n_279 ,in7[5]);
  xnor mul_84_22_g3698(mul_84_22_n_362 ,mul_84_22_n_146 ,in7[7]);
  xnor mul_84_22_g3699(mul_84_22_n_361 ,mul_84_22_n_124 ,in7[1]);
  xnor mul_84_22_g3700(mul_84_22_n_360 ,mul_84_22_n_102 ,in7[1]);
  xnor mul_84_22_g3701(mul_84_22_n_359 ,mul_84_22_n_124 ,in7[7]);
  xnor mul_84_22_g3702(mul_84_22_n_358 ,mul_84_22_n_114 ,in7[7]);
  xnor mul_84_22_g3703(mul_84_22_n_357 ,mul_84_22_n_98 ,in7[1]);
  xnor mul_84_22_g3704(mul_84_22_n_356 ,mul_84_22_n_118 ,in7[7]);
  xnor mul_84_22_g3705(mul_84_22_n_355 ,mul_84_22_n_108 ,in7[1]);
  xnor mul_84_22_g3706(mul_84_22_n_354 ,mul_84_22_n_108 ,in7[7]);
  xnor mul_84_22_g3707(mul_84_22_n_353 ,mul_84_22_n_106 ,in7[1]);
  xnor mul_84_22_g3708(mul_84_22_n_352 ,mul_84_22_n_96 ,in7[1]);
  xnor mul_84_22_g3709(mul_84_22_n_351 ,mul_84_22_n_118 ,in7[1]);
  xnor mul_84_22_g3710(mul_84_22_n_350 ,mul_84_22_n_104 ,in7[1]);
  xnor mul_84_22_g3711(mul_84_22_n_349 ,mul_84_22_n_116 ,in7[7]);
  xnor mul_84_22_g3712(mul_84_22_n_348 ,mul_84_22_n_146 ,in7[1]);
  xnor mul_84_22_g3713(mul_84_22_n_347 ,mul_84_22_n_267 ,in7[1]);
  xnor mul_84_22_g3714(mul_84_22_n_346 ,mul_84_22_n_122 ,in7[7]);
  xnor mul_84_22_g3715(mul_84_22_n_345 ,mul_84_22_n_130 ,in7[7]);
  xnor mul_84_22_g3716(mul_84_22_n_344 ,mul_84_22_n_104 ,in7[7]);
  xnor mul_84_22_g3717(mul_84_22_n_343 ,mul_84_22_n_102 ,in7[7]);
  xnor mul_84_22_g3718(mul_84_22_n_342 ,mul_84_22_n_96 ,in7[7]);
  xnor mul_84_22_g3719(mul_84_22_n_341 ,mul_84_22_n_106 ,in7[7]);
  xnor mul_84_22_g3720(mul_84_22_n_340 ,mul_84_22_n_116 ,in7[1]);
  xnor mul_84_22_g3721(mul_84_22_n_339 ,mul_84_22_n_130 ,in7[3]);
  xnor mul_84_22_g3722(mul_84_22_n_338 ,mul_84_22_n_112 ,in7[1]);
  xnor mul_84_22_g3723(mul_84_22_n_337 ,mul_84_22_n_100 ,in7[1]);
  xnor mul_84_22_g3724(mul_84_22_n_334 ,in7[8] ,in7[7]);
  xnor mul_84_22_g3725(mul_84_22_n_331 ,mul_84_22_n_202 ,in7[2]);
  nor mul_84_22_g3726(mul_84_22_n_327 ,mul_84_22_n_70 ,mul_84_22_n_163);
  nor mul_84_22_g3727(mul_84_22_n_326 ,mul_84_22_n_166 ,in7[4]);
  not mul_84_22_g3728(mul_84_22_n_325 ,mul_84_22_n_324);
  and mul_84_22_g3729(mul_84_22_n_324 ,in7[1] ,in7[0]);
  or mul_84_22_g3730(mul_84_22_n_323 ,mul_84_22_n_159 ,mul_84_22_n_313);
  or mul_84_22_g3731(mul_84_22_n_322 ,mul_84_22_n_160 ,mul_84_22_n_318);
  nor mul_84_22_g3732(mul_84_22_n_321 ,mul_84_22_n_19 ,in7[2]);
  nor mul_84_22_g3733(mul_84_22_n_320 ,mul_84_22_n_168 ,in7[6]);
  or mul_84_22_g3734(mul_84_22_n_319 ,mul_84_22_n_160 ,mul_84_22_n_314);
  not mul_84_22_g3735(mul_84_22_n_318 ,in7[2]);
  not mul_84_22_g3736(mul_84_22_n_317 ,in7[0]);
  not mul_84_22_g3737(mul_84_22_n_316 ,in7[3]);
  not mul_84_22_g3738(mul_84_22_n_315 ,in7[5]);
  not mul_84_22_g3739(mul_84_22_n_314 ,in7[6]);
  not mul_84_22_g3740(mul_84_22_n_313 ,in7[4]);
  not mul_84_22_g3741(mul_84_22_n_312 ,mul_84_22_n_165);
  not mul_84_22_g3742(mul_84_22_n_311 ,in7[1]);
  not mul_84_22_g3743(mul_84_22_n_310 ,in7[7]);
  not mul_84_22_drc_bufs3784(mul_84_22_n_297 ,mul_84_22_n_295);
  not mul_84_22_drc_bufs3785(mul_84_22_n_296 ,mul_84_22_n_295);
  not mul_84_22_drc_bufs3786(mul_84_22_n_295 ,n_191);
  not mul_84_22_drc_bufs3814(mul_84_22_n_294 ,mul_84_22_n_292);
  not mul_84_22_drc_bufs3815(mul_84_22_n_293 ,mul_84_22_n_292);
  not mul_84_22_drc_bufs3816(mul_84_22_n_292 ,n_194);
  not mul_84_22_drc_bufs3818(mul_84_22_n_291 ,mul_84_22_n_289);
  not mul_84_22_drc_bufs3819(mul_84_22_n_290 ,mul_84_22_n_289);
  not mul_84_22_drc_bufs3820(mul_84_22_n_289 ,n_192);
  not mul_84_22_drc_bufs3822(mul_84_22_n_288 ,mul_84_22_n_286);
  not mul_84_22_drc_bufs3823(mul_84_22_n_287 ,mul_84_22_n_286);
  not mul_84_22_drc_bufs3824(mul_84_22_n_286 ,n_198);
  not mul_84_22_drc_bufs3826(mul_84_22_n_285 ,mul_84_22_n_283);
  not mul_84_22_drc_bufs3827(mul_84_22_n_284 ,mul_84_22_n_283);
  not mul_84_22_drc_bufs3828(mul_84_22_n_283 ,n_199);
  not mul_84_22_drc_bufs3830(mul_84_22_n_282 ,mul_84_22_n_280);
  not mul_84_22_drc_bufs3831(mul_84_22_n_281 ,mul_84_22_n_280);
  not mul_84_22_drc_bufs3832(mul_84_22_n_280 ,n_195);
  not mul_84_22_drc_bufs3834(mul_84_22_n_279 ,mul_84_22_n_277);
  not mul_84_22_drc_bufs3835(mul_84_22_n_278 ,mul_84_22_n_277);
  not mul_84_22_drc_bufs3836(mul_84_22_n_277 ,n_200);
  not mul_84_22_drc_bufs3838(mul_84_22_n_276 ,mul_84_22_n_274);
  not mul_84_22_drc_bufs3839(mul_84_22_n_275 ,mul_84_22_n_274);
  not mul_84_22_drc_bufs3840(mul_84_22_n_274 ,n_201);
  not mul_84_22_drc_bufs3842(mul_84_22_n_273 ,mul_84_22_n_271);
  not mul_84_22_drc_bufs3843(mul_84_22_n_272 ,mul_84_22_n_271);
  not mul_84_22_drc_bufs3844(mul_84_22_n_271 ,n_196);
  not mul_84_22_drc_bufs3846(mul_84_22_n_270 ,mul_84_22_n_268);
  not mul_84_22_drc_bufs3847(mul_84_22_n_269 ,mul_84_22_n_268);
  not mul_84_22_drc_bufs3848(mul_84_22_n_268 ,n_202);
  not mul_84_22_drc_bufs3850(mul_84_22_n_267 ,mul_84_22_n_265);
  not mul_84_22_drc_bufs3851(mul_84_22_n_266 ,mul_84_22_n_265);
  not mul_84_22_drc_bufs3852(mul_84_22_n_265 ,n_193);
  not mul_84_22_drc_bufs3854(mul_84_22_n_264 ,mul_84_22_n_262);
  not mul_84_22_drc_bufs3855(mul_84_22_n_263 ,mul_84_22_n_262);
  not mul_84_22_drc_bufs3856(mul_84_22_n_262 ,n_203);
  not mul_84_22_drc_bufs3858(mul_84_22_n_261 ,mul_84_22_n_259);
  not mul_84_22_drc_bufs3859(mul_84_22_n_260 ,mul_84_22_n_259);
  not mul_84_22_drc_bufs3860(mul_84_22_n_259 ,n_197);
  not mul_84_22_drc_bufs3862(mul_84_22_n_258 ,mul_84_22_n_256);
  not mul_84_22_drc_bufs3863(mul_84_22_n_257 ,mul_84_22_n_256);
  not mul_84_22_drc_bufs3864(mul_84_22_n_256 ,n_204);
  not mul_84_22_drc_bufs3866(mul_84_22_n_255 ,mul_84_22_n_253);
  not mul_84_22_drc_bufs3867(mul_84_22_n_254 ,mul_84_22_n_253);
  not mul_84_22_drc_bufs3868(mul_84_22_n_253 ,n_205);
  not mul_84_22_drc_bufs3870(mul_84_22_n_252 ,mul_84_22_n_250);
  not mul_84_22_drc_bufs3871(mul_84_22_n_251 ,mul_84_22_n_250);
  not mul_84_22_drc_bufs3872(mul_84_22_n_250 ,n_206);
  not mul_84_22_drc_bufs3874(mul_84_22_n_249 ,mul_84_22_n_247);
  not mul_84_22_drc_bufs3875(mul_84_22_n_248 ,mul_84_22_n_247);
  not mul_84_22_drc_bufs3876(mul_84_22_n_247 ,mul_84_22_n_303);
  not mul_84_22_drc_bufs3878(mul_84_22_n_246 ,mul_84_22_n_244);
  not mul_84_22_drc_bufs3879(mul_84_22_n_245 ,mul_84_22_n_244);
  not mul_84_22_drc_bufs3880(mul_84_22_n_244 ,mul_84_22_n_335);
  not mul_84_22_drc_bufs3882(mul_84_22_n_243 ,mul_84_22_n_241);
  not mul_84_22_drc_bufs3883(mul_84_22_n_242 ,mul_84_22_n_241);
  not mul_84_22_drc_bufs3884(mul_84_22_n_241 ,mul_84_22_n_299);
  not mul_84_22_drc_bufs3886(mul_84_22_n_240 ,mul_84_22_n_238);
  not mul_84_22_drc_bufs3887(mul_84_22_n_239 ,mul_84_22_n_238);
  not mul_84_22_drc_bufs3888(mul_84_22_n_238 ,mul_84_22_n_298);
  not mul_84_22_drc_bufs3890(mul_84_22_n_237 ,mul_84_22_n_235);
  not mul_84_22_drc_bufs3891(mul_84_22_n_236 ,mul_84_22_n_235);
  not mul_84_22_drc_bufs3892(mul_84_22_n_235 ,mul_84_22_n_336);
  not mul_84_22_drc_bufs3894(mul_84_22_n_234 ,mul_84_22_n_232);
  not mul_84_22_drc_bufs3895(mul_84_22_n_233 ,mul_84_22_n_232);
  not mul_84_22_drc_bufs3896(mul_84_22_n_232 ,mul_84_22_n_383);
  not mul_84_22_drc_bufs3898(mul_84_22_n_231 ,mul_84_22_n_229);
  not mul_84_22_drc_bufs3899(mul_84_22_n_230 ,mul_84_22_n_229);
  not mul_84_22_drc_bufs3900(mul_84_22_n_229 ,mul_84_22_n_382);
  not mul_84_22_drc_bufs3902(mul_84_22_n_228 ,mul_84_22_n_226);
  not mul_84_22_drc_bufs3903(mul_84_22_n_227 ,mul_84_22_n_226);
  not mul_84_22_drc_bufs3904(mul_84_22_n_226 ,mul_84_22_n_305);
  not mul_84_22_drc_bufs3906(mul_84_22_n_225 ,mul_84_22_n_223);
  not mul_84_22_drc_bufs3907(mul_84_22_n_224 ,mul_84_22_n_223);
  not mul_84_22_drc_bufs3908(mul_84_22_n_223 ,mul_84_22_n_304);
  not mul_84_22_drc_bufs3910(mul_84_22_n_222 ,mul_84_22_n_220);
  not mul_84_22_drc_bufs3911(mul_84_22_n_221 ,mul_84_22_n_220);
  not mul_84_22_drc_bufs3912(mul_84_22_n_220 ,mul_84_22_n_379);
  not mul_84_22_drc_bufs3914(mul_84_22_n_219 ,mul_84_22_n_217);
  not mul_84_22_drc_bufs3915(mul_84_22_n_218 ,mul_84_22_n_217);
  not mul_84_22_drc_bufs3916(mul_84_22_n_217 ,mul_84_22_n_380);
  not mul_84_22_drc_bufs3918(mul_84_22_n_216 ,mul_84_22_n_214);
  not mul_84_22_drc_bufs3919(mul_84_22_n_215 ,mul_84_22_n_214);
  not mul_84_22_drc_bufs3920(mul_84_22_n_214 ,mul_84_22_n_302);
  not mul_84_22_drc_bufs3922(mul_84_22_n_213 ,mul_84_22_n_211);
  not mul_84_22_drc_bufs3923(mul_84_22_n_212 ,mul_84_22_n_211);
  not mul_84_22_drc_bufs3924(mul_84_22_n_211 ,mul_84_22_n_332);
  not mul_84_22_drc_bufs3926(mul_84_22_n_210 ,mul_84_22_n_208);
  not mul_84_22_drc_bufs3927(mul_84_22_n_209 ,mul_84_22_n_208);
  not mul_84_22_drc_bufs3928(mul_84_22_n_208 ,mul_84_22_n_300);
  not mul_84_22_drc_bufs3930(mul_84_22_n_207 ,mul_84_22_n_205);
  not mul_84_22_drc_bufs3931(mul_84_22_n_206 ,mul_84_22_n_205);
  not mul_84_22_drc_bufs3932(mul_84_22_n_205 ,mul_84_22_n_333);
  not mul_84_22_drc_bufs3934(mul_84_22_n_204 ,mul_84_22_n_649);
  not mul_84_22_drc_bufs3935(mul_84_22_n_203 ,mul_84_22_n_649);
  not mul_84_22_drc_bufs3940(mul_84_22_n_307 ,mul_84_22_n_650);
  not mul_84_22_drc_bufs3943(mul_84_22_n_202 ,mul_84_22_n_201);
  not mul_84_22_drc_bufs3944(mul_84_22_n_201 ,mul_84_22_n_311);
  not mul_84_22_drc_bufs3946(mul_84_22_n_200 ,mul_84_22_n_198);
  not mul_84_22_drc_bufs3947(mul_84_22_n_199 ,mul_84_22_n_198);
  not mul_84_22_drc_bufs3948(mul_84_22_n_198 ,mul_84_22_n_301);
  buf mul_84_22_drc_bufs3957(n_184 ,mul_84_22_n_1140);
  buf mul_84_22_drc_bufs3958(n_185 ,mul_84_22_n_1143);
  buf mul_84_22_drc_bufs3959(n_178 ,mul_84_22_n_1121);
  buf mul_84_22_drc_bufs3960(n_180 ,mul_84_22_n_1127);
  buf mul_84_22_drc_bufs3961(n_181 ,mul_84_22_n_1130);
  buf mul_84_22_drc_bufs3962(n_188 ,mul_84_22_n_1153);
  buf mul_84_22_drc_bufs3963(n_183 ,mul_84_22_n_1137);
  buf mul_84_22_drc_bufs3964(n_182 ,mul_84_22_n_1134);
  buf mul_84_22_drc_bufs3965(n_179 ,mul_84_22_n_1124);
  buf mul_84_22_drc_bufs3966(n_189 ,mul_84_22_n_1156);
  buf mul_84_22_drc_bufs3967(n_186 ,mul_84_22_n_1147);
  buf mul_84_22_drc_bufs3968(n_187 ,mul_84_22_n_1150);
  buf mul_84_22_drc_bufs3969(n_175 ,mul_84_22_n_1112);
  buf mul_84_22_drc_bufs3970(n_176 ,mul_84_22_n_1115);
  buf mul_84_22_drc_bufs3971(n_177 ,mul_84_22_n_1118);
  not mul_84_22_drc_bufs3973(mul_84_22_n_182 ,mul_84_22_n_308);
  not mul_84_22_drc_bufs3974(mul_84_22_n_308 ,mul_84_22_n_885);
  not mul_84_22_drc_bufs3996(mul_84_22_n_181 ,mul_84_22_n_180);
  not mul_84_22_drc_bufs3998(mul_84_22_n_180 ,mul_84_22_n_446);
  not mul_84_22_drc_bufs4001(mul_84_22_n_179 ,mul_84_22_n_178);
  not mul_84_22_drc_bufs4003(mul_84_22_n_178 ,mul_84_22_n_444);
  not mul_84_22_drc_bufs4006(mul_84_22_n_177 ,mul_84_22_n_176);
  not mul_84_22_drc_bufs4008(mul_84_22_n_176 ,mul_84_22_n_447);
  not mul_84_22_drc_bufs4011(mul_84_22_n_175 ,mul_84_22_n_174);
  not mul_84_22_drc_bufs4013(mul_84_22_n_174 ,mul_84_22_n_445);
  not mul_84_22_drc_bufs4021(mul_84_22_n_173 ,mul_84_22_n_172);
  not mul_84_22_drc_bufs4023(mul_84_22_n_172 ,mul_84_22_n_317);
  not mul_84_22_drc_bufs4031(mul_84_22_n_171 ,mul_84_22_n_169);
  not mul_84_22_drc_bufs4032(mul_84_22_n_170 ,mul_84_22_n_169);
  not mul_84_22_drc_bufs4033(mul_84_22_n_169 ,mul_84_22_n_448);
  not mul_84_22_drc_bufs4036(mul_84_22_n_168 ,mul_84_22_n_167);
  not mul_84_22_drc_bufs4037(mul_84_22_n_167 ,mul_84_22_n_297);
  not mul_84_22_drc_bufs4039(mul_84_22_n_166 ,mul_84_22_n_164);
  not mul_84_22_drc_bufs4040(mul_84_22_n_165 ,mul_84_22_n_164);
  not mul_84_22_drc_bufs4041(mul_84_22_n_164 ,mul_84_22_n_296);
  not mul_84_22_drc_bufs4043(mul_84_22_n_163 ,mul_84_22_n_161);
  not mul_84_22_drc_bufs4044(mul_84_22_n_162 ,mul_84_22_n_161);
  not mul_84_22_drc_bufs4045(mul_84_22_n_161 ,mul_84_22_n_312);
  not mul_84_22_drc_bufs4047(mul_84_22_n_160 ,mul_84_22_n_158);
  not mul_84_22_drc_bufs4048(mul_84_22_n_159 ,mul_84_22_n_158);
  not mul_84_22_drc_bufs4049(mul_84_22_n_158 ,mul_84_22_n_312);
  not mul_84_22_drc_bufs4051(mul_84_22_n_157 ,mul_84_22_n_306);
  not mul_84_22_drc_bufs4053(mul_84_22_n_306 ,mul_84_22_n_648);
  not mul_84_22_drc_bufs4056(mul_84_22_n_156 ,mul_84_22_n_155);
  not mul_84_22_drc_bufs4057(mul_84_22_n_155 ,mul_84_22_n_648);
  not mul_84_22_drc_bufs4059(mul_84_22_n_154 ,mul_84_22_n_299);
  not mul_84_22_drc_bufs4061(mul_84_22_n_299 ,mul_84_22_n_331);
  not mul_84_22_drc_bufs4063(mul_84_22_n_153 ,mul_84_22_n_298);
  not mul_84_22_drc_bufs4065(mul_84_22_n_298 ,mul_84_22_n_331);
  not mul_84_22_drc_bufs4067(mul_84_22_n_152 ,mul_84_22_n_305);
  not mul_84_22_drc_bufs4069(mul_84_22_n_305 ,mul_84_22_n_381);
  not mul_84_22_drc_bufs4071(mul_84_22_n_151 ,mul_84_22_n_304);
  not mul_84_22_drc_bufs4073(mul_84_22_n_304 ,mul_84_22_n_381);
  not mul_84_22_drc_bufs4075(mul_84_22_n_150 ,mul_84_22_n_303);
  not mul_84_22_drc_bufs4077(mul_84_22_n_303 ,mul_84_22_n_378);
  not mul_84_22_drc_bufs4079(mul_84_22_n_149 ,mul_84_22_n_302);
  not mul_84_22_drc_bufs4081(mul_84_22_n_302 ,mul_84_22_n_378);
  not mul_84_22_drc_bufs4083(mul_84_22_n_148 ,mul_84_22_n_301);
  not mul_84_22_drc_bufs4085(mul_84_22_n_301 ,mul_84_22_n_334);
  not mul_84_22_drc_bufs4087(mul_84_22_n_147 ,mul_84_22_n_300);
  not mul_84_22_drc_bufs4089(mul_84_22_n_300 ,mul_84_22_n_334);
  not mul_84_22_drc_bufs4091(mul_84_22_n_146 ,mul_84_22_n_145);
  not mul_84_22_drc_bufs4093(mul_84_22_n_145 ,mul_84_22_n_281);
  not mul_84_22_drc_bufs4095(mul_84_22_n_144 ,mul_84_22_n_143);
  not mul_84_22_drc_bufs4097(mul_84_22_n_143 ,mul_84_22_n_291);
  not mul_84_22_drc_bufs4099(mul_84_22_n_142 ,mul_84_22_n_141);
  not mul_84_22_drc_bufs4101(mul_84_22_n_141 ,mul_84_22_n_273);
  not mul_84_22_drc_bufs4103(mul_84_22_n_140 ,mul_84_22_n_139);
  not mul_84_22_drc_bufs4105(mul_84_22_n_139 ,mul_84_22_n_294);
  not mul_84_22_drc_bufs4107(mul_84_22_n_138 ,mul_84_22_n_137);
  not mul_84_22_drc_bufs4109(mul_84_22_n_137 ,mul_84_22_n_255);
  not mul_84_22_drc_bufs4111(mul_84_22_n_136 ,mul_84_22_n_135);
  not mul_84_22_drc_bufs4113(mul_84_22_n_135 ,mul_84_22_n_282);
  not mul_84_22_drc_bufs4115(mul_84_22_n_134 ,mul_84_22_n_133);
  not mul_84_22_drc_bufs4117(mul_84_22_n_133 ,mul_84_22_n_261);
  not mul_84_22_drc_bufs4119(mul_84_22_n_132 ,mul_84_22_n_131);
  not mul_84_22_drc_bufs4121(mul_84_22_n_131 ,mul_84_22_n_264);
  not mul_84_22_drc_bufs4123(mul_84_22_n_130 ,mul_84_22_n_129);
  not mul_84_22_drc_bufs4125(mul_84_22_n_129 ,mul_84_22_n_266);
  not mul_84_22_drc_bufs4127(mul_84_22_n_128 ,mul_84_22_n_127);
  not mul_84_22_drc_bufs4129(mul_84_22_n_127 ,mul_84_22_n_276);
  not mul_84_22_drc_bufs4131(mul_84_22_n_126 ,mul_84_22_n_125);
  not mul_84_22_drc_bufs4133(mul_84_22_n_125 ,mul_84_22_n_258);
  not mul_84_22_drc_bufs4135(mul_84_22_n_124 ,mul_84_22_n_123);
  not mul_84_22_drc_bufs4137(mul_84_22_n_123 ,mul_84_22_n_260);
  not mul_84_22_drc_bufs4139(mul_84_22_n_122 ,mul_84_22_n_121);
  not mul_84_22_drc_bufs4141(mul_84_22_n_121 ,mul_84_22_n_252);
  not mul_84_22_drc_bufs4143(mul_84_22_n_120 ,mul_84_22_n_119);
  not mul_84_22_drc_bufs4145(mul_84_22_n_119 ,mul_84_22_n_270);
  not mul_84_22_drc_bufs4147(mul_84_22_n_118 ,mul_84_22_n_117);
  not mul_84_22_drc_bufs4149(mul_84_22_n_117 ,mul_84_22_n_254);
  not mul_84_22_drc_bufs4151(mul_84_22_n_116 ,mul_84_22_n_115);
  not mul_84_22_drc_bufs4153(mul_84_22_n_115 ,mul_84_22_n_263);
  not mul_84_22_drc_bufs4155(mul_84_22_n_114 ,mul_84_22_n_113);
  not mul_84_22_drc_bufs4157(mul_84_22_n_113 ,mul_84_22_n_290);
  not mul_84_22_drc_bufs4159(mul_84_22_n_112 ,mul_84_22_n_111);
  not mul_84_22_drc_bufs4161(mul_84_22_n_111 ,mul_84_22_n_293);
  not mul_84_22_drc_bufs4163(mul_84_22_n_110 ,mul_84_22_n_109);
  not mul_84_22_drc_bufs4165(mul_84_22_n_109 ,mul_84_22_n_267);
  not mul_84_22_drc_bufs4167(mul_84_22_n_108 ,mul_84_22_n_107);
  not mul_84_22_drc_bufs4169(mul_84_22_n_107 ,mul_84_22_n_284);
  not mul_84_22_drc_bufs4171(mul_84_22_n_106 ,mul_84_22_n_105);
  not mul_84_22_drc_bufs4173(mul_84_22_n_105 ,mul_84_22_n_269);
  not mul_84_22_drc_bufs4175(mul_84_22_n_104 ,mul_84_22_n_103);
  not mul_84_22_drc_bufs4177(mul_84_22_n_103 ,mul_84_22_n_278);
  not mul_84_22_drc_bufs4179(mul_84_22_n_102 ,mul_84_22_n_101);
  not mul_84_22_drc_bufs4181(mul_84_22_n_101 ,mul_84_22_n_275);
  not mul_84_22_drc_bufs4183(mul_84_22_n_100 ,mul_84_22_n_99);
  not mul_84_22_drc_bufs4185(mul_84_22_n_99 ,mul_84_22_n_257);
  not mul_84_22_drc_bufs4187(mul_84_22_n_98 ,mul_84_22_n_97);
  not mul_84_22_drc_bufs4189(mul_84_22_n_97 ,mul_84_22_n_272);
  not mul_84_22_drc_bufs4191(mul_84_22_n_96 ,mul_84_22_n_95);
  not mul_84_22_drc_bufs4193(mul_84_22_n_95 ,mul_84_22_n_287);
  not mul_84_22_drc_bufs4195(mul_84_22_n_94 ,mul_84_22_n_93);
  not mul_84_22_drc_bufs4197(mul_84_22_n_93 ,mul_84_22_n_285);
  not mul_84_22_drc_bufs4199(mul_84_22_n_92 ,mul_84_22_n_91);
  not mul_84_22_drc_bufs4201(mul_84_22_n_91 ,mul_84_22_n_279);
  not mul_84_22_drc_bufs4203(mul_84_22_n_90 ,mul_84_22_n_89);
  not mul_84_22_drc_bufs4205(mul_84_22_n_89 ,mul_84_22_n_288);
  not mul_84_22_drc_bufs4207(mul_84_22_n_88 ,mul_84_22_n_86);
  not mul_84_22_drc_bufs4208(mul_84_22_n_87 ,mul_84_22_n_86);
  not mul_84_22_drc_bufs4209(mul_84_22_n_86 ,mul_84_22_n_446);
  not mul_84_22_drc_bufs4211(mul_84_22_n_85 ,mul_84_22_n_83);
  not mul_84_22_drc_bufs4212(mul_84_22_n_84 ,mul_84_22_n_83);
  not mul_84_22_drc_bufs4213(mul_84_22_n_83 ,mul_84_22_n_444);
  not mul_84_22_drc_bufs4215(mul_84_22_n_82 ,mul_84_22_n_80);
  not mul_84_22_drc_bufs4216(mul_84_22_n_81 ,mul_84_22_n_80);
  not mul_84_22_drc_bufs4217(mul_84_22_n_80 ,mul_84_22_n_445);
  not mul_84_22_drc_bufs4219(mul_84_22_n_79 ,mul_84_22_n_77);
  not mul_84_22_drc_bufs4220(mul_84_22_n_78 ,mul_84_22_n_77);
  not mul_84_22_drc_bufs4221(mul_84_22_n_77 ,mul_84_22_n_447);
  not mul_84_22_drc_bufs4223(mul_84_22_n_76 ,mul_84_22_n_74);
  not mul_84_22_drc_bufs4224(mul_84_22_n_75 ,mul_84_22_n_74);
  not mul_84_22_drc_bufs4225(mul_84_22_n_74 ,mul_84_22_n_181);
  not mul_84_22_drc_bufs4227(mul_84_22_n_73 ,mul_84_22_n_71);
  not mul_84_22_drc_bufs4228(mul_84_22_n_72 ,mul_84_22_n_71);
  not mul_84_22_drc_bufs4229(mul_84_22_n_71 ,mul_84_22_n_317);
  not mul_84_22_drc_bufs4231(mul_84_22_n_70 ,mul_84_22_n_68);
  not mul_84_22_drc_bufs4232(mul_84_22_n_69 ,mul_84_22_n_68);
  not mul_84_22_drc_bufs4233(mul_84_22_n_68 ,mul_84_22_n_173);
  not mul_84_22_drc_bufs4235(mul_84_22_n_67 ,mul_84_22_n_65);
  not mul_84_22_drc_bufs4236(mul_84_22_n_66 ,mul_84_22_n_65);
  not mul_84_22_drc_bufs4237(mul_84_22_n_65 ,mul_84_22_n_446);
  not mul_84_22_drc_bufs4239(mul_84_22_n_64 ,mul_84_22_n_62);
  not mul_84_22_drc_bufs4240(mul_84_22_n_63 ,mul_84_22_n_62);
  not mul_84_22_drc_bufs4241(mul_84_22_n_62 ,mul_84_22_n_179);
  not mul_84_22_drc_bufs4243(mul_84_22_n_61 ,mul_84_22_n_59);
  not mul_84_22_drc_bufs4244(mul_84_22_n_60 ,mul_84_22_n_59);
  not mul_84_22_drc_bufs4245(mul_84_22_n_59 ,mul_84_22_n_177);
  not mul_84_22_drc_bufs4247(mul_84_22_n_58 ,mul_84_22_n_56);
  not mul_84_22_drc_bufs4248(mul_84_22_n_57 ,mul_84_22_n_56);
  not mul_84_22_drc_bufs4249(mul_84_22_n_56 ,mul_84_22_n_175);
  not mul_84_22_drc_bufs4251(mul_84_22_n_55 ,mul_84_22_n_53);
  not mul_84_22_drc_bufs4252(mul_84_22_n_54 ,mul_84_22_n_53);
  not mul_84_22_drc_bufs4253(mul_84_22_n_53 ,mul_84_22_n_317);
  not mul_84_22_drc_bufs4255(mul_84_22_n_52 ,mul_84_22_n_50);
  not mul_84_22_drc_bufs4256(mul_84_22_n_51 ,mul_84_22_n_50);
  not mul_84_22_drc_bufs4257(mul_84_22_n_50 ,mul_84_22_n_177);
  not mul_84_22_drc_bufs4259(mul_84_22_n_49 ,mul_84_22_n_47);
  not mul_84_22_drc_bufs4260(mul_84_22_n_48 ,mul_84_22_n_47);
  not mul_84_22_drc_bufs4261(mul_84_22_n_47 ,mul_84_22_n_444);
  not mul_84_22_drc_bufs4263(mul_84_22_n_46 ,mul_84_22_n_44);
  not mul_84_22_drc_bufs4264(mul_84_22_n_45 ,mul_84_22_n_44);
  not mul_84_22_drc_bufs4265(mul_84_22_n_44 ,mul_84_22_n_448);
  not mul_84_22_drc_bufs4267(mul_84_22_n_43 ,mul_84_22_n_41);
  not mul_84_22_drc_bufs4268(mul_84_22_n_42 ,mul_84_22_n_41);
  not mul_84_22_drc_bufs4269(mul_84_22_n_41 ,mul_84_22_n_173);
  not mul_84_22_drc_bufs4271(mul_84_22_n_40 ,mul_84_22_n_38);
  not mul_84_22_drc_bufs4272(mul_84_22_n_39 ,mul_84_22_n_38);
  not mul_84_22_drc_bufs4273(mul_84_22_n_38 ,mul_84_22_n_181);
  not mul_84_22_drc_bufs4275(mul_84_22_n_37 ,mul_84_22_n_35);
  not mul_84_22_drc_bufs4276(mul_84_22_n_36 ,mul_84_22_n_35);
  not mul_84_22_drc_bufs4277(mul_84_22_n_35 ,mul_84_22_n_175);
  not mul_84_22_drc_bufs4279(mul_84_22_n_34 ,mul_84_22_n_32);
  not mul_84_22_drc_bufs4280(mul_84_22_n_33 ,mul_84_22_n_32);
  not mul_84_22_drc_bufs4281(mul_84_22_n_32 ,mul_84_22_n_448);
  not mul_84_22_drc_bufs4283(mul_84_22_n_31 ,mul_84_22_n_29);
  not mul_84_22_drc_bufs4284(mul_84_22_n_30 ,mul_84_22_n_29);
  not mul_84_22_drc_bufs4285(mul_84_22_n_29 ,mul_84_22_n_447);
  not mul_84_22_drc_bufs4287(mul_84_22_n_28 ,mul_84_22_n_26);
  not mul_84_22_drc_bufs4288(mul_84_22_n_27 ,mul_84_22_n_26);
  not mul_84_22_drc_bufs4289(mul_84_22_n_26 ,mul_84_22_n_179);
  not mul_84_22_drc_bufs4291(mul_84_22_n_25 ,mul_84_22_n_23);
  not mul_84_22_drc_bufs4292(mul_84_22_n_24 ,mul_84_22_n_23);
  not mul_84_22_drc_bufs4293(mul_84_22_n_23 ,mul_84_22_n_445);
  not mul_84_22_drc_bufs4295(mul_84_22_n_22 ,mul_84_22_n_20);
  not mul_84_22_drc_bufs4296(mul_84_22_n_21 ,mul_84_22_n_20);
  not mul_84_22_drc_bufs4297(mul_84_22_n_20 ,mul_84_22_n_171);
  not mul_84_22_drc_bufs4299(mul_84_22_n_19 ,mul_84_22_n_17);
  not mul_84_22_drc_bufs4300(mul_84_22_n_18 ,mul_84_22_n_17);
  not mul_84_22_drc_bufs4301(mul_84_22_n_17 ,mul_84_22_n_297);
  not mul_84_22_drc_bufs4303(mul_84_22_n_16 ,mul_84_22_n_15);
  not mul_84_22_drc_bufs4305(mul_84_22_n_15 ,mul_84_22_n_170);
  not mul_84_22_drc_bufs4307(mul_84_22_n_14 ,mul_84_22_n_13);
  not mul_84_22_drc_bufs4309(mul_84_22_n_13 ,mul_84_22_n_88);
  not mul_84_22_drc_bufs4311(mul_84_22_n_12 ,mul_84_22_n_11);
  not mul_84_22_drc_bufs4313(mul_84_22_n_11 ,mul_84_22_n_79);
  not mul_84_22_drc_bufs4315(mul_84_22_n_10 ,mul_84_22_n_9);
  not mul_84_22_drc_bufs4317(mul_84_22_n_9 ,mul_84_22_n_82);
  not mul_84_22_drc_bufs4319(mul_84_22_n_8 ,mul_84_22_n_7);
  not mul_84_22_drc_bufs4321(mul_84_22_n_7 ,mul_84_22_n_85);
  and mul_84_22_g2(mul_84_22_n_6 ,mul_84_22_n_982 ,mul_84_22_n_996);
  and mul_84_22_g4323(mul_84_22_n_5 ,mul_84_22_n_913 ,mul_84_22_n_966);
  xor mul_84_22_g4324(mul_84_22_n_4 ,mul_84_22_n_882 ,mul_84_22_n_963);
  xor mul_84_22_g4325(mul_84_22_n_3 ,mul_84_22_n_889 ,mul_84_22_n_960);
  xor mul_84_22_g4326(mul_84_22_n_2 ,mul_84_22_n_890 ,mul_84_22_n_930);
  xor mul_84_22_g4327(mul_84_22_n_1 ,mul_84_22_n_599 ,mul_84_22_n_847);
  xor mul_84_22_g4328(mul_84_22_n_0 ,mul_84_22_n_801 ,mul_84_22_n_307);
  xnor mul_90_22_g2868(n_158 ,mul_90_22_n_984 ,mul_90_22_n_1157);
  nor mul_90_22_g2869(mul_90_22_n_1157 ,mul_90_22_n_1026 ,mul_90_22_n_1155);
  xnor mul_90_22_g2870(mul_90_22_n_1156 ,mul_90_22_n_1154 ,mul_90_22_n_1040);
  and mul_90_22_g2871(mul_90_22_n_1155 ,mul_90_22_n_1027 ,mul_90_22_n_1154);
  or mul_90_22_g2872(mul_90_22_n_1154 ,mul_90_22_n_1050 ,mul_90_22_n_1152);
  xnor mul_90_22_g2873(mul_90_22_n_1153 ,mul_90_22_n_1151 ,mul_90_22_n_1061);
  and mul_90_22_g2874(mul_90_22_n_1152 ,mul_90_22_n_1051 ,mul_90_22_n_1151);
  or mul_90_22_g2875(mul_90_22_n_1151 ,mul_90_22_n_1079 ,mul_90_22_n_1149);
  xnor mul_90_22_g2876(mul_90_22_n_1150 ,mul_90_22_n_1148 ,mul_90_22_n_1081);
  nor mul_90_22_g2877(mul_90_22_n_1149 ,mul_90_22_n_1072 ,mul_90_22_n_1148);
  and mul_90_22_g2878(mul_90_22_n_1148 ,mul_90_22_n_1094 ,mul_90_22_n_1146);
  xnor mul_90_22_g2879(mul_90_22_n_1147 ,mul_90_22_n_1144 ,mul_90_22_n_1106);
  or mul_90_22_g2880(mul_90_22_n_1146 ,mul_90_22_n_1093 ,mul_90_22_n_1145);
  not mul_90_22_g2881(mul_90_22_n_1145 ,mul_90_22_n_1144);
  or mul_90_22_g2882(mul_90_22_n_1144 ,mul_90_22_n_1073 ,mul_90_22_n_1142);
  xnor mul_90_22_g2883(mul_90_22_n_1143 ,mul_90_22_n_1141 ,mul_90_22_n_1082);
  and mul_90_22_g2884(mul_90_22_n_1142 ,mul_90_22_n_1080 ,mul_90_22_n_1141);
  or mul_90_22_g2885(mul_90_22_n_1141 ,mul_90_22_n_1087 ,mul_90_22_n_1139);
  xnor mul_90_22_g2886(mul_90_22_n_1140 ,mul_90_22_n_1138 ,mul_90_22_n_1105);
  and mul_90_22_g2887(mul_90_22_n_1139 ,mul_90_22_n_1086 ,mul_90_22_n_1138);
  or mul_90_22_g2888(mul_90_22_n_1138 ,mul_90_22_n_1085 ,mul_90_22_n_1136);
  xnor mul_90_22_g2889(mul_90_22_n_1137 ,mul_90_22_n_1135 ,mul_90_22_n_1104);
  nor mul_90_22_g2890(mul_90_22_n_1136 ,mul_90_22_n_1135 ,mul_90_22_n_1099);
  and mul_90_22_g2891(mul_90_22_n_1135 ,mul_90_22_n_1092 ,mul_90_22_n_1133);
  xnor mul_90_22_g2892(mul_90_22_n_1134 ,mul_90_22_n_1131 ,mul_90_22_n_1103);
  or mul_90_22_g2893(mul_90_22_n_1133 ,mul_90_22_n_1090 ,mul_90_22_n_1132);
  not mul_90_22_g2894(mul_90_22_n_1132 ,mul_90_22_n_1131);
  or mul_90_22_g2895(mul_90_22_n_1131 ,mul_90_22_n_1089 ,mul_90_22_n_1129);
  xnor mul_90_22_g2896(mul_90_22_n_1130 ,mul_90_22_n_1128 ,mul_90_22_n_1102);
  and mul_90_22_g2897(mul_90_22_n_1129 ,mul_90_22_n_1088 ,mul_90_22_n_1128);
  or mul_90_22_g2898(mul_90_22_n_1128 ,mul_90_22_n_1075 ,mul_90_22_n_1126);
  xnor mul_90_22_g2899(mul_90_22_n_1127 ,mul_90_22_n_1125 ,mul_90_22_n_1084);
  and mul_90_22_g2900(mul_90_22_n_1126 ,mul_90_22_n_1074 ,mul_90_22_n_1125);
  or mul_90_22_g2901(mul_90_22_n_1125 ,mul_90_22_n_1098 ,mul_90_22_n_1123);
  xnor mul_90_22_g2902(mul_90_22_n_1124 ,mul_90_22_n_1122 ,mul_90_22_n_1101);
  and mul_90_22_g2903(mul_90_22_n_1123 ,mul_90_22_n_1097 ,mul_90_22_n_1122);
  or mul_90_22_g2904(mul_90_22_n_1122 ,mul_90_22_n_1078 ,mul_90_22_n_1120);
  xnor mul_90_22_g2905(mul_90_22_n_1121 ,mul_90_22_n_1119 ,mul_90_22_n_1083);
  and mul_90_22_g2906(mul_90_22_n_1120 ,mul_90_22_n_1077 ,mul_90_22_n_1119);
  or mul_90_22_g2907(mul_90_22_n_1119 ,mul_90_22_n_1096 ,mul_90_22_n_1117);
  xnor mul_90_22_g2908(mul_90_22_n_1118 ,mul_90_22_n_1116 ,mul_90_22_n_1100);
  and mul_90_22_g2909(mul_90_22_n_1117 ,mul_90_22_n_1095 ,mul_90_22_n_1116);
  or mul_90_22_g2910(mul_90_22_n_1116 ,mul_90_22_n_1041 ,mul_90_22_n_1114);
  xnor mul_90_22_g2911(mul_90_22_n_1115 ,mul_90_22_n_1113 ,mul_90_22_n_1060);
  and mul_90_22_g2912(mul_90_22_n_1114 ,mul_90_22_n_1042 ,mul_90_22_n_1113);
  or mul_90_22_g2913(mul_90_22_n_1113 ,mul_90_22_n_1043 ,mul_90_22_n_1111);
  xnor mul_90_22_g2914(mul_90_22_n_1112 ,mul_90_22_n_1110 ,mul_90_22_n_1059);
  and mul_90_22_g2915(mul_90_22_n_1111 ,mul_90_22_n_1044 ,mul_90_22_n_1110);
  or mul_90_22_g2916(mul_90_22_n_1110 ,mul_90_22_n_6 ,mul_90_22_n_1109);
  nor mul_90_22_g2917(mul_90_22_n_1109 ,mul_90_22_n_1016 ,mul_90_22_n_1108);
  nor mul_90_22_g2918(mul_90_22_n_1108 ,mul_90_22_n_5 ,mul_90_22_n_1107);
  nor mul_90_22_g2919(mul_90_22_n_1107 ,mul_90_22_n_1003 ,mul_90_22_n_1091);
  xnor mul_90_22_g2920(mul_90_22_n_1106 ,mul_90_22_n_1062 ,mul_90_22_n_1039);
  xnor mul_90_22_g2921(mul_90_22_n_1105 ,mul_90_22_n_1019 ,mul_90_22_n_1063);
  xnor mul_90_22_g2922(mul_90_22_n_1104 ,mul_90_22_n_1038 ,mul_90_22_n_1070);
  xnor mul_90_22_g2923(mul_90_22_n_1103 ,mul_90_22_n_1037 ,mul_90_22_n_1069);
  xnor mul_90_22_g2924(mul_90_22_n_1102 ,mul_90_22_n_1055 ,mul_90_22_n_1066);
  xnor mul_90_22_g2925(mul_90_22_n_1101 ,mul_90_22_n_1065 ,mul_90_22_n_1058);
  xnor mul_90_22_g2926(mul_90_22_n_1100 ,mul_90_22_n_1035 ,mul_90_22_n_1067);
  and mul_90_22_g2927(mul_90_22_n_1099 ,mul_90_22_n_1038 ,mul_90_22_n_1071);
  nor mul_90_22_g2928(mul_90_22_n_1098 ,mul_90_22_n_1058 ,mul_90_22_n_1065);
  or mul_90_22_g2929(mul_90_22_n_1097 ,mul_90_22_n_1057 ,mul_90_22_n_1064);
  and mul_90_22_g2930(mul_90_22_n_1096 ,mul_90_22_n_1035 ,mul_90_22_n_1067);
  or mul_90_22_g2931(mul_90_22_n_1095 ,mul_90_22_n_1035 ,mul_90_22_n_1067);
  or mul_90_22_g2932(mul_90_22_n_1094 ,mul_90_22_n_1039 ,mul_90_22_n_1062);
  and mul_90_22_g2933(mul_90_22_n_1093 ,mul_90_22_n_1039 ,mul_90_22_n_1062);
  or mul_90_22_g2934(mul_90_22_n_1092 ,mul_90_22_n_1036 ,mul_90_22_n_1068);
  nor mul_90_22_g2935(mul_90_22_n_1091 ,mul_90_22_n_1000 ,mul_90_22_n_1076);
  nor mul_90_22_g2936(mul_90_22_n_1090 ,mul_90_22_n_1037 ,mul_90_22_n_1069);
  and mul_90_22_g2937(mul_90_22_n_1089 ,mul_90_22_n_1055 ,mul_90_22_n_1066);
  or mul_90_22_g2938(mul_90_22_n_1088 ,mul_90_22_n_1055 ,mul_90_22_n_1066);
  and mul_90_22_g2939(mul_90_22_n_1087 ,mul_90_22_n_1019 ,mul_90_22_n_1063);
  or mul_90_22_g2940(mul_90_22_n_1086 ,mul_90_22_n_1019 ,mul_90_22_n_1063);
  nor mul_90_22_g2941(mul_90_22_n_1085 ,mul_90_22_n_1038 ,mul_90_22_n_1071);
  xnor mul_90_22_g2942(mul_90_22_n_1084 ,mul_90_22_n_1056 ,mul_90_22_n_1045);
  xnor mul_90_22_g2943(mul_90_22_n_1083 ,mul_90_22_n_1047 ,mul_90_22_n_1053);
  xnor mul_90_22_g2944(mul_90_22_n_1082 ,mul_90_22_n_1034 ,mul_90_22_n_1048);
  xnor mul_90_22_g2945(mul_90_22_n_1081 ,mul_90_22_n_1054 ,mul_90_22_n_1017);
  or mul_90_22_g2946(mul_90_22_n_1080 ,mul_90_22_n_1034 ,mul_90_22_n_1048);
  nor mul_90_22_g2947(mul_90_22_n_1079 ,mul_90_22_n_1054 ,mul_90_22_n_1018);
  nor mul_90_22_g2948(mul_90_22_n_1078 ,mul_90_22_n_1053 ,mul_90_22_n_1047);
  or mul_90_22_g2949(mul_90_22_n_1077 ,mul_90_22_n_1052 ,mul_90_22_n_1046);
  nor mul_90_22_g2950(mul_90_22_n_1076 ,mul_90_22_n_999 ,mul_90_22_n_1049);
  and mul_90_22_g2951(mul_90_22_n_1075 ,mul_90_22_n_1056 ,mul_90_22_n_1045);
  or mul_90_22_g2952(mul_90_22_n_1074 ,mul_90_22_n_1056 ,mul_90_22_n_1045);
  and mul_90_22_g2953(mul_90_22_n_1073 ,mul_90_22_n_1034 ,mul_90_22_n_1048);
  and mul_90_22_g2954(mul_90_22_n_1072 ,mul_90_22_n_1054 ,mul_90_22_n_1018);
  not mul_90_22_g2955(mul_90_22_n_1071 ,mul_90_22_n_1070);
  not mul_90_22_g2956(mul_90_22_n_1069 ,mul_90_22_n_1068);
  not mul_90_22_g2957(mul_90_22_n_1065 ,mul_90_22_n_1064);
  xnor mul_90_22_g2958(mul_90_22_n_1061 ,mul_90_22_n_1023 ,mul_90_22_n_1033);
  xnor mul_90_22_g2959(mul_90_22_n_1060 ,mul_90_22_n_1009 ,mul_90_22_n_1021);
  xnor mul_90_22_g2960(mul_90_22_n_1059 ,mul_90_22_n_1010 ,mul_90_22_n_1020);
  xnor mul_90_22_g2961(mul_90_22_n_1070 ,mul_90_22_n_941 ,mul_90_22_n_1011);
  xnor mul_90_22_g2962(mul_90_22_n_1068 ,mul_90_22_n_925 ,mul_90_22_n_4);
  xnor mul_90_22_g2963(mul_90_22_n_1067 ,mul_90_22_n_945 ,mul_90_22_n_1014);
  xnor mul_90_22_g2964(mul_90_22_n_1066 ,mul_90_22_n_942 ,mul_90_22_n_3);
  xnor mul_90_22_g2965(mul_90_22_n_1064 ,mul_90_22_n_912 ,mul_90_22_n_1012);
  xnor mul_90_22_g2966(mul_90_22_n_1063 ,mul_90_22_n_939 ,mul_90_22_n_1013);
  xnor mul_90_22_g2967(mul_90_22_n_1062 ,mul_90_22_n_944 ,mul_90_22_n_1015);
  not mul_90_22_g2968(mul_90_22_n_1057 ,mul_90_22_n_1058);
  not mul_90_22_g2969(mul_90_22_n_1052 ,mul_90_22_n_1053);
  or mul_90_22_g2970(mul_90_22_n_1051 ,mul_90_22_n_1032 ,mul_90_22_n_1022);
  nor mul_90_22_g2971(mul_90_22_n_1050 ,mul_90_22_n_1033 ,mul_90_22_n_1023);
  nor mul_90_22_g2972(mul_90_22_n_1049 ,mul_90_22_n_921 ,mul_90_22_n_1031);
  and mul_90_22_g2973(mul_90_22_n_1058 ,mul_90_22_n_993 ,mul_90_22_n_1024);
  or mul_90_22_g2974(mul_90_22_n_1056 ,mul_90_22_n_1005 ,mul_90_22_n_1030);
  or mul_90_22_g2975(mul_90_22_n_1055 ,mul_90_22_n_997 ,mul_90_22_n_1025);
  and mul_90_22_g2976(mul_90_22_n_1054 ,mul_90_22_n_1007 ,mul_90_22_n_1029);
  and mul_90_22_g2977(mul_90_22_n_1053 ,mul_90_22_n_991 ,mul_90_22_n_1028);
  not mul_90_22_g2978(mul_90_22_n_1047 ,mul_90_22_n_1046);
  or mul_90_22_g2979(mul_90_22_n_1044 ,mul_90_22_n_1010 ,mul_90_22_n_1020);
  and mul_90_22_g2980(mul_90_22_n_1043 ,mul_90_22_n_1010 ,mul_90_22_n_1020);
  or mul_90_22_g2981(mul_90_22_n_1042 ,mul_90_22_n_1009 ,mul_90_22_n_1021);
  and mul_90_22_g2982(mul_90_22_n_1041 ,mul_90_22_n_1009 ,mul_90_22_n_1021);
  xnor mul_90_22_g2983(mul_90_22_n_1040 ,mul_90_22_n_927 ,mul_90_22_n_995);
  xnor mul_90_22_g2984(mul_90_22_n_1048 ,mul_90_22_n_940 ,mul_90_22_n_2);
  xnor mul_90_22_g2985(mul_90_22_n_1046 ,mul_90_22_n_956 ,mul_90_22_n_983);
  xnor mul_90_22_g2986(mul_90_22_n_1045 ,mul_90_22_n_952 ,mul_90_22_n_985);
  not mul_90_22_g2987(mul_90_22_n_1037 ,mul_90_22_n_1036);
  not mul_90_22_g2988(mul_90_22_n_1033 ,mul_90_22_n_1032);
  nor mul_90_22_g2989(mul_90_22_n_1031 ,mul_90_22_n_920 ,mul_90_22_n_1002);
  and mul_90_22_g2990(mul_90_22_n_1030 ,mul_90_22_n_912 ,mul_90_22_n_987);
  or mul_90_22_g2991(mul_90_22_n_1029 ,mul_90_22_n_944 ,mul_90_22_n_1004);
  or mul_90_22_g2992(mul_90_22_n_1028 ,mul_90_22_n_945 ,mul_90_22_n_990);
  or mul_90_22_g2993(mul_90_22_n_1027 ,mul_90_22_n_927 ,mul_90_22_n_995);
  and mul_90_22_g2994(mul_90_22_n_1026 ,mul_90_22_n_927 ,mul_90_22_n_995);
  nor mul_90_22_g2995(mul_90_22_n_1025 ,mul_90_22_n_943 ,mul_90_22_n_1001);
  or mul_90_22_g2996(mul_90_22_n_1024 ,mul_90_22_n_929 ,mul_90_22_n_992);
  and mul_90_22_g2997(mul_90_22_n_1039 ,mul_90_22_n_973 ,mul_90_22_n_994);
  and mul_90_22_g2998(mul_90_22_n_1038 ,mul_90_22_n_969 ,mul_90_22_n_989);
  and mul_90_22_g2999(mul_90_22_n_1036 ,mul_90_22_n_971 ,mul_90_22_n_998);
  or mul_90_22_g3000(mul_90_22_n_1035 ,mul_90_22_n_976 ,mul_90_22_n_986);
  or mul_90_22_g3001(mul_90_22_n_1034 ,mul_90_22_n_978 ,mul_90_22_n_1006);
  or mul_90_22_g3002(mul_90_22_n_1032 ,mul_90_22_n_937 ,mul_90_22_n_1008);
  not mul_90_22_g3003(mul_90_22_n_1022 ,mul_90_22_n_1023);
  not mul_90_22_g3004(mul_90_22_n_1018 ,mul_90_22_n_1017);
  nor mul_90_22_g3006(mul_90_22_n_1016 ,mul_90_22_n_982 ,mul_90_22_n_996);
  xnor mul_90_22_g3007(mul_90_22_n_1015 ,mul_90_22_n_959 ,mul_90_22_n_862);
  xnor mul_90_22_g3008(mul_90_22_n_1014 ,mul_90_22_n_794 ,mul_90_22_n_954);
  xnor mul_90_22_g3009(mul_90_22_n_1013 ,mul_90_22_n_878 ,mul_90_22_n_962);
  xnor mul_90_22_g3010(mul_90_22_n_1012 ,mul_90_22_n_958 ,mul_90_22_n_885);
  xnor mul_90_22_g3011(mul_90_22_n_1011 ,mul_90_22_n_906 ,mul_90_22_n_961);
  xnor mul_90_22_g3014(mul_90_22_n_1023 ,mul_90_22_n_842 ,mul_90_22_n_947);
  xnor mul_90_22_g3015(mul_90_22_n_1021 ,mul_90_22_n_926 ,mul_90_22_n_946);
  xnor mul_90_22_g3016(mul_90_22_n_1020 ,mul_90_22_n_928 ,mul_90_22_n_948);
  or mul_90_22_g3017(mul_90_22_n_1019 ,mul_90_22_n_951 ,mul_90_22_n_988);
  xnor mul_90_22_g3018(mul_90_22_n_1017 ,mul_90_22_n_981 ,mul_90_22_n_949);
  and mul_90_22_g3020(mul_90_22_n_1008 ,mul_90_22_n_981 ,mul_90_22_n_931);
  or mul_90_22_g3021(mul_90_22_n_1007 ,mul_90_22_n_862 ,mul_90_22_n_959);
  and mul_90_22_g3022(mul_90_22_n_1006 ,mul_90_22_n_962 ,mul_90_22_n_977);
  nor mul_90_22_g3023(mul_90_22_n_1005 ,mul_90_22_n_182 ,mul_90_22_n_958);
  and mul_90_22_g3024(mul_90_22_n_1004 ,mul_90_22_n_862 ,mul_90_22_n_959);
  nor mul_90_22_g3025(mul_90_22_n_1003 ,mul_90_22_n_913 ,mul_90_22_n_966);
  nor mul_90_22_g3026(mul_90_22_n_1002 ,mul_90_22_n_935 ,mul_90_22_n_979);
  and mul_90_22_g3027(mul_90_22_n_1001 ,mul_90_22_n_886 ,mul_90_22_n_952);
  nor mul_90_22_g3028(mul_90_22_n_1000 ,mul_90_22_n_848 ,mul_90_22_n_965);
  nor mul_90_22_g3029(mul_90_22_n_999 ,mul_90_22_n_849 ,mul_90_22_n_964);
  or mul_90_22_g3030(mul_90_22_n_998 ,mul_90_22_n_970 ,mul_90_22_n_960);
  nor mul_90_22_g3031(mul_90_22_n_997 ,mul_90_22_n_886 ,mul_90_22_n_952);
  or mul_90_22_g3032(mul_90_22_n_1010 ,mul_90_22_n_923 ,mul_90_22_n_972);
  or mul_90_22_g3033(mul_90_22_n_1009 ,mul_90_22_n_918 ,mul_90_22_n_974);
  or mul_90_22_g3035(mul_90_22_n_994 ,mul_90_22_n_930 ,mul_90_22_n_980);
  or mul_90_22_g3036(mul_90_22_n_993 ,mul_90_22_n_884 ,mul_90_22_n_955);
  nor mul_90_22_g3037(mul_90_22_n_992 ,mul_90_22_n_883 ,mul_90_22_n_956);
  or mul_90_22_g3038(mul_90_22_n_991 ,mul_90_22_n_794 ,mul_90_22_n_953);
  nor mul_90_22_g3039(mul_90_22_n_990 ,mul_90_22_n_793 ,mul_90_22_n_954);
  or mul_90_22_g3040(mul_90_22_n_989 ,mul_90_22_n_968 ,mul_90_22_n_963);
  nor mul_90_22_g3041(mul_90_22_n_988 ,mul_90_22_n_950 ,mul_90_22_n_961);
  or mul_90_22_g3042(mul_90_22_n_987 ,mul_90_22_n_308 ,mul_90_22_n_957);
  nor mul_90_22_g3043(mul_90_22_n_986 ,mul_90_22_n_840 ,mul_90_22_n_975);
  xor mul_90_22_g3044(mul_90_22_n_985 ,mul_90_22_n_943 ,mul_90_22_n_886);
  xnor mul_90_22_g3046(mul_90_22_n_984 ,mul_90_22_n_0 ,mul_90_22_n_916);
  xnor mul_90_22_g3047(mul_90_22_n_996 ,mul_90_22_n_876 ,mul_90_22_n_1);
  xnor mul_90_22_g3048(mul_90_22_n_983 ,mul_90_22_n_929 ,mul_90_22_n_884);
  or mul_90_22_g3049(mul_90_22_n_995 ,mul_90_22_n_933 ,mul_90_22_n_967);
  and mul_90_22_g3051(mul_90_22_n_980 ,mul_90_22_n_890 ,mul_90_22_n_940);
  and mul_90_22_g3052(mul_90_22_n_979 ,mul_90_22_n_802 ,mul_90_22_n_934);
  nor mul_90_22_g3053(mul_90_22_n_978 ,mul_90_22_n_878 ,mul_90_22_n_939);
  or mul_90_22_g3054(mul_90_22_n_977 ,mul_90_22_n_877 ,mul_90_22_n_938);
  nor mul_90_22_g3055(mul_90_22_n_976 ,mul_90_22_n_905 ,mul_90_22_n_926);
  and mul_90_22_g3056(mul_90_22_n_975 ,mul_90_22_n_905 ,mul_90_22_n_926);
  and mul_90_22_g3057(mul_90_22_n_974 ,mul_90_22_n_928 ,mul_90_22_n_917);
  or mul_90_22_g3058(mul_90_22_n_973 ,mul_90_22_n_890 ,mul_90_22_n_940);
  nor mul_90_22_g3059(mul_90_22_n_972 ,mul_90_22_n_847 ,mul_90_22_n_919);
  or mul_90_22_g3060(mul_90_22_n_971 ,mul_90_22_n_889 ,mul_90_22_n_942);
  and mul_90_22_g3061(mul_90_22_n_970 ,mul_90_22_n_889 ,mul_90_22_n_942);
  or mul_90_22_g3062(mul_90_22_n_969 ,mul_90_22_n_882 ,mul_90_22_n_924);
  nor mul_90_22_g3063(mul_90_22_n_968 ,mul_90_22_n_881 ,mul_90_22_n_925);
  and mul_90_22_g3064(mul_90_22_n_967 ,mul_90_22_n_842 ,mul_90_22_n_936);
  or mul_90_22_g3065(mul_90_22_n_982 ,mul_90_22_n_705 ,mul_90_22_n_922);
  or mul_90_22_g3066(mul_90_22_n_981 ,mul_90_22_n_746 ,mul_90_22_n_932);
  not mul_90_22_g3068(mul_90_22_n_965 ,mul_90_22_n_964);
  not mul_90_22_g3071(mul_90_22_n_958 ,mul_90_22_n_957);
  not mul_90_22_g3072(mul_90_22_n_956 ,mul_90_22_n_955);
  not mul_90_22_g3073(mul_90_22_n_953 ,mul_90_22_n_954);
  nor mul_90_22_g3074(mul_90_22_n_951 ,mul_90_22_n_907 ,mul_90_22_n_941);
  and mul_90_22_g3075(mul_90_22_n_950 ,mul_90_22_n_907 ,mul_90_22_n_941);
  xnor mul_90_22_g3076(mul_90_22_n_966 ,mul_90_22_n_910 ,mul_90_22_n_780);
  xnor mul_90_22_g3077(mul_90_22_n_964 ,mul_90_22_n_602 ,mul_90_22_n_875);
  xnor mul_90_22_g3078(mul_90_22_n_949 ,mul_90_22_n_888 ,mul_90_22_n_839);
  xnor mul_90_22_g3079(mul_90_22_n_948 ,mul_90_22_n_880 ,mul_90_22_n_909);
  xnor mul_90_22_g3080(mul_90_22_n_947 ,mul_90_22_n_904 ,mul_90_22_n_649);
  xor mul_90_22_g3081(mul_90_22_n_946 ,mul_90_22_n_905 ,mul_90_22_n_840);
  xnor mul_90_22_g3082(mul_90_22_n_963 ,mul_90_22_n_841 ,mul_90_22_n_868);
  xnor mul_90_22_g3083(mul_90_22_n_962 ,mul_90_22_n_867 ,mul_90_22_n_870);
  xnor mul_90_22_g3084(mul_90_22_n_961 ,mul_90_22_n_866 ,mul_90_22_n_869);
  xnor mul_90_22_g3085(mul_90_22_n_960 ,mul_90_22_n_845 ,mul_90_22_n_874);
  xnor mul_90_22_g3086(mul_90_22_n_959 ,mul_90_22_n_911 ,mul_90_22_n_787);
  xnor mul_90_22_g3087(mul_90_22_n_957 ,mul_90_22_n_865 ,mul_90_22_n_872);
  xnor mul_90_22_g3088(mul_90_22_n_955 ,mul_90_22_n_762 ,mul_90_22_n_871);
  xnor mul_90_22_g3089(mul_90_22_n_954 ,mul_90_22_n_843 ,mul_90_22_n_893);
  xnor mul_90_22_g3090(mul_90_22_n_952 ,mul_90_22_n_864 ,mul_90_22_n_873);
  not mul_90_22_g3091(mul_90_22_n_939 ,mul_90_22_n_938);
  nor mul_90_22_g3092(mul_90_22_n_937 ,mul_90_22_n_839 ,mul_90_22_n_888);
  or mul_90_22_g3093(mul_90_22_n_936 ,mul_90_22_n_204 ,mul_90_22_n_904);
  nor mul_90_22_g3094(mul_90_22_n_935 ,mul_90_22_n_643 ,mul_90_22_n_914);
  or mul_90_22_g3095(mul_90_22_n_934 ,mul_90_22_n_644 ,mul_90_22_n_915);
  and mul_90_22_g3096(mul_90_22_n_933 ,mul_90_22_n_203 ,mul_90_22_n_904);
  and mul_90_22_g3097(mul_90_22_n_932 ,mul_90_22_n_755 ,mul_90_22_n_911);
  or mul_90_22_g3098(mul_90_22_n_931 ,mul_90_22_n_838 ,mul_90_22_n_887);
  and mul_90_22_g3099(mul_90_22_n_945 ,mul_90_22_n_754 ,mul_90_22_n_899);
  and mul_90_22_g3100(mul_90_22_n_944 ,mul_90_22_n_804 ,mul_90_22_n_897);
  and mul_90_22_g3101(mul_90_22_n_943 ,mul_90_22_n_857 ,mul_90_22_n_901);
  and mul_90_22_g3102(mul_90_22_n_942 ,mul_90_22_n_861 ,mul_90_22_n_902);
  and mul_90_22_g3103(mul_90_22_n_941 ,mul_90_22_n_832 ,mul_90_22_n_898);
  and mul_90_22_g3104(mul_90_22_n_940 ,mul_90_22_n_855 ,mul_90_22_n_903);
  or mul_90_22_g3105(mul_90_22_n_938 ,mul_90_22_n_854 ,mul_90_22_n_900);
  not mul_90_22_g3107(mul_90_22_n_924 ,mul_90_22_n_925);
  nor mul_90_22_g3108(mul_90_22_n_923 ,mul_90_22_n_599 ,mul_90_22_n_876);
  and mul_90_22_g3109(mul_90_22_n_922 ,mul_90_22_n_704 ,mul_90_22_n_910);
  nor mul_90_22_g3110(mul_90_22_n_921 ,mul_90_22_n_769 ,mul_90_22_n_891);
  nor mul_90_22_g3111(mul_90_22_n_920 ,mul_90_22_n_768 ,mul_90_22_n_892);
  and mul_90_22_g3112(mul_90_22_n_919 ,mul_90_22_n_599 ,mul_90_22_n_876);
  nor mul_90_22_g3113(mul_90_22_n_918 ,mul_90_22_n_909 ,mul_90_22_n_880);
  or mul_90_22_g3114(mul_90_22_n_917 ,mul_90_22_n_908 ,mul_90_22_n_879);
  or mul_90_22_g3116(mul_90_22_n_916 ,mul_90_22_n_719 ,mul_90_22_n_894);
  xnor mul_90_22_g3117(mul_90_22_n_930 ,mul_90_22_n_844 ,mul_90_22_n_830);
  and mul_90_22_g3118(mul_90_22_n_929 ,mul_90_22_n_851 ,mul_90_22_n_895);
  xnor mul_90_22_g3119(mul_90_22_n_928 ,mul_90_22_n_606 ,mul_90_22_n_831);
  xnor mul_90_22_g3120(mul_90_22_n_927 ,mul_90_22_n_863 ,mul_90_22_n_782);
  xnor mul_90_22_g3121(mul_90_22_n_926 ,mul_90_22_n_846 ,mul_90_22_n_783);
  or mul_90_22_g3122(mul_90_22_n_925 ,mul_90_22_n_835 ,mul_90_22_n_896);
  not mul_90_22_g3123(mul_90_22_n_915 ,mul_90_22_n_914);
  not mul_90_22_g3125(mul_90_22_n_908 ,mul_90_22_n_909);
  not mul_90_22_g3126(mul_90_22_n_907 ,mul_90_22_n_906);
  or mul_90_22_g3127(mul_90_22_n_903 ,mul_90_22_n_858 ,mul_90_22_n_867);
  or mul_90_22_g3128(mul_90_22_n_902 ,mul_90_22_n_860 ,mul_90_22_n_864);
  or mul_90_22_g3129(mul_90_22_n_901 ,mul_90_22_n_856 ,mul_90_22_n_865);
  nor mul_90_22_g3130(mul_90_22_n_900 ,mul_90_22_n_852 ,mul_90_22_n_866);
  or mul_90_22_g3131(mul_90_22_n_899 ,mul_90_22_n_726 ,mul_90_22_n_846);
  or mul_90_22_g3132(mul_90_22_n_898 ,mul_90_22_n_837 ,mul_90_22_n_841);
  or mul_90_22_g3133(mul_90_22_n_897 ,mul_90_22_n_803 ,mul_90_22_n_844);
  nor mul_90_22_g3134(mul_90_22_n_896 ,mul_90_22_n_834 ,mul_90_22_n_845);
  or mul_90_22_g3135(mul_90_22_n_895 ,mul_90_22_n_843 ,mul_90_22_n_850);
  and mul_90_22_g3136(mul_90_22_n_894 ,mul_90_22_n_720 ,mul_90_22_n_863);
  and mul_90_22_g3137(mul_90_22_n_914 ,mul_90_22_n_753 ,mul_90_22_n_859);
  xnor mul_90_22_g3138(mul_90_22_n_893 ,mul_90_22_n_663 ,mul_90_22_n_792);
  xnor mul_90_22_g3139(mul_90_22_n_913 ,mul_90_22_n_731 ,mul_90_22_n_774);
  or mul_90_22_g3140(mul_90_22_n_912 ,mul_90_22_n_816 ,mul_90_22_n_853);
  xnor mul_90_22_g3141(mul_90_22_n_911 ,mul_90_22_n_692 ,mul_90_22_n_800);
  or mul_90_22_g3142(mul_90_22_n_910 ,mul_90_22_n_703 ,mul_90_22_n_833);
  and mul_90_22_g3143(mul_90_22_n_909 ,mul_90_22_n_713 ,mul_90_22_n_836);
  xnor mul_90_22_g3144(mul_90_22_n_906 ,mul_90_22_n_672 ,mul_90_22_n_785);
  xnor mul_90_22_g3145(mul_90_22_n_905 ,mul_90_22_n_661 ,mul_90_22_n_779);
  xnor mul_90_22_g3146(mul_90_22_n_904 ,mul_90_22_n_687 ,mul_90_22_n_777);
  not mul_90_22_g3147(mul_90_22_n_892 ,mul_90_22_n_891);
  not mul_90_22_g3148(mul_90_22_n_888 ,mul_90_22_n_887);
  not mul_90_22_g3150(mul_90_22_n_883 ,mul_90_22_n_884);
  not mul_90_22_g3151(mul_90_22_n_881 ,mul_90_22_n_882);
  not mul_90_22_g3152(mul_90_22_n_879 ,mul_90_22_n_880);
  not mul_90_22_g3153(mul_90_22_n_877 ,mul_90_22_n_878);
  xnor mul_90_22_g3154(mul_90_22_n_875 ,mul_90_22_n_618 ,mul_90_22_n_797);
  xnor mul_90_22_g3155(mul_90_22_n_874 ,mul_90_22_n_758 ,mul_90_22_n_796);
  xnor mul_90_22_g3156(mul_90_22_n_873 ,mul_90_22_n_764 ,mul_90_22_n_829);
  xnor mul_90_22_g3157(mul_90_22_n_872 ,mul_90_22_n_760 ,mul_90_22_n_827);
  xnor mul_90_22_g3158(mul_90_22_n_871 ,mul_90_22_n_767 ,mul_90_22_n_799);
  xnor mul_90_22_g3159(mul_90_22_n_870 ,mul_90_22_n_757 ,mul_90_22_n_825);
  xnor mul_90_22_g3160(mul_90_22_n_869 ,mul_90_22_n_765 ,mul_90_22_n_795);
  xnor mul_90_22_g3161(mul_90_22_n_868 ,mul_90_22_n_730 ,mul_90_22_n_790);
  xnor mul_90_22_g3162(mul_90_22_n_891 ,mul_90_22_n_641 ,mul_90_22_n_775);
  xnor mul_90_22_g3164(mul_90_22_n_890 ,mul_90_22_n_697 ,mul_90_22_n_781);
  xnor mul_90_22_g3165(mul_90_22_n_889 ,mul_90_22_n_608 ,mul_90_22_n_778);
  xnor mul_90_22_g3166(mul_90_22_n_887 ,mul_90_22_n_786 ,mul_90_22_n_204);
  xnor mul_90_22_g3167(mul_90_22_n_886 ,mul_90_22_n_621 ,mul_90_22_n_773);
  xnor mul_90_22_g3168(mul_90_22_n_885 ,mul_90_22_n_632 ,mul_90_22_n_771);
  xnor mul_90_22_g3169(mul_90_22_n_884 ,mul_90_22_n_627 ,mul_90_22_n_770);
  xnor mul_90_22_g3170(mul_90_22_n_882 ,mul_90_22_n_664 ,mul_90_22_n_788);
  xnor mul_90_22_g3171(mul_90_22_n_880 ,mul_90_22_n_631 ,mul_90_22_n_776);
  xnor mul_90_22_g3172(mul_90_22_n_878 ,mul_90_22_n_633 ,mul_90_22_n_772);
  xnor mul_90_22_g3173(mul_90_22_n_876 ,mul_90_22_n_798 ,mul_90_22_n_784);
  or mul_90_22_g3174(mul_90_22_n_861 ,mul_90_22_n_763 ,mul_90_22_n_828);
  nor mul_90_22_g3175(mul_90_22_n_860 ,mul_90_22_n_764 ,mul_90_22_n_829);
  or mul_90_22_g3176(mul_90_22_n_859 ,mul_90_22_n_821 ,mul_90_22_n_751);
  nor mul_90_22_g3177(mul_90_22_n_858 ,mul_90_22_n_757 ,mul_90_22_n_824);
  or mul_90_22_g3178(mul_90_22_n_857 ,mul_90_22_n_760 ,mul_90_22_n_826);
  nor mul_90_22_g3179(mul_90_22_n_856 ,mul_90_22_n_759 ,mul_90_22_n_827);
  or mul_90_22_g3180(mul_90_22_n_855 ,mul_90_22_n_756 ,mul_90_22_n_825);
  and mul_90_22_g3181(mul_90_22_n_854 ,mul_90_22_n_765 ,mul_90_22_n_795);
  and mul_90_22_g3182(mul_90_22_n_853 ,mul_90_22_n_799 ,mul_90_22_n_815);
  nor mul_90_22_g3183(mul_90_22_n_852 ,mul_90_22_n_765 ,mul_90_22_n_795);
  or mul_90_22_g3184(mul_90_22_n_851 ,mul_90_22_n_663 ,mul_90_22_n_791);
  nor mul_90_22_g3185(mul_90_22_n_850 ,mul_90_22_n_662 ,mul_90_22_n_792);
  and mul_90_22_g3186(mul_90_22_n_867 ,mul_90_22_n_715 ,mul_90_22_n_820);
  and mul_90_22_g3187(mul_90_22_n_866 ,mul_90_22_n_736 ,mul_90_22_n_814);
  and mul_90_22_g3188(mul_90_22_n_865 ,mul_90_22_n_743 ,mul_90_22_n_817);
  and mul_90_22_g3189(mul_90_22_n_864 ,mul_90_22_n_752 ,mul_90_22_n_819);
  or mul_90_22_g3190(mul_90_22_n_863 ,mul_90_22_n_741 ,mul_90_22_n_818);
  and mul_90_22_g3191(mul_90_22_n_862 ,mul_90_22_n_737 ,mul_90_22_n_813);
  not mul_90_22_g3192(mul_90_22_n_849 ,mul_90_22_n_848);
  not mul_90_22_g3193(mul_90_22_n_838 ,mul_90_22_n_839);
  nor mul_90_22_g3194(mul_90_22_n_837 ,mul_90_22_n_730 ,mul_90_22_n_790);
  or mul_90_22_g3195(mul_90_22_n_836 ,mul_90_22_n_711 ,mul_90_22_n_798);
  and mul_90_22_g3196(mul_90_22_n_835 ,mul_90_22_n_758 ,mul_90_22_n_796);
  nor mul_90_22_g3197(mul_90_22_n_834 ,mul_90_22_n_758 ,mul_90_22_n_796);
  and mul_90_22_g3198(mul_90_22_n_833 ,mul_90_22_n_750 ,mul_90_22_n_797);
  or mul_90_22_g3199(mul_90_22_n_832 ,mul_90_22_n_729 ,mul_90_22_n_789);
  and mul_90_22_g3200(mul_90_22_n_848 ,mul_90_22_n_747 ,mul_90_22_n_822);
  xnor mul_90_22_g3201(mul_90_22_n_831 ,mul_90_22_n_598 ,mul_90_22_n_733);
  xnor mul_90_22_g3202(mul_90_22_n_830 ,mul_90_22_n_728 ,mul_90_22_n_648);
  and mul_90_22_g3203(mul_90_22_n_847 ,mul_90_22_n_709 ,mul_90_22_n_809);
  and mul_90_22_g3204(mul_90_22_n_846 ,mul_90_22_n_735 ,mul_90_22_n_812);
  and mul_90_22_g3205(mul_90_22_n_845 ,mul_90_22_n_710 ,mul_90_22_n_808);
  and mul_90_22_g3206(mul_90_22_n_844 ,mul_90_22_n_745 ,mul_90_22_n_807);
  and mul_90_22_g3207(mul_90_22_n_843 ,mul_90_22_n_738 ,mul_90_22_n_806);
  or mul_90_22_g3208(mul_90_22_n_842 ,mul_90_22_n_725 ,mul_90_22_n_805);
  and mul_90_22_g3209(mul_90_22_n_841 ,mul_90_22_n_722 ,mul_90_22_n_811);
  and mul_90_22_g3210(mul_90_22_n_840 ,mul_90_22_n_721 ,mul_90_22_n_810);
  and mul_90_22_g3211(mul_90_22_n_839 ,mul_90_22_n_706 ,mul_90_22_n_823);
  not mul_90_22_g3212(mul_90_22_n_828 ,mul_90_22_n_829);
  not mul_90_22_g3213(mul_90_22_n_826 ,mul_90_22_n_827);
  not mul_90_22_g3214(mul_90_22_n_824 ,mul_90_22_n_825);
  or mul_90_22_g3215(mul_90_22_n_823 ,mul_90_22_n_692 ,mul_90_22_n_749);
  or mul_90_22_g3216(mul_90_22_n_822 ,mul_90_22_n_641 ,mul_90_22_n_716);
  or mul_90_22_g3217(mul_90_22_n_821 ,mul_90_22_n_327 ,mul_90_22_n_727);
  or mul_90_22_g3218(mul_90_22_n_820 ,mul_90_22_n_630 ,mul_90_22_n_744);
  or mul_90_22_g3219(mul_90_22_n_819 ,mul_90_22_n_632 ,mul_90_22_n_718);
  and mul_90_22_g3220(mul_90_22_n_818 ,mul_90_22_n_687 ,mul_90_22_n_748);
  or mul_90_22_g3221(mul_90_22_n_817 ,mul_90_22_n_627 ,mul_90_22_n_742);
  nor mul_90_22_g3222(mul_90_22_n_816 ,mul_90_22_n_767 ,mul_90_22_n_761);
  or mul_90_22_g3223(mul_90_22_n_815 ,mul_90_22_n_766 ,mul_90_22_n_762);
  or mul_90_22_g3224(mul_90_22_n_814 ,mul_90_22_n_624 ,mul_90_22_n_739);
  or mul_90_22_g3225(mul_90_22_n_813 ,mul_90_22_n_697 ,mul_90_22_n_723);
  or mul_90_22_g3226(mul_90_22_n_812 ,mul_90_22_n_631 ,mul_90_22_n_724);
  or mul_90_22_g3227(mul_90_22_n_811 ,mul_90_22_n_622 ,mul_90_22_n_714);
  or mul_90_22_g3228(mul_90_22_n_810 ,mul_90_22_n_734 ,mul_90_22_n_717);
  or mul_90_22_g3229(mul_90_22_n_809 ,mul_90_22_n_708 ,mul_90_22_n_732);
  or mul_90_22_g3230(mul_90_22_n_808 ,mul_90_22_n_621 ,mul_90_22_n_707);
  or mul_90_22_g3231(mul_90_22_n_807 ,mul_90_22_n_633 ,mul_90_22_n_702);
  or mul_90_22_g3232(mul_90_22_n_806 ,mul_90_22_n_623 ,mul_90_22_n_740);
  nor mul_90_22_g3233(mul_90_22_n_805 ,mul_90_22_n_203 ,mul_90_22_n_712);
  or mul_90_22_g3234(mul_90_22_n_804 ,mul_90_22_n_156 ,mul_90_22_n_728);
  and mul_90_22_g3235(mul_90_22_n_803 ,mul_90_22_n_157 ,mul_90_22_n_728);
  xnor mul_90_22_g3236(mul_90_22_n_802 ,mul_90_22_n_698 ,mul_90_22_n_547);
  xnor mul_90_22_g3237(mul_90_22_n_801 ,mul_90_22_n_647 ,mul_90_22_n_646);
  xnor mul_90_22_g3238(mul_90_22_n_800 ,mul_90_22_n_604 ,mul_90_22_n_656);
  xnor mul_90_22_g3239(mul_90_22_n_829 ,mul_90_22_n_628 ,mul_90_22_n_636);
  xnor mul_90_22_g3240(mul_90_22_n_827 ,mul_90_22_n_679 ,mul_90_22_n_696);
  xnor mul_90_22_g3241(mul_90_22_n_825 ,mul_90_22_n_645 ,mul_90_22_n_700);
  not mul_90_22_g3242(mul_90_22_n_793 ,mul_90_22_n_794);
  not mul_90_22_g3243(mul_90_22_n_791 ,mul_90_22_n_792);
  not mul_90_22_g3244(mul_90_22_n_789 ,mul_90_22_n_790);
  xnor mul_90_22_g3245(mul_90_22_n_788 ,mul_90_22_n_667 ,mul_90_22_n_624);
  xnor mul_90_22_g3246(mul_90_22_n_787 ,mul_90_22_n_677 ,mul_90_22_n_157);
  xnor mul_90_22_g3247(mul_90_22_n_786 ,mul_90_22_n_670 ,mul_90_22_n_611);
  xor mul_90_22_g3248(mul_90_22_n_785 ,mul_90_22_n_666 ,mul_90_22_n_630);
  xnor mul_90_22_g3249(mul_90_22_n_784 ,mul_90_22_n_609 ,mul_90_22_n_669);
  xnor mul_90_22_g3250(mul_90_22_n_783 ,mul_90_22_n_674 ,mul_90_22_n_654);
  xnor mul_90_22_g3251(mul_90_22_n_782 ,mul_90_22_n_614 ,mul_90_22_n_650);
  xnor mul_90_22_g3252(mul_90_22_n_781 ,mul_90_22_n_657 ,mul_90_22_n_612);
  xnor mul_90_22_g3253(mul_90_22_n_780 ,mul_90_22_n_594 ,mul_90_22_n_596);
  xor mul_90_22_g3254(mul_90_22_n_779 ,mul_90_22_n_659 ,mul_90_22_n_623);
  xnor mul_90_22_g3255(mul_90_22_n_778 ,mul_90_22_n_600 ,mul_90_22_n_622);
  xnor mul_90_22_g3256(mul_90_22_n_777 ,mul_90_22_n_616 ,mul_90_22_n_653);
  xnor mul_90_22_g3257(mul_90_22_n_776 ,mul_90_22_n_449 ,mul_90_22_n_673);
  xnor mul_90_22_g3258(mul_90_22_n_775 ,mul_90_22_n_451 ,mul_90_22_n_651);
  xnor mul_90_22_g3259(mul_90_22_n_774 ,mul_90_22_n_450 ,mul_90_22_n_605);
  xnor mul_90_22_g3260(mul_90_22_n_773 ,mul_90_22_n_592 ,mul_90_22_n_597);
  xnor mul_90_22_g3261(mul_90_22_n_772 ,mul_90_22_n_607 ,mul_90_22_n_665);
  xnor mul_90_22_g3262(mul_90_22_n_771 ,mul_90_22_n_610 ,mul_90_22_n_668);
  xnor mul_90_22_g3263(mul_90_22_n_770 ,mul_90_22_n_678 ,mul_90_22_n_675);
  xnor mul_90_22_g3264(mul_90_22_n_799 ,mul_90_22_n_684 ,mul_90_22_n_682);
  xnor mul_90_22_g3265(mul_90_22_n_798 ,mul_90_22_n_639 ,mul_90_22_n_544);
  xnor mul_90_22_g3266(mul_90_22_n_797 ,mul_90_22_n_546 ,mul_90_22_n_634);
  xnor mul_90_22_g3267(mul_90_22_n_796 ,mul_90_22_n_619 ,mul_90_22_n_629);
  xnor mul_90_22_g3268(mul_90_22_n_795 ,mul_90_22_n_694 ,mul_90_22_n_693);
  xnor mul_90_22_g3269(mul_90_22_n_794 ,mul_90_22_n_690 ,mul_90_22_n_625);
  xnor mul_90_22_g3270(mul_90_22_n_792 ,mul_90_22_n_681 ,mul_90_22_n_685);
  xnor mul_90_22_g3271(mul_90_22_n_790 ,mul_90_22_n_638 ,mul_90_22_n_688);
  not mul_90_22_g3272(mul_90_22_n_769 ,mul_90_22_n_768);
  not mul_90_22_g3273(mul_90_22_n_767 ,mul_90_22_n_766);
  not mul_90_22_g3274(mul_90_22_n_764 ,mul_90_22_n_763);
  not mul_90_22_g3275(mul_90_22_n_761 ,mul_90_22_n_762);
  not mul_90_22_g3276(mul_90_22_n_760 ,mul_90_22_n_759);
  not mul_90_22_g3277(mul_90_22_n_757 ,mul_90_22_n_756);
  or mul_90_22_g3278(mul_90_22_n_755 ,mul_90_22_n_156 ,mul_90_22_n_676);
  or mul_90_22_g3279(mul_90_22_n_754 ,mul_90_22_n_654 ,mul_90_22_n_674);
  or mul_90_22_g3280(mul_90_22_n_753 ,mul_90_22_n_456 ,mul_90_22_n_642);
  or mul_90_22_g3281(mul_90_22_n_752 ,mul_90_22_n_668 ,mul_90_22_n_610);
  and mul_90_22_g3282(mul_90_22_n_751 ,mul_90_22_n_456 ,mul_90_22_n_642);
  or mul_90_22_g3283(mul_90_22_n_750 ,mul_90_22_n_601 ,mul_90_22_n_617);
  nor mul_90_22_g3284(mul_90_22_n_749 ,mul_90_22_n_604 ,mul_90_22_n_655);
  or mul_90_22_g3285(mul_90_22_n_748 ,mul_90_22_n_652 ,mul_90_22_n_615);
  or mul_90_22_g3286(mul_90_22_n_747 ,mul_90_22_n_451 ,mul_90_22_n_651);
  nor mul_90_22_g3287(mul_90_22_n_746 ,mul_90_22_n_306 ,mul_90_22_n_677);
  or mul_90_22_g3288(mul_90_22_n_745 ,mul_90_22_n_665 ,mul_90_22_n_607);
  and mul_90_22_g3289(mul_90_22_n_744 ,mul_90_22_n_672 ,mul_90_22_n_666);
  or mul_90_22_g3290(mul_90_22_n_743 ,mul_90_22_n_675 ,mul_90_22_n_678);
  and mul_90_22_g3291(mul_90_22_n_742 ,mul_90_22_n_675 ,mul_90_22_n_678);
  nor mul_90_22_g3292(mul_90_22_n_741 ,mul_90_22_n_653 ,mul_90_22_n_616);
  nor mul_90_22_g3293(mul_90_22_n_740 ,mul_90_22_n_661 ,mul_90_22_n_658);
  and mul_90_22_g3294(mul_90_22_n_739 ,mul_90_22_n_667 ,mul_90_22_n_664);
  or mul_90_22_g3295(mul_90_22_n_738 ,mul_90_22_n_660 ,mul_90_22_n_659);
  or mul_90_22_g3296(mul_90_22_n_737 ,mul_90_22_n_612 ,mul_90_22_n_657);
  or mul_90_22_g3297(mul_90_22_n_736 ,mul_90_22_n_667 ,mul_90_22_n_664);
  or mul_90_22_g3298(mul_90_22_n_735 ,mul_90_22_n_449 ,mul_90_22_n_673);
  and mul_90_22_g3299(mul_90_22_n_768 ,mul_90_22_n_547 ,mul_90_22_n_699);
  and mul_90_22_g3300(mul_90_22_n_766 ,mul_90_22_n_681 ,mul_90_22_n_686);
  and mul_90_22_g3301(mul_90_22_n_765 ,mul_90_22_n_638 ,mul_90_22_n_689);
  or mul_90_22_g3302(mul_90_22_n_763 ,mul_90_22_n_680 ,mul_90_22_n_696);
  and mul_90_22_g3303(mul_90_22_n_762 ,mul_90_22_n_626 ,mul_90_22_n_691);
  and mul_90_22_g3304(mul_90_22_n_759 ,mul_90_22_n_684 ,mul_90_22_n_683);
  and mul_90_22_g3305(mul_90_22_n_758 ,mul_90_22_n_628 ,mul_90_22_n_637);
  or mul_90_22_g3306(mul_90_22_n_756 ,mul_90_22_n_695 ,mul_90_22_n_693);
  not mul_90_22_g3307(mul_90_22_n_734 ,mul_90_22_n_733);
  not mul_90_22_g3308(mul_90_22_n_732 ,mul_90_22_n_731);
  not mul_90_22_g3309(mul_90_22_n_730 ,mul_90_22_n_729);
  or mul_90_22_g3310(mul_90_22_n_727 ,mul_90_22_n_311 ,mul_90_22_n_591);
  and mul_90_22_g3311(mul_90_22_n_726 ,mul_90_22_n_654 ,mul_90_22_n_674);
  nor mul_90_22_g3312(mul_90_22_n_725 ,mul_90_22_n_671 ,mul_90_22_n_611);
  and mul_90_22_g3313(mul_90_22_n_724 ,mul_90_22_n_449 ,mul_90_22_n_673);
  and mul_90_22_g3314(mul_90_22_n_723 ,mul_90_22_n_612 ,mul_90_22_n_657);
  or mul_90_22_g3315(mul_90_22_n_722 ,mul_90_22_n_600 ,mul_90_22_n_608);
  or mul_90_22_g3316(mul_90_22_n_721 ,mul_90_22_n_598 ,mul_90_22_n_606);
  or mul_90_22_g3317(mul_90_22_n_720 ,mul_90_22_n_307 ,mul_90_22_n_613);
  nor mul_90_22_g3318(mul_90_22_n_719 ,mul_90_22_n_650 ,mul_90_22_n_614);
  and mul_90_22_g3319(mul_90_22_n_718 ,mul_90_22_n_668 ,mul_90_22_n_610);
  and mul_90_22_g3320(mul_90_22_n_717 ,mul_90_22_n_598 ,mul_90_22_n_606);
  and mul_90_22_g3321(mul_90_22_n_716 ,mul_90_22_n_451 ,mul_90_22_n_651);
  or mul_90_22_g3322(mul_90_22_n_715 ,mul_90_22_n_672 ,mul_90_22_n_666);
  and mul_90_22_g3323(mul_90_22_n_714 ,mul_90_22_n_600 ,mul_90_22_n_608);
  or mul_90_22_g3324(mul_90_22_n_713 ,mul_90_22_n_669 ,mul_90_22_n_609);
  and mul_90_22_g3325(mul_90_22_n_712 ,mul_90_22_n_671 ,mul_90_22_n_611);
  and mul_90_22_g3326(mul_90_22_n_711 ,mul_90_22_n_669 ,mul_90_22_n_609);
  or mul_90_22_g3327(mul_90_22_n_710 ,mul_90_22_n_597 ,mul_90_22_n_592);
  or mul_90_22_g3328(mul_90_22_n_709 ,mul_90_22_n_450 ,mul_90_22_n_605);
  and mul_90_22_g3329(mul_90_22_n_708 ,mul_90_22_n_450 ,mul_90_22_n_605);
  and mul_90_22_g3330(mul_90_22_n_707 ,mul_90_22_n_597 ,mul_90_22_n_592);
  or mul_90_22_g3331(mul_90_22_n_706 ,mul_90_22_n_603 ,mul_90_22_n_656);
  nor mul_90_22_g3332(mul_90_22_n_705 ,mul_90_22_n_596 ,mul_90_22_n_594);
  or mul_90_22_g3333(mul_90_22_n_704 ,mul_90_22_n_595 ,mul_90_22_n_593);
  nor mul_90_22_g3334(mul_90_22_n_703 ,mul_90_22_n_602 ,mul_90_22_n_618);
  and mul_90_22_g3335(mul_90_22_n_702 ,mul_90_22_n_665 ,mul_90_22_n_607);
  and mul_90_22_g3336(mul_90_22_n_733 ,mul_90_22_n_545 ,mul_90_22_n_640);
  and mul_90_22_g3337(mul_90_22_n_731 ,mul_90_22_n_546 ,mul_90_22_n_635);
  or mul_90_22_g3338(mul_90_22_n_729 ,mul_90_22_n_620 ,mul_90_22_n_629);
  and mul_90_22_g3339(mul_90_22_n_728 ,mul_90_22_n_645 ,mul_90_22_n_701);
  not mul_90_22_g3340(mul_90_22_n_701 ,mul_90_22_n_700);
  not mul_90_22_g3341(mul_90_22_n_699 ,mul_90_22_n_698);
  not mul_90_22_g3342(mul_90_22_n_695 ,mul_90_22_n_694);
  not mul_90_22_g3343(mul_90_22_n_691 ,mul_90_22_n_690);
  not mul_90_22_g3344(mul_90_22_n_689 ,mul_90_22_n_688);
  not mul_90_22_g3345(mul_90_22_n_686 ,mul_90_22_n_685);
  not mul_90_22_g3346(mul_90_22_n_683 ,mul_90_22_n_682);
  not mul_90_22_g3347(mul_90_22_n_680 ,mul_90_22_n_679);
  not mul_90_22_g3348(mul_90_22_n_676 ,mul_90_22_n_677);
  not mul_90_22_g3349(mul_90_22_n_671 ,mul_90_22_n_670);
  not mul_90_22_g3350(mul_90_22_n_662 ,mul_90_22_n_663);
  not mul_90_22_g3351(mul_90_22_n_660 ,mul_90_22_n_661);
  not mul_90_22_g3352(mul_90_22_n_658 ,mul_90_22_n_659);
  not mul_90_22_g3353(mul_90_22_n_655 ,mul_90_22_n_656);
  not mul_90_22_g3354(mul_90_22_n_652 ,mul_90_22_n_653);
  or mul_90_22_g3358(mul_90_22_n_700 ,mul_90_22_n_502 ,mul_90_22_n_578);
  and mul_90_22_g3359(mul_90_22_n_698 ,mul_90_22_n_422 ,mul_90_22_n_536);
  or mul_90_22_g3360(mul_90_22_n_647 ,mul_90_22_n_457 ,mul_90_22_n_506);
  or mul_90_22_g3361(mul_90_22_n_646 ,mul_90_22_n_497 ,mul_90_22_n_580);
  and mul_90_22_g3362(mul_90_22_n_697 ,mul_90_22_n_429 ,mul_90_22_n_565);
  and mul_90_22_g3363(mul_90_22_n_696 ,mul_90_22_n_460 ,mul_90_22_n_561);
  or mul_90_22_g3364(mul_90_22_n_694 ,mul_90_22_n_500 ,mul_90_22_n_588);
  and mul_90_22_g3365(mul_90_22_n_693 ,mul_90_22_n_466 ,mul_90_22_n_573);
  and mul_90_22_g3366(mul_90_22_n_692 ,mul_90_22_n_461 ,mul_90_22_n_517);
  and mul_90_22_g3367(mul_90_22_n_690 ,mul_90_22_n_470 ,mul_90_22_n_526);
  and mul_90_22_g3368(mul_90_22_n_688 ,mul_90_22_n_472 ,mul_90_22_n_562);
  or mul_90_22_g3369(mul_90_22_n_687 ,mul_90_22_n_495 ,mul_90_22_n_587);
  and mul_90_22_g3370(mul_90_22_n_685 ,mul_90_22_n_412 ,mul_90_22_n_563);
  or mul_90_22_g3371(mul_90_22_n_684 ,mul_90_22_n_499 ,mul_90_22_n_585);
  and mul_90_22_g3372(mul_90_22_n_682 ,mul_90_22_n_441 ,mul_90_22_n_568);
  or mul_90_22_g3373(mul_90_22_n_681 ,mul_90_22_n_491 ,mul_90_22_n_582);
  or mul_90_22_g3374(mul_90_22_n_679 ,mul_90_22_n_501 ,mul_90_22_n_589);
  and mul_90_22_g3375(mul_90_22_n_678 ,mul_90_22_n_471 ,mul_90_22_n_528);
  and mul_90_22_g3376(mul_90_22_n_677 ,mul_90_22_n_440 ,mul_90_22_n_567);
  and mul_90_22_g3377(mul_90_22_n_675 ,mul_90_22_n_464 ,mul_90_22_n_529);
  and mul_90_22_g3378(mul_90_22_n_674 ,mul_90_22_n_467 ,mul_90_22_n_538);
  and mul_90_22_g3379(mul_90_22_n_673 ,mul_90_22_n_443 ,mul_90_22_n_555);
  and mul_90_22_g3380(mul_90_22_n_672 ,mul_90_22_n_459 ,mul_90_22_n_521);
  or mul_90_22_g3381(mul_90_22_n_670 ,mul_90_22_n_492 ,mul_90_22_n_579);
  and mul_90_22_g3382(mul_90_22_n_669 ,mul_90_22_n_434 ,mul_90_22_n_514);
  and mul_90_22_g3383(mul_90_22_n_668 ,mul_90_22_n_462 ,mul_90_22_n_535);
  and mul_90_22_g3384(mul_90_22_n_667 ,mul_90_22_n_473 ,mul_90_22_n_524);
  and mul_90_22_g3385(mul_90_22_n_666 ,mul_90_22_n_436 ,mul_90_22_n_533);
  and mul_90_22_g3386(mul_90_22_n_665 ,mul_90_22_n_432 ,mul_90_22_n_552);
  and mul_90_22_g3387(mul_90_22_n_664 ,mul_90_22_n_423 ,mul_90_22_n_523);
  and mul_90_22_g3388(mul_90_22_n_663 ,mul_90_22_n_426 ,mul_90_22_n_518);
  or mul_90_22_g3389(mul_90_22_n_661 ,mul_90_22_n_494 ,mul_90_22_n_540);
  and mul_90_22_g3390(mul_90_22_n_659 ,mul_90_22_n_433 ,mul_90_22_n_558);
  and mul_90_22_g3391(mul_90_22_n_657 ,mul_90_22_n_431 ,mul_90_22_n_531);
  or mul_90_22_g3392(mul_90_22_n_656 ,mul_90_22_n_454 ,mul_90_22_n_504);
  and mul_90_22_g3393(mul_90_22_n_654 ,mul_90_22_n_418 ,mul_90_22_n_527);
  or mul_90_22_g3394(mul_90_22_n_653 ,mul_90_22_n_452 ,mul_90_22_n_505);
  and mul_90_22_g3395(mul_90_22_n_651 ,mul_90_22_n_413 ,mul_90_22_n_532);
  or mul_90_22_g3396(mul_90_22_n_650 ,mul_90_22_n_493 ,mul_90_22_n_577);
  and mul_90_22_g3397(mul_90_22_n_649 ,mul_90_22_n_425 ,mul_90_22_n_559);
  or mul_90_22_g3398(mul_90_22_n_648 ,mul_90_22_n_498 ,mul_90_22_n_584);
  not mul_90_22_g3399(mul_90_22_n_644 ,mul_90_22_n_643);
  not mul_90_22_g3400(mul_90_22_n_640 ,mul_90_22_n_639);
  not mul_90_22_g3401(mul_90_22_n_637 ,mul_90_22_n_636);
  not mul_90_22_g3402(mul_90_22_n_635 ,mul_90_22_n_634);
  not mul_90_22_g3403(mul_90_22_n_626 ,mul_90_22_n_625);
  not mul_90_22_g3404(mul_90_22_n_620 ,mul_90_22_n_619);
  not mul_90_22_g3405(mul_90_22_n_617 ,mul_90_22_n_618);
  not mul_90_22_g3406(mul_90_22_n_615 ,mul_90_22_n_616);
  not mul_90_22_g3407(mul_90_22_n_613 ,mul_90_22_n_614);
  not mul_90_22_g3408(mul_90_22_n_603 ,mul_90_22_n_604);
  not mul_90_22_g3409(mul_90_22_n_601 ,mul_90_22_n_602);
  not mul_90_22_g3411(mul_90_22_n_595 ,mul_90_22_n_596);
  not mul_90_22_g3412(mul_90_22_n_593 ,mul_90_22_n_594);
  nor mul_90_22_g3413(mul_90_22_n_591 ,mul_90_22_n_486 ,mul_90_22_n_574);
  or mul_90_22_g3414(mul_90_22_n_645 ,mul_90_22_n_324 ,mul_90_22_n_507);
  and mul_90_22_g3415(mul_90_22_n_643 ,mul_90_22_n_488 ,mul_90_22_n_571);
  and mul_90_22_g3416(mul_90_22_n_642 ,mul_90_22_n_478 ,mul_90_22_n_570);
  and mul_90_22_g3417(mul_90_22_n_641 ,mul_90_22_n_481 ,mul_90_22_n_572);
  and mul_90_22_g3418(mul_90_22_n_639 ,mul_90_22_n_421 ,mul_90_22_n_575);
  or mul_90_22_g3419(mul_90_22_n_638 ,mul_90_22_n_490 ,mul_90_22_n_581);
  and mul_90_22_g3420(mul_90_22_n_636 ,mul_90_22_n_428 ,mul_90_22_n_512);
  and mul_90_22_g3421(mul_90_22_n_634 ,mul_90_22_n_468 ,mul_90_22_n_539);
  and mul_90_22_g3422(mul_90_22_n_633 ,mul_90_22_n_430 ,mul_90_22_n_509);
  and mul_90_22_g3423(mul_90_22_n_632 ,mul_90_22_n_484 ,mul_90_22_n_590);
  and mul_90_22_g3424(mul_90_22_n_631 ,mul_90_22_n_437 ,mul_90_22_n_520);
  and mul_90_22_g3425(mul_90_22_n_630 ,mul_90_22_n_325 ,mul_90_22_n_556);
  and mul_90_22_g3426(mul_90_22_n_629 ,mul_90_22_n_427 ,mul_90_22_n_519);
  or mul_90_22_g3427(mul_90_22_n_628 ,mul_90_22_n_496 ,mul_90_22_n_569);
  and mul_90_22_g3428(mul_90_22_n_627 ,mul_90_22_n_482 ,mul_90_22_n_566);
  and mul_90_22_g3429(mul_90_22_n_625 ,mul_90_22_n_479 ,mul_90_22_n_560);
  and mul_90_22_g3430(mul_90_22_n_624 ,mul_90_22_n_477 ,mul_90_22_n_576);
  and mul_90_22_g3431(mul_90_22_n_623 ,mul_90_22_n_475 ,mul_90_22_n_557);
  and mul_90_22_g3432(mul_90_22_n_622 ,mul_90_22_n_474 ,mul_90_22_n_553);
  and mul_90_22_g3433(mul_90_22_n_621 ,mul_90_22_n_487 ,mul_90_22_n_541);
  or mul_90_22_g3434(mul_90_22_n_619 ,mul_90_22_n_503 ,mul_90_22_n_583);
  and mul_90_22_g3435(mul_90_22_n_618 ,mul_90_22_n_416 ,mul_90_22_n_530);
  and mul_90_22_g3436(mul_90_22_n_616 ,mul_90_22_n_420 ,mul_90_22_n_542);
  and mul_90_22_g3437(mul_90_22_n_614 ,mul_90_22_n_458 ,mul_90_22_n_564);
  and mul_90_22_g3438(mul_90_22_n_612 ,mul_90_22_n_455 ,mul_90_22_n_543);
  and mul_90_22_g3439(mul_90_22_n_611 ,mul_90_22_n_453 ,mul_90_22_n_515);
  and mul_90_22_g3440(mul_90_22_n_610 ,mul_90_22_n_438 ,mul_90_22_n_534);
  and mul_90_22_g3441(mul_90_22_n_609 ,mul_90_22_n_469 ,mul_90_22_n_513);
  and mul_90_22_g3442(mul_90_22_n_608 ,mul_90_22_n_442 ,mul_90_22_n_537);
  and mul_90_22_g3443(mul_90_22_n_607 ,mul_90_22_n_419 ,mul_90_22_n_510);
  and mul_90_22_g3444(mul_90_22_n_606 ,mul_90_22_n_463 ,mul_90_22_n_516);
  and mul_90_22_g3445(mul_90_22_n_605 ,mul_90_22_n_465 ,mul_90_22_n_511);
  or mul_90_22_g3446(mul_90_22_n_604 ,mul_90_22_n_489 ,mul_90_22_n_586);
  and mul_90_22_g3447(mul_90_22_n_602 ,mul_90_22_n_485 ,mul_90_22_n_522);
  and mul_90_22_g3448(mul_90_22_n_600 ,mul_90_22_n_435 ,mul_90_22_n_548);
  and mul_90_22_g3449(mul_90_22_n_599 ,mul_90_22_n_483 ,mul_90_22_n_551);
  and mul_90_22_g3450(mul_90_22_n_598 ,mul_90_22_n_476 ,mul_90_22_n_554);
  and mul_90_22_g3451(mul_90_22_n_597 ,mul_90_22_n_417 ,mul_90_22_n_550);
  and mul_90_22_g3452(mul_90_22_n_596 ,mul_90_22_n_480 ,mul_90_22_n_549);
  and mul_90_22_g3453(mul_90_22_n_594 ,mul_90_22_n_411 ,mul_90_22_n_525);
  and mul_90_22_g3454(mul_90_22_n_592 ,mul_90_22_n_414 ,mul_90_22_n_508);
  or mul_90_22_g3455(mul_90_22_n_590 ,mul_90_22_n_353 ,mul_90_22_n_66);
  and mul_90_22_g3456(mul_90_22_n_589 ,mul_90_22_n_140 ,mul_90_22_n_33);
  and mul_90_22_g3457(mul_90_22_n_588 ,mul_90_22_n_90 ,mul_90_22_n_45);
  and mul_90_22_g3458(mul_90_22_n_587 ,mul_90_22_n_132 ,mul_90_22_n_16);
  and mul_90_22_g3459(mul_90_22_n_586 ,mul_90_22_n_128 ,mul_90_22_n_33);
  and mul_90_22_g3460(mul_90_22_n_585 ,mul_90_22_n_110 ,mul_90_22_n_34);
  and mul_90_22_g3461(mul_90_22_n_584 ,mul_90_22_n_92 ,mul_90_22_n_46);
  and mul_90_22_g3462(mul_90_22_n_583 ,mul_90_22_n_142 ,mul_90_22_n_22);
  and mul_90_22_g3463(mul_90_22_n_582 ,mul_90_22_n_144 ,mul_90_22_n_21);
  and mul_90_22_g3464(mul_90_22_n_581 ,mul_90_22_n_134 ,mul_90_22_n_34);
  and mul_90_22_g3465(mul_90_22_n_580 ,mul_90_22_n_138 ,mul_90_22_n_21);
  and mul_90_22_g3466(mul_90_22_n_579 ,mul_90_22_n_120 ,mul_90_22_n_46);
  and mul_90_22_g3467(mul_90_22_n_578 ,mul_90_22_n_94 ,mul_90_22_n_45);
  and mul_90_22_g3468(mul_90_22_n_577 ,mul_90_22_n_126 ,mul_90_22_n_170);
  or mul_90_22_g3469(mul_90_22_n_576 ,mul_90_22_n_351 ,mul_90_22_n_76);
  or mul_90_22_g3470(mul_90_22_n_575 ,mul_90_22_n_328 ,mul_90_22_n_25);
  nor mul_90_22_g3471(mul_90_22_n_574 ,mul_90_22_n_76 ,mul_90_22_n_330);
  or mul_90_22_g3472(mul_90_22_n_573 ,mul_90_22_n_344 ,mul_90_22_n_58);
  or mul_90_22_g3473(mul_90_22_n_572 ,mul_90_22_n_338 ,mul_90_22_n_75);
  or mul_90_22_g3474(mul_90_22_n_571 ,mul_90_22_n_347 ,mul_90_22_n_40);
  or mul_90_22_g3475(mul_90_22_n_570 ,mul_90_22_n_365 ,mul_90_22_n_39);
  and mul_90_22_g3476(mul_90_22_n_569 ,mul_90_22_n_136 ,mul_90_22_n_22);
  or mul_90_22_g3477(mul_90_22_n_568 ,mul_90_22_n_362 ,mul_90_22_n_37);
  or mul_90_22_g3478(mul_90_22_n_567 ,mul_90_22_n_349 ,mul_90_22_n_57);
  or mul_90_22_g3479(mul_90_22_n_566 ,mul_90_22_n_360 ,mul_90_22_n_40);
  or mul_90_22_g3480(mul_90_22_n_565 ,mul_90_22_n_341 ,mul_90_22_n_81);
  or mul_90_22_g3481(mul_90_22_n_564 ,mul_90_22_n_346 ,mul_90_22_n_36);
  or mul_90_22_g3482(mul_90_22_n_563 ,mul_90_22_n_366 ,mul_90_22_n_25);
  or mul_90_22_g3483(mul_90_22_n_562 ,mul_90_22_n_354 ,mul_90_22_n_24);
  or mul_90_22_g3484(mul_90_22_n_561 ,mul_90_22_n_369 ,mul_90_22_n_24);
  or mul_90_22_g3485(mul_90_22_n_560 ,mul_90_22_n_350 ,mul_90_22_n_14);
  or mul_90_22_g3486(mul_90_22_n_559 ,mul_90_22_n_368 ,mul_90_22_n_37);
  or mul_90_22_g3487(mul_90_22_n_558 ,mul_90_22_n_345 ,mul_90_22_n_57);
  or mul_90_22_g3488(mul_90_22_n_557 ,mul_90_22_n_355 ,mul_90_22_n_88);
  or mul_90_22_g3489(mul_90_22_n_556 ,mul_90_22_n_364 ,mul_90_22_n_39);
  or mul_90_22_g3490(mul_90_22_n_555 ,mul_90_22_n_358 ,mul_90_22_n_81);
  or mul_90_22_g3491(mul_90_22_n_554 ,mul_90_22_n_352 ,mul_90_22_n_66);
  or mul_90_22_g3492(mul_90_22_n_553 ,mul_90_22_n_337 ,mul_90_22_n_75);
  or mul_90_22_g3493(mul_90_22_n_552 ,mul_90_22_n_343 ,mul_90_22_n_36);
  or mul_90_22_g3494(mul_90_22_n_551 ,mul_90_22_n_361 ,mul_90_22_n_67);
  or mul_90_22_g3495(mul_90_22_n_550 ,mul_90_22_n_359 ,mul_90_22_n_10);
  or mul_90_22_g3496(mul_90_22_n_549 ,mul_90_22_n_357 ,mul_90_22_n_87);
  or mul_90_22_g3497(mul_90_22_n_548 ,mul_90_22_n_342 ,mul_90_22_n_10);
  not mul_90_22_g3498(mul_90_22_n_545 ,mul_90_22_n_544);
  or mul_90_22_g3499(mul_90_22_n_543 ,mul_90_22_n_392 ,mul_90_22_n_49);
  or mul_90_22_g3500(mul_90_22_n_542 ,mul_90_22_n_356 ,mul_90_22_n_82);
  or mul_90_22_g3501(mul_90_22_n_541 ,mul_90_22_n_340 ,mul_90_22_n_87);
  and mul_90_22_g3502(mul_90_22_n_540 ,mul_90_22_n_165 ,mul_90_22_n_16);
  or mul_90_22_g3503(mul_90_22_n_539 ,mul_90_22_n_377 ,mul_90_22_n_31);
  or mul_90_22_g3504(mul_90_22_n_538 ,mul_90_22_n_388 ,mul_90_22_n_64);
  or mul_90_22_g3505(mul_90_22_n_537 ,mul_90_22_n_407 ,mul_90_22_n_28);
  or mul_90_22_g3506(mul_90_22_n_536 ,mul_90_22_n_370 ,mul_90_22_n_63);
  or mul_90_22_g3507(mul_90_22_n_535 ,mul_90_22_n_405 ,mul_90_22_n_61);
  or mul_90_22_g3508(mul_90_22_n_534 ,mul_90_22_n_404 ,mul_90_22_n_84);
  or mul_90_22_g3509(mul_90_22_n_533 ,mul_90_22_n_386 ,mul_90_22_n_27);
  or mul_90_22_g3510(mul_90_22_n_532 ,mul_90_22_n_399 ,mul_90_22_n_49);
  or mul_90_22_g3511(mul_90_22_n_531 ,mul_90_22_n_390 ,mul_90_22_n_52);
  or mul_90_22_g3512(mul_90_22_n_530 ,mul_90_22_n_339 ,mul_90_22_n_48);
  or mul_90_22_g3513(mul_90_22_n_529 ,mul_90_22_n_410 ,mul_90_22_n_60);
  or mul_90_22_g3514(mul_90_22_n_528 ,mul_90_22_n_385 ,mul_90_22_n_48);
  or mul_90_22_g3515(mul_90_22_n_527 ,mul_90_22_n_389 ,mul_90_22_n_78);
  or mul_90_22_g3516(mul_90_22_n_526 ,mul_90_22_n_408 ,mul_90_22_n_28);
  or mul_90_22_g3517(mul_90_22_n_525 ,mul_90_22_n_397 ,mul_90_22_n_63);
  or mul_90_22_g3518(mul_90_22_n_524 ,mul_90_22_n_395 ,mul_90_22_n_51);
  or mul_90_22_g3519(mul_90_22_n_523 ,mul_90_22_n_403 ,mul_90_22_n_84);
  or mul_90_22_g3520(mul_90_22_n_522 ,mul_90_22_n_348 ,mul_90_22_n_14);
  or mul_90_22_g3521(mul_90_22_n_521 ,mul_90_22_n_406 ,mul_90_22_n_31);
  or mul_90_22_g3522(mul_90_22_n_520 ,mul_90_22_n_396 ,mul_90_22_n_30);
  or mul_90_22_g3523(mul_90_22_n_519 ,mul_90_22_n_363 ,mul_90_22_n_30);
  or mul_90_22_g3524(mul_90_22_n_518 ,mul_90_22_n_391 ,mul_90_22_n_52);
  or mul_90_22_g3525(mul_90_22_n_517 ,mul_90_22_n_394 ,mul_90_22_n_60);
  or mul_90_22_g3526(mul_90_22_n_516 ,mul_90_22_n_400 ,mul_90_22_n_27);
  or mul_90_22_g3527(mul_90_22_n_515 ,mul_90_22_n_387 ,mul_90_22_n_78);
  or mul_90_22_g3528(mul_90_22_n_514 ,mul_90_22_n_384 ,mul_90_22_n_51);
  or mul_90_22_g3529(mul_90_22_n_513 ,mul_90_22_n_409 ,mul_90_22_n_8);
  or mul_90_22_g3530(mul_90_22_n_512 ,mul_90_22_n_393 ,mul_90_22_n_12);
  or mul_90_22_g3531(mul_90_22_n_511 ,mul_90_22_n_401 ,mul_90_22_n_12);
  or mul_90_22_g3532(mul_90_22_n_510 ,mul_90_22_n_367 ,mul_90_22_n_79);
  or mul_90_22_g3533(mul_90_22_n_509 ,mul_90_22_n_402 ,mul_90_22_n_8);
  or mul_90_22_g3534(mul_90_22_n_508 ,mul_90_22_n_398 ,mul_90_22_n_85);
  nor mul_90_22_g3535(mul_90_22_n_507 ,mul_90_22_n_67 ,mul_90_22_n_311);
  nor mul_90_22_g3536(mul_90_22_n_506 ,mul_90_22_n_58 ,mul_90_22_n_310);
  nor mul_90_22_g3537(mul_90_22_n_505 ,mul_90_22_n_61 ,mul_90_22_n_315);
  nor mul_90_22_g3538(mul_90_22_n_504 ,mul_90_22_n_64 ,mul_90_22_n_316);
  and mul_90_22_g3539(mul_90_22_n_547 ,in12[3] ,mul_90_22_n_439);
  and mul_90_22_g3540(mul_90_22_n_546 ,in12[5] ,mul_90_22_n_415);
  or mul_90_22_g3541(mul_90_22_n_544 ,mul_90_22_n_310 ,mul_90_22_n_424);
  and mul_90_22_g3542(mul_90_22_n_503 ,mul_90_22_n_134 ,mul_90_22_n_246);
  and mul_90_22_g3543(mul_90_22_n_502 ,mul_90_22_n_92 ,mul_90_22_n_236);
  and mul_90_22_g3544(mul_90_22_n_501 ,mul_90_22_n_136 ,mul_90_22_n_209);
  and mul_90_22_g3545(mul_90_22_n_500 ,mul_90_22_n_94 ,mul_90_22_n_237);
  and mul_90_22_g3546(mul_90_22_n_499 ,mul_90_22_n_140 ,mul_90_22_n_209);
  and mul_90_22_g3547(mul_90_22_n_498 ,mul_90_22_n_128 ,mul_90_22_n_210);
  and mul_90_22_g3548(mul_90_22_n_497 ,mul_90_22_n_252 ,mul_90_22_n_210);
  and mul_90_22_g3549(mul_90_22_n_496 ,mul_90_22_n_142 ,mul_90_22_n_237);
  and mul_90_22_g3550(mul_90_22_n_495 ,mul_90_22_n_126 ,mul_90_22_n_200);
  and mul_90_22_g3551(mul_90_22_n_494 ,mul_90_22_n_144 ,mul_90_22_n_199);
  and mul_90_22_g3552(mul_90_22_n_493 ,mul_90_22_n_138 ,mul_90_22_n_236);
  and mul_90_22_g3553(mul_90_22_n_492 ,mul_90_22_n_132 ,mul_90_22_n_246);
  and mul_90_22_g3554(mul_90_22_n_491 ,mul_90_22_n_110 ,mul_90_22_n_200);
  and mul_90_22_g3555(mul_90_22_n_490 ,mul_90_22_n_90 ,mul_90_22_n_245);
  and mul_90_22_g3556(mul_90_22_n_489 ,mul_90_22_n_120 ,mul_90_22_n_245);
  or mul_90_22_g3557(mul_90_22_n_488 ,mul_90_22_n_70 ,mul_90_22_n_338);
  or mul_90_22_g3558(mul_90_22_n_487 ,mul_90_22_n_42 ,mul_90_22_n_337);
  nor mul_90_22_g3559(mul_90_22_n_486 ,mul_90_22_n_73 ,mul_90_22_n_365);
  or mul_90_22_g3560(mul_90_22_n_485 ,mul_90_22_n_54 ,mul_90_22_n_357);
  or mul_90_22_g3561(mul_90_22_n_484 ,mul_90_22_n_72 ,mul_90_22_n_340);
  or mul_90_22_g3562(mul_90_22_n_483 ,mul_90_22_n_69 ,mul_90_22_n_352);
  or mul_90_22_g3563(mul_90_22_n_482 ,mul_90_22_n_43 ,mul_90_22_n_353);
  or mul_90_22_g3564(mul_90_22_n_481 ,mul_90_22_n_55 ,mul_90_22_n_348);
  or mul_90_22_g3565(mul_90_22_n_480 ,mul_90_22_n_72 ,mul_90_22_n_361);
  or mul_90_22_g3566(mul_90_22_n_479 ,mul_90_22_n_69 ,mul_90_22_n_360);
  or mul_90_22_g3567(mul_90_22_n_478 ,mul_90_22_n_42 ,mul_90_22_n_347);
  or mul_90_22_g3568(mul_90_22_n_477 ,mul_90_22_n_54 ,mul_90_22_n_364);
  or mul_90_22_g3569(mul_90_22_n_476 ,mul_90_22_n_55 ,mul_90_22_n_355);
  or mul_90_22_g3570(mul_90_22_n_475 ,mul_90_22_n_43 ,mul_90_22_n_350);
  or mul_90_22_g3571(mul_90_22_n_474 ,mul_90_22_n_73 ,mul_90_22_n_351);
  or mul_90_22_g3572(mul_90_22_n_473 ,mul_90_22_n_406 ,mul_90_22_n_224);
  or mul_90_22_g3573(mul_90_22_n_472 ,mul_90_22_n_344 ,mul_90_22_n_215);
  or mul_90_22_g3574(mul_90_22_n_471 ,mul_90_22_n_404 ,mul_90_22_n_239);
  or mul_90_22_g3575(mul_90_22_n_470 ,mul_90_22_n_385 ,mul_90_22_n_206);
  or mul_90_22_g3576(mul_90_22_n_469 ,mul_90_22_n_400 ,mul_90_22_n_206);
  or mul_90_22_g3577(mul_90_22_n_468 ,mul_90_22_n_401 ,mul_90_22_n_233);
  or mul_90_22_g3578(mul_90_22_n_467 ,mul_90_22_n_408 ,mul_90_22_n_240);
  or mul_90_22_g3579(mul_90_22_n_466 ,mul_90_22_n_343 ,mul_90_22_n_218);
  or mul_90_22_g3580(mul_90_22_n_465 ,mul_90_22_n_384 ,mul_90_22_n_233);
  or mul_90_22_g3581(mul_90_22_n_464 ,mul_90_22_n_405 ,mul_90_22_n_225);
  or mul_90_22_g3582(mul_90_22_n_463 ,mul_90_22_n_388 ,mul_90_22_n_243);
  or mul_90_22_g3583(mul_90_22_n_462 ,mul_90_22_n_393 ,mul_90_22_n_228);
  or mul_90_22_g3584(mul_90_22_n_461 ,mul_90_22_n_387 ,mul_90_22_n_224);
  or mul_90_22_g3585(mul_90_22_n_460 ,mul_90_22_n_359 ,mul_90_22_n_218);
  or mul_90_22_g3586(mul_90_22_n_459 ,mul_90_22_n_367 ,mul_90_22_n_227);
  not mul_90_22_g3587(mul_90_22_n_458 ,mul_90_22_n_457);
  not mul_90_22_g3588(mul_90_22_n_455 ,mul_90_22_n_454);
  not mul_90_22_g3589(mul_90_22_n_453 ,mul_90_22_n_452);
  or mul_90_22_g3590(mul_90_22_n_443 ,mul_90_22_n_345 ,mul_90_22_n_216);
  or mul_90_22_g3591(mul_90_22_n_442 ,mul_90_22_n_403 ,mul_90_22_n_239);
  or mul_90_22_g3592(mul_90_22_n_441 ,mul_90_22_n_369 ,mul_90_22_n_249);
  or mul_90_22_g3593(mul_90_22_n_440 ,mul_90_22_n_368 ,mul_90_22_n_215);
  or mul_90_22_g3594(mul_90_22_n_439 ,mul_90_22_n_321 ,mul_90_22_n_376);
  or mul_90_22_g3595(mul_90_22_n_438 ,mul_90_22_n_398 ,mul_90_22_n_242);
  or mul_90_22_g3596(mul_90_22_n_437 ,mul_90_22_n_389 ,mul_90_22_n_230);
  or mul_90_22_g3597(mul_90_22_n_436 ,mul_90_22_n_402 ,mul_90_22_n_212);
  or mul_90_22_g3598(mul_90_22_n_435 ,mul_90_22_n_354 ,mul_90_22_n_248);
  or mul_90_22_g3599(mul_90_22_n_434 ,mul_90_22_n_396 ,mul_90_22_n_230);
  or mul_90_22_g3600(mul_90_22_n_433 ,mul_90_22_n_366 ,mul_90_22_n_221);
  or mul_90_22_g3601(mul_90_22_n_432 ,mul_90_22_n_341 ,mul_90_22_n_221);
  or mul_90_22_g3602(mul_90_22_n_431 ,mul_90_22_n_394 ,mul_90_22_n_227);
  or mul_90_22_g3603(mul_90_22_n_430 ,mul_90_22_n_392 ,mul_90_22_n_212);
  or mul_90_22_g3604(mul_90_22_n_429 ,mul_90_22_n_349 ,mul_90_22_n_248);
  or mul_90_22_g3605(mul_90_22_n_428 ,mul_90_22_n_363 ,mul_90_22_n_234);
  or mul_90_22_g3606(mul_90_22_n_427 ,mul_90_22_n_395 ,mul_90_22_n_228);
  or mul_90_22_g3607(mul_90_22_n_426 ,mul_90_22_n_410 ,mul_90_22_n_231);
  or mul_90_22_g3608(mul_90_22_n_425 ,mul_90_22_n_356 ,mul_90_22_n_219);
  nor mul_90_22_g3609(mul_90_22_n_424 ,mul_90_22_n_320 ,mul_90_22_n_374);
  or mul_90_22_g3610(mul_90_22_n_423 ,mul_90_22_n_386 ,mul_90_22_n_242);
  or mul_90_22_g3611(mul_90_22_n_422 ,mul_90_22_n_399 ,mul_90_22_n_207);
  or mul_90_22_g3612(mul_90_22_n_421 ,mul_90_22_n_358 ,mul_90_22_n_249);
  or mul_90_22_g3613(mul_90_22_n_420 ,mul_90_22_n_346 ,mul_90_22_n_222);
  or mul_90_22_g3614(mul_90_22_n_419 ,mul_90_22_n_390 ,mul_90_22_n_225);
  or mul_90_22_g3615(mul_90_22_n_418 ,mul_90_22_n_391 ,mul_90_22_n_234);
  or mul_90_22_g3616(mul_90_22_n_417 ,mul_90_22_n_342 ,mul_90_22_n_216);
  or mul_90_22_g3617(mul_90_22_n_416 ,mul_90_22_n_397 ,mul_90_22_n_243);
  or mul_90_22_g3618(mul_90_22_n_415 ,mul_90_22_n_326 ,mul_90_22_n_373);
  or mul_90_22_g3619(mul_90_22_n_414 ,mul_90_22_n_407 ,mul_90_22_n_213);
  or mul_90_22_g3620(mul_90_22_n_413 ,mul_90_22_n_339 ,mul_90_22_n_240);
  or mul_90_22_g3621(mul_90_22_n_412 ,mul_90_22_n_362 ,mul_90_22_n_219);
  or mul_90_22_g3622(mul_90_22_n_411 ,mul_90_22_n_409 ,mul_90_22_n_207);
  and mul_90_22_g3623(mul_90_22_n_457 ,in12[7] ,mul_90_22_n_150);
  or mul_90_22_g3624(mul_90_22_n_456 ,mul_90_22_n_159 ,mul_90_22_n_213);
  and mul_90_22_g3625(mul_90_22_n_454 ,in12[3] ,mul_90_22_n_154);
  and mul_90_22_g3626(mul_90_22_n_452 ,in12[5] ,mul_90_22_n_152);
  or mul_90_22_g3627(mul_90_22_n_451 ,mul_90_22_n_163 ,mul_90_22_n_231);
  or mul_90_22_g3628(mul_90_22_n_450 ,mul_90_22_n_162 ,mul_90_22_n_222);
  or mul_90_22_g3629(mul_90_22_n_449 ,mul_90_22_n_162 ,mul_90_22_n_148);
  and mul_90_22_g3630(mul_90_22_n_448 ,in12[8] ,mul_90_22_n_147);
  or mul_90_22_g3631(mul_90_22_n_447 ,mul_90_22_n_371 ,mul_90_22_n_151);
  or mul_90_22_g3632(mul_90_22_n_446 ,in12[0] ,mul_90_22_n_375);
  or mul_90_22_g3633(mul_90_22_n_445 ,mul_90_22_n_329 ,mul_90_22_n_149);
  or mul_90_22_g3634(mul_90_22_n_444 ,mul_90_22_n_372 ,mul_90_22_n_153);
  not mul_90_22_g3635(mul_90_22_n_383 ,mul_90_22_n_152);
  not mul_90_22_g3636(mul_90_22_n_382 ,mul_90_22_n_151);
  not mul_90_22_g3639(mul_90_22_n_380 ,mul_90_22_n_150);
  not mul_90_22_g3640(mul_90_22_n_379 ,mul_90_22_n_149);
  xnor mul_90_22_g3643(mul_90_22_n_377 ,mul_90_22_n_18 ,in12[5]);
  and mul_90_22_g3644(mul_90_22_n_376 ,mul_90_22_n_202 ,mul_90_22_n_322);
  and mul_90_22_g3646(mul_90_22_n_374 ,mul_90_22_n_315 ,mul_90_22_n_319);
  and mul_90_22_g3647(mul_90_22_n_373 ,mul_90_22_n_316 ,mul_90_22_n_323);
  xnor mul_90_22_g3648(mul_90_22_n_372 ,in12[3] ,in12[2]);
  xnor mul_90_22_g3649(mul_90_22_n_371 ,in12[5] ,in12[4]);
  xnor mul_90_22_g3650(mul_90_22_n_370 ,mul_90_22_n_18 ,in12[3]);
  xnor mul_90_22_g3651(mul_90_22_n_410 ,mul_90_22_n_260 ,in12[5]);
  xnor mul_90_22_g3652(mul_90_22_n_409 ,mul_90_22_n_281 ,in12[3]);
  xnor mul_90_22_g3653(mul_90_22_n_408 ,mul_90_22_n_287 ,in12[3]);
  xnor mul_90_22_g3654(mul_90_22_n_407 ,mul_90_22_n_269 ,in12[3]);
  xnor mul_90_22_g3655(mul_90_22_n_406 ,mul_90_22_n_270 ,in12[5]);
  xnor mul_90_22_g3656(mul_90_22_n_405 ,mul_90_22_n_288 ,in12[5]);
  xnor mul_90_22_g3657(mul_90_22_n_404 ,mul_90_22_n_278 ,in12[3]);
  xnor mul_90_22_g3658(mul_90_22_n_403 ,mul_90_22_n_263 ,in12[3]);
  xnor mul_90_22_g3659(mul_90_22_n_402 ,mul_90_22_n_254 ,in12[3]);
  xnor mul_90_22_g3660(mul_90_22_n_401 ,mul_90_22_n_290 ,in12[5]);
  xnor mul_90_22_g3661(mul_90_22_n_400 ,mul_90_22_n_272 ,in12[3]);
  xnor mul_90_22_g3662(mul_90_22_n_399 ,mul_90_22_n_291 ,in12[3]);
  xnor mul_90_22_g3663(mul_90_22_n_398 ,mul_90_22_n_275 ,in12[3]);
  xnor mul_90_22_g3664(mul_90_22_n_397 ,mul_90_22_n_293 ,in12[3]);
  xnor mul_90_22_g3665(mul_90_22_n_396 ,mul_90_22_n_294 ,in12[5]);
  xnor mul_90_22_g3666(mul_90_22_n_395 ,mul_90_22_n_276 ,in12[5]);
  xnor mul_90_22_g3667(mul_90_22_n_394 ,mul_90_22_n_255 ,in12[5]);
  xnor mul_90_22_g3668(mul_90_22_n_393 ,mul_90_22_n_284 ,in12[5]);
  xnor mul_90_22_g3669(mul_90_22_n_392 ,mul_90_22_n_251 ,in12[3]);
  xnor mul_90_22_g3670(mul_90_22_n_391 ,mul_90_22_n_273 ,in12[5]);
  xnor mul_90_22_g3671(mul_90_22_n_390 ,mul_90_22_n_257 ,in12[5]);
  xnor mul_90_22_g3672(mul_90_22_n_389 ,mul_90_22_n_282 ,in12[5]);
  xnor mul_90_22_g3673(mul_90_22_n_388 ,mul_90_22_n_261 ,in12[3]);
  xnor mul_90_22_g3674(mul_90_22_n_387 ,mul_90_22_n_122 ,in12[5]);
  xnor mul_90_22_g3675(mul_90_22_n_386 ,mul_90_22_n_258 ,in12[3]);
  xnor mul_90_22_g3676(mul_90_22_n_385 ,mul_90_22_n_285 ,in12[3]);
  xnor mul_90_22_g3677(mul_90_22_n_384 ,mul_90_22_n_266 ,in12[5]);
  xnor mul_90_22_g3678(mul_90_22_n_381 ,mul_90_22_n_316 ,in12[4]);
  xnor mul_90_22_g3679(mul_90_22_n_378 ,mul_90_22_n_315 ,in12[6]);
  not mul_90_22_g3680(mul_90_22_n_336 ,mul_90_22_n_148);
  not mul_90_22_g3681(mul_90_22_n_335 ,mul_90_22_n_147);
  not mul_90_22_g3684(mul_90_22_n_333 ,mul_90_22_n_154);
  not mul_90_22_g3685(mul_90_22_n_332 ,mul_90_22_n_153);
  xnor mul_90_22_g3689(mul_90_22_n_329 ,in12[7] ,in12[6]);
  xnor mul_90_22_g3690(mul_90_22_n_328 ,mul_90_22_n_168 ,in12[7]);
  xnor mul_90_22_g3691(mul_90_22_n_369 ,mul_90_22_n_98 ,in12[7]);
  xnor mul_90_22_g3692(mul_90_22_n_368 ,mul_90_22_n_100 ,in12[7]);
  xnor mul_90_22_g3693(mul_90_22_n_367 ,mul_90_22_n_264 ,in12[5]);
  xnor mul_90_22_g3694(mul_90_22_n_366 ,mul_90_22_n_112 ,in12[7]);
  xnor mul_90_22_g3695(mul_90_22_n_365 ,mul_90_22_n_114 ,in12[1]);
  xnor mul_90_22_g3696(mul_90_22_n_364 ,mul_90_22_n_251 ,in12[1]);
  xnor mul_90_22_g3697(mul_90_22_n_363 ,mul_90_22_n_279 ,in12[5]);
  xnor mul_90_22_g3698(mul_90_22_n_362 ,mul_90_22_n_146 ,in12[7]);
  xnor mul_90_22_g3699(mul_90_22_n_361 ,mul_90_22_n_124 ,in12[1]);
  xnor mul_90_22_g3700(mul_90_22_n_360 ,mul_90_22_n_102 ,in12[1]);
  xnor mul_90_22_g3701(mul_90_22_n_359 ,mul_90_22_n_124 ,in12[7]);
  xnor mul_90_22_g3702(mul_90_22_n_358 ,mul_90_22_n_114 ,in12[7]);
  xnor mul_90_22_g3703(mul_90_22_n_357 ,mul_90_22_n_98 ,in12[1]);
  xnor mul_90_22_g3704(mul_90_22_n_356 ,mul_90_22_n_118 ,in12[7]);
  xnor mul_90_22_g3705(mul_90_22_n_355 ,mul_90_22_n_108 ,in12[1]);
  xnor mul_90_22_g3706(mul_90_22_n_354 ,mul_90_22_n_108 ,in12[7]);
  xnor mul_90_22_g3707(mul_90_22_n_353 ,mul_90_22_n_106 ,in12[1]);
  xnor mul_90_22_g3708(mul_90_22_n_352 ,mul_90_22_n_96 ,in12[1]);
  xnor mul_90_22_g3709(mul_90_22_n_351 ,mul_90_22_n_118 ,in12[1]);
  xnor mul_90_22_g3710(mul_90_22_n_350 ,mul_90_22_n_104 ,in12[1]);
  xnor mul_90_22_g3711(mul_90_22_n_349 ,mul_90_22_n_116 ,in12[7]);
  xnor mul_90_22_g3712(mul_90_22_n_348 ,mul_90_22_n_146 ,in12[1]);
  xnor mul_90_22_g3713(mul_90_22_n_347 ,mul_90_22_n_267 ,in12[1]);
  xnor mul_90_22_g3714(mul_90_22_n_346 ,mul_90_22_n_122 ,in12[7]);
  xnor mul_90_22_g3715(mul_90_22_n_345 ,mul_90_22_n_130 ,in12[7]);
  xnor mul_90_22_g3716(mul_90_22_n_344 ,mul_90_22_n_104 ,in12[7]);
  xnor mul_90_22_g3717(mul_90_22_n_343 ,mul_90_22_n_102 ,in12[7]);
  xnor mul_90_22_g3718(mul_90_22_n_342 ,mul_90_22_n_96 ,in12[7]);
  xnor mul_90_22_g3719(mul_90_22_n_341 ,mul_90_22_n_106 ,in12[7]);
  xnor mul_90_22_g3720(mul_90_22_n_340 ,mul_90_22_n_116 ,in12[1]);
  xnor mul_90_22_g3721(mul_90_22_n_339 ,mul_90_22_n_130 ,in12[3]);
  xnor mul_90_22_g3722(mul_90_22_n_338 ,mul_90_22_n_112 ,in12[1]);
  xnor mul_90_22_g3723(mul_90_22_n_337 ,mul_90_22_n_100 ,in12[1]);
  xnor mul_90_22_g3724(mul_90_22_n_334 ,in12[8] ,in12[7]);
  xnor mul_90_22_g3725(mul_90_22_n_331 ,mul_90_22_n_202 ,in12[2]);
  nor mul_90_22_g3726(mul_90_22_n_327 ,mul_90_22_n_70 ,mul_90_22_n_163);
  nor mul_90_22_g3727(mul_90_22_n_326 ,mul_90_22_n_166 ,in12[4]);
  not mul_90_22_g3728(mul_90_22_n_325 ,mul_90_22_n_324);
  and mul_90_22_g3729(mul_90_22_n_324 ,in12[1] ,in12[0]);
  or mul_90_22_g3730(mul_90_22_n_323 ,mul_90_22_n_159 ,mul_90_22_n_313);
  or mul_90_22_g3731(mul_90_22_n_322 ,mul_90_22_n_160 ,mul_90_22_n_318);
  nor mul_90_22_g3732(mul_90_22_n_321 ,mul_90_22_n_19 ,in12[2]);
  nor mul_90_22_g3733(mul_90_22_n_320 ,mul_90_22_n_168 ,in12[6]);
  or mul_90_22_g3734(mul_90_22_n_319 ,mul_90_22_n_160 ,mul_90_22_n_314);
  not mul_90_22_g3735(mul_90_22_n_318 ,in12[2]);
  not mul_90_22_g3736(mul_90_22_n_317 ,in12[0]);
  not mul_90_22_g3737(mul_90_22_n_316 ,in12[3]);
  not mul_90_22_g3738(mul_90_22_n_315 ,in12[5]);
  not mul_90_22_g3739(mul_90_22_n_314 ,in12[6]);
  not mul_90_22_g3740(mul_90_22_n_313 ,in12[4]);
  not mul_90_22_g3741(mul_90_22_n_312 ,mul_90_22_n_165);
  not mul_90_22_g3742(mul_90_22_n_311 ,in12[1]);
  not mul_90_22_g3743(mul_90_22_n_310 ,in12[7]);
  not mul_90_22_drc_bufs3784(mul_90_22_n_297 ,mul_90_22_n_295);
  not mul_90_22_drc_bufs3785(mul_90_22_n_296 ,mul_90_22_n_295);
  not mul_90_22_drc_bufs3786(mul_90_22_n_295 ,n_159);
  not mul_90_22_drc_bufs3814(mul_90_22_n_294 ,mul_90_22_n_292);
  not mul_90_22_drc_bufs3815(mul_90_22_n_293 ,mul_90_22_n_292);
  not mul_90_22_drc_bufs3816(mul_90_22_n_292 ,n_162);
  not mul_90_22_drc_bufs3818(mul_90_22_n_291 ,mul_90_22_n_289);
  not mul_90_22_drc_bufs3819(mul_90_22_n_290 ,mul_90_22_n_289);
  not mul_90_22_drc_bufs3820(mul_90_22_n_289 ,n_160);
  not mul_90_22_drc_bufs3822(mul_90_22_n_288 ,mul_90_22_n_286);
  not mul_90_22_drc_bufs3823(mul_90_22_n_287 ,mul_90_22_n_286);
  not mul_90_22_drc_bufs3824(mul_90_22_n_286 ,n_166);
  not mul_90_22_drc_bufs3826(mul_90_22_n_285 ,mul_90_22_n_283);
  not mul_90_22_drc_bufs3827(mul_90_22_n_284 ,mul_90_22_n_283);
  not mul_90_22_drc_bufs3828(mul_90_22_n_283 ,n_167);
  not mul_90_22_drc_bufs3830(mul_90_22_n_282 ,mul_90_22_n_280);
  not mul_90_22_drc_bufs3831(mul_90_22_n_281 ,mul_90_22_n_280);
  not mul_90_22_drc_bufs3832(mul_90_22_n_280 ,n_163);
  not mul_90_22_drc_bufs3834(mul_90_22_n_279 ,mul_90_22_n_277);
  not mul_90_22_drc_bufs3835(mul_90_22_n_278 ,mul_90_22_n_277);
  not mul_90_22_drc_bufs3836(mul_90_22_n_277 ,n_168);
  not mul_90_22_drc_bufs3838(mul_90_22_n_276 ,mul_90_22_n_274);
  not mul_90_22_drc_bufs3839(mul_90_22_n_275 ,mul_90_22_n_274);
  not mul_90_22_drc_bufs3840(mul_90_22_n_274 ,n_169);
  not mul_90_22_drc_bufs3842(mul_90_22_n_273 ,mul_90_22_n_271);
  not mul_90_22_drc_bufs3843(mul_90_22_n_272 ,mul_90_22_n_271);
  not mul_90_22_drc_bufs3844(mul_90_22_n_271 ,n_164);
  not mul_90_22_drc_bufs3846(mul_90_22_n_270 ,mul_90_22_n_268);
  not mul_90_22_drc_bufs3847(mul_90_22_n_269 ,mul_90_22_n_268);
  not mul_90_22_drc_bufs3848(mul_90_22_n_268 ,n_170);
  not mul_90_22_drc_bufs3850(mul_90_22_n_267 ,mul_90_22_n_265);
  not mul_90_22_drc_bufs3851(mul_90_22_n_266 ,mul_90_22_n_265);
  not mul_90_22_drc_bufs3852(mul_90_22_n_265 ,n_161);
  not mul_90_22_drc_bufs3854(mul_90_22_n_264 ,mul_90_22_n_262);
  not mul_90_22_drc_bufs3855(mul_90_22_n_263 ,mul_90_22_n_262);
  not mul_90_22_drc_bufs3856(mul_90_22_n_262 ,n_171);
  not mul_90_22_drc_bufs3858(mul_90_22_n_261 ,mul_90_22_n_259);
  not mul_90_22_drc_bufs3859(mul_90_22_n_260 ,mul_90_22_n_259);
  not mul_90_22_drc_bufs3860(mul_90_22_n_259 ,n_165);
  not mul_90_22_drc_bufs3862(mul_90_22_n_258 ,mul_90_22_n_256);
  not mul_90_22_drc_bufs3863(mul_90_22_n_257 ,mul_90_22_n_256);
  not mul_90_22_drc_bufs3864(mul_90_22_n_256 ,n_172);
  not mul_90_22_drc_bufs3866(mul_90_22_n_255 ,mul_90_22_n_253);
  not mul_90_22_drc_bufs3867(mul_90_22_n_254 ,mul_90_22_n_253);
  not mul_90_22_drc_bufs3868(mul_90_22_n_253 ,n_173);
  not mul_90_22_drc_bufs3870(mul_90_22_n_252 ,mul_90_22_n_250);
  not mul_90_22_drc_bufs3871(mul_90_22_n_251 ,mul_90_22_n_250);
  not mul_90_22_drc_bufs3872(mul_90_22_n_250 ,n_174);
  not mul_90_22_drc_bufs3874(mul_90_22_n_249 ,mul_90_22_n_247);
  not mul_90_22_drc_bufs3875(mul_90_22_n_248 ,mul_90_22_n_247);
  not mul_90_22_drc_bufs3876(mul_90_22_n_247 ,mul_90_22_n_303);
  not mul_90_22_drc_bufs3878(mul_90_22_n_246 ,mul_90_22_n_244);
  not mul_90_22_drc_bufs3879(mul_90_22_n_245 ,mul_90_22_n_244);
  not mul_90_22_drc_bufs3880(mul_90_22_n_244 ,mul_90_22_n_335);
  not mul_90_22_drc_bufs3882(mul_90_22_n_243 ,mul_90_22_n_241);
  not mul_90_22_drc_bufs3883(mul_90_22_n_242 ,mul_90_22_n_241);
  not mul_90_22_drc_bufs3884(mul_90_22_n_241 ,mul_90_22_n_299);
  not mul_90_22_drc_bufs3886(mul_90_22_n_240 ,mul_90_22_n_238);
  not mul_90_22_drc_bufs3887(mul_90_22_n_239 ,mul_90_22_n_238);
  not mul_90_22_drc_bufs3888(mul_90_22_n_238 ,mul_90_22_n_298);
  not mul_90_22_drc_bufs3890(mul_90_22_n_237 ,mul_90_22_n_235);
  not mul_90_22_drc_bufs3891(mul_90_22_n_236 ,mul_90_22_n_235);
  not mul_90_22_drc_bufs3892(mul_90_22_n_235 ,mul_90_22_n_336);
  not mul_90_22_drc_bufs3894(mul_90_22_n_234 ,mul_90_22_n_232);
  not mul_90_22_drc_bufs3895(mul_90_22_n_233 ,mul_90_22_n_232);
  not mul_90_22_drc_bufs3896(mul_90_22_n_232 ,mul_90_22_n_383);
  not mul_90_22_drc_bufs3898(mul_90_22_n_231 ,mul_90_22_n_229);
  not mul_90_22_drc_bufs3899(mul_90_22_n_230 ,mul_90_22_n_229);
  not mul_90_22_drc_bufs3900(mul_90_22_n_229 ,mul_90_22_n_382);
  not mul_90_22_drc_bufs3902(mul_90_22_n_228 ,mul_90_22_n_226);
  not mul_90_22_drc_bufs3903(mul_90_22_n_227 ,mul_90_22_n_226);
  not mul_90_22_drc_bufs3904(mul_90_22_n_226 ,mul_90_22_n_305);
  not mul_90_22_drc_bufs3906(mul_90_22_n_225 ,mul_90_22_n_223);
  not mul_90_22_drc_bufs3907(mul_90_22_n_224 ,mul_90_22_n_223);
  not mul_90_22_drc_bufs3908(mul_90_22_n_223 ,mul_90_22_n_304);
  not mul_90_22_drc_bufs3910(mul_90_22_n_222 ,mul_90_22_n_220);
  not mul_90_22_drc_bufs3911(mul_90_22_n_221 ,mul_90_22_n_220);
  not mul_90_22_drc_bufs3912(mul_90_22_n_220 ,mul_90_22_n_379);
  not mul_90_22_drc_bufs3914(mul_90_22_n_219 ,mul_90_22_n_217);
  not mul_90_22_drc_bufs3915(mul_90_22_n_218 ,mul_90_22_n_217);
  not mul_90_22_drc_bufs3916(mul_90_22_n_217 ,mul_90_22_n_380);
  not mul_90_22_drc_bufs3918(mul_90_22_n_216 ,mul_90_22_n_214);
  not mul_90_22_drc_bufs3919(mul_90_22_n_215 ,mul_90_22_n_214);
  not mul_90_22_drc_bufs3920(mul_90_22_n_214 ,mul_90_22_n_302);
  not mul_90_22_drc_bufs3922(mul_90_22_n_213 ,mul_90_22_n_211);
  not mul_90_22_drc_bufs3923(mul_90_22_n_212 ,mul_90_22_n_211);
  not mul_90_22_drc_bufs3924(mul_90_22_n_211 ,mul_90_22_n_332);
  not mul_90_22_drc_bufs3926(mul_90_22_n_210 ,mul_90_22_n_208);
  not mul_90_22_drc_bufs3927(mul_90_22_n_209 ,mul_90_22_n_208);
  not mul_90_22_drc_bufs3928(mul_90_22_n_208 ,mul_90_22_n_300);
  not mul_90_22_drc_bufs3930(mul_90_22_n_207 ,mul_90_22_n_205);
  not mul_90_22_drc_bufs3931(mul_90_22_n_206 ,mul_90_22_n_205);
  not mul_90_22_drc_bufs3932(mul_90_22_n_205 ,mul_90_22_n_333);
  not mul_90_22_drc_bufs3934(mul_90_22_n_204 ,mul_90_22_n_649);
  not mul_90_22_drc_bufs3935(mul_90_22_n_203 ,mul_90_22_n_649);
  not mul_90_22_drc_bufs3940(mul_90_22_n_307 ,mul_90_22_n_650);
  not mul_90_22_drc_bufs3943(mul_90_22_n_202 ,mul_90_22_n_201);
  not mul_90_22_drc_bufs3944(mul_90_22_n_201 ,mul_90_22_n_311);
  not mul_90_22_drc_bufs3946(mul_90_22_n_200 ,mul_90_22_n_198);
  not mul_90_22_drc_bufs3947(mul_90_22_n_199 ,mul_90_22_n_198);
  not mul_90_22_drc_bufs3948(mul_90_22_n_198 ,mul_90_22_n_301);
  buf mul_90_22_drc_bufs3957(n_152 ,mul_90_22_n_1140);
  buf mul_90_22_drc_bufs3958(n_153 ,mul_90_22_n_1143);
  buf mul_90_22_drc_bufs3959(n_146 ,mul_90_22_n_1121);
  buf mul_90_22_drc_bufs3960(n_148 ,mul_90_22_n_1127);
  buf mul_90_22_drc_bufs3961(n_149 ,mul_90_22_n_1130);
  buf mul_90_22_drc_bufs3962(n_156 ,mul_90_22_n_1153);
  buf mul_90_22_drc_bufs3963(n_151 ,mul_90_22_n_1137);
  buf mul_90_22_drc_bufs3964(n_150 ,mul_90_22_n_1134);
  buf mul_90_22_drc_bufs3965(n_147 ,mul_90_22_n_1124);
  buf mul_90_22_drc_bufs3966(n_157 ,mul_90_22_n_1156);
  buf mul_90_22_drc_bufs3967(n_154 ,mul_90_22_n_1147);
  buf mul_90_22_drc_bufs3968(n_155 ,mul_90_22_n_1150);
  buf mul_90_22_drc_bufs3969(n_143 ,mul_90_22_n_1112);
  buf mul_90_22_drc_bufs3970(n_144 ,mul_90_22_n_1115);
  buf mul_90_22_drc_bufs3971(n_145 ,mul_90_22_n_1118);
  not mul_90_22_drc_bufs3973(mul_90_22_n_182 ,mul_90_22_n_308);
  not mul_90_22_drc_bufs3974(mul_90_22_n_308 ,mul_90_22_n_885);
  not mul_90_22_drc_bufs3996(mul_90_22_n_181 ,mul_90_22_n_180);
  not mul_90_22_drc_bufs3998(mul_90_22_n_180 ,mul_90_22_n_446);
  not mul_90_22_drc_bufs4001(mul_90_22_n_179 ,mul_90_22_n_178);
  not mul_90_22_drc_bufs4003(mul_90_22_n_178 ,mul_90_22_n_444);
  not mul_90_22_drc_bufs4006(mul_90_22_n_177 ,mul_90_22_n_176);
  not mul_90_22_drc_bufs4008(mul_90_22_n_176 ,mul_90_22_n_447);
  not mul_90_22_drc_bufs4011(mul_90_22_n_175 ,mul_90_22_n_174);
  not mul_90_22_drc_bufs4013(mul_90_22_n_174 ,mul_90_22_n_445);
  not mul_90_22_drc_bufs4021(mul_90_22_n_173 ,mul_90_22_n_172);
  not mul_90_22_drc_bufs4023(mul_90_22_n_172 ,mul_90_22_n_317);
  not mul_90_22_drc_bufs4031(mul_90_22_n_171 ,mul_90_22_n_169);
  not mul_90_22_drc_bufs4032(mul_90_22_n_170 ,mul_90_22_n_169);
  not mul_90_22_drc_bufs4033(mul_90_22_n_169 ,mul_90_22_n_448);
  not mul_90_22_drc_bufs4036(mul_90_22_n_168 ,mul_90_22_n_167);
  not mul_90_22_drc_bufs4037(mul_90_22_n_167 ,mul_90_22_n_297);
  not mul_90_22_drc_bufs4039(mul_90_22_n_166 ,mul_90_22_n_164);
  not mul_90_22_drc_bufs4040(mul_90_22_n_165 ,mul_90_22_n_164);
  not mul_90_22_drc_bufs4041(mul_90_22_n_164 ,mul_90_22_n_296);
  not mul_90_22_drc_bufs4043(mul_90_22_n_163 ,mul_90_22_n_161);
  not mul_90_22_drc_bufs4044(mul_90_22_n_162 ,mul_90_22_n_161);
  not mul_90_22_drc_bufs4045(mul_90_22_n_161 ,mul_90_22_n_312);
  not mul_90_22_drc_bufs4047(mul_90_22_n_160 ,mul_90_22_n_158);
  not mul_90_22_drc_bufs4048(mul_90_22_n_159 ,mul_90_22_n_158);
  not mul_90_22_drc_bufs4049(mul_90_22_n_158 ,mul_90_22_n_312);
  not mul_90_22_drc_bufs4051(mul_90_22_n_157 ,mul_90_22_n_306);
  not mul_90_22_drc_bufs4053(mul_90_22_n_306 ,mul_90_22_n_648);
  not mul_90_22_drc_bufs4056(mul_90_22_n_156 ,mul_90_22_n_155);
  not mul_90_22_drc_bufs4057(mul_90_22_n_155 ,mul_90_22_n_648);
  not mul_90_22_drc_bufs4059(mul_90_22_n_154 ,mul_90_22_n_299);
  not mul_90_22_drc_bufs4061(mul_90_22_n_299 ,mul_90_22_n_331);
  not mul_90_22_drc_bufs4063(mul_90_22_n_153 ,mul_90_22_n_298);
  not mul_90_22_drc_bufs4065(mul_90_22_n_298 ,mul_90_22_n_331);
  not mul_90_22_drc_bufs4067(mul_90_22_n_152 ,mul_90_22_n_305);
  not mul_90_22_drc_bufs4069(mul_90_22_n_305 ,mul_90_22_n_381);
  not mul_90_22_drc_bufs4071(mul_90_22_n_151 ,mul_90_22_n_304);
  not mul_90_22_drc_bufs4073(mul_90_22_n_304 ,mul_90_22_n_381);
  not mul_90_22_drc_bufs4075(mul_90_22_n_150 ,mul_90_22_n_303);
  not mul_90_22_drc_bufs4077(mul_90_22_n_303 ,mul_90_22_n_378);
  not mul_90_22_drc_bufs4079(mul_90_22_n_149 ,mul_90_22_n_302);
  not mul_90_22_drc_bufs4081(mul_90_22_n_302 ,mul_90_22_n_378);
  not mul_90_22_drc_bufs4083(mul_90_22_n_148 ,mul_90_22_n_301);
  not mul_90_22_drc_bufs4085(mul_90_22_n_301 ,mul_90_22_n_334);
  not mul_90_22_drc_bufs4087(mul_90_22_n_147 ,mul_90_22_n_300);
  not mul_90_22_drc_bufs4089(mul_90_22_n_300 ,mul_90_22_n_334);
  not mul_90_22_drc_bufs4091(mul_90_22_n_146 ,mul_90_22_n_145);
  not mul_90_22_drc_bufs4093(mul_90_22_n_145 ,mul_90_22_n_281);
  not mul_90_22_drc_bufs4095(mul_90_22_n_144 ,mul_90_22_n_143);
  not mul_90_22_drc_bufs4097(mul_90_22_n_143 ,mul_90_22_n_291);
  not mul_90_22_drc_bufs4099(mul_90_22_n_142 ,mul_90_22_n_141);
  not mul_90_22_drc_bufs4101(mul_90_22_n_141 ,mul_90_22_n_273);
  not mul_90_22_drc_bufs4103(mul_90_22_n_140 ,mul_90_22_n_139);
  not mul_90_22_drc_bufs4105(mul_90_22_n_139 ,mul_90_22_n_294);
  not mul_90_22_drc_bufs4107(mul_90_22_n_138 ,mul_90_22_n_137);
  not mul_90_22_drc_bufs4109(mul_90_22_n_137 ,mul_90_22_n_255);
  not mul_90_22_drc_bufs4111(mul_90_22_n_136 ,mul_90_22_n_135);
  not mul_90_22_drc_bufs4113(mul_90_22_n_135 ,mul_90_22_n_282);
  not mul_90_22_drc_bufs4115(mul_90_22_n_134 ,mul_90_22_n_133);
  not mul_90_22_drc_bufs4117(mul_90_22_n_133 ,mul_90_22_n_261);
  not mul_90_22_drc_bufs4119(mul_90_22_n_132 ,mul_90_22_n_131);
  not mul_90_22_drc_bufs4121(mul_90_22_n_131 ,mul_90_22_n_264);
  not mul_90_22_drc_bufs4123(mul_90_22_n_130 ,mul_90_22_n_129);
  not mul_90_22_drc_bufs4125(mul_90_22_n_129 ,mul_90_22_n_266);
  not mul_90_22_drc_bufs4127(mul_90_22_n_128 ,mul_90_22_n_127);
  not mul_90_22_drc_bufs4129(mul_90_22_n_127 ,mul_90_22_n_276);
  not mul_90_22_drc_bufs4131(mul_90_22_n_126 ,mul_90_22_n_125);
  not mul_90_22_drc_bufs4133(mul_90_22_n_125 ,mul_90_22_n_258);
  not mul_90_22_drc_bufs4135(mul_90_22_n_124 ,mul_90_22_n_123);
  not mul_90_22_drc_bufs4137(mul_90_22_n_123 ,mul_90_22_n_260);
  not mul_90_22_drc_bufs4139(mul_90_22_n_122 ,mul_90_22_n_121);
  not mul_90_22_drc_bufs4141(mul_90_22_n_121 ,mul_90_22_n_252);
  not mul_90_22_drc_bufs4143(mul_90_22_n_120 ,mul_90_22_n_119);
  not mul_90_22_drc_bufs4145(mul_90_22_n_119 ,mul_90_22_n_270);
  not mul_90_22_drc_bufs4147(mul_90_22_n_118 ,mul_90_22_n_117);
  not mul_90_22_drc_bufs4149(mul_90_22_n_117 ,mul_90_22_n_254);
  not mul_90_22_drc_bufs4151(mul_90_22_n_116 ,mul_90_22_n_115);
  not mul_90_22_drc_bufs4153(mul_90_22_n_115 ,mul_90_22_n_263);
  not mul_90_22_drc_bufs4155(mul_90_22_n_114 ,mul_90_22_n_113);
  not mul_90_22_drc_bufs4157(mul_90_22_n_113 ,mul_90_22_n_290);
  not mul_90_22_drc_bufs4159(mul_90_22_n_112 ,mul_90_22_n_111);
  not mul_90_22_drc_bufs4161(mul_90_22_n_111 ,mul_90_22_n_293);
  not mul_90_22_drc_bufs4163(mul_90_22_n_110 ,mul_90_22_n_109);
  not mul_90_22_drc_bufs4165(mul_90_22_n_109 ,mul_90_22_n_267);
  not mul_90_22_drc_bufs4167(mul_90_22_n_108 ,mul_90_22_n_107);
  not mul_90_22_drc_bufs4169(mul_90_22_n_107 ,mul_90_22_n_284);
  not mul_90_22_drc_bufs4171(mul_90_22_n_106 ,mul_90_22_n_105);
  not mul_90_22_drc_bufs4173(mul_90_22_n_105 ,mul_90_22_n_269);
  not mul_90_22_drc_bufs4175(mul_90_22_n_104 ,mul_90_22_n_103);
  not mul_90_22_drc_bufs4177(mul_90_22_n_103 ,mul_90_22_n_278);
  not mul_90_22_drc_bufs4179(mul_90_22_n_102 ,mul_90_22_n_101);
  not mul_90_22_drc_bufs4181(mul_90_22_n_101 ,mul_90_22_n_275);
  not mul_90_22_drc_bufs4183(mul_90_22_n_100 ,mul_90_22_n_99);
  not mul_90_22_drc_bufs4185(mul_90_22_n_99 ,mul_90_22_n_257);
  not mul_90_22_drc_bufs4187(mul_90_22_n_98 ,mul_90_22_n_97);
  not mul_90_22_drc_bufs4189(mul_90_22_n_97 ,mul_90_22_n_272);
  not mul_90_22_drc_bufs4191(mul_90_22_n_96 ,mul_90_22_n_95);
  not mul_90_22_drc_bufs4193(mul_90_22_n_95 ,mul_90_22_n_287);
  not mul_90_22_drc_bufs4195(mul_90_22_n_94 ,mul_90_22_n_93);
  not mul_90_22_drc_bufs4197(mul_90_22_n_93 ,mul_90_22_n_285);
  not mul_90_22_drc_bufs4199(mul_90_22_n_92 ,mul_90_22_n_91);
  not mul_90_22_drc_bufs4201(mul_90_22_n_91 ,mul_90_22_n_279);
  not mul_90_22_drc_bufs4203(mul_90_22_n_90 ,mul_90_22_n_89);
  not mul_90_22_drc_bufs4205(mul_90_22_n_89 ,mul_90_22_n_288);
  not mul_90_22_drc_bufs4207(mul_90_22_n_88 ,mul_90_22_n_86);
  not mul_90_22_drc_bufs4208(mul_90_22_n_87 ,mul_90_22_n_86);
  not mul_90_22_drc_bufs4209(mul_90_22_n_86 ,mul_90_22_n_446);
  not mul_90_22_drc_bufs4211(mul_90_22_n_85 ,mul_90_22_n_83);
  not mul_90_22_drc_bufs4212(mul_90_22_n_84 ,mul_90_22_n_83);
  not mul_90_22_drc_bufs4213(mul_90_22_n_83 ,mul_90_22_n_444);
  not mul_90_22_drc_bufs4215(mul_90_22_n_82 ,mul_90_22_n_80);
  not mul_90_22_drc_bufs4216(mul_90_22_n_81 ,mul_90_22_n_80);
  not mul_90_22_drc_bufs4217(mul_90_22_n_80 ,mul_90_22_n_445);
  not mul_90_22_drc_bufs4219(mul_90_22_n_79 ,mul_90_22_n_77);
  not mul_90_22_drc_bufs4220(mul_90_22_n_78 ,mul_90_22_n_77);
  not mul_90_22_drc_bufs4221(mul_90_22_n_77 ,mul_90_22_n_447);
  not mul_90_22_drc_bufs4223(mul_90_22_n_76 ,mul_90_22_n_74);
  not mul_90_22_drc_bufs4224(mul_90_22_n_75 ,mul_90_22_n_74);
  not mul_90_22_drc_bufs4225(mul_90_22_n_74 ,mul_90_22_n_181);
  not mul_90_22_drc_bufs4227(mul_90_22_n_73 ,mul_90_22_n_71);
  not mul_90_22_drc_bufs4228(mul_90_22_n_72 ,mul_90_22_n_71);
  not mul_90_22_drc_bufs4229(mul_90_22_n_71 ,mul_90_22_n_317);
  not mul_90_22_drc_bufs4231(mul_90_22_n_70 ,mul_90_22_n_68);
  not mul_90_22_drc_bufs4232(mul_90_22_n_69 ,mul_90_22_n_68);
  not mul_90_22_drc_bufs4233(mul_90_22_n_68 ,mul_90_22_n_173);
  not mul_90_22_drc_bufs4235(mul_90_22_n_67 ,mul_90_22_n_65);
  not mul_90_22_drc_bufs4236(mul_90_22_n_66 ,mul_90_22_n_65);
  not mul_90_22_drc_bufs4237(mul_90_22_n_65 ,mul_90_22_n_446);
  not mul_90_22_drc_bufs4239(mul_90_22_n_64 ,mul_90_22_n_62);
  not mul_90_22_drc_bufs4240(mul_90_22_n_63 ,mul_90_22_n_62);
  not mul_90_22_drc_bufs4241(mul_90_22_n_62 ,mul_90_22_n_179);
  not mul_90_22_drc_bufs4243(mul_90_22_n_61 ,mul_90_22_n_59);
  not mul_90_22_drc_bufs4244(mul_90_22_n_60 ,mul_90_22_n_59);
  not mul_90_22_drc_bufs4245(mul_90_22_n_59 ,mul_90_22_n_177);
  not mul_90_22_drc_bufs4247(mul_90_22_n_58 ,mul_90_22_n_56);
  not mul_90_22_drc_bufs4248(mul_90_22_n_57 ,mul_90_22_n_56);
  not mul_90_22_drc_bufs4249(mul_90_22_n_56 ,mul_90_22_n_175);
  not mul_90_22_drc_bufs4251(mul_90_22_n_55 ,mul_90_22_n_53);
  not mul_90_22_drc_bufs4252(mul_90_22_n_54 ,mul_90_22_n_53);
  not mul_90_22_drc_bufs4253(mul_90_22_n_53 ,mul_90_22_n_317);
  not mul_90_22_drc_bufs4255(mul_90_22_n_52 ,mul_90_22_n_50);
  not mul_90_22_drc_bufs4256(mul_90_22_n_51 ,mul_90_22_n_50);
  not mul_90_22_drc_bufs4257(mul_90_22_n_50 ,mul_90_22_n_177);
  not mul_90_22_drc_bufs4259(mul_90_22_n_49 ,mul_90_22_n_47);
  not mul_90_22_drc_bufs4260(mul_90_22_n_48 ,mul_90_22_n_47);
  not mul_90_22_drc_bufs4261(mul_90_22_n_47 ,mul_90_22_n_444);
  not mul_90_22_drc_bufs4263(mul_90_22_n_46 ,mul_90_22_n_44);
  not mul_90_22_drc_bufs4264(mul_90_22_n_45 ,mul_90_22_n_44);
  not mul_90_22_drc_bufs4265(mul_90_22_n_44 ,mul_90_22_n_448);
  not mul_90_22_drc_bufs4267(mul_90_22_n_43 ,mul_90_22_n_41);
  not mul_90_22_drc_bufs4268(mul_90_22_n_42 ,mul_90_22_n_41);
  not mul_90_22_drc_bufs4269(mul_90_22_n_41 ,mul_90_22_n_173);
  not mul_90_22_drc_bufs4271(mul_90_22_n_40 ,mul_90_22_n_38);
  not mul_90_22_drc_bufs4272(mul_90_22_n_39 ,mul_90_22_n_38);
  not mul_90_22_drc_bufs4273(mul_90_22_n_38 ,mul_90_22_n_181);
  not mul_90_22_drc_bufs4275(mul_90_22_n_37 ,mul_90_22_n_35);
  not mul_90_22_drc_bufs4276(mul_90_22_n_36 ,mul_90_22_n_35);
  not mul_90_22_drc_bufs4277(mul_90_22_n_35 ,mul_90_22_n_175);
  not mul_90_22_drc_bufs4279(mul_90_22_n_34 ,mul_90_22_n_32);
  not mul_90_22_drc_bufs4280(mul_90_22_n_33 ,mul_90_22_n_32);
  not mul_90_22_drc_bufs4281(mul_90_22_n_32 ,mul_90_22_n_448);
  not mul_90_22_drc_bufs4283(mul_90_22_n_31 ,mul_90_22_n_29);
  not mul_90_22_drc_bufs4284(mul_90_22_n_30 ,mul_90_22_n_29);
  not mul_90_22_drc_bufs4285(mul_90_22_n_29 ,mul_90_22_n_447);
  not mul_90_22_drc_bufs4287(mul_90_22_n_28 ,mul_90_22_n_26);
  not mul_90_22_drc_bufs4288(mul_90_22_n_27 ,mul_90_22_n_26);
  not mul_90_22_drc_bufs4289(mul_90_22_n_26 ,mul_90_22_n_179);
  not mul_90_22_drc_bufs4291(mul_90_22_n_25 ,mul_90_22_n_23);
  not mul_90_22_drc_bufs4292(mul_90_22_n_24 ,mul_90_22_n_23);
  not mul_90_22_drc_bufs4293(mul_90_22_n_23 ,mul_90_22_n_445);
  not mul_90_22_drc_bufs4295(mul_90_22_n_22 ,mul_90_22_n_20);
  not mul_90_22_drc_bufs4296(mul_90_22_n_21 ,mul_90_22_n_20);
  not mul_90_22_drc_bufs4297(mul_90_22_n_20 ,mul_90_22_n_171);
  not mul_90_22_drc_bufs4299(mul_90_22_n_19 ,mul_90_22_n_17);
  not mul_90_22_drc_bufs4300(mul_90_22_n_18 ,mul_90_22_n_17);
  not mul_90_22_drc_bufs4301(mul_90_22_n_17 ,mul_90_22_n_297);
  not mul_90_22_drc_bufs4303(mul_90_22_n_16 ,mul_90_22_n_15);
  not mul_90_22_drc_bufs4305(mul_90_22_n_15 ,mul_90_22_n_170);
  not mul_90_22_drc_bufs4307(mul_90_22_n_14 ,mul_90_22_n_13);
  not mul_90_22_drc_bufs4309(mul_90_22_n_13 ,mul_90_22_n_88);
  not mul_90_22_drc_bufs4311(mul_90_22_n_12 ,mul_90_22_n_11);
  not mul_90_22_drc_bufs4313(mul_90_22_n_11 ,mul_90_22_n_79);
  not mul_90_22_drc_bufs4315(mul_90_22_n_10 ,mul_90_22_n_9);
  not mul_90_22_drc_bufs4317(mul_90_22_n_9 ,mul_90_22_n_82);
  not mul_90_22_drc_bufs4319(mul_90_22_n_8 ,mul_90_22_n_7);
  not mul_90_22_drc_bufs4321(mul_90_22_n_7 ,mul_90_22_n_85);
  and mul_90_22_g2(mul_90_22_n_6 ,mul_90_22_n_982 ,mul_90_22_n_996);
  and mul_90_22_g4323(mul_90_22_n_5 ,mul_90_22_n_913 ,mul_90_22_n_966);
  xor mul_90_22_g4324(mul_90_22_n_4 ,mul_90_22_n_882 ,mul_90_22_n_963);
  xor mul_90_22_g4325(mul_90_22_n_3 ,mul_90_22_n_889 ,mul_90_22_n_960);
  xor mul_90_22_g4326(mul_90_22_n_2 ,mul_90_22_n_890 ,mul_90_22_n_930);
  xor mul_90_22_g4327(mul_90_22_n_1 ,mul_90_22_n_599 ,mul_90_22_n_847);
  xor mul_90_22_g4328(mul_90_22_n_0 ,mul_90_22_n_801 ,mul_90_22_n_307);
  xnor mul_102_22_g2868(n_222 ,mul_102_22_n_984 ,mul_102_22_n_1157);
  nor mul_102_22_g2869(mul_102_22_n_1157 ,mul_102_22_n_1026 ,mul_102_22_n_1155);
  xnor mul_102_22_g2870(mul_102_22_n_1156 ,mul_102_22_n_1154 ,mul_102_22_n_1040);
  and mul_102_22_g2871(mul_102_22_n_1155 ,mul_102_22_n_1027 ,mul_102_22_n_1154);
  or mul_102_22_g2872(mul_102_22_n_1154 ,mul_102_22_n_1050 ,mul_102_22_n_1152);
  xnor mul_102_22_g2873(mul_102_22_n_1153 ,mul_102_22_n_1151 ,mul_102_22_n_1061);
  and mul_102_22_g2874(mul_102_22_n_1152 ,mul_102_22_n_1051 ,mul_102_22_n_1151);
  or mul_102_22_g2875(mul_102_22_n_1151 ,mul_102_22_n_1079 ,mul_102_22_n_1149);
  xnor mul_102_22_g2876(mul_102_22_n_1150 ,mul_102_22_n_1148 ,mul_102_22_n_1081);
  nor mul_102_22_g2877(mul_102_22_n_1149 ,mul_102_22_n_1072 ,mul_102_22_n_1148);
  and mul_102_22_g2878(mul_102_22_n_1148 ,mul_102_22_n_1094 ,mul_102_22_n_1146);
  xnor mul_102_22_g2879(mul_102_22_n_1147 ,mul_102_22_n_1144 ,mul_102_22_n_1106);
  or mul_102_22_g2880(mul_102_22_n_1146 ,mul_102_22_n_1093 ,mul_102_22_n_1145);
  not mul_102_22_g2881(mul_102_22_n_1145 ,mul_102_22_n_1144);
  or mul_102_22_g2882(mul_102_22_n_1144 ,mul_102_22_n_1073 ,mul_102_22_n_1142);
  xnor mul_102_22_g2883(mul_102_22_n_1143 ,mul_102_22_n_1141 ,mul_102_22_n_1082);
  and mul_102_22_g2884(mul_102_22_n_1142 ,mul_102_22_n_1080 ,mul_102_22_n_1141);
  or mul_102_22_g2885(mul_102_22_n_1141 ,mul_102_22_n_1087 ,mul_102_22_n_1139);
  xnor mul_102_22_g2886(mul_102_22_n_1140 ,mul_102_22_n_1138 ,mul_102_22_n_1105);
  and mul_102_22_g2887(mul_102_22_n_1139 ,mul_102_22_n_1086 ,mul_102_22_n_1138);
  or mul_102_22_g2888(mul_102_22_n_1138 ,mul_102_22_n_1085 ,mul_102_22_n_1136);
  xnor mul_102_22_g2889(mul_102_22_n_1137 ,mul_102_22_n_1135 ,mul_102_22_n_1104);
  nor mul_102_22_g2890(mul_102_22_n_1136 ,mul_102_22_n_1135 ,mul_102_22_n_1099);
  and mul_102_22_g2891(mul_102_22_n_1135 ,mul_102_22_n_1092 ,mul_102_22_n_1133);
  xnor mul_102_22_g2892(mul_102_22_n_1134 ,mul_102_22_n_1131 ,mul_102_22_n_1103);
  or mul_102_22_g2893(mul_102_22_n_1133 ,mul_102_22_n_1090 ,mul_102_22_n_1132);
  not mul_102_22_g2894(mul_102_22_n_1132 ,mul_102_22_n_1131);
  or mul_102_22_g2895(mul_102_22_n_1131 ,mul_102_22_n_1089 ,mul_102_22_n_1129);
  xnor mul_102_22_g2896(mul_102_22_n_1130 ,mul_102_22_n_1128 ,mul_102_22_n_1102);
  and mul_102_22_g2897(mul_102_22_n_1129 ,mul_102_22_n_1088 ,mul_102_22_n_1128);
  or mul_102_22_g2898(mul_102_22_n_1128 ,mul_102_22_n_1075 ,mul_102_22_n_1126);
  xnor mul_102_22_g2899(mul_102_22_n_1127 ,mul_102_22_n_1125 ,mul_102_22_n_1084);
  and mul_102_22_g2900(mul_102_22_n_1126 ,mul_102_22_n_1074 ,mul_102_22_n_1125);
  or mul_102_22_g2901(mul_102_22_n_1125 ,mul_102_22_n_1098 ,mul_102_22_n_1123);
  xnor mul_102_22_g2902(mul_102_22_n_1124 ,mul_102_22_n_1122 ,mul_102_22_n_1101);
  and mul_102_22_g2903(mul_102_22_n_1123 ,mul_102_22_n_1097 ,mul_102_22_n_1122);
  or mul_102_22_g2904(mul_102_22_n_1122 ,mul_102_22_n_1078 ,mul_102_22_n_1120);
  xnor mul_102_22_g2905(mul_102_22_n_1121 ,mul_102_22_n_1119 ,mul_102_22_n_1083);
  and mul_102_22_g2906(mul_102_22_n_1120 ,mul_102_22_n_1077 ,mul_102_22_n_1119);
  or mul_102_22_g2907(mul_102_22_n_1119 ,mul_102_22_n_1096 ,mul_102_22_n_1117);
  xnor mul_102_22_g2908(mul_102_22_n_1118 ,mul_102_22_n_1116 ,mul_102_22_n_1100);
  and mul_102_22_g2909(mul_102_22_n_1117 ,mul_102_22_n_1095 ,mul_102_22_n_1116);
  or mul_102_22_g2910(mul_102_22_n_1116 ,mul_102_22_n_1041 ,mul_102_22_n_1114);
  xnor mul_102_22_g2911(mul_102_22_n_1115 ,mul_102_22_n_1113 ,mul_102_22_n_1060);
  and mul_102_22_g2912(mul_102_22_n_1114 ,mul_102_22_n_1042 ,mul_102_22_n_1113);
  or mul_102_22_g2913(mul_102_22_n_1113 ,mul_102_22_n_1043 ,mul_102_22_n_1111);
  xnor mul_102_22_g2914(mul_102_22_n_1112 ,mul_102_22_n_1110 ,mul_102_22_n_1059);
  and mul_102_22_g2915(mul_102_22_n_1111 ,mul_102_22_n_1044 ,mul_102_22_n_1110);
  or mul_102_22_g2916(mul_102_22_n_1110 ,mul_102_22_n_6 ,mul_102_22_n_1109);
  nor mul_102_22_g2917(mul_102_22_n_1109 ,mul_102_22_n_1016 ,mul_102_22_n_1108);
  nor mul_102_22_g2918(mul_102_22_n_1108 ,mul_102_22_n_5 ,mul_102_22_n_1107);
  nor mul_102_22_g2919(mul_102_22_n_1107 ,mul_102_22_n_1003 ,mul_102_22_n_1091);
  xnor mul_102_22_g2920(mul_102_22_n_1106 ,mul_102_22_n_1062 ,mul_102_22_n_1039);
  xnor mul_102_22_g2921(mul_102_22_n_1105 ,mul_102_22_n_1019 ,mul_102_22_n_1063);
  xnor mul_102_22_g2922(mul_102_22_n_1104 ,mul_102_22_n_1038 ,mul_102_22_n_1070);
  xnor mul_102_22_g2923(mul_102_22_n_1103 ,mul_102_22_n_1037 ,mul_102_22_n_1069);
  xnor mul_102_22_g2924(mul_102_22_n_1102 ,mul_102_22_n_1055 ,mul_102_22_n_1066);
  xnor mul_102_22_g2925(mul_102_22_n_1101 ,mul_102_22_n_1065 ,mul_102_22_n_1058);
  xnor mul_102_22_g2926(mul_102_22_n_1100 ,mul_102_22_n_1035 ,mul_102_22_n_1067);
  and mul_102_22_g2927(mul_102_22_n_1099 ,mul_102_22_n_1038 ,mul_102_22_n_1071);
  nor mul_102_22_g2928(mul_102_22_n_1098 ,mul_102_22_n_1058 ,mul_102_22_n_1065);
  or mul_102_22_g2929(mul_102_22_n_1097 ,mul_102_22_n_1057 ,mul_102_22_n_1064);
  and mul_102_22_g2930(mul_102_22_n_1096 ,mul_102_22_n_1035 ,mul_102_22_n_1067);
  or mul_102_22_g2931(mul_102_22_n_1095 ,mul_102_22_n_1035 ,mul_102_22_n_1067);
  or mul_102_22_g2932(mul_102_22_n_1094 ,mul_102_22_n_1039 ,mul_102_22_n_1062);
  and mul_102_22_g2933(mul_102_22_n_1093 ,mul_102_22_n_1039 ,mul_102_22_n_1062);
  or mul_102_22_g2934(mul_102_22_n_1092 ,mul_102_22_n_1036 ,mul_102_22_n_1068);
  nor mul_102_22_g2935(mul_102_22_n_1091 ,mul_102_22_n_1000 ,mul_102_22_n_1076);
  nor mul_102_22_g2936(mul_102_22_n_1090 ,mul_102_22_n_1037 ,mul_102_22_n_1069);
  and mul_102_22_g2937(mul_102_22_n_1089 ,mul_102_22_n_1055 ,mul_102_22_n_1066);
  or mul_102_22_g2938(mul_102_22_n_1088 ,mul_102_22_n_1055 ,mul_102_22_n_1066);
  and mul_102_22_g2939(mul_102_22_n_1087 ,mul_102_22_n_1019 ,mul_102_22_n_1063);
  or mul_102_22_g2940(mul_102_22_n_1086 ,mul_102_22_n_1019 ,mul_102_22_n_1063);
  nor mul_102_22_g2941(mul_102_22_n_1085 ,mul_102_22_n_1038 ,mul_102_22_n_1071);
  xnor mul_102_22_g2942(mul_102_22_n_1084 ,mul_102_22_n_1056 ,mul_102_22_n_1045);
  xnor mul_102_22_g2943(mul_102_22_n_1083 ,mul_102_22_n_1047 ,mul_102_22_n_1053);
  xnor mul_102_22_g2944(mul_102_22_n_1082 ,mul_102_22_n_1034 ,mul_102_22_n_1048);
  xnor mul_102_22_g2945(mul_102_22_n_1081 ,mul_102_22_n_1054 ,mul_102_22_n_1017);
  or mul_102_22_g2946(mul_102_22_n_1080 ,mul_102_22_n_1034 ,mul_102_22_n_1048);
  nor mul_102_22_g2947(mul_102_22_n_1079 ,mul_102_22_n_1054 ,mul_102_22_n_1018);
  nor mul_102_22_g2948(mul_102_22_n_1078 ,mul_102_22_n_1053 ,mul_102_22_n_1047);
  or mul_102_22_g2949(mul_102_22_n_1077 ,mul_102_22_n_1052 ,mul_102_22_n_1046);
  nor mul_102_22_g2950(mul_102_22_n_1076 ,mul_102_22_n_999 ,mul_102_22_n_1049);
  and mul_102_22_g2951(mul_102_22_n_1075 ,mul_102_22_n_1056 ,mul_102_22_n_1045);
  or mul_102_22_g2952(mul_102_22_n_1074 ,mul_102_22_n_1056 ,mul_102_22_n_1045);
  and mul_102_22_g2953(mul_102_22_n_1073 ,mul_102_22_n_1034 ,mul_102_22_n_1048);
  and mul_102_22_g2954(mul_102_22_n_1072 ,mul_102_22_n_1054 ,mul_102_22_n_1018);
  not mul_102_22_g2955(mul_102_22_n_1071 ,mul_102_22_n_1070);
  not mul_102_22_g2956(mul_102_22_n_1069 ,mul_102_22_n_1068);
  not mul_102_22_g2957(mul_102_22_n_1065 ,mul_102_22_n_1064);
  xnor mul_102_22_g2958(mul_102_22_n_1061 ,mul_102_22_n_1023 ,mul_102_22_n_1033);
  xnor mul_102_22_g2959(mul_102_22_n_1060 ,mul_102_22_n_1009 ,mul_102_22_n_1021);
  xnor mul_102_22_g2960(mul_102_22_n_1059 ,mul_102_22_n_1010 ,mul_102_22_n_1020);
  xnor mul_102_22_g2961(mul_102_22_n_1070 ,mul_102_22_n_941 ,mul_102_22_n_1011);
  xnor mul_102_22_g2962(mul_102_22_n_1068 ,mul_102_22_n_925 ,mul_102_22_n_4);
  xnor mul_102_22_g2963(mul_102_22_n_1067 ,mul_102_22_n_945 ,mul_102_22_n_1014);
  xnor mul_102_22_g2964(mul_102_22_n_1066 ,mul_102_22_n_942 ,mul_102_22_n_3);
  xnor mul_102_22_g2965(mul_102_22_n_1064 ,mul_102_22_n_912 ,mul_102_22_n_1012);
  xnor mul_102_22_g2966(mul_102_22_n_1063 ,mul_102_22_n_939 ,mul_102_22_n_1013);
  xnor mul_102_22_g2967(mul_102_22_n_1062 ,mul_102_22_n_944 ,mul_102_22_n_1015);
  not mul_102_22_g2968(mul_102_22_n_1057 ,mul_102_22_n_1058);
  not mul_102_22_g2969(mul_102_22_n_1052 ,mul_102_22_n_1053);
  or mul_102_22_g2970(mul_102_22_n_1051 ,mul_102_22_n_1032 ,mul_102_22_n_1022);
  nor mul_102_22_g2971(mul_102_22_n_1050 ,mul_102_22_n_1033 ,mul_102_22_n_1023);
  nor mul_102_22_g2972(mul_102_22_n_1049 ,mul_102_22_n_921 ,mul_102_22_n_1031);
  and mul_102_22_g2973(mul_102_22_n_1058 ,mul_102_22_n_993 ,mul_102_22_n_1024);
  or mul_102_22_g2974(mul_102_22_n_1056 ,mul_102_22_n_1005 ,mul_102_22_n_1030);
  or mul_102_22_g2975(mul_102_22_n_1055 ,mul_102_22_n_997 ,mul_102_22_n_1025);
  and mul_102_22_g2976(mul_102_22_n_1054 ,mul_102_22_n_1007 ,mul_102_22_n_1029);
  and mul_102_22_g2977(mul_102_22_n_1053 ,mul_102_22_n_991 ,mul_102_22_n_1028);
  not mul_102_22_g2978(mul_102_22_n_1047 ,mul_102_22_n_1046);
  or mul_102_22_g2979(mul_102_22_n_1044 ,mul_102_22_n_1010 ,mul_102_22_n_1020);
  and mul_102_22_g2980(mul_102_22_n_1043 ,mul_102_22_n_1010 ,mul_102_22_n_1020);
  or mul_102_22_g2981(mul_102_22_n_1042 ,mul_102_22_n_1009 ,mul_102_22_n_1021);
  and mul_102_22_g2982(mul_102_22_n_1041 ,mul_102_22_n_1009 ,mul_102_22_n_1021);
  xnor mul_102_22_g2983(mul_102_22_n_1040 ,mul_102_22_n_927 ,mul_102_22_n_995);
  xnor mul_102_22_g2984(mul_102_22_n_1048 ,mul_102_22_n_940 ,mul_102_22_n_2);
  xnor mul_102_22_g2985(mul_102_22_n_1046 ,mul_102_22_n_956 ,mul_102_22_n_983);
  xnor mul_102_22_g2986(mul_102_22_n_1045 ,mul_102_22_n_952 ,mul_102_22_n_985);
  not mul_102_22_g2987(mul_102_22_n_1037 ,mul_102_22_n_1036);
  not mul_102_22_g2988(mul_102_22_n_1033 ,mul_102_22_n_1032);
  nor mul_102_22_g2989(mul_102_22_n_1031 ,mul_102_22_n_920 ,mul_102_22_n_1002);
  and mul_102_22_g2990(mul_102_22_n_1030 ,mul_102_22_n_912 ,mul_102_22_n_987);
  or mul_102_22_g2991(mul_102_22_n_1029 ,mul_102_22_n_944 ,mul_102_22_n_1004);
  or mul_102_22_g2992(mul_102_22_n_1028 ,mul_102_22_n_945 ,mul_102_22_n_990);
  or mul_102_22_g2993(mul_102_22_n_1027 ,mul_102_22_n_927 ,mul_102_22_n_995);
  and mul_102_22_g2994(mul_102_22_n_1026 ,mul_102_22_n_927 ,mul_102_22_n_995);
  nor mul_102_22_g2995(mul_102_22_n_1025 ,mul_102_22_n_943 ,mul_102_22_n_1001);
  or mul_102_22_g2996(mul_102_22_n_1024 ,mul_102_22_n_929 ,mul_102_22_n_992);
  and mul_102_22_g2997(mul_102_22_n_1039 ,mul_102_22_n_973 ,mul_102_22_n_994);
  and mul_102_22_g2998(mul_102_22_n_1038 ,mul_102_22_n_969 ,mul_102_22_n_989);
  and mul_102_22_g2999(mul_102_22_n_1036 ,mul_102_22_n_971 ,mul_102_22_n_998);
  or mul_102_22_g3000(mul_102_22_n_1035 ,mul_102_22_n_976 ,mul_102_22_n_986);
  or mul_102_22_g3001(mul_102_22_n_1034 ,mul_102_22_n_978 ,mul_102_22_n_1006);
  or mul_102_22_g3002(mul_102_22_n_1032 ,mul_102_22_n_937 ,mul_102_22_n_1008);
  not mul_102_22_g3003(mul_102_22_n_1022 ,mul_102_22_n_1023);
  not mul_102_22_g3004(mul_102_22_n_1018 ,mul_102_22_n_1017);
  nor mul_102_22_g3006(mul_102_22_n_1016 ,mul_102_22_n_982 ,mul_102_22_n_996);
  xnor mul_102_22_g3007(mul_102_22_n_1015 ,mul_102_22_n_959 ,mul_102_22_n_862);
  xnor mul_102_22_g3008(mul_102_22_n_1014 ,mul_102_22_n_794 ,mul_102_22_n_954);
  xnor mul_102_22_g3009(mul_102_22_n_1013 ,mul_102_22_n_878 ,mul_102_22_n_962);
  xnor mul_102_22_g3010(mul_102_22_n_1012 ,mul_102_22_n_958 ,mul_102_22_n_885);
  xnor mul_102_22_g3011(mul_102_22_n_1011 ,mul_102_22_n_906 ,mul_102_22_n_961);
  xnor mul_102_22_g3014(mul_102_22_n_1023 ,mul_102_22_n_842 ,mul_102_22_n_947);
  xnor mul_102_22_g3015(mul_102_22_n_1021 ,mul_102_22_n_926 ,mul_102_22_n_946);
  xnor mul_102_22_g3016(mul_102_22_n_1020 ,mul_102_22_n_928 ,mul_102_22_n_948);
  or mul_102_22_g3017(mul_102_22_n_1019 ,mul_102_22_n_951 ,mul_102_22_n_988);
  xnor mul_102_22_g3018(mul_102_22_n_1017 ,mul_102_22_n_981 ,mul_102_22_n_949);
  and mul_102_22_g3020(mul_102_22_n_1008 ,mul_102_22_n_981 ,mul_102_22_n_931);
  or mul_102_22_g3021(mul_102_22_n_1007 ,mul_102_22_n_862 ,mul_102_22_n_959);
  and mul_102_22_g3022(mul_102_22_n_1006 ,mul_102_22_n_962 ,mul_102_22_n_977);
  nor mul_102_22_g3023(mul_102_22_n_1005 ,mul_102_22_n_182 ,mul_102_22_n_958);
  and mul_102_22_g3024(mul_102_22_n_1004 ,mul_102_22_n_862 ,mul_102_22_n_959);
  nor mul_102_22_g3025(mul_102_22_n_1003 ,mul_102_22_n_913 ,mul_102_22_n_966);
  nor mul_102_22_g3026(mul_102_22_n_1002 ,mul_102_22_n_935 ,mul_102_22_n_979);
  and mul_102_22_g3027(mul_102_22_n_1001 ,mul_102_22_n_886 ,mul_102_22_n_952);
  nor mul_102_22_g3028(mul_102_22_n_1000 ,mul_102_22_n_848 ,mul_102_22_n_965);
  nor mul_102_22_g3029(mul_102_22_n_999 ,mul_102_22_n_849 ,mul_102_22_n_964);
  or mul_102_22_g3030(mul_102_22_n_998 ,mul_102_22_n_970 ,mul_102_22_n_960);
  nor mul_102_22_g3031(mul_102_22_n_997 ,mul_102_22_n_886 ,mul_102_22_n_952);
  or mul_102_22_g3032(mul_102_22_n_1010 ,mul_102_22_n_923 ,mul_102_22_n_972);
  or mul_102_22_g3033(mul_102_22_n_1009 ,mul_102_22_n_918 ,mul_102_22_n_974);
  or mul_102_22_g3035(mul_102_22_n_994 ,mul_102_22_n_930 ,mul_102_22_n_980);
  or mul_102_22_g3036(mul_102_22_n_993 ,mul_102_22_n_884 ,mul_102_22_n_955);
  nor mul_102_22_g3037(mul_102_22_n_992 ,mul_102_22_n_883 ,mul_102_22_n_956);
  or mul_102_22_g3038(mul_102_22_n_991 ,mul_102_22_n_794 ,mul_102_22_n_953);
  nor mul_102_22_g3039(mul_102_22_n_990 ,mul_102_22_n_793 ,mul_102_22_n_954);
  or mul_102_22_g3040(mul_102_22_n_989 ,mul_102_22_n_968 ,mul_102_22_n_963);
  nor mul_102_22_g3041(mul_102_22_n_988 ,mul_102_22_n_950 ,mul_102_22_n_961);
  or mul_102_22_g3042(mul_102_22_n_987 ,mul_102_22_n_308 ,mul_102_22_n_957);
  nor mul_102_22_g3043(mul_102_22_n_986 ,mul_102_22_n_840 ,mul_102_22_n_975);
  xor mul_102_22_g3044(mul_102_22_n_985 ,mul_102_22_n_943 ,mul_102_22_n_886);
  xnor mul_102_22_g3046(mul_102_22_n_984 ,mul_102_22_n_0 ,mul_102_22_n_916);
  xnor mul_102_22_g3047(mul_102_22_n_996 ,mul_102_22_n_876 ,mul_102_22_n_1);
  xnor mul_102_22_g3048(mul_102_22_n_983 ,mul_102_22_n_929 ,mul_102_22_n_884);
  or mul_102_22_g3049(mul_102_22_n_995 ,mul_102_22_n_933 ,mul_102_22_n_967);
  and mul_102_22_g3051(mul_102_22_n_980 ,mul_102_22_n_890 ,mul_102_22_n_940);
  and mul_102_22_g3052(mul_102_22_n_979 ,mul_102_22_n_802 ,mul_102_22_n_934);
  nor mul_102_22_g3053(mul_102_22_n_978 ,mul_102_22_n_878 ,mul_102_22_n_939);
  or mul_102_22_g3054(mul_102_22_n_977 ,mul_102_22_n_877 ,mul_102_22_n_938);
  nor mul_102_22_g3055(mul_102_22_n_976 ,mul_102_22_n_905 ,mul_102_22_n_926);
  and mul_102_22_g3056(mul_102_22_n_975 ,mul_102_22_n_905 ,mul_102_22_n_926);
  and mul_102_22_g3057(mul_102_22_n_974 ,mul_102_22_n_928 ,mul_102_22_n_917);
  or mul_102_22_g3058(mul_102_22_n_973 ,mul_102_22_n_890 ,mul_102_22_n_940);
  nor mul_102_22_g3059(mul_102_22_n_972 ,mul_102_22_n_847 ,mul_102_22_n_919);
  or mul_102_22_g3060(mul_102_22_n_971 ,mul_102_22_n_889 ,mul_102_22_n_942);
  and mul_102_22_g3061(mul_102_22_n_970 ,mul_102_22_n_889 ,mul_102_22_n_942);
  or mul_102_22_g3062(mul_102_22_n_969 ,mul_102_22_n_882 ,mul_102_22_n_924);
  nor mul_102_22_g3063(mul_102_22_n_968 ,mul_102_22_n_881 ,mul_102_22_n_925);
  and mul_102_22_g3064(mul_102_22_n_967 ,mul_102_22_n_842 ,mul_102_22_n_936);
  or mul_102_22_g3065(mul_102_22_n_982 ,mul_102_22_n_705 ,mul_102_22_n_922);
  or mul_102_22_g3066(mul_102_22_n_981 ,mul_102_22_n_746 ,mul_102_22_n_932);
  not mul_102_22_g3068(mul_102_22_n_965 ,mul_102_22_n_964);
  not mul_102_22_g3071(mul_102_22_n_958 ,mul_102_22_n_957);
  not mul_102_22_g3072(mul_102_22_n_956 ,mul_102_22_n_955);
  not mul_102_22_g3073(mul_102_22_n_953 ,mul_102_22_n_954);
  nor mul_102_22_g3074(mul_102_22_n_951 ,mul_102_22_n_907 ,mul_102_22_n_941);
  and mul_102_22_g3075(mul_102_22_n_950 ,mul_102_22_n_907 ,mul_102_22_n_941);
  xnor mul_102_22_g3076(mul_102_22_n_966 ,mul_102_22_n_910 ,mul_102_22_n_780);
  xnor mul_102_22_g3077(mul_102_22_n_964 ,mul_102_22_n_602 ,mul_102_22_n_875);
  xnor mul_102_22_g3078(mul_102_22_n_949 ,mul_102_22_n_888 ,mul_102_22_n_839);
  xnor mul_102_22_g3079(mul_102_22_n_948 ,mul_102_22_n_880 ,mul_102_22_n_909);
  xnor mul_102_22_g3080(mul_102_22_n_947 ,mul_102_22_n_904 ,mul_102_22_n_649);
  xor mul_102_22_g3081(mul_102_22_n_946 ,mul_102_22_n_905 ,mul_102_22_n_840);
  xnor mul_102_22_g3082(mul_102_22_n_963 ,mul_102_22_n_841 ,mul_102_22_n_868);
  xnor mul_102_22_g3083(mul_102_22_n_962 ,mul_102_22_n_867 ,mul_102_22_n_870);
  xnor mul_102_22_g3084(mul_102_22_n_961 ,mul_102_22_n_866 ,mul_102_22_n_869);
  xnor mul_102_22_g3085(mul_102_22_n_960 ,mul_102_22_n_845 ,mul_102_22_n_874);
  xnor mul_102_22_g3086(mul_102_22_n_959 ,mul_102_22_n_911 ,mul_102_22_n_787);
  xnor mul_102_22_g3087(mul_102_22_n_957 ,mul_102_22_n_865 ,mul_102_22_n_872);
  xnor mul_102_22_g3088(mul_102_22_n_955 ,mul_102_22_n_762 ,mul_102_22_n_871);
  xnor mul_102_22_g3089(mul_102_22_n_954 ,mul_102_22_n_843 ,mul_102_22_n_893);
  xnor mul_102_22_g3090(mul_102_22_n_952 ,mul_102_22_n_864 ,mul_102_22_n_873);
  not mul_102_22_g3091(mul_102_22_n_939 ,mul_102_22_n_938);
  nor mul_102_22_g3092(mul_102_22_n_937 ,mul_102_22_n_839 ,mul_102_22_n_888);
  or mul_102_22_g3093(mul_102_22_n_936 ,mul_102_22_n_204 ,mul_102_22_n_904);
  nor mul_102_22_g3094(mul_102_22_n_935 ,mul_102_22_n_643 ,mul_102_22_n_914);
  or mul_102_22_g3095(mul_102_22_n_934 ,mul_102_22_n_644 ,mul_102_22_n_915);
  and mul_102_22_g3096(mul_102_22_n_933 ,mul_102_22_n_203 ,mul_102_22_n_904);
  and mul_102_22_g3097(mul_102_22_n_932 ,mul_102_22_n_755 ,mul_102_22_n_911);
  or mul_102_22_g3098(mul_102_22_n_931 ,mul_102_22_n_838 ,mul_102_22_n_887);
  and mul_102_22_g3099(mul_102_22_n_945 ,mul_102_22_n_754 ,mul_102_22_n_899);
  and mul_102_22_g3100(mul_102_22_n_944 ,mul_102_22_n_804 ,mul_102_22_n_897);
  and mul_102_22_g3101(mul_102_22_n_943 ,mul_102_22_n_857 ,mul_102_22_n_901);
  and mul_102_22_g3102(mul_102_22_n_942 ,mul_102_22_n_861 ,mul_102_22_n_902);
  and mul_102_22_g3103(mul_102_22_n_941 ,mul_102_22_n_832 ,mul_102_22_n_898);
  and mul_102_22_g3104(mul_102_22_n_940 ,mul_102_22_n_855 ,mul_102_22_n_903);
  or mul_102_22_g3105(mul_102_22_n_938 ,mul_102_22_n_854 ,mul_102_22_n_900);
  not mul_102_22_g3107(mul_102_22_n_924 ,mul_102_22_n_925);
  nor mul_102_22_g3108(mul_102_22_n_923 ,mul_102_22_n_599 ,mul_102_22_n_876);
  and mul_102_22_g3109(mul_102_22_n_922 ,mul_102_22_n_704 ,mul_102_22_n_910);
  nor mul_102_22_g3110(mul_102_22_n_921 ,mul_102_22_n_769 ,mul_102_22_n_891);
  nor mul_102_22_g3111(mul_102_22_n_920 ,mul_102_22_n_768 ,mul_102_22_n_892);
  and mul_102_22_g3112(mul_102_22_n_919 ,mul_102_22_n_599 ,mul_102_22_n_876);
  nor mul_102_22_g3113(mul_102_22_n_918 ,mul_102_22_n_909 ,mul_102_22_n_880);
  or mul_102_22_g3114(mul_102_22_n_917 ,mul_102_22_n_908 ,mul_102_22_n_879);
  or mul_102_22_g3116(mul_102_22_n_916 ,mul_102_22_n_719 ,mul_102_22_n_894);
  xnor mul_102_22_g3117(mul_102_22_n_930 ,mul_102_22_n_844 ,mul_102_22_n_830);
  and mul_102_22_g3118(mul_102_22_n_929 ,mul_102_22_n_851 ,mul_102_22_n_895);
  xnor mul_102_22_g3119(mul_102_22_n_928 ,mul_102_22_n_606 ,mul_102_22_n_831);
  xnor mul_102_22_g3120(mul_102_22_n_927 ,mul_102_22_n_863 ,mul_102_22_n_782);
  xnor mul_102_22_g3121(mul_102_22_n_926 ,mul_102_22_n_846 ,mul_102_22_n_783);
  or mul_102_22_g3122(mul_102_22_n_925 ,mul_102_22_n_835 ,mul_102_22_n_896);
  not mul_102_22_g3123(mul_102_22_n_915 ,mul_102_22_n_914);
  not mul_102_22_g3125(mul_102_22_n_908 ,mul_102_22_n_909);
  not mul_102_22_g3126(mul_102_22_n_907 ,mul_102_22_n_906);
  or mul_102_22_g3127(mul_102_22_n_903 ,mul_102_22_n_858 ,mul_102_22_n_867);
  or mul_102_22_g3128(mul_102_22_n_902 ,mul_102_22_n_860 ,mul_102_22_n_864);
  or mul_102_22_g3129(mul_102_22_n_901 ,mul_102_22_n_856 ,mul_102_22_n_865);
  nor mul_102_22_g3130(mul_102_22_n_900 ,mul_102_22_n_852 ,mul_102_22_n_866);
  or mul_102_22_g3131(mul_102_22_n_899 ,mul_102_22_n_726 ,mul_102_22_n_846);
  or mul_102_22_g3132(mul_102_22_n_898 ,mul_102_22_n_837 ,mul_102_22_n_841);
  or mul_102_22_g3133(mul_102_22_n_897 ,mul_102_22_n_803 ,mul_102_22_n_844);
  nor mul_102_22_g3134(mul_102_22_n_896 ,mul_102_22_n_834 ,mul_102_22_n_845);
  or mul_102_22_g3135(mul_102_22_n_895 ,mul_102_22_n_843 ,mul_102_22_n_850);
  and mul_102_22_g3136(mul_102_22_n_894 ,mul_102_22_n_720 ,mul_102_22_n_863);
  and mul_102_22_g3137(mul_102_22_n_914 ,mul_102_22_n_753 ,mul_102_22_n_859);
  xnor mul_102_22_g3138(mul_102_22_n_893 ,mul_102_22_n_663 ,mul_102_22_n_792);
  xnor mul_102_22_g3139(mul_102_22_n_913 ,mul_102_22_n_731 ,mul_102_22_n_774);
  or mul_102_22_g3140(mul_102_22_n_912 ,mul_102_22_n_816 ,mul_102_22_n_853);
  xnor mul_102_22_g3141(mul_102_22_n_911 ,mul_102_22_n_692 ,mul_102_22_n_800);
  or mul_102_22_g3142(mul_102_22_n_910 ,mul_102_22_n_703 ,mul_102_22_n_833);
  and mul_102_22_g3143(mul_102_22_n_909 ,mul_102_22_n_713 ,mul_102_22_n_836);
  xnor mul_102_22_g3144(mul_102_22_n_906 ,mul_102_22_n_672 ,mul_102_22_n_785);
  xnor mul_102_22_g3145(mul_102_22_n_905 ,mul_102_22_n_661 ,mul_102_22_n_779);
  xnor mul_102_22_g3146(mul_102_22_n_904 ,mul_102_22_n_687 ,mul_102_22_n_777);
  not mul_102_22_g3147(mul_102_22_n_892 ,mul_102_22_n_891);
  not mul_102_22_g3148(mul_102_22_n_888 ,mul_102_22_n_887);
  not mul_102_22_g3150(mul_102_22_n_883 ,mul_102_22_n_884);
  not mul_102_22_g3151(mul_102_22_n_881 ,mul_102_22_n_882);
  not mul_102_22_g3152(mul_102_22_n_879 ,mul_102_22_n_880);
  not mul_102_22_g3153(mul_102_22_n_877 ,mul_102_22_n_878);
  xnor mul_102_22_g3154(mul_102_22_n_875 ,mul_102_22_n_618 ,mul_102_22_n_797);
  xnor mul_102_22_g3155(mul_102_22_n_874 ,mul_102_22_n_758 ,mul_102_22_n_796);
  xnor mul_102_22_g3156(mul_102_22_n_873 ,mul_102_22_n_764 ,mul_102_22_n_829);
  xnor mul_102_22_g3157(mul_102_22_n_872 ,mul_102_22_n_760 ,mul_102_22_n_827);
  xnor mul_102_22_g3158(mul_102_22_n_871 ,mul_102_22_n_767 ,mul_102_22_n_799);
  xnor mul_102_22_g3159(mul_102_22_n_870 ,mul_102_22_n_757 ,mul_102_22_n_825);
  xnor mul_102_22_g3160(mul_102_22_n_869 ,mul_102_22_n_765 ,mul_102_22_n_795);
  xnor mul_102_22_g3161(mul_102_22_n_868 ,mul_102_22_n_730 ,mul_102_22_n_790);
  xnor mul_102_22_g3162(mul_102_22_n_891 ,mul_102_22_n_641 ,mul_102_22_n_775);
  xnor mul_102_22_g3164(mul_102_22_n_890 ,mul_102_22_n_697 ,mul_102_22_n_781);
  xnor mul_102_22_g3165(mul_102_22_n_889 ,mul_102_22_n_608 ,mul_102_22_n_778);
  xnor mul_102_22_g3166(mul_102_22_n_887 ,mul_102_22_n_786 ,mul_102_22_n_204);
  xnor mul_102_22_g3167(mul_102_22_n_886 ,mul_102_22_n_621 ,mul_102_22_n_773);
  xnor mul_102_22_g3168(mul_102_22_n_885 ,mul_102_22_n_632 ,mul_102_22_n_771);
  xnor mul_102_22_g3169(mul_102_22_n_884 ,mul_102_22_n_627 ,mul_102_22_n_770);
  xnor mul_102_22_g3170(mul_102_22_n_882 ,mul_102_22_n_664 ,mul_102_22_n_788);
  xnor mul_102_22_g3171(mul_102_22_n_880 ,mul_102_22_n_631 ,mul_102_22_n_776);
  xnor mul_102_22_g3172(mul_102_22_n_878 ,mul_102_22_n_633 ,mul_102_22_n_772);
  xnor mul_102_22_g3173(mul_102_22_n_876 ,mul_102_22_n_798 ,mul_102_22_n_784);
  or mul_102_22_g3174(mul_102_22_n_861 ,mul_102_22_n_763 ,mul_102_22_n_828);
  nor mul_102_22_g3175(mul_102_22_n_860 ,mul_102_22_n_764 ,mul_102_22_n_829);
  or mul_102_22_g3176(mul_102_22_n_859 ,mul_102_22_n_821 ,mul_102_22_n_751);
  nor mul_102_22_g3177(mul_102_22_n_858 ,mul_102_22_n_757 ,mul_102_22_n_824);
  or mul_102_22_g3178(mul_102_22_n_857 ,mul_102_22_n_760 ,mul_102_22_n_826);
  nor mul_102_22_g3179(mul_102_22_n_856 ,mul_102_22_n_759 ,mul_102_22_n_827);
  or mul_102_22_g3180(mul_102_22_n_855 ,mul_102_22_n_756 ,mul_102_22_n_825);
  and mul_102_22_g3181(mul_102_22_n_854 ,mul_102_22_n_765 ,mul_102_22_n_795);
  and mul_102_22_g3182(mul_102_22_n_853 ,mul_102_22_n_799 ,mul_102_22_n_815);
  nor mul_102_22_g3183(mul_102_22_n_852 ,mul_102_22_n_765 ,mul_102_22_n_795);
  or mul_102_22_g3184(mul_102_22_n_851 ,mul_102_22_n_663 ,mul_102_22_n_791);
  nor mul_102_22_g3185(mul_102_22_n_850 ,mul_102_22_n_662 ,mul_102_22_n_792);
  and mul_102_22_g3186(mul_102_22_n_867 ,mul_102_22_n_715 ,mul_102_22_n_820);
  and mul_102_22_g3187(mul_102_22_n_866 ,mul_102_22_n_736 ,mul_102_22_n_814);
  and mul_102_22_g3188(mul_102_22_n_865 ,mul_102_22_n_743 ,mul_102_22_n_817);
  and mul_102_22_g3189(mul_102_22_n_864 ,mul_102_22_n_752 ,mul_102_22_n_819);
  or mul_102_22_g3190(mul_102_22_n_863 ,mul_102_22_n_741 ,mul_102_22_n_818);
  and mul_102_22_g3191(mul_102_22_n_862 ,mul_102_22_n_737 ,mul_102_22_n_813);
  not mul_102_22_g3192(mul_102_22_n_849 ,mul_102_22_n_848);
  not mul_102_22_g3193(mul_102_22_n_838 ,mul_102_22_n_839);
  nor mul_102_22_g3194(mul_102_22_n_837 ,mul_102_22_n_730 ,mul_102_22_n_790);
  or mul_102_22_g3195(mul_102_22_n_836 ,mul_102_22_n_711 ,mul_102_22_n_798);
  and mul_102_22_g3196(mul_102_22_n_835 ,mul_102_22_n_758 ,mul_102_22_n_796);
  nor mul_102_22_g3197(mul_102_22_n_834 ,mul_102_22_n_758 ,mul_102_22_n_796);
  and mul_102_22_g3198(mul_102_22_n_833 ,mul_102_22_n_750 ,mul_102_22_n_797);
  or mul_102_22_g3199(mul_102_22_n_832 ,mul_102_22_n_729 ,mul_102_22_n_789);
  and mul_102_22_g3200(mul_102_22_n_848 ,mul_102_22_n_747 ,mul_102_22_n_822);
  xnor mul_102_22_g3201(mul_102_22_n_831 ,mul_102_22_n_598 ,mul_102_22_n_733);
  xnor mul_102_22_g3202(mul_102_22_n_830 ,mul_102_22_n_728 ,mul_102_22_n_648);
  and mul_102_22_g3203(mul_102_22_n_847 ,mul_102_22_n_709 ,mul_102_22_n_809);
  and mul_102_22_g3204(mul_102_22_n_846 ,mul_102_22_n_735 ,mul_102_22_n_812);
  and mul_102_22_g3205(mul_102_22_n_845 ,mul_102_22_n_710 ,mul_102_22_n_808);
  and mul_102_22_g3206(mul_102_22_n_844 ,mul_102_22_n_745 ,mul_102_22_n_807);
  and mul_102_22_g3207(mul_102_22_n_843 ,mul_102_22_n_738 ,mul_102_22_n_806);
  or mul_102_22_g3208(mul_102_22_n_842 ,mul_102_22_n_725 ,mul_102_22_n_805);
  and mul_102_22_g3209(mul_102_22_n_841 ,mul_102_22_n_722 ,mul_102_22_n_811);
  and mul_102_22_g3210(mul_102_22_n_840 ,mul_102_22_n_721 ,mul_102_22_n_810);
  and mul_102_22_g3211(mul_102_22_n_839 ,mul_102_22_n_706 ,mul_102_22_n_823);
  not mul_102_22_g3212(mul_102_22_n_828 ,mul_102_22_n_829);
  not mul_102_22_g3213(mul_102_22_n_826 ,mul_102_22_n_827);
  not mul_102_22_g3214(mul_102_22_n_824 ,mul_102_22_n_825);
  or mul_102_22_g3215(mul_102_22_n_823 ,mul_102_22_n_692 ,mul_102_22_n_749);
  or mul_102_22_g3216(mul_102_22_n_822 ,mul_102_22_n_641 ,mul_102_22_n_716);
  or mul_102_22_g3217(mul_102_22_n_821 ,mul_102_22_n_327 ,mul_102_22_n_727);
  or mul_102_22_g3218(mul_102_22_n_820 ,mul_102_22_n_630 ,mul_102_22_n_744);
  or mul_102_22_g3219(mul_102_22_n_819 ,mul_102_22_n_632 ,mul_102_22_n_718);
  and mul_102_22_g3220(mul_102_22_n_818 ,mul_102_22_n_687 ,mul_102_22_n_748);
  or mul_102_22_g3221(mul_102_22_n_817 ,mul_102_22_n_627 ,mul_102_22_n_742);
  nor mul_102_22_g3222(mul_102_22_n_816 ,mul_102_22_n_767 ,mul_102_22_n_761);
  or mul_102_22_g3223(mul_102_22_n_815 ,mul_102_22_n_766 ,mul_102_22_n_762);
  or mul_102_22_g3224(mul_102_22_n_814 ,mul_102_22_n_624 ,mul_102_22_n_739);
  or mul_102_22_g3225(mul_102_22_n_813 ,mul_102_22_n_697 ,mul_102_22_n_723);
  or mul_102_22_g3226(mul_102_22_n_812 ,mul_102_22_n_631 ,mul_102_22_n_724);
  or mul_102_22_g3227(mul_102_22_n_811 ,mul_102_22_n_622 ,mul_102_22_n_714);
  or mul_102_22_g3228(mul_102_22_n_810 ,mul_102_22_n_734 ,mul_102_22_n_717);
  or mul_102_22_g3229(mul_102_22_n_809 ,mul_102_22_n_708 ,mul_102_22_n_732);
  or mul_102_22_g3230(mul_102_22_n_808 ,mul_102_22_n_621 ,mul_102_22_n_707);
  or mul_102_22_g3231(mul_102_22_n_807 ,mul_102_22_n_633 ,mul_102_22_n_702);
  or mul_102_22_g3232(mul_102_22_n_806 ,mul_102_22_n_623 ,mul_102_22_n_740);
  nor mul_102_22_g3233(mul_102_22_n_805 ,mul_102_22_n_203 ,mul_102_22_n_712);
  or mul_102_22_g3234(mul_102_22_n_804 ,mul_102_22_n_156 ,mul_102_22_n_728);
  and mul_102_22_g3235(mul_102_22_n_803 ,mul_102_22_n_157 ,mul_102_22_n_728);
  xnor mul_102_22_g3236(mul_102_22_n_802 ,mul_102_22_n_698 ,mul_102_22_n_547);
  xnor mul_102_22_g3237(mul_102_22_n_801 ,mul_102_22_n_647 ,mul_102_22_n_646);
  xnor mul_102_22_g3238(mul_102_22_n_800 ,mul_102_22_n_604 ,mul_102_22_n_656);
  xnor mul_102_22_g3239(mul_102_22_n_829 ,mul_102_22_n_628 ,mul_102_22_n_636);
  xnor mul_102_22_g3240(mul_102_22_n_827 ,mul_102_22_n_679 ,mul_102_22_n_696);
  xnor mul_102_22_g3241(mul_102_22_n_825 ,mul_102_22_n_645 ,mul_102_22_n_700);
  not mul_102_22_g3242(mul_102_22_n_793 ,mul_102_22_n_794);
  not mul_102_22_g3243(mul_102_22_n_791 ,mul_102_22_n_792);
  not mul_102_22_g3244(mul_102_22_n_789 ,mul_102_22_n_790);
  xnor mul_102_22_g3245(mul_102_22_n_788 ,mul_102_22_n_667 ,mul_102_22_n_624);
  xnor mul_102_22_g3246(mul_102_22_n_787 ,mul_102_22_n_677 ,mul_102_22_n_157);
  xnor mul_102_22_g3247(mul_102_22_n_786 ,mul_102_22_n_670 ,mul_102_22_n_611);
  xor mul_102_22_g3248(mul_102_22_n_785 ,mul_102_22_n_666 ,mul_102_22_n_630);
  xnor mul_102_22_g3249(mul_102_22_n_784 ,mul_102_22_n_609 ,mul_102_22_n_669);
  xnor mul_102_22_g3250(mul_102_22_n_783 ,mul_102_22_n_674 ,mul_102_22_n_654);
  xnor mul_102_22_g3251(mul_102_22_n_782 ,mul_102_22_n_614 ,mul_102_22_n_650);
  xnor mul_102_22_g3252(mul_102_22_n_781 ,mul_102_22_n_657 ,mul_102_22_n_612);
  xnor mul_102_22_g3253(mul_102_22_n_780 ,mul_102_22_n_594 ,mul_102_22_n_596);
  xor mul_102_22_g3254(mul_102_22_n_779 ,mul_102_22_n_659 ,mul_102_22_n_623);
  xnor mul_102_22_g3255(mul_102_22_n_778 ,mul_102_22_n_600 ,mul_102_22_n_622);
  xnor mul_102_22_g3256(mul_102_22_n_777 ,mul_102_22_n_616 ,mul_102_22_n_653);
  xnor mul_102_22_g3257(mul_102_22_n_776 ,mul_102_22_n_449 ,mul_102_22_n_673);
  xnor mul_102_22_g3258(mul_102_22_n_775 ,mul_102_22_n_451 ,mul_102_22_n_651);
  xnor mul_102_22_g3259(mul_102_22_n_774 ,mul_102_22_n_450 ,mul_102_22_n_605);
  xnor mul_102_22_g3260(mul_102_22_n_773 ,mul_102_22_n_592 ,mul_102_22_n_597);
  xnor mul_102_22_g3261(mul_102_22_n_772 ,mul_102_22_n_607 ,mul_102_22_n_665);
  xnor mul_102_22_g3262(mul_102_22_n_771 ,mul_102_22_n_610 ,mul_102_22_n_668);
  xnor mul_102_22_g3263(mul_102_22_n_770 ,mul_102_22_n_678 ,mul_102_22_n_675);
  xnor mul_102_22_g3264(mul_102_22_n_799 ,mul_102_22_n_684 ,mul_102_22_n_682);
  xnor mul_102_22_g3265(mul_102_22_n_798 ,mul_102_22_n_639 ,mul_102_22_n_544);
  xnor mul_102_22_g3266(mul_102_22_n_797 ,mul_102_22_n_546 ,mul_102_22_n_634);
  xnor mul_102_22_g3267(mul_102_22_n_796 ,mul_102_22_n_619 ,mul_102_22_n_629);
  xnor mul_102_22_g3268(mul_102_22_n_795 ,mul_102_22_n_694 ,mul_102_22_n_693);
  xnor mul_102_22_g3269(mul_102_22_n_794 ,mul_102_22_n_690 ,mul_102_22_n_625);
  xnor mul_102_22_g3270(mul_102_22_n_792 ,mul_102_22_n_681 ,mul_102_22_n_685);
  xnor mul_102_22_g3271(mul_102_22_n_790 ,mul_102_22_n_638 ,mul_102_22_n_688);
  not mul_102_22_g3272(mul_102_22_n_769 ,mul_102_22_n_768);
  not mul_102_22_g3273(mul_102_22_n_767 ,mul_102_22_n_766);
  not mul_102_22_g3274(mul_102_22_n_764 ,mul_102_22_n_763);
  not mul_102_22_g3275(mul_102_22_n_761 ,mul_102_22_n_762);
  not mul_102_22_g3276(mul_102_22_n_760 ,mul_102_22_n_759);
  not mul_102_22_g3277(mul_102_22_n_757 ,mul_102_22_n_756);
  or mul_102_22_g3278(mul_102_22_n_755 ,mul_102_22_n_156 ,mul_102_22_n_676);
  or mul_102_22_g3279(mul_102_22_n_754 ,mul_102_22_n_654 ,mul_102_22_n_674);
  or mul_102_22_g3280(mul_102_22_n_753 ,mul_102_22_n_456 ,mul_102_22_n_642);
  or mul_102_22_g3281(mul_102_22_n_752 ,mul_102_22_n_668 ,mul_102_22_n_610);
  and mul_102_22_g3282(mul_102_22_n_751 ,mul_102_22_n_456 ,mul_102_22_n_642);
  or mul_102_22_g3283(mul_102_22_n_750 ,mul_102_22_n_601 ,mul_102_22_n_617);
  nor mul_102_22_g3284(mul_102_22_n_749 ,mul_102_22_n_604 ,mul_102_22_n_655);
  or mul_102_22_g3285(mul_102_22_n_748 ,mul_102_22_n_652 ,mul_102_22_n_615);
  or mul_102_22_g3286(mul_102_22_n_747 ,mul_102_22_n_451 ,mul_102_22_n_651);
  nor mul_102_22_g3287(mul_102_22_n_746 ,mul_102_22_n_306 ,mul_102_22_n_677);
  or mul_102_22_g3288(mul_102_22_n_745 ,mul_102_22_n_665 ,mul_102_22_n_607);
  and mul_102_22_g3289(mul_102_22_n_744 ,mul_102_22_n_672 ,mul_102_22_n_666);
  or mul_102_22_g3290(mul_102_22_n_743 ,mul_102_22_n_675 ,mul_102_22_n_678);
  and mul_102_22_g3291(mul_102_22_n_742 ,mul_102_22_n_675 ,mul_102_22_n_678);
  nor mul_102_22_g3292(mul_102_22_n_741 ,mul_102_22_n_653 ,mul_102_22_n_616);
  nor mul_102_22_g3293(mul_102_22_n_740 ,mul_102_22_n_661 ,mul_102_22_n_658);
  and mul_102_22_g3294(mul_102_22_n_739 ,mul_102_22_n_667 ,mul_102_22_n_664);
  or mul_102_22_g3295(mul_102_22_n_738 ,mul_102_22_n_660 ,mul_102_22_n_659);
  or mul_102_22_g3296(mul_102_22_n_737 ,mul_102_22_n_612 ,mul_102_22_n_657);
  or mul_102_22_g3297(mul_102_22_n_736 ,mul_102_22_n_667 ,mul_102_22_n_664);
  or mul_102_22_g3298(mul_102_22_n_735 ,mul_102_22_n_449 ,mul_102_22_n_673);
  and mul_102_22_g3299(mul_102_22_n_768 ,mul_102_22_n_547 ,mul_102_22_n_699);
  and mul_102_22_g3300(mul_102_22_n_766 ,mul_102_22_n_681 ,mul_102_22_n_686);
  and mul_102_22_g3301(mul_102_22_n_765 ,mul_102_22_n_638 ,mul_102_22_n_689);
  or mul_102_22_g3302(mul_102_22_n_763 ,mul_102_22_n_680 ,mul_102_22_n_696);
  and mul_102_22_g3303(mul_102_22_n_762 ,mul_102_22_n_626 ,mul_102_22_n_691);
  and mul_102_22_g3304(mul_102_22_n_759 ,mul_102_22_n_684 ,mul_102_22_n_683);
  and mul_102_22_g3305(mul_102_22_n_758 ,mul_102_22_n_628 ,mul_102_22_n_637);
  or mul_102_22_g3306(mul_102_22_n_756 ,mul_102_22_n_695 ,mul_102_22_n_693);
  not mul_102_22_g3307(mul_102_22_n_734 ,mul_102_22_n_733);
  not mul_102_22_g3308(mul_102_22_n_732 ,mul_102_22_n_731);
  not mul_102_22_g3309(mul_102_22_n_730 ,mul_102_22_n_729);
  or mul_102_22_g3310(mul_102_22_n_727 ,mul_102_22_n_311 ,mul_102_22_n_591);
  and mul_102_22_g3311(mul_102_22_n_726 ,mul_102_22_n_654 ,mul_102_22_n_674);
  nor mul_102_22_g3312(mul_102_22_n_725 ,mul_102_22_n_671 ,mul_102_22_n_611);
  and mul_102_22_g3313(mul_102_22_n_724 ,mul_102_22_n_449 ,mul_102_22_n_673);
  and mul_102_22_g3314(mul_102_22_n_723 ,mul_102_22_n_612 ,mul_102_22_n_657);
  or mul_102_22_g3315(mul_102_22_n_722 ,mul_102_22_n_600 ,mul_102_22_n_608);
  or mul_102_22_g3316(mul_102_22_n_721 ,mul_102_22_n_598 ,mul_102_22_n_606);
  or mul_102_22_g3317(mul_102_22_n_720 ,mul_102_22_n_307 ,mul_102_22_n_613);
  nor mul_102_22_g3318(mul_102_22_n_719 ,mul_102_22_n_650 ,mul_102_22_n_614);
  and mul_102_22_g3319(mul_102_22_n_718 ,mul_102_22_n_668 ,mul_102_22_n_610);
  and mul_102_22_g3320(mul_102_22_n_717 ,mul_102_22_n_598 ,mul_102_22_n_606);
  and mul_102_22_g3321(mul_102_22_n_716 ,mul_102_22_n_451 ,mul_102_22_n_651);
  or mul_102_22_g3322(mul_102_22_n_715 ,mul_102_22_n_672 ,mul_102_22_n_666);
  and mul_102_22_g3323(mul_102_22_n_714 ,mul_102_22_n_600 ,mul_102_22_n_608);
  or mul_102_22_g3324(mul_102_22_n_713 ,mul_102_22_n_669 ,mul_102_22_n_609);
  and mul_102_22_g3325(mul_102_22_n_712 ,mul_102_22_n_671 ,mul_102_22_n_611);
  and mul_102_22_g3326(mul_102_22_n_711 ,mul_102_22_n_669 ,mul_102_22_n_609);
  or mul_102_22_g3327(mul_102_22_n_710 ,mul_102_22_n_597 ,mul_102_22_n_592);
  or mul_102_22_g3328(mul_102_22_n_709 ,mul_102_22_n_450 ,mul_102_22_n_605);
  and mul_102_22_g3329(mul_102_22_n_708 ,mul_102_22_n_450 ,mul_102_22_n_605);
  and mul_102_22_g3330(mul_102_22_n_707 ,mul_102_22_n_597 ,mul_102_22_n_592);
  or mul_102_22_g3331(mul_102_22_n_706 ,mul_102_22_n_603 ,mul_102_22_n_656);
  nor mul_102_22_g3332(mul_102_22_n_705 ,mul_102_22_n_596 ,mul_102_22_n_594);
  or mul_102_22_g3333(mul_102_22_n_704 ,mul_102_22_n_595 ,mul_102_22_n_593);
  nor mul_102_22_g3334(mul_102_22_n_703 ,mul_102_22_n_602 ,mul_102_22_n_618);
  and mul_102_22_g3335(mul_102_22_n_702 ,mul_102_22_n_665 ,mul_102_22_n_607);
  and mul_102_22_g3336(mul_102_22_n_733 ,mul_102_22_n_545 ,mul_102_22_n_640);
  and mul_102_22_g3337(mul_102_22_n_731 ,mul_102_22_n_546 ,mul_102_22_n_635);
  or mul_102_22_g3338(mul_102_22_n_729 ,mul_102_22_n_620 ,mul_102_22_n_629);
  and mul_102_22_g3339(mul_102_22_n_728 ,mul_102_22_n_645 ,mul_102_22_n_701);
  not mul_102_22_g3340(mul_102_22_n_701 ,mul_102_22_n_700);
  not mul_102_22_g3341(mul_102_22_n_699 ,mul_102_22_n_698);
  not mul_102_22_g3342(mul_102_22_n_695 ,mul_102_22_n_694);
  not mul_102_22_g3343(mul_102_22_n_691 ,mul_102_22_n_690);
  not mul_102_22_g3344(mul_102_22_n_689 ,mul_102_22_n_688);
  not mul_102_22_g3345(mul_102_22_n_686 ,mul_102_22_n_685);
  not mul_102_22_g3346(mul_102_22_n_683 ,mul_102_22_n_682);
  not mul_102_22_g3347(mul_102_22_n_680 ,mul_102_22_n_679);
  not mul_102_22_g3348(mul_102_22_n_676 ,mul_102_22_n_677);
  not mul_102_22_g3349(mul_102_22_n_671 ,mul_102_22_n_670);
  not mul_102_22_g3350(mul_102_22_n_662 ,mul_102_22_n_663);
  not mul_102_22_g3351(mul_102_22_n_660 ,mul_102_22_n_661);
  not mul_102_22_g3352(mul_102_22_n_658 ,mul_102_22_n_659);
  not mul_102_22_g3353(mul_102_22_n_655 ,mul_102_22_n_656);
  not mul_102_22_g3354(mul_102_22_n_652 ,mul_102_22_n_653);
  or mul_102_22_g3358(mul_102_22_n_700 ,mul_102_22_n_502 ,mul_102_22_n_578);
  and mul_102_22_g3359(mul_102_22_n_698 ,mul_102_22_n_422 ,mul_102_22_n_536);
  or mul_102_22_g3360(mul_102_22_n_647 ,mul_102_22_n_457 ,mul_102_22_n_506);
  or mul_102_22_g3361(mul_102_22_n_646 ,mul_102_22_n_497 ,mul_102_22_n_580);
  and mul_102_22_g3362(mul_102_22_n_697 ,mul_102_22_n_429 ,mul_102_22_n_565);
  and mul_102_22_g3363(mul_102_22_n_696 ,mul_102_22_n_460 ,mul_102_22_n_561);
  or mul_102_22_g3364(mul_102_22_n_694 ,mul_102_22_n_500 ,mul_102_22_n_588);
  and mul_102_22_g3365(mul_102_22_n_693 ,mul_102_22_n_466 ,mul_102_22_n_573);
  and mul_102_22_g3366(mul_102_22_n_692 ,mul_102_22_n_461 ,mul_102_22_n_517);
  and mul_102_22_g3367(mul_102_22_n_690 ,mul_102_22_n_470 ,mul_102_22_n_526);
  and mul_102_22_g3368(mul_102_22_n_688 ,mul_102_22_n_472 ,mul_102_22_n_562);
  or mul_102_22_g3369(mul_102_22_n_687 ,mul_102_22_n_495 ,mul_102_22_n_587);
  and mul_102_22_g3370(mul_102_22_n_685 ,mul_102_22_n_412 ,mul_102_22_n_563);
  or mul_102_22_g3371(mul_102_22_n_684 ,mul_102_22_n_499 ,mul_102_22_n_585);
  and mul_102_22_g3372(mul_102_22_n_682 ,mul_102_22_n_441 ,mul_102_22_n_568);
  or mul_102_22_g3373(mul_102_22_n_681 ,mul_102_22_n_491 ,mul_102_22_n_582);
  or mul_102_22_g3374(mul_102_22_n_679 ,mul_102_22_n_501 ,mul_102_22_n_589);
  and mul_102_22_g3375(mul_102_22_n_678 ,mul_102_22_n_471 ,mul_102_22_n_528);
  and mul_102_22_g3376(mul_102_22_n_677 ,mul_102_22_n_440 ,mul_102_22_n_567);
  and mul_102_22_g3377(mul_102_22_n_675 ,mul_102_22_n_464 ,mul_102_22_n_529);
  and mul_102_22_g3378(mul_102_22_n_674 ,mul_102_22_n_467 ,mul_102_22_n_538);
  and mul_102_22_g3379(mul_102_22_n_673 ,mul_102_22_n_443 ,mul_102_22_n_555);
  and mul_102_22_g3380(mul_102_22_n_672 ,mul_102_22_n_459 ,mul_102_22_n_521);
  or mul_102_22_g3381(mul_102_22_n_670 ,mul_102_22_n_492 ,mul_102_22_n_579);
  and mul_102_22_g3382(mul_102_22_n_669 ,mul_102_22_n_434 ,mul_102_22_n_514);
  and mul_102_22_g3383(mul_102_22_n_668 ,mul_102_22_n_462 ,mul_102_22_n_535);
  and mul_102_22_g3384(mul_102_22_n_667 ,mul_102_22_n_473 ,mul_102_22_n_524);
  and mul_102_22_g3385(mul_102_22_n_666 ,mul_102_22_n_436 ,mul_102_22_n_533);
  and mul_102_22_g3386(mul_102_22_n_665 ,mul_102_22_n_432 ,mul_102_22_n_552);
  and mul_102_22_g3387(mul_102_22_n_664 ,mul_102_22_n_423 ,mul_102_22_n_523);
  and mul_102_22_g3388(mul_102_22_n_663 ,mul_102_22_n_426 ,mul_102_22_n_518);
  or mul_102_22_g3389(mul_102_22_n_661 ,mul_102_22_n_494 ,mul_102_22_n_540);
  and mul_102_22_g3390(mul_102_22_n_659 ,mul_102_22_n_433 ,mul_102_22_n_558);
  and mul_102_22_g3391(mul_102_22_n_657 ,mul_102_22_n_431 ,mul_102_22_n_531);
  or mul_102_22_g3392(mul_102_22_n_656 ,mul_102_22_n_454 ,mul_102_22_n_504);
  and mul_102_22_g3393(mul_102_22_n_654 ,mul_102_22_n_418 ,mul_102_22_n_527);
  or mul_102_22_g3394(mul_102_22_n_653 ,mul_102_22_n_452 ,mul_102_22_n_505);
  and mul_102_22_g3395(mul_102_22_n_651 ,mul_102_22_n_413 ,mul_102_22_n_532);
  or mul_102_22_g3396(mul_102_22_n_650 ,mul_102_22_n_493 ,mul_102_22_n_577);
  and mul_102_22_g3397(mul_102_22_n_649 ,mul_102_22_n_425 ,mul_102_22_n_559);
  or mul_102_22_g3398(mul_102_22_n_648 ,mul_102_22_n_498 ,mul_102_22_n_584);
  not mul_102_22_g3399(mul_102_22_n_644 ,mul_102_22_n_643);
  not mul_102_22_g3400(mul_102_22_n_640 ,mul_102_22_n_639);
  not mul_102_22_g3401(mul_102_22_n_637 ,mul_102_22_n_636);
  not mul_102_22_g3402(mul_102_22_n_635 ,mul_102_22_n_634);
  not mul_102_22_g3403(mul_102_22_n_626 ,mul_102_22_n_625);
  not mul_102_22_g3404(mul_102_22_n_620 ,mul_102_22_n_619);
  not mul_102_22_g3405(mul_102_22_n_617 ,mul_102_22_n_618);
  not mul_102_22_g3406(mul_102_22_n_615 ,mul_102_22_n_616);
  not mul_102_22_g3407(mul_102_22_n_613 ,mul_102_22_n_614);
  not mul_102_22_g3408(mul_102_22_n_603 ,mul_102_22_n_604);
  not mul_102_22_g3409(mul_102_22_n_601 ,mul_102_22_n_602);
  not mul_102_22_g3411(mul_102_22_n_595 ,mul_102_22_n_596);
  not mul_102_22_g3412(mul_102_22_n_593 ,mul_102_22_n_594);
  nor mul_102_22_g3413(mul_102_22_n_591 ,mul_102_22_n_486 ,mul_102_22_n_574);
  or mul_102_22_g3414(mul_102_22_n_645 ,mul_102_22_n_324 ,mul_102_22_n_507);
  and mul_102_22_g3415(mul_102_22_n_643 ,mul_102_22_n_488 ,mul_102_22_n_571);
  and mul_102_22_g3416(mul_102_22_n_642 ,mul_102_22_n_478 ,mul_102_22_n_570);
  and mul_102_22_g3417(mul_102_22_n_641 ,mul_102_22_n_481 ,mul_102_22_n_572);
  and mul_102_22_g3418(mul_102_22_n_639 ,mul_102_22_n_421 ,mul_102_22_n_575);
  or mul_102_22_g3419(mul_102_22_n_638 ,mul_102_22_n_490 ,mul_102_22_n_581);
  and mul_102_22_g3420(mul_102_22_n_636 ,mul_102_22_n_428 ,mul_102_22_n_512);
  and mul_102_22_g3421(mul_102_22_n_634 ,mul_102_22_n_468 ,mul_102_22_n_539);
  and mul_102_22_g3422(mul_102_22_n_633 ,mul_102_22_n_430 ,mul_102_22_n_509);
  and mul_102_22_g3423(mul_102_22_n_632 ,mul_102_22_n_484 ,mul_102_22_n_590);
  and mul_102_22_g3424(mul_102_22_n_631 ,mul_102_22_n_437 ,mul_102_22_n_520);
  and mul_102_22_g3425(mul_102_22_n_630 ,mul_102_22_n_325 ,mul_102_22_n_556);
  and mul_102_22_g3426(mul_102_22_n_629 ,mul_102_22_n_427 ,mul_102_22_n_519);
  or mul_102_22_g3427(mul_102_22_n_628 ,mul_102_22_n_496 ,mul_102_22_n_569);
  and mul_102_22_g3428(mul_102_22_n_627 ,mul_102_22_n_482 ,mul_102_22_n_566);
  and mul_102_22_g3429(mul_102_22_n_625 ,mul_102_22_n_479 ,mul_102_22_n_560);
  and mul_102_22_g3430(mul_102_22_n_624 ,mul_102_22_n_477 ,mul_102_22_n_576);
  and mul_102_22_g3431(mul_102_22_n_623 ,mul_102_22_n_475 ,mul_102_22_n_557);
  and mul_102_22_g3432(mul_102_22_n_622 ,mul_102_22_n_474 ,mul_102_22_n_553);
  and mul_102_22_g3433(mul_102_22_n_621 ,mul_102_22_n_487 ,mul_102_22_n_541);
  or mul_102_22_g3434(mul_102_22_n_619 ,mul_102_22_n_503 ,mul_102_22_n_583);
  and mul_102_22_g3435(mul_102_22_n_618 ,mul_102_22_n_416 ,mul_102_22_n_530);
  and mul_102_22_g3436(mul_102_22_n_616 ,mul_102_22_n_420 ,mul_102_22_n_542);
  and mul_102_22_g3437(mul_102_22_n_614 ,mul_102_22_n_458 ,mul_102_22_n_564);
  and mul_102_22_g3438(mul_102_22_n_612 ,mul_102_22_n_455 ,mul_102_22_n_543);
  and mul_102_22_g3439(mul_102_22_n_611 ,mul_102_22_n_453 ,mul_102_22_n_515);
  and mul_102_22_g3440(mul_102_22_n_610 ,mul_102_22_n_438 ,mul_102_22_n_534);
  and mul_102_22_g3441(mul_102_22_n_609 ,mul_102_22_n_469 ,mul_102_22_n_513);
  and mul_102_22_g3442(mul_102_22_n_608 ,mul_102_22_n_442 ,mul_102_22_n_537);
  and mul_102_22_g3443(mul_102_22_n_607 ,mul_102_22_n_419 ,mul_102_22_n_510);
  and mul_102_22_g3444(mul_102_22_n_606 ,mul_102_22_n_463 ,mul_102_22_n_516);
  and mul_102_22_g3445(mul_102_22_n_605 ,mul_102_22_n_465 ,mul_102_22_n_511);
  or mul_102_22_g3446(mul_102_22_n_604 ,mul_102_22_n_489 ,mul_102_22_n_586);
  and mul_102_22_g3447(mul_102_22_n_602 ,mul_102_22_n_485 ,mul_102_22_n_522);
  and mul_102_22_g3448(mul_102_22_n_600 ,mul_102_22_n_435 ,mul_102_22_n_548);
  and mul_102_22_g3449(mul_102_22_n_599 ,mul_102_22_n_483 ,mul_102_22_n_551);
  and mul_102_22_g3450(mul_102_22_n_598 ,mul_102_22_n_476 ,mul_102_22_n_554);
  and mul_102_22_g3451(mul_102_22_n_597 ,mul_102_22_n_417 ,mul_102_22_n_550);
  and mul_102_22_g3452(mul_102_22_n_596 ,mul_102_22_n_480 ,mul_102_22_n_549);
  and mul_102_22_g3453(mul_102_22_n_594 ,mul_102_22_n_411 ,mul_102_22_n_525);
  and mul_102_22_g3454(mul_102_22_n_592 ,mul_102_22_n_414 ,mul_102_22_n_508);
  or mul_102_22_g3455(mul_102_22_n_590 ,mul_102_22_n_353 ,mul_102_22_n_66);
  and mul_102_22_g3456(mul_102_22_n_589 ,mul_102_22_n_140 ,mul_102_22_n_33);
  and mul_102_22_g3457(mul_102_22_n_588 ,mul_102_22_n_90 ,mul_102_22_n_45);
  and mul_102_22_g3458(mul_102_22_n_587 ,mul_102_22_n_132 ,mul_102_22_n_16);
  and mul_102_22_g3459(mul_102_22_n_586 ,mul_102_22_n_128 ,mul_102_22_n_33);
  and mul_102_22_g3460(mul_102_22_n_585 ,mul_102_22_n_110 ,mul_102_22_n_34);
  and mul_102_22_g3461(mul_102_22_n_584 ,mul_102_22_n_92 ,mul_102_22_n_46);
  and mul_102_22_g3462(mul_102_22_n_583 ,mul_102_22_n_142 ,mul_102_22_n_22);
  and mul_102_22_g3463(mul_102_22_n_582 ,mul_102_22_n_144 ,mul_102_22_n_21);
  and mul_102_22_g3464(mul_102_22_n_581 ,mul_102_22_n_134 ,mul_102_22_n_34);
  and mul_102_22_g3465(mul_102_22_n_580 ,mul_102_22_n_138 ,mul_102_22_n_21);
  and mul_102_22_g3466(mul_102_22_n_579 ,mul_102_22_n_120 ,mul_102_22_n_46);
  and mul_102_22_g3467(mul_102_22_n_578 ,mul_102_22_n_94 ,mul_102_22_n_45);
  and mul_102_22_g3468(mul_102_22_n_577 ,mul_102_22_n_126 ,mul_102_22_n_170);
  or mul_102_22_g3469(mul_102_22_n_576 ,mul_102_22_n_351 ,mul_102_22_n_76);
  or mul_102_22_g3470(mul_102_22_n_575 ,mul_102_22_n_328 ,mul_102_22_n_25);
  nor mul_102_22_g3471(mul_102_22_n_574 ,mul_102_22_n_76 ,mul_102_22_n_330);
  or mul_102_22_g3472(mul_102_22_n_573 ,mul_102_22_n_344 ,mul_102_22_n_58);
  or mul_102_22_g3473(mul_102_22_n_572 ,mul_102_22_n_338 ,mul_102_22_n_75);
  or mul_102_22_g3474(mul_102_22_n_571 ,mul_102_22_n_347 ,mul_102_22_n_40);
  or mul_102_22_g3475(mul_102_22_n_570 ,mul_102_22_n_365 ,mul_102_22_n_39);
  and mul_102_22_g3476(mul_102_22_n_569 ,mul_102_22_n_136 ,mul_102_22_n_22);
  or mul_102_22_g3477(mul_102_22_n_568 ,mul_102_22_n_362 ,mul_102_22_n_37);
  or mul_102_22_g3478(mul_102_22_n_567 ,mul_102_22_n_349 ,mul_102_22_n_57);
  or mul_102_22_g3479(mul_102_22_n_566 ,mul_102_22_n_360 ,mul_102_22_n_40);
  or mul_102_22_g3480(mul_102_22_n_565 ,mul_102_22_n_341 ,mul_102_22_n_81);
  or mul_102_22_g3481(mul_102_22_n_564 ,mul_102_22_n_346 ,mul_102_22_n_36);
  or mul_102_22_g3482(mul_102_22_n_563 ,mul_102_22_n_366 ,mul_102_22_n_25);
  or mul_102_22_g3483(mul_102_22_n_562 ,mul_102_22_n_354 ,mul_102_22_n_24);
  or mul_102_22_g3484(mul_102_22_n_561 ,mul_102_22_n_369 ,mul_102_22_n_24);
  or mul_102_22_g3485(mul_102_22_n_560 ,mul_102_22_n_350 ,mul_102_22_n_14);
  or mul_102_22_g3486(mul_102_22_n_559 ,mul_102_22_n_368 ,mul_102_22_n_37);
  or mul_102_22_g3487(mul_102_22_n_558 ,mul_102_22_n_345 ,mul_102_22_n_57);
  or mul_102_22_g3488(mul_102_22_n_557 ,mul_102_22_n_355 ,mul_102_22_n_88);
  or mul_102_22_g3489(mul_102_22_n_556 ,mul_102_22_n_364 ,mul_102_22_n_39);
  or mul_102_22_g3490(mul_102_22_n_555 ,mul_102_22_n_358 ,mul_102_22_n_81);
  or mul_102_22_g3491(mul_102_22_n_554 ,mul_102_22_n_352 ,mul_102_22_n_66);
  or mul_102_22_g3492(mul_102_22_n_553 ,mul_102_22_n_337 ,mul_102_22_n_75);
  or mul_102_22_g3493(mul_102_22_n_552 ,mul_102_22_n_343 ,mul_102_22_n_36);
  or mul_102_22_g3494(mul_102_22_n_551 ,mul_102_22_n_361 ,mul_102_22_n_67);
  or mul_102_22_g3495(mul_102_22_n_550 ,mul_102_22_n_359 ,mul_102_22_n_10);
  or mul_102_22_g3496(mul_102_22_n_549 ,mul_102_22_n_357 ,mul_102_22_n_87);
  or mul_102_22_g3497(mul_102_22_n_548 ,mul_102_22_n_342 ,mul_102_22_n_10);
  not mul_102_22_g3498(mul_102_22_n_545 ,mul_102_22_n_544);
  or mul_102_22_g3499(mul_102_22_n_543 ,mul_102_22_n_392 ,mul_102_22_n_49);
  or mul_102_22_g3500(mul_102_22_n_542 ,mul_102_22_n_356 ,mul_102_22_n_82);
  or mul_102_22_g3501(mul_102_22_n_541 ,mul_102_22_n_340 ,mul_102_22_n_87);
  and mul_102_22_g3502(mul_102_22_n_540 ,mul_102_22_n_165 ,mul_102_22_n_16);
  or mul_102_22_g3503(mul_102_22_n_539 ,mul_102_22_n_377 ,mul_102_22_n_31);
  or mul_102_22_g3504(mul_102_22_n_538 ,mul_102_22_n_388 ,mul_102_22_n_64);
  or mul_102_22_g3505(mul_102_22_n_537 ,mul_102_22_n_407 ,mul_102_22_n_28);
  or mul_102_22_g3506(mul_102_22_n_536 ,mul_102_22_n_370 ,mul_102_22_n_63);
  or mul_102_22_g3507(mul_102_22_n_535 ,mul_102_22_n_405 ,mul_102_22_n_61);
  or mul_102_22_g3508(mul_102_22_n_534 ,mul_102_22_n_404 ,mul_102_22_n_84);
  or mul_102_22_g3509(mul_102_22_n_533 ,mul_102_22_n_386 ,mul_102_22_n_27);
  or mul_102_22_g3510(mul_102_22_n_532 ,mul_102_22_n_399 ,mul_102_22_n_49);
  or mul_102_22_g3511(mul_102_22_n_531 ,mul_102_22_n_390 ,mul_102_22_n_52);
  or mul_102_22_g3512(mul_102_22_n_530 ,mul_102_22_n_339 ,mul_102_22_n_48);
  or mul_102_22_g3513(mul_102_22_n_529 ,mul_102_22_n_410 ,mul_102_22_n_60);
  or mul_102_22_g3514(mul_102_22_n_528 ,mul_102_22_n_385 ,mul_102_22_n_48);
  or mul_102_22_g3515(mul_102_22_n_527 ,mul_102_22_n_389 ,mul_102_22_n_78);
  or mul_102_22_g3516(mul_102_22_n_526 ,mul_102_22_n_408 ,mul_102_22_n_28);
  or mul_102_22_g3517(mul_102_22_n_525 ,mul_102_22_n_397 ,mul_102_22_n_63);
  or mul_102_22_g3518(mul_102_22_n_524 ,mul_102_22_n_395 ,mul_102_22_n_51);
  or mul_102_22_g3519(mul_102_22_n_523 ,mul_102_22_n_403 ,mul_102_22_n_84);
  or mul_102_22_g3520(mul_102_22_n_522 ,mul_102_22_n_348 ,mul_102_22_n_14);
  or mul_102_22_g3521(mul_102_22_n_521 ,mul_102_22_n_406 ,mul_102_22_n_31);
  or mul_102_22_g3522(mul_102_22_n_520 ,mul_102_22_n_396 ,mul_102_22_n_30);
  or mul_102_22_g3523(mul_102_22_n_519 ,mul_102_22_n_363 ,mul_102_22_n_30);
  or mul_102_22_g3524(mul_102_22_n_518 ,mul_102_22_n_391 ,mul_102_22_n_52);
  or mul_102_22_g3525(mul_102_22_n_517 ,mul_102_22_n_394 ,mul_102_22_n_60);
  or mul_102_22_g3526(mul_102_22_n_516 ,mul_102_22_n_400 ,mul_102_22_n_27);
  or mul_102_22_g3527(mul_102_22_n_515 ,mul_102_22_n_387 ,mul_102_22_n_78);
  or mul_102_22_g3528(mul_102_22_n_514 ,mul_102_22_n_384 ,mul_102_22_n_51);
  or mul_102_22_g3529(mul_102_22_n_513 ,mul_102_22_n_409 ,mul_102_22_n_8);
  or mul_102_22_g3530(mul_102_22_n_512 ,mul_102_22_n_393 ,mul_102_22_n_12);
  or mul_102_22_g3531(mul_102_22_n_511 ,mul_102_22_n_401 ,mul_102_22_n_12);
  or mul_102_22_g3532(mul_102_22_n_510 ,mul_102_22_n_367 ,mul_102_22_n_79);
  or mul_102_22_g3533(mul_102_22_n_509 ,mul_102_22_n_402 ,mul_102_22_n_8);
  or mul_102_22_g3534(mul_102_22_n_508 ,mul_102_22_n_398 ,mul_102_22_n_85);
  nor mul_102_22_g3535(mul_102_22_n_507 ,mul_102_22_n_67 ,mul_102_22_n_311);
  nor mul_102_22_g3536(mul_102_22_n_506 ,mul_102_22_n_58 ,mul_102_22_n_310);
  nor mul_102_22_g3537(mul_102_22_n_505 ,mul_102_22_n_61 ,mul_102_22_n_315);
  nor mul_102_22_g3538(mul_102_22_n_504 ,mul_102_22_n_64 ,mul_102_22_n_316);
  and mul_102_22_g3539(mul_102_22_n_547 ,in20[3] ,mul_102_22_n_439);
  and mul_102_22_g3540(mul_102_22_n_546 ,in20[5] ,mul_102_22_n_415);
  or mul_102_22_g3541(mul_102_22_n_544 ,mul_102_22_n_310 ,mul_102_22_n_424);
  and mul_102_22_g3542(mul_102_22_n_503 ,mul_102_22_n_134 ,mul_102_22_n_246);
  and mul_102_22_g3543(mul_102_22_n_502 ,mul_102_22_n_92 ,mul_102_22_n_236);
  and mul_102_22_g3544(mul_102_22_n_501 ,mul_102_22_n_136 ,mul_102_22_n_209);
  and mul_102_22_g3545(mul_102_22_n_500 ,mul_102_22_n_94 ,mul_102_22_n_237);
  and mul_102_22_g3546(mul_102_22_n_499 ,mul_102_22_n_140 ,mul_102_22_n_209);
  and mul_102_22_g3547(mul_102_22_n_498 ,mul_102_22_n_128 ,mul_102_22_n_210);
  and mul_102_22_g3548(mul_102_22_n_497 ,mul_102_22_n_252 ,mul_102_22_n_210);
  and mul_102_22_g3549(mul_102_22_n_496 ,mul_102_22_n_142 ,mul_102_22_n_237);
  and mul_102_22_g3550(mul_102_22_n_495 ,mul_102_22_n_126 ,mul_102_22_n_200);
  and mul_102_22_g3551(mul_102_22_n_494 ,mul_102_22_n_144 ,mul_102_22_n_199);
  and mul_102_22_g3552(mul_102_22_n_493 ,mul_102_22_n_138 ,mul_102_22_n_236);
  and mul_102_22_g3553(mul_102_22_n_492 ,mul_102_22_n_132 ,mul_102_22_n_246);
  and mul_102_22_g3554(mul_102_22_n_491 ,mul_102_22_n_110 ,mul_102_22_n_200);
  and mul_102_22_g3555(mul_102_22_n_490 ,mul_102_22_n_90 ,mul_102_22_n_245);
  and mul_102_22_g3556(mul_102_22_n_489 ,mul_102_22_n_120 ,mul_102_22_n_245);
  or mul_102_22_g3557(mul_102_22_n_488 ,mul_102_22_n_70 ,mul_102_22_n_338);
  or mul_102_22_g3558(mul_102_22_n_487 ,mul_102_22_n_42 ,mul_102_22_n_337);
  nor mul_102_22_g3559(mul_102_22_n_486 ,mul_102_22_n_73 ,mul_102_22_n_365);
  or mul_102_22_g3560(mul_102_22_n_485 ,mul_102_22_n_54 ,mul_102_22_n_357);
  or mul_102_22_g3561(mul_102_22_n_484 ,mul_102_22_n_72 ,mul_102_22_n_340);
  or mul_102_22_g3562(mul_102_22_n_483 ,mul_102_22_n_69 ,mul_102_22_n_352);
  or mul_102_22_g3563(mul_102_22_n_482 ,mul_102_22_n_43 ,mul_102_22_n_353);
  or mul_102_22_g3564(mul_102_22_n_481 ,mul_102_22_n_55 ,mul_102_22_n_348);
  or mul_102_22_g3565(mul_102_22_n_480 ,mul_102_22_n_72 ,mul_102_22_n_361);
  or mul_102_22_g3566(mul_102_22_n_479 ,mul_102_22_n_69 ,mul_102_22_n_360);
  or mul_102_22_g3567(mul_102_22_n_478 ,mul_102_22_n_42 ,mul_102_22_n_347);
  or mul_102_22_g3568(mul_102_22_n_477 ,mul_102_22_n_54 ,mul_102_22_n_364);
  or mul_102_22_g3569(mul_102_22_n_476 ,mul_102_22_n_55 ,mul_102_22_n_355);
  or mul_102_22_g3570(mul_102_22_n_475 ,mul_102_22_n_43 ,mul_102_22_n_350);
  or mul_102_22_g3571(mul_102_22_n_474 ,mul_102_22_n_73 ,mul_102_22_n_351);
  or mul_102_22_g3572(mul_102_22_n_473 ,mul_102_22_n_406 ,mul_102_22_n_224);
  or mul_102_22_g3573(mul_102_22_n_472 ,mul_102_22_n_344 ,mul_102_22_n_215);
  or mul_102_22_g3574(mul_102_22_n_471 ,mul_102_22_n_404 ,mul_102_22_n_239);
  or mul_102_22_g3575(mul_102_22_n_470 ,mul_102_22_n_385 ,mul_102_22_n_206);
  or mul_102_22_g3576(mul_102_22_n_469 ,mul_102_22_n_400 ,mul_102_22_n_206);
  or mul_102_22_g3577(mul_102_22_n_468 ,mul_102_22_n_401 ,mul_102_22_n_233);
  or mul_102_22_g3578(mul_102_22_n_467 ,mul_102_22_n_408 ,mul_102_22_n_240);
  or mul_102_22_g3579(mul_102_22_n_466 ,mul_102_22_n_343 ,mul_102_22_n_218);
  or mul_102_22_g3580(mul_102_22_n_465 ,mul_102_22_n_384 ,mul_102_22_n_233);
  or mul_102_22_g3581(mul_102_22_n_464 ,mul_102_22_n_405 ,mul_102_22_n_225);
  or mul_102_22_g3582(mul_102_22_n_463 ,mul_102_22_n_388 ,mul_102_22_n_243);
  or mul_102_22_g3583(mul_102_22_n_462 ,mul_102_22_n_393 ,mul_102_22_n_228);
  or mul_102_22_g3584(mul_102_22_n_461 ,mul_102_22_n_387 ,mul_102_22_n_224);
  or mul_102_22_g3585(mul_102_22_n_460 ,mul_102_22_n_359 ,mul_102_22_n_218);
  or mul_102_22_g3586(mul_102_22_n_459 ,mul_102_22_n_367 ,mul_102_22_n_227);
  not mul_102_22_g3587(mul_102_22_n_458 ,mul_102_22_n_457);
  not mul_102_22_g3588(mul_102_22_n_455 ,mul_102_22_n_454);
  not mul_102_22_g3589(mul_102_22_n_453 ,mul_102_22_n_452);
  or mul_102_22_g3590(mul_102_22_n_443 ,mul_102_22_n_345 ,mul_102_22_n_216);
  or mul_102_22_g3591(mul_102_22_n_442 ,mul_102_22_n_403 ,mul_102_22_n_239);
  or mul_102_22_g3592(mul_102_22_n_441 ,mul_102_22_n_369 ,mul_102_22_n_249);
  or mul_102_22_g3593(mul_102_22_n_440 ,mul_102_22_n_368 ,mul_102_22_n_215);
  or mul_102_22_g3594(mul_102_22_n_439 ,mul_102_22_n_321 ,mul_102_22_n_376);
  or mul_102_22_g3595(mul_102_22_n_438 ,mul_102_22_n_398 ,mul_102_22_n_242);
  or mul_102_22_g3596(mul_102_22_n_437 ,mul_102_22_n_389 ,mul_102_22_n_230);
  or mul_102_22_g3597(mul_102_22_n_436 ,mul_102_22_n_402 ,mul_102_22_n_212);
  or mul_102_22_g3598(mul_102_22_n_435 ,mul_102_22_n_354 ,mul_102_22_n_248);
  or mul_102_22_g3599(mul_102_22_n_434 ,mul_102_22_n_396 ,mul_102_22_n_230);
  or mul_102_22_g3600(mul_102_22_n_433 ,mul_102_22_n_366 ,mul_102_22_n_221);
  or mul_102_22_g3601(mul_102_22_n_432 ,mul_102_22_n_341 ,mul_102_22_n_221);
  or mul_102_22_g3602(mul_102_22_n_431 ,mul_102_22_n_394 ,mul_102_22_n_227);
  or mul_102_22_g3603(mul_102_22_n_430 ,mul_102_22_n_392 ,mul_102_22_n_212);
  or mul_102_22_g3604(mul_102_22_n_429 ,mul_102_22_n_349 ,mul_102_22_n_248);
  or mul_102_22_g3605(mul_102_22_n_428 ,mul_102_22_n_363 ,mul_102_22_n_234);
  or mul_102_22_g3606(mul_102_22_n_427 ,mul_102_22_n_395 ,mul_102_22_n_228);
  or mul_102_22_g3607(mul_102_22_n_426 ,mul_102_22_n_410 ,mul_102_22_n_231);
  or mul_102_22_g3608(mul_102_22_n_425 ,mul_102_22_n_356 ,mul_102_22_n_219);
  nor mul_102_22_g3609(mul_102_22_n_424 ,mul_102_22_n_320 ,mul_102_22_n_374);
  or mul_102_22_g3610(mul_102_22_n_423 ,mul_102_22_n_386 ,mul_102_22_n_242);
  or mul_102_22_g3611(mul_102_22_n_422 ,mul_102_22_n_399 ,mul_102_22_n_207);
  or mul_102_22_g3612(mul_102_22_n_421 ,mul_102_22_n_358 ,mul_102_22_n_249);
  or mul_102_22_g3613(mul_102_22_n_420 ,mul_102_22_n_346 ,mul_102_22_n_222);
  or mul_102_22_g3614(mul_102_22_n_419 ,mul_102_22_n_390 ,mul_102_22_n_225);
  or mul_102_22_g3615(mul_102_22_n_418 ,mul_102_22_n_391 ,mul_102_22_n_234);
  or mul_102_22_g3616(mul_102_22_n_417 ,mul_102_22_n_342 ,mul_102_22_n_216);
  or mul_102_22_g3617(mul_102_22_n_416 ,mul_102_22_n_397 ,mul_102_22_n_243);
  or mul_102_22_g3618(mul_102_22_n_415 ,mul_102_22_n_326 ,mul_102_22_n_373);
  or mul_102_22_g3619(mul_102_22_n_414 ,mul_102_22_n_407 ,mul_102_22_n_213);
  or mul_102_22_g3620(mul_102_22_n_413 ,mul_102_22_n_339 ,mul_102_22_n_240);
  or mul_102_22_g3621(mul_102_22_n_412 ,mul_102_22_n_362 ,mul_102_22_n_219);
  or mul_102_22_g3622(mul_102_22_n_411 ,mul_102_22_n_409 ,mul_102_22_n_207);
  and mul_102_22_g3623(mul_102_22_n_457 ,in20[7] ,mul_102_22_n_150);
  or mul_102_22_g3624(mul_102_22_n_456 ,mul_102_22_n_159 ,mul_102_22_n_213);
  and mul_102_22_g3625(mul_102_22_n_454 ,in20[3] ,mul_102_22_n_154);
  and mul_102_22_g3626(mul_102_22_n_452 ,in20[5] ,mul_102_22_n_152);
  or mul_102_22_g3627(mul_102_22_n_451 ,mul_102_22_n_163 ,mul_102_22_n_231);
  or mul_102_22_g3628(mul_102_22_n_450 ,mul_102_22_n_162 ,mul_102_22_n_222);
  or mul_102_22_g3629(mul_102_22_n_449 ,mul_102_22_n_162 ,mul_102_22_n_148);
  and mul_102_22_g3630(mul_102_22_n_448 ,in20[8] ,mul_102_22_n_147);
  or mul_102_22_g3631(mul_102_22_n_447 ,mul_102_22_n_371 ,mul_102_22_n_151);
  or mul_102_22_g3632(mul_102_22_n_446 ,in20[0] ,mul_102_22_n_375);
  or mul_102_22_g3633(mul_102_22_n_445 ,mul_102_22_n_329 ,mul_102_22_n_149);
  or mul_102_22_g3634(mul_102_22_n_444 ,mul_102_22_n_372 ,mul_102_22_n_153);
  not mul_102_22_g3635(mul_102_22_n_383 ,mul_102_22_n_152);
  not mul_102_22_g3636(mul_102_22_n_382 ,mul_102_22_n_151);
  not mul_102_22_g3639(mul_102_22_n_380 ,mul_102_22_n_150);
  not mul_102_22_g3640(mul_102_22_n_379 ,mul_102_22_n_149);
  xnor mul_102_22_g3643(mul_102_22_n_377 ,mul_102_22_n_18 ,in20[5]);
  and mul_102_22_g3644(mul_102_22_n_376 ,mul_102_22_n_202 ,mul_102_22_n_322);
  and mul_102_22_g3646(mul_102_22_n_374 ,mul_102_22_n_315 ,mul_102_22_n_319);
  and mul_102_22_g3647(mul_102_22_n_373 ,mul_102_22_n_316 ,mul_102_22_n_323);
  xnor mul_102_22_g3648(mul_102_22_n_372 ,in20[3] ,in20[2]);
  xnor mul_102_22_g3649(mul_102_22_n_371 ,in20[5] ,in20[4]);
  xnor mul_102_22_g3650(mul_102_22_n_370 ,mul_102_22_n_18 ,in20[3]);
  xnor mul_102_22_g3651(mul_102_22_n_410 ,mul_102_22_n_260 ,in20[5]);
  xnor mul_102_22_g3652(mul_102_22_n_409 ,mul_102_22_n_281 ,in20[3]);
  xnor mul_102_22_g3653(mul_102_22_n_408 ,mul_102_22_n_287 ,in20[3]);
  xnor mul_102_22_g3654(mul_102_22_n_407 ,mul_102_22_n_269 ,in20[3]);
  xnor mul_102_22_g3655(mul_102_22_n_406 ,mul_102_22_n_270 ,in20[5]);
  xnor mul_102_22_g3656(mul_102_22_n_405 ,mul_102_22_n_288 ,in20[5]);
  xnor mul_102_22_g3657(mul_102_22_n_404 ,mul_102_22_n_278 ,in20[3]);
  xnor mul_102_22_g3658(mul_102_22_n_403 ,mul_102_22_n_263 ,in20[3]);
  xnor mul_102_22_g3659(mul_102_22_n_402 ,mul_102_22_n_254 ,in20[3]);
  xnor mul_102_22_g3660(mul_102_22_n_401 ,mul_102_22_n_290 ,in20[5]);
  xnor mul_102_22_g3661(mul_102_22_n_400 ,mul_102_22_n_272 ,in20[3]);
  xnor mul_102_22_g3662(mul_102_22_n_399 ,mul_102_22_n_291 ,in20[3]);
  xnor mul_102_22_g3663(mul_102_22_n_398 ,mul_102_22_n_275 ,in20[3]);
  xnor mul_102_22_g3664(mul_102_22_n_397 ,mul_102_22_n_293 ,in20[3]);
  xnor mul_102_22_g3665(mul_102_22_n_396 ,mul_102_22_n_294 ,in20[5]);
  xnor mul_102_22_g3666(mul_102_22_n_395 ,mul_102_22_n_276 ,in20[5]);
  xnor mul_102_22_g3667(mul_102_22_n_394 ,mul_102_22_n_255 ,in20[5]);
  xnor mul_102_22_g3668(mul_102_22_n_393 ,mul_102_22_n_284 ,in20[5]);
  xnor mul_102_22_g3669(mul_102_22_n_392 ,mul_102_22_n_251 ,in20[3]);
  xnor mul_102_22_g3670(mul_102_22_n_391 ,mul_102_22_n_273 ,in20[5]);
  xnor mul_102_22_g3671(mul_102_22_n_390 ,mul_102_22_n_257 ,in20[5]);
  xnor mul_102_22_g3672(mul_102_22_n_389 ,mul_102_22_n_282 ,in20[5]);
  xnor mul_102_22_g3673(mul_102_22_n_388 ,mul_102_22_n_261 ,in20[3]);
  xnor mul_102_22_g3674(mul_102_22_n_387 ,mul_102_22_n_122 ,in20[5]);
  xnor mul_102_22_g3675(mul_102_22_n_386 ,mul_102_22_n_258 ,in20[3]);
  xnor mul_102_22_g3676(mul_102_22_n_385 ,mul_102_22_n_285 ,in20[3]);
  xnor mul_102_22_g3677(mul_102_22_n_384 ,mul_102_22_n_266 ,in20[5]);
  xnor mul_102_22_g3678(mul_102_22_n_381 ,mul_102_22_n_316 ,in20[4]);
  xnor mul_102_22_g3679(mul_102_22_n_378 ,mul_102_22_n_315 ,in20[6]);
  not mul_102_22_g3680(mul_102_22_n_336 ,mul_102_22_n_148);
  not mul_102_22_g3681(mul_102_22_n_335 ,mul_102_22_n_147);
  not mul_102_22_g3684(mul_102_22_n_333 ,mul_102_22_n_154);
  not mul_102_22_g3685(mul_102_22_n_332 ,mul_102_22_n_153);
  xnor mul_102_22_g3689(mul_102_22_n_329 ,in20[7] ,in20[6]);
  xnor mul_102_22_g3690(mul_102_22_n_328 ,mul_102_22_n_168 ,in20[7]);
  xnor mul_102_22_g3691(mul_102_22_n_369 ,mul_102_22_n_98 ,in20[7]);
  xnor mul_102_22_g3692(mul_102_22_n_368 ,mul_102_22_n_100 ,in20[7]);
  xnor mul_102_22_g3693(mul_102_22_n_367 ,mul_102_22_n_264 ,in20[5]);
  xnor mul_102_22_g3694(mul_102_22_n_366 ,mul_102_22_n_112 ,in20[7]);
  xnor mul_102_22_g3695(mul_102_22_n_365 ,mul_102_22_n_114 ,in20[1]);
  xnor mul_102_22_g3696(mul_102_22_n_364 ,mul_102_22_n_251 ,in20[1]);
  xnor mul_102_22_g3697(mul_102_22_n_363 ,mul_102_22_n_279 ,in20[5]);
  xnor mul_102_22_g3698(mul_102_22_n_362 ,mul_102_22_n_146 ,in20[7]);
  xnor mul_102_22_g3699(mul_102_22_n_361 ,mul_102_22_n_124 ,in20[1]);
  xnor mul_102_22_g3700(mul_102_22_n_360 ,mul_102_22_n_102 ,in20[1]);
  xnor mul_102_22_g3701(mul_102_22_n_359 ,mul_102_22_n_124 ,in20[7]);
  xnor mul_102_22_g3702(mul_102_22_n_358 ,mul_102_22_n_114 ,in20[7]);
  xnor mul_102_22_g3703(mul_102_22_n_357 ,mul_102_22_n_98 ,in20[1]);
  xnor mul_102_22_g3704(mul_102_22_n_356 ,mul_102_22_n_118 ,in20[7]);
  xnor mul_102_22_g3705(mul_102_22_n_355 ,mul_102_22_n_108 ,in20[1]);
  xnor mul_102_22_g3706(mul_102_22_n_354 ,mul_102_22_n_108 ,in20[7]);
  xnor mul_102_22_g3707(mul_102_22_n_353 ,mul_102_22_n_106 ,in20[1]);
  xnor mul_102_22_g3708(mul_102_22_n_352 ,mul_102_22_n_96 ,in20[1]);
  xnor mul_102_22_g3709(mul_102_22_n_351 ,mul_102_22_n_118 ,in20[1]);
  xnor mul_102_22_g3710(mul_102_22_n_350 ,mul_102_22_n_104 ,in20[1]);
  xnor mul_102_22_g3711(mul_102_22_n_349 ,mul_102_22_n_116 ,in20[7]);
  xnor mul_102_22_g3712(mul_102_22_n_348 ,mul_102_22_n_146 ,in20[1]);
  xnor mul_102_22_g3713(mul_102_22_n_347 ,mul_102_22_n_267 ,in20[1]);
  xnor mul_102_22_g3714(mul_102_22_n_346 ,mul_102_22_n_122 ,in20[7]);
  xnor mul_102_22_g3715(mul_102_22_n_345 ,mul_102_22_n_130 ,in20[7]);
  xnor mul_102_22_g3716(mul_102_22_n_344 ,mul_102_22_n_104 ,in20[7]);
  xnor mul_102_22_g3717(mul_102_22_n_343 ,mul_102_22_n_102 ,in20[7]);
  xnor mul_102_22_g3718(mul_102_22_n_342 ,mul_102_22_n_96 ,in20[7]);
  xnor mul_102_22_g3719(mul_102_22_n_341 ,mul_102_22_n_106 ,in20[7]);
  xnor mul_102_22_g3720(mul_102_22_n_340 ,mul_102_22_n_116 ,in20[1]);
  xnor mul_102_22_g3721(mul_102_22_n_339 ,mul_102_22_n_130 ,in20[3]);
  xnor mul_102_22_g3722(mul_102_22_n_338 ,mul_102_22_n_112 ,in20[1]);
  xnor mul_102_22_g3723(mul_102_22_n_337 ,mul_102_22_n_100 ,in20[1]);
  xnor mul_102_22_g3724(mul_102_22_n_334 ,in20[8] ,in20[7]);
  xnor mul_102_22_g3725(mul_102_22_n_331 ,mul_102_22_n_202 ,in20[2]);
  nor mul_102_22_g3726(mul_102_22_n_327 ,mul_102_22_n_70 ,mul_102_22_n_163);
  nor mul_102_22_g3727(mul_102_22_n_326 ,mul_102_22_n_166 ,in20[4]);
  not mul_102_22_g3728(mul_102_22_n_325 ,mul_102_22_n_324);
  and mul_102_22_g3729(mul_102_22_n_324 ,in20[1] ,in20[0]);
  or mul_102_22_g3730(mul_102_22_n_323 ,mul_102_22_n_159 ,mul_102_22_n_313);
  or mul_102_22_g3731(mul_102_22_n_322 ,mul_102_22_n_160 ,mul_102_22_n_318);
  nor mul_102_22_g3732(mul_102_22_n_321 ,mul_102_22_n_19 ,in20[2]);
  nor mul_102_22_g3733(mul_102_22_n_320 ,mul_102_22_n_168 ,in20[6]);
  or mul_102_22_g3734(mul_102_22_n_319 ,mul_102_22_n_160 ,mul_102_22_n_314);
  not mul_102_22_g3735(mul_102_22_n_318 ,in20[2]);
  not mul_102_22_g3736(mul_102_22_n_317 ,in20[0]);
  not mul_102_22_g3737(mul_102_22_n_316 ,in20[3]);
  not mul_102_22_g3738(mul_102_22_n_315 ,in20[5]);
  not mul_102_22_g3739(mul_102_22_n_314 ,in20[6]);
  not mul_102_22_g3740(mul_102_22_n_313 ,in20[4]);
  not mul_102_22_g3741(mul_102_22_n_312 ,mul_102_22_n_165);
  not mul_102_22_g3742(mul_102_22_n_311 ,in20[1]);
  not mul_102_22_g3743(mul_102_22_n_310 ,in20[7]);
  not mul_102_22_drc_bufs3784(mul_102_22_n_297 ,mul_102_22_n_295);
  not mul_102_22_drc_bufs3785(mul_102_22_n_296 ,mul_102_22_n_295);
  not mul_102_22_drc_bufs3786(mul_102_22_n_295 ,n_223);
  not mul_102_22_drc_bufs3814(mul_102_22_n_294 ,mul_102_22_n_292);
  not mul_102_22_drc_bufs3815(mul_102_22_n_293 ,mul_102_22_n_292);
  not mul_102_22_drc_bufs3816(mul_102_22_n_292 ,n_226);
  not mul_102_22_drc_bufs3818(mul_102_22_n_291 ,mul_102_22_n_289);
  not mul_102_22_drc_bufs3819(mul_102_22_n_290 ,mul_102_22_n_289);
  not mul_102_22_drc_bufs3820(mul_102_22_n_289 ,n_224);
  not mul_102_22_drc_bufs3822(mul_102_22_n_288 ,mul_102_22_n_286);
  not mul_102_22_drc_bufs3823(mul_102_22_n_287 ,mul_102_22_n_286);
  not mul_102_22_drc_bufs3824(mul_102_22_n_286 ,n_230);
  not mul_102_22_drc_bufs3826(mul_102_22_n_285 ,mul_102_22_n_283);
  not mul_102_22_drc_bufs3827(mul_102_22_n_284 ,mul_102_22_n_283);
  not mul_102_22_drc_bufs3828(mul_102_22_n_283 ,n_231);
  not mul_102_22_drc_bufs3830(mul_102_22_n_282 ,mul_102_22_n_280);
  not mul_102_22_drc_bufs3831(mul_102_22_n_281 ,mul_102_22_n_280);
  not mul_102_22_drc_bufs3832(mul_102_22_n_280 ,n_227);
  not mul_102_22_drc_bufs3834(mul_102_22_n_279 ,mul_102_22_n_277);
  not mul_102_22_drc_bufs3835(mul_102_22_n_278 ,mul_102_22_n_277);
  not mul_102_22_drc_bufs3836(mul_102_22_n_277 ,n_232);
  not mul_102_22_drc_bufs3838(mul_102_22_n_276 ,mul_102_22_n_274);
  not mul_102_22_drc_bufs3839(mul_102_22_n_275 ,mul_102_22_n_274);
  not mul_102_22_drc_bufs3840(mul_102_22_n_274 ,n_233);
  not mul_102_22_drc_bufs3842(mul_102_22_n_273 ,mul_102_22_n_271);
  not mul_102_22_drc_bufs3843(mul_102_22_n_272 ,mul_102_22_n_271);
  not mul_102_22_drc_bufs3844(mul_102_22_n_271 ,n_228);
  not mul_102_22_drc_bufs3846(mul_102_22_n_270 ,mul_102_22_n_268);
  not mul_102_22_drc_bufs3847(mul_102_22_n_269 ,mul_102_22_n_268);
  not mul_102_22_drc_bufs3848(mul_102_22_n_268 ,n_234);
  not mul_102_22_drc_bufs3850(mul_102_22_n_267 ,mul_102_22_n_265);
  not mul_102_22_drc_bufs3851(mul_102_22_n_266 ,mul_102_22_n_265);
  not mul_102_22_drc_bufs3852(mul_102_22_n_265 ,n_225);
  not mul_102_22_drc_bufs3854(mul_102_22_n_264 ,mul_102_22_n_262);
  not mul_102_22_drc_bufs3855(mul_102_22_n_263 ,mul_102_22_n_262);
  not mul_102_22_drc_bufs3856(mul_102_22_n_262 ,n_235);
  not mul_102_22_drc_bufs3858(mul_102_22_n_261 ,mul_102_22_n_259);
  not mul_102_22_drc_bufs3859(mul_102_22_n_260 ,mul_102_22_n_259);
  not mul_102_22_drc_bufs3860(mul_102_22_n_259 ,n_229);
  not mul_102_22_drc_bufs3862(mul_102_22_n_258 ,mul_102_22_n_256);
  not mul_102_22_drc_bufs3863(mul_102_22_n_257 ,mul_102_22_n_256);
  not mul_102_22_drc_bufs3864(mul_102_22_n_256 ,n_236);
  not mul_102_22_drc_bufs3866(mul_102_22_n_255 ,mul_102_22_n_253);
  not mul_102_22_drc_bufs3867(mul_102_22_n_254 ,mul_102_22_n_253);
  not mul_102_22_drc_bufs3868(mul_102_22_n_253 ,n_237);
  not mul_102_22_drc_bufs3870(mul_102_22_n_252 ,mul_102_22_n_250);
  not mul_102_22_drc_bufs3871(mul_102_22_n_251 ,mul_102_22_n_250);
  not mul_102_22_drc_bufs3872(mul_102_22_n_250 ,n_238);
  not mul_102_22_drc_bufs3874(mul_102_22_n_249 ,mul_102_22_n_247);
  not mul_102_22_drc_bufs3875(mul_102_22_n_248 ,mul_102_22_n_247);
  not mul_102_22_drc_bufs3876(mul_102_22_n_247 ,mul_102_22_n_303);
  not mul_102_22_drc_bufs3878(mul_102_22_n_246 ,mul_102_22_n_244);
  not mul_102_22_drc_bufs3879(mul_102_22_n_245 ,mul_102_22_n_244);
  not mul_102_22_drc_bufs3880(mul_102_22_n_244 ,mul_102_22_n_335);
  not mul_102_22_drc_bufs3882(mul_102_22_n_243 ,mul_102_22_n_241);
  not mul_102_22_drc_bufs3883(mul_102_22_n_242 ,mul_102_22_n_241);
  not mul_102_22_drc_bufs3884(mul_102_22_n_241 ,mul_102_22_n_299);
  not mul_102_22_drc_bufs3886(mul_102_22_n_240 ,mul_102_22_n_238);
  not mul_102_22_drc_bufs3887(mul_102_22_n_239 ,mul_102_22_n_238);
  not mul_102_22_drc_bufs3888(mul_102_22_n_238 ,mul_102_22_n_298);
  not mul_102_22_drc_bufs3890(mul_102_22_n_237 ,mul_102_22_n_235);
  not mul_102_22_drc_bufs3891(mul_102_22_n_236 ,mul_102_22_n_235);
  not mul_102_22_drc_bufs3892(mul_102_22_n_235 ,mul_102_22_n_336);
  not mul_102_22_drc_bufs3894(mul_102_22_n_234 ,mul_102_22_n_232);
  not mul_102_22_drc_bufs3895(mul_102_22_n_233 ,mul_102_22_n_232);
  not mul_102_22_drc_bufs3896(mul_102_22_n_232 ,mul_102_22_n_383);
  not mul_102_22_drc_bufs3898(mul_102_22_n_231 ,mul_102_22_n_229);
  not mul_102_22_drc_bufs3899(mul_102_22_n_230 ,mul_102_22_n_229);
  not mul_102_22_drc_bufs3900(mul_102_22_n_229 ,mul_102_22_n_382);
  not mul_102_22_drc_bufs3902(mul_102_22_n_228 ,mul_102_22_n_226);
  not mul_102_22_drc_bufs3903(mul_102_22_n_227 ,mul_102_22_n_226);
  not mul_102_22_drc_bufs3904(mul_102_22_n_226 ,mul_102_22_n_305);
  not mul_102_22_drc_bufs3906(mul_102_22_n_225 ,mul_102_22_n_223);
  not mul_102_22_drc_bufs3907(mul_102_22_n_224 ,mul_102_22_n_223);
  not mul_102_22_drc_bufs3908(mul_102_22_n_223 ,mul_102_22_n_304);
  not mul_102_22_drc_bufs3910(mul_102_22_n_222 ,mul_102_22_n_220);
  not mul_102_22_drc_bufs3911(mul_102_22_n_221 ,mul_102_22_n_220);
  not mul_102_22_drc_bufs3912(mul_102_22_n_220 ,mul_102_22_n_379);
  not mul_102_22_drc_bufs3914(mul_102_22_n_219 ,mul_102_22_n_217);
  not mul_102_22_drc_bufs3915(mul_102_22_n_218 ,mul_102_22_n_217);
  not mul_102_22_drc_bufs3916(mul_102_22_n_217 ,mul_102_22_n_380);
  not mul_102_22_drc_bufs3918(mul_102_22_n_216 ,mul_102_22_n_214);
  not mul_102_22_drc_bufs3919(mul_102_22_n_215 ,mul_102_22_n_214);
  not mul_102_22_drc_bufs3920(mul_102_22_n_214 ,mul_102_22_n_302);
  not mul_102_22_drc_bufs3922(mul_102_22_n_213 ,mul_102_22_n_211);
  not mul_102_22_drc_bufs3923(mul_102_22_n_212 ,mul_102_22_n_211);
  not mul_102_22_drc_bufs3924(mul_102_22_n_211 ,mul_102_22_n_332);
  not mul_102_22_drc_bufs3926(mul_102_22_n_210 ,mul_102_22_n_208);
  not mul_102_22_drc_bufs3927(mul_102_22_n_209 ,mul_102_22_n_208);
  not mul_102_22_drc_bufs3928(mul_102_22_n_208 ,mul_102_22_n_300);
  not mul_102_22_drc_bufs3930(mul_102_22_n_207 ,mul_102_22_n_205);
  not mul_102_22_drc_bufs3931(mul_102_22_n_206 ,mul_102_22_n_205);
  not mul_102_22_drc_bufs3932(mul_102_22_n_205 ,mul_102_22_n_333);
  not mul_102_22_drc_bufs3934(mul_102_22_n_204 ,mul_102_22_n_649);
  not mul_102_22_drc_bufs3935(mul_102_22_n_203 ,mul_102_22_n_649);
  not mul_102_22_drc_bufs3940(mul_102_22_n_307 ,mul_102_22_n_650);
  not mul_102_22_drc_bufs3943(mul_102_22_n_202 ,mul_102_22_n_201);
  not mul_102_22_drc_bufs3944(mul_102_22_n_201 ,mul_102_22_n_311);
  not mul_102_22_drc_bufs3946(mul_102_22_n_200 ,mul_102_22_n_198);
  not mul_102_22_drc_bufs3947(mul_102_22_n_199 ,mul_102_22_n_198);
  not mul_102_22_drc_bufs3948(mul_102_22_n_198 ,mul_102_22_n_301);
  buf mul_102_22_drc_bufs3957(n_216 ,mul_102_22_n_1140);
  buf mul_102_22_drc_bufs3958(n_217 ,mul_102_22_n_1143);
  buf mul_102_22_drc_bufs3959(n_210 ,mul_102_22_n_1121);
  buf mul_102_22_drc_bufs3960(n_212 ,mul_102_22_n_1127);
  buf mul_102_22_drc_bufs3961(n_213 ,mul_102_22_n_1130);
  buf mul_102_22_drc_bufs3962(n_220 ,mul_102_22_n_1153);
  buf mul_102_22_drc_bufs3963(n_215 ,mul_102_22_n_1137);
  buf mul_102_22_drc_bufs3964(n_214 ,mul_102_22_n_1134);
  buf mul_102_22_drc_bufs3965(n_211 ,mul_102_22_n_1124);
  buf mul_102_22_drc_bufs3966(n_221 ,mul_102_22_n_1156);
  buf mul_102_22_drc_bufs3967(n_218 ,mul_102_22_n_1147);
  buf mul_102_22_drc_bufs3968(n_219 ,mul_102_22_n_1150);
  buf mul_102_22_drc_bufs3969(n_207 ,mul_102_22_n_1112);
  buf mul_102_22_drc_bufs3970(n_208 ,mul_102_22_n_1115);
  buf mul_102_22_drc_bufs3971(n_209 ,mul_102_22_n_1118);
  not mul_102_22_drc_bufs3973(mul_102_22_n_182 ,mul_102_22_n_308);
  not mul_102_22_drc_bufs3974(mul_102_22_n_308 ,mul_102_22_n_885);
  not mul_102_22_drc_bufs3996(mul_102_22_n_181 ,mul_102_22_n_180);
  not mul_102_22_drc_bufs3998(mul_102_22_n_180 ,mul_102_22_n_446);
  not mul_102_22_drc_bufs4001(mul_102_22_n_179 ,mul_102_22_n_178);
  not mul_102_22_drc_bufs4003(mul_102_22_n_178 ,mul_102_22_n_444);
  not mul_102_22_drc_bufs4006(mul_102_22_n_177 ,mul_102_22_n_176);
  not mul_102_22_drc_bufs4008(mul_102_22_n_176 ,mul_102_22_n_447);
  not mul_102_22_drc_bufs4011(mul_102_22_n_175 ,mul_102_22_n_174);
  not mul_102_22_drc_bufs4013(mul_102_22_n_174 ,mul_102_22_n_445);
  not mul_102_22_drc_bufs4021(mul_102_22_n_173 ,mul_102_22_n_172);
  not mul_102_22_drc_bufs4023(mul_102_22_n_172 ,mul_102_22_n_317);
  not mul_102_22_drc_bufs4031(mul_102_22_n_171 ,mul_102_22_n_169);
  not mul_102_22_drc_bufs4032(mul_102_22_n_170 ,mul_102_22_n_169);
  not mul_102_22_drc_bufs4033(mul_102_22_n_169 ,mul_102_22_n_448);
  not mul_102_22_drc_bufs4036(mul_102_22_n_168 ,mul_102_22_n_167);
  not mul_102_22_drc_bufs4037(mul_102_22_n_167 ,mul_102_22_n_297);
  not mul_102_22_drc_bufs4039(mul_102_22_n_166 ,mul_102_22_n_164);
  not mul_102_22_drc_bufs4040(mul_102_22_n_165 ,mul_102_22_n_164);
  not mul_102_22_drc_bufs4041(mul_102_22_n_164 ,mul_102_22_n_296);
  not mul_102_22_drc_bufs4043(mul_102_22_n_163 ,mul_102_22_n_161);
  not mul_102_22_drc_bufs4044(mul_102_22_n_162 ,mul_102_22_n_161);
  not mul_102_22_drc_bufs4045(mul_102_22_n_161 ,mul_102_22_n_312);
  not mul_102_22_drc_bufs4047(mul_102_22_n_160 ,mul_102_22_n_158);
  not mul_102_22_drc_bufs4048(mul_102_22_n_159 ,mul_102_22_n_158);
  not mul_102_22_drc_bufs4049(mul_102_22_n_158 ,mul_102_22_n_312);
  not mul_102_22_drc_bufs4051(mul_102_22_n_157 ,mul_102_22_n_306);
  not mul_102_22_drc_bufs4053(mul_102_22_n_306 ,mul_102_22_n_648);
  not mul_102_22_drc_bufs4056(mul_102_22_n_156 ,mul_102_22_n_155);
  not mul_102_22_drc_bufs4057(mul_102_22_n_155 ,mul_102_22_n_648);
  not mul_102_22_drc_bufs4059(mul_102_22_n_154 ,mul_102_22_n_299);
  not mul_102_22_drc_bufs4061(mul_102_22_n_299 ,mul_102_22_n_331);
  not mul_102_22_drc_bufs4063(mul_102_22_n_153 ,mul_102_22_n_298);
  not mul_102_22_drc_bufs4065(mul_102_22_n_298 ,mul_102_22_n_331);
  not mul_102_22_drc_bufs4067(mul_102_22_n_152 ,mul_102_22_n_305);
  not mul_102_22_drc_bufs4069(mul_102_22_n_305 ,mul_102_22_n_381);
  not mul_102_22_drc_bufs4071(mul_102_22_n_151 ,mul_102_22_n_304);
  not mul_102_22_drc_bufs4073(mul_102_22_n_304 ,mul_102_22_n_381);
  not mul_102_22_drc_bufs4075(mul_102_22_n_150 ,mul_102_22_n_303);
  not mul_102_22_drc_bufs4077(mul_102_22_n_303 ,mul_102_22_n_378);
  not mul_102_22_drc_bufs4079(mul_102_22_n_149 ,mul_102_22_n_302);
  not mul_102_22_drc_bufs4081(mul_102_22_n_302 ,mul_102_22_n_378);
  not mul_102_22_drc_bufs4083(mul_102_22_n_148 ,mul_102_22_n_301);
  not mul_102_22_drc_bufs4085(mul_102_22_n_301 ,mul_102_22_n_334);
  not mul_102_22_drc_bufs4087(mul_102_22_n_147 ,mul_102_22_n_300);
  not mul_102_22_drc_bufs4089(mul_102_22_n_300 ,mul_102_22_n_334);
  not mul_102_22_drc_bufs4091(mul_102_22_n_146 ,mul_102_22_n_145);
  not mul_102_22_drc_bufs4093(mul_102_22_n_145 ,mul_102_22_n_281);
  not mul_102_22_drc_bufs4095(mul_102_22_n_144 ,mul_102_22_n_143);
  not mul_102_22_drc_bufs4097(mul_102_22_n_143 ,mul_102_22_n_291);
  not mul_102_22_drc_bufs4099(mul_102_22_n_142 ,mul_102_22_n_141);
  not mul_102_22_drc_bufs4101(mul_102_22_n_141 ,mul_102_22_n_273);
  not mul_102_22_drc_bufs4103(mul_102_22_n_140 ,mul_102_22_n_139);
  not mul_102_22_drc_bufs4105(mul_102_22_n_139 ,mul_102_22_n_294);
  not mul_102_22_drc_bufs4107(mul_102_22_n_138 ,mul_102_22_n_137);
  not mul_102_22_drc_bufs4109(mul_102_22_n_137 ,mul_102_22_n_255);
  not mul_102_22_drc_bufs4111(mul_102_22_n_136 ,mul_102_22_n_135);
  not mul_102_22_drc_bufs4113(mul_102_22_n_135 ,mul_102_22_n_282);
  not mul_102_22_drc_bufs4115(mul_102_22_n_134 ,mul_102_22_n_133);
  not mul_102_22_drc_bufs4117(mul_102_22_n_133 ,mul_102_22_n_261);
  not mul_102_22_drc_bufs4119(mul_102_22_n_132 ,mul_102_22_n_131);
  not mul_102_22_drc_bufs4121(mul_102_22_n_131 ,mul_102_22_n_264);
  not mul_102_22_drc_bufs4123(mul_102_22_n_130 ,mul_102_22_n_129);
  not mul_102_22_drc_bufs4125(mul_102_22_n_129 ,mul_102_22_n_266);
  not mul_102_22_drc_bufs4127(mul_102_22_n_128 ,mul_102_22_n_127);
  not mul_102_22_drc_bufs4129(mul_102_22_n_127 ,mul_102_22_n_276);
  not mul_102_22_drc_bufs4131(mul_102_22_n_126 ,mul_102_22_n_125);
  not mul_102_22_drc_bufs4133(mul_102_22_n_125 ,mul_102_22_n_258);
  not mul_102_22_drc_bufs4135(mul_102_22_n_124 ,mul_102_22_n_123);
  not mul_102_22_drc_bufs4137(mul_102_22_n_123 ,mul_102_22_n_260);
  not mul_102_22_drc_bufs4139(mul_102_22_n_122 ,mul_102_22_n_121);
  not mul_102_22_drc_bufs4141(mul_102_22_n_121 ,mul_102_22_n_252);
  not mul_102_22_drc_bufs4143(mul_102_22_n_120 ,mul_102_22_n_119);
  not mul_102_22_drc_bufs4145(mul_102_22_n_119 ,mul_102_22_n_270);
  not mul_102_22_drc_bufs4147(mul_102_22_n_118 ,mul_102_22_n_117);
  not mul_102_22_drc_bufs4149(mul_102_22_n_117 ,mul_102_22_n_254);
  not mul_102_22_drc_bufs4151(mul_102_22_n_116 ,mul_102_22_n_115);
  not mul_102_22_drc_bufs4153(mul_102_22_n_115 ,mul_102_22_n_263);
  not mul_102_22_drc_bufs4155(mul_102_22_n_114 ,mul_102_22_n_113);
  not mul_102_22_drc_bufs4157(mul_102_22_n_113 ,mul_102_22_n_290);
  not mul_102_22_drc_bufs4159(mul_102_22_n_112 ,mul_102_22_n_111);
  not mul_102_22_drc_bufs4161(mul_102_22_n_111 ,mul_102_22_n_293);
  not mul_102_22_drc_bufs4163(mul_102_22_n_110 ,mul_102_22_n_109);
  not mul_102_22_drc_bufs4165(mul_102_22_n_109 ,mul_102_22_n_267);
  not mul_102_22_drc_bufs4167(mul_102_22_n_108 ,mul_102_22_n_107);
  not mul_102_22_drc_bufs4169(mul_102_22_n_107 ,mul_102_22_n_284);
  not mul_102_22_drc_bufs4171(mul_102_22_n_106 ,mul_102_22_n_105);
  not mul_102_22_drc_bufs4173(mul_102_22_n_105 ,mul_102_22_n_269);
  not mul_102_22_drc_bufs4175(mul_102_22_n_104 ,mul_102_22_n_103);
  not mul_102_22_drc_bufs4177(mul_102_22_n_103 ,mul_102_22_n_278);
  not mul_102_22_drc_bufs4179(mul_102_22_n_102 ,mul_102_22_n_101);
  not mul_102_22_drc_bufs4181(mul_102_22_n_101 ,mul_102_22_n_275);
  not mul_102_22_drc_bufs4183(mul_102_22_n_100 ,mul_102_22_n_99);
  not mul_102_22_drc_bufs4185(mul_102_22_n_99 ,mul_102_22_n_257);
  not mul_102_22_drc_bufs4187(mul_102_22_n_98 ,mul_102_22_n_97);
  not mul_102_22_drc_bufs4189(mul_102_22_n_97 ,mul_102_22_n_272);
  not mul_102_22_drc_bufs4191(mul_102_22_n_96 ,mul_102_22_n_95);
  not mul_102_22_drc_bufs4193(mul_102_22_n_95 ,mul_102_22_n_287);
  not mul_102_22_drc_bufs4195(mul_102_22_n_94 ,mul_102_22_n_93);
  not mul_102_22_drc_bufs4197(mul_102_22_n_93 ,mul_102_22_n_285);
  not mul_102_22_drc_bufs4199(mul_102_22_n_92 ,mul_102_22_n_91);
  not mul_102_22_drc_bufs4201(mul_102_22_n_91 ,mul_102_22_n_279);
  not mul_102_22_drc_bufs4203(mul_102_22_n_90 ,mul_102_22_n_89);
  not mul_102_22_drc_bufs4205(mul_102_22_n_89 ,mul_102_22_n_288);
  not mul_102_22_drc_bufs4207(mul_102_22_n_88 ,mul_102_22_n_86);
  not mul_102_22_drc_bufs4208(mul_102_22_n_87 ,mul_102_22_n_86);
  not mul_102_22_drc_bufs4209(mul_102_22_n_86 ,mul_102_22_n_446);
  not mul_102_22_drc_bufs4211(mul_102_22_n_85 ,mul_102_22_n_83);
  not mul_102_22_drc_bufs4212(mul_102_22_n_84 ,mul_102_22_n_83);
  not mul_102_22_drc_bufs4213(mul_102_22_n_83 ,mul_102_22_n_444);
  not mul_102_22_drc_bufs4215(mul_102_22_n_82 ,mul_102_22_n_80);
  not mul_102_22_drc_bufs4216(mul_102_22_n_81 ,mul_102_22_n_80);
  not mul_102_22_drc_bufs4217(mul_102_22_n_80 ,mul_102_22_n_445);
  not mul_102_22_drc_bufs4219(mul_102_22_n_79 ,mul_102_22_n_77);
  not mul_102_22_drc_bufs4220(mul_102_22_n_78 ,mul_102_22_n_77);
  not mul_102_22_drc_bufs4221(mul_102_22_n_77 ,mul_102_22_n_447);
  not mul_102_22_drc_bufs4223(mul_102_22_n_76 ,mul_102_22_n_74);
  not mul_102_22_drc_bufs4224(mul_102_22_n_75 ,mul_102_22_n_74);
  not mul_102_22_drc_bufs4225(mul_102_22_n_74 ,mul_102_22_n_181);
  not mul_102_22_drc_bufs4227(mul_102_22_n_73 ,mul_102_22_n_71);
  not mul_102_22_drc_bufs4228(mul_102_22_n_72 ,mul_102_22_n_71);
  not mul_102_22_drc_bufs4229(mul_102_22_n_71 ,mul_102_22_n_317);
  not mul_102_22_drc_bufs4231(mul_102_22_n_70 ,mul_102_22_n_68);
  not mul_102_22_drc_bufs4232(mul_102_22_n_69 ,mul_102_22_n_68);
  not mul_102_22_drc_bufs4233(mul_102_22_n_68 ,mul_102_22_n_173);
  not mul_102_22_drc_bufs4235(mul_102_22_n_67 ,mul_102_22_n_65);
  not mul_102_22_drc_bufs4236(mul_102_22_n_66 ,mul_102_22_n_65);
  not mul_102_22_drc_bufs4237(mul_102_22_n_65 ,mul_102_22_n_446);
  not mul_102_22_drc_bufs4239(mul_102_22_n_64 ,mul_102_22_n_62);
  not mul_102_22_drc_bufs4240(mul_102_22_n_63 ,mul_102_22_n_62);
  not mul_102_22_drc_bufs4241(mul_102_22_n_62 ,mul_102_22_n_179);
  not mul_102_22_drc_bufs4243(mul_102_22_n_61 ,mul_102_22_n_59);
  not mul_102_22_drc_bufs4244(mul_102_22_n_60 ,mul_102_22_n_59);
  not mul_102_22_drc_bufs4245(mul_102_22_n_59 ,mul_102_22_n_177);
  not mul_102_22_drc_bufs4247(mul_102_22_n_58 ,mul_102_22_n_56);
  not mul_102_22_drc_bufs4248(mul_102_22_n_57 ,mul_102_22_n_56);
  not mul_102_22_drc_bufs4249(mul_102_22_n_56 ,mul_102_22_n_175);
  not mul_102_22_drc_bufs4251(mul_102_22_n_55 ,mul_102_22_n_53);
  not mul_102_22_drc_bufs4252(mul_102_22_n_54 ,mul_102_22_n_53);
  not mul_102_22_drc_bufs4253(mul_102_22_n_53 ,mul_102_22_n_317);
  not mul_102_22_drc_bufs4255(mul_102_22_n_52 ,mul_102_22_n_50);
  not mul_102_22_drc_bufs4256(mul_102_22_n_51 ,mul_102_22_n_50);
  not mul_102_22_drc_bufs4257(mul_102_22_n_50 ,mul_102_22_n_177);
  not mul_102_22_drc_bufs4259(mul_102_22_n_49 ,mul_102_22_n_47);
  not mul_102_22_drc_bufs4260(mul_102_22_n_48 ,mul_102_22_n_47);
  not mul_102_22_drc_bufs4261(mul_102_22_n_47 ,mul_102_22_n_444);
  not mul_102_22_drc_bufs4263(mul_102_22_n_46 ,mul_102_22_n_44);
  not mul_102_22_drc_bufs4264(mul_102_22_n_45 ,mul_102_22_n_44);
  not mul_102_22_drc_bufs4265(mul_102_22_n_44 ,mul_102_22_n_448);
  not mul_102_22_drc_bufs4267(mul_102_22_n_43 ,mul_102_22_n_41);
  not mul_102_22_drc_bufs4268(mul_102_22_n_42 ,mul_102_22_n_41);
  not mul_102_22_drc_bufs4269(mul_102_22_n_41 ,mul_102_22_n_173);
  not mul_102_22_drc_bufs4271(mul_102_22_n_40 ,mul_102_22_n_38);
  not mul_102_22_drc_bufs4272(mul_102_22_n_39 ,mul_102_22_n_38);
  not mul_102_22_drc_bufs4273(mul_102_22_n_38 ,mul_102_22_n_181);
  not mul_102_22_drc_bufs4275(mul_102_22_n_37 ,mul_102_22_n_35);
  not mul_102_22_drc_bufs4276(mul_102_22_n_36 ,mul_102_22_n_35);
  not mul_102_22_drc_bufs4277(mul_102_22_n_35 ,mul_102_22_n_175);
  not mul_102_22_drc_bufs4279(mul_102_22_n_34 ,mul_102_22_n_32);
  not mul_102_22_drc_bufs4280(mul_102_22_n_33 ,mul_102_22_n_32);
  not mul_102_22_drc_bufs4281(mul_102_22_n_32 ,mul_102_22_n_448);
  not mul_102_22_drc_bufs4283(mul_102_22_n_31 ,mul_102_22_n_29);
  not mul_102_22_drc_bufs4284(mul_102_22_n_30 ,mul_102_22_n_29);
  not mul_102_22_drc_bufs4285(mul_102_22_n_29 ,mul_102_22_n_447);
  not mul_102_22_drc_bufs4287(mul_102_22_n_28 ,mul_102_22_n_26);
  not mul_102_22_drc_bufs4288(mul_102_22_n_27 ,mul_102_22_n_26);
  not mul_102_22_drc_bufs4289(mul_102_22_n_26 ,mul_102_22_n_179);
  not mul_102_22_drc_bufs4291(mul_102_22_n_25 ,mul_102_22_n_23);
  not mul_102_22_drc_bufs4292(mul_102_22_n_24 ,mul_102_22_n_23);
  not mul_102_22_drc_bufs4293(mul_102_22_n_23 ,mul_102_22_n_445);
  not mul_102_22_drc_bufs4295(mul_102_22_n_22 ,mul_102_22_n_20);
  not mul_102_22_drc_bufs4296(mul_102_22_n_21 ,mul_102_22_n_20);
  not mul_102_22_drc_bufs4297(mul_102_22_n_20 ,mul_102_22_n_171);
  not mul_102_22_drc_bufs4299(mul_102_22_n_19 ,mul_102_22_n_17);
  not mul_102_22_drc_bufs4300(mul_102_22_n_18 ,mul_102_22_n_17);
  not mul_102_22_drc_bufs4301(mul_102_22_n_17 ,mul_102_22_n_297);
  not mul_102_22_drc_bufs4303(mul_102_22_n_16 ,mul_102_22_n_15);
  not mul_102_22_drc_bufs4305(mul_102_22_n_15 ,mul_102_22_n_170);
  not mul_102_22_drc_bufs4307(mul_102_22_n_14 ,mul_102_22_n_13);
  not mul_102_22_drc_bufs4309(mul_102_22_n_13 ,mul_102_22_n_88);
  not mul_102_22_drc_bufs4311(mul_102_22_n_12 ,mul_102_22_n_11);
  not mul_102_22_drc_bufs4313(mul_102_22_n_11 ,mul_102_22_n_79);
  not mul_102_22_drc_bufs4315(mul_102_22_n_10 ,mul_102_22_n_9);
  not mul_102_22_drc_bufs4317(mul_102_22_n_9 ,mul_102_22_n_82);
  not mul_102_22_drc_bufs4319(mul_102_22_n_8 ,mul_102_22_n_7);
  not mul_102_22_drc_bufs4321(mul_102_22_n_7 ,mul_102_22_n_85);
  and mul_102_22_g2(mul_102_22_n_6 ,mul_102_22_n_982 ,mul_102_22_n_996);
  and mul_102_22_g4323(mul_102_22_n_5 ,mul_102_22_n_913 ,mul_102_22_n_966);
  xor mul_102_22_g4324(mul_102_22_n_4 ,mul_102_22_n_882 ,mul_102_22_n_963);
  xor mul_102_22_g4325(mul_102_22_n_3 ,mul_102_22_n_889 ,mul_102_22_n_960);
  xor mul_102_22_g4326(mul_102_22_n_2 ,mul_102_22_n_890 ,mul_102_22_n_930);
  xor mul_102_22_g4327(mul_102_22_n_1 ,mul_102_22_n_599 ,mul_102_22_n_847);
  xor mul_102_22_g4328(mul_102_22_n_0 ,mul_102_22_n_801 ,mul_102_22_n_307);
  xnor mul_108_22_g2868(n_254 ,mul_108_22_n_984 ,mul_108_22_n_1157);
  nor mul_108_22_g2869(mul_108_22_n_1157 ,mul_108_22_n_1026 ,mul_108_22_n_1155);
  xnor mul_108_22_g2870(mul_108_22_n_1156 ,mul_108_22_n_1154 ,mul_108_22_n_1040);
  and mul_108_22_g2871(mul_108_22_n_1155 ,mul_108_22_n_1027 ,mul_108_22_n_1154);
  or mul_108_22_g2872(mul_108_22_n_1154 ,mul_108_22_n_1050 ,mul_108_22_n_1152);
  xnor mul_108_22_g2873(mul_108_22_n_1153 ,mul_108_22_n_1151 ,mul_108_22_n_1061);
  and mul_108_22_g2874(mul_108_22_n_1152 ,mul_108_22_n_1051 ,mul_108_22_n_1151);
  or mul_108_22_g2875(mul_108_22_n_1151 ,mul_108_22_n_1079 ,mul_108_22_n_1149);
  xnor mul_108_22_g2876(mul_108_22_n_1150 ,mul_108_22_n_1148 ,mul_108_22_n_1081);
  nor mul_108_22_g2877(mul_108_22_n_1149 ,mul_108_22_n_1072 ,mul_108_22_n_1148);
  and mul_108_22_g2878(mul_108_22_n_1148 ,mul_108_22_n_1094 ,mul_108_22_n_1146);
  xnor mul_108_22_g2879(mul_108_22_n_1147 ,mul_108_22_n_1144 ,mul_108_22_n_1106);
  or mul_108_22_g2880(mul_108_22_n_1146 ,mul_108_22_n_1093 ,mul_108_22_n_1145);
  not mul_108_22_g2881(mul_108_22_n_1145 ,mul_108_22_n_1144);
  or mul_108_22_g2882(mul_108_22_n_1144 ,mul_108_22_n_1073 ,mul_108_22_n_1142);
  xnor mul_108_22_g2883(mul_108_22_n_1143 ,mul_108_22_n_1141 ,mul_108_22_n_1082);
  and mul_108_22_g2884(mul_108_22_n_1142 ,mul_108_22_n_1080 ,mul_108_22_n_1141);
  or mul_108_22_g2885(mul_108_22_n_1141 ,mul_108_22_n_1087 ,mul_108_22_n_1139);
  xnor mul_108_22_g2886(mul_108_22_n_1140 ,mul_108_22_n_1138 ,mul_108_22_n_1105);
  and mul_108_22_g2887(mul_108_22_n_1139 ,mul_108_22_n_1086 ,mul_108_22_n_1138);
  or mul_108_22_g2888(mul_108_22_n_1138 ,mul_108_22_n_1085 ,mul_108_22_n_1136);
  xnor mul_108_22_g2889(mul_108_22_n_1137 ,mul_108_22_n_1135 ,mul_108_22_n_1104);
  nor mul_108_22_g2890(mul_108_22_n_1136 ,mul_108_22_n_1135 ,mul_108_22_n_1099);
  and mul_108_22_g2891(mul_108_22_n_1135 ,mul_108_22_n_1092 ,mul_108_22_n_1133);
  xnor mul_108_22_g2892(mul_108_22_n_1134 ,mul_108_22_n_1131 ,mul_108_22_n_1103);
  or mul_108_22_g2893(mul_108_22_n_1133 ,mul_108_22_n_1090 ,mul_108_22_n_1132);
  not mul_108_22_g2894(mul_108_22_n_1132 ,mul_108_22_n_1131);
  or mul_108_22_g2895(mul_108_22_n_1131 ,mul_108_22_n_1089 ,mul_108_22_n_1129);
  xnor mul_108_22_g2896(mul_108_22_n_1130 ,mul_108_22_n_1128 ,mul_108_22_n_1102);
  and mul_108_22_g2897(mul_108_22_n_1129 ,mul_108_22_n_1088 ,mul_108_22_n_1128);
  or mul_108_22_g2898(mul_108_22_n_1128 ,mul_108_22_n_1075 ,mul_108_22_n_1126);
  xnor mul_108_22_g2899(mul_108_22_n_1127 ,mul_108_22_n_1125 ,mul_108_22_n_1084);
  and mul_108_22_g2900(mul_108_22_n_1126 ,mul_108_22_n_1074 ,mul_108_22_n_1125);
  or mul_108_22_g2901(mul_108_22_n_1125 ,mul_108_22_n_1098 ,mul_108_22_n_1123);
  xnor mul_108_22_g2902(mul_108_22_n_1124 ,mul_108_22_n_1122 ,mul_108_22_n_1101);
  and mul_108_22_g2903(mul_108_22_n_1123 ,mul_108_22_n_1097 ,mul_108_22_n_1122);
  or mul_108_22_g2904(mul_108_22_n_1122 ,mul_108_22_n_1078 ,mul_108_22_n_1120);
  xnor mul_108_22_g2905(mul_108_22_n_1121 ,mul_108_22_n_1119 ,mul_108_22_n_1083);
  and mul_108_22_g2906(mul_108_22_n_1120 ,mul_108_22_n_1077 ,mul_108_22_n_1119);
  or mul_108_22_g2907(mul_108_22_n_1119 ,mul_108_22_n_1096 ,mul_108_22_n_1117);
  xnor mul_108_22_g2908(mul_108_22_n_1118 ,mul_108_22_n_1116 ,mul_108_22_n_1100);
  and mul_108_22_g2909(mul_108_22_n_1117 ,mul_108_22_n_1095 ,mul_108_22_n_1116);
  or mul_108_22_g2910(mul_108_22_n_1116 ,mul_108_22_n_1041 ,mul_108_22_n_1114);
  xnor mul_108_22_g2911(mul_108_22_n_1115 ,mul_108_22_n_1113 ,mul_108_22_n_1060);
  and mul_108_22_g2912(mul_108_22_n_1114 ,mul_108_22_n_1042 ,mul_108_22_n_1113);
  or mul_108_22_g2913(mul_108_22_n_1113 ,mul_108_22_n_1043 ,mul_108_22_n_1111);
  xnor mul_108_22_g2914(mul_108_22_n_1112 ,mul_108_22_n_1110 ,mul_108_22_n_1059);
  and mul_108_22_g2915(mul_108_22_n_1111 ,mul_108_22_n_1044 ,mul_108_22_n_1110);
  or mul_108_22_g2916(mul_108_22_n_1110 ,mul_108_22_n_6 ,mul_108_22_n_1109);
  nor mul_108_22_g2917(mul_108_22_n_1109 ,mul_108_22_n_1016 ,mul_108_22_n_1108);
  nor mul_108_22_g2918(mul_108_22_n_1108 ,mul_108_22_n_5 ,mul_108_22_n_1107);
  nor mul_108_22_g2919(mul_108_22_n_1107 ,mul_108_22_n_1003 ,mul_108_22_n_1091);
  xnor mul_108_22_g2920(mul_108_22_n_1106 ,mul_108_22_n_1062 ,mul_108_22_n_1039);
  xnor mul_108_22_g2921(mul_108_22_n_1105 ,mul_108_22_n_1019 ,mul_108_22_n_1063);
  xnor mul_108_22_g2922(mul_108_22_n_1104 ,mul_108_22_n_1038 ,mul_108_22_n_1070);
  xnor mul_108_22_g2923(mul_108_22_n_1103 ,mul_108_22_n_1037 ,mul_108_22_n_1069);
  xnor mul_108_22_g2924(mul_108_22_n_1102 ,mul_108_22_n_1055 ,mul_108_22_n_1066);
  xnor mul_108_22_g2925(mul_108_22_n_1101 ,mul_108_22_n_1065 ,mul_108_22_n_1058);
  xnor mul_108_22_g2926(mul_108_22_n_1100 ,mul_108_22_n_1035 ,mul_108_22_n_1067);
  and mul_108_22_g2927(mul_108_22_n_1099 ,mul_108_22_n_1038 ,mul_108_22_n_1071);
  nor mul_108_22_g2928(mul_108_22_n_1098 ,mul_108_22_n_1058 ,mul_108_22_n_1065);
  or mul_108_22_g2929(mul_108_22_n_1097 ,mul_108_22_n_1057 ,mul_108_22_n_1064);
  and mul_108_22_g2930(mul_108_22_n_1096 ,mul_108_22_n_1035 ,mul_108_22_n_1067);
  or mul_108_22_g2931(mul_108_22_n_1095 ,mul_108_22_n_1035 ,mul_108_22_n_1067);
  or mul_108_22_g2932(mul_108_22_n_1094 ,mul_108_22_n_1039 ,mul_108_22_n_1062);
  and mul_108_22_g2933(mul_108_22_n_1093 ,mul_108_22_n_1039 ,mul_108_22_n_1062);
  or mul_108_22_g2934(mul_108_22_n_1092 ,mul_108_22_n_1036 ,mul_108_22_n_1068);
  nor mul_108_22_g2935(mul_108_22_n_1091 ,mul_108_22_n_1000 ,mul_108_22_n_1076);
  nor mul_108_22_g2936(mul_108_22_n_1090 ,mul_108_22_n_1037 ,mul_108_22_n_1069);
  and mul_108_22_g2937(mul_108_22_n_1089 ,mul_108_22_n_1055 ,mul_108_22_n_1066);
  or mul_108_22_g2938(mul_108_22_n_1088 ,mul_108_22_n_1055 ,mul_108_22_n_1066);
  and mul_108_22_g2939(mul_108_22_n_1087 ,mul_108_22_n_1019 ,mul_108_22_n_1063);
  or mul_108_22_g2940(mul_108_22_n_1086 ,mul_108_22_n_1019 ,mul_108_22_n_1063);
  nor mul_108_22_g2941(mul_108_22_n_1085 ,mul_108_22_n_1038 ,mul_108_22_n_1071);
  xnor mul_108_22_g2942(mul_108_22_n_1084 ,mul_108_22_n_1056 ,mul_108_22_n_1045);
  xnor mul_108_22_g2943(mul_108_22_n_1083 ,mul_108_22_n_1047 ,mul_108_22_n_1053);
  xnor mul_108_22_g2944(mul_108_22_n_1082 ,mul_108_22_n_1034 ,mul_108_22_n_1048);
  xnor mul_108_22_g2945(mul_108_22_n_1081 ,mul_108_22_n_1054 ,mul_108_22_n_1017);
  or mul_108_22_g2946(mul_108_22_n_1080 ,mul_108_22_n_1034 ,mul_108_22_n_1048);
  nor mul_108_22_g2947(mul_108_22_n_1079 ,mul_108_22_n_1054 ,mul_108_22_n_1018);
  nor mul_108_22_g2948(mul_108_22_n_1078 ,mul_108_22_n_1053 ,mul_108_22_n_1047);
  or mul_108_22_g2949(mul_108_22_n_1077 ,mul_108_22_n_1052 ,mul_108_22_n_1046);
  nor mul_108_22_g2950(mul_108_22_n_1076 ,mul_108_22_n_999 ,mul_108_22_n_1049);
  and mul_108_22_g2951(mul_108_22_n_1075 ,mul_108_22_n_1056 ,mul_108_22_n_1045);
  or mul_108_22_g2952(mul_108_22_n_1074 ,mul_108_22_n_1056 ,mul_108_22_n_1045);
  and mul_108_22_g2953(mul_108_22_n_1073 ,mul_108_22_n_1034 ,mul_108_22_n_1048);
  and mul_108_22_g2954(mul_108_22_n_1072 ,mul_108_22_n_1054 ,mul_108_22_n_1018);
  not mul_108_22_g2955(mul_108_22_n_1071 ,mul_108_22_n_1070);
  not mul_108_22_g2956(mul_108_22_n_1069 ,mul_108_22_n_1068);
  not mul_108_22_g2957(mul_108_22_n_1065 ,mul_108_22_n_1064);
  xnor mul_108_22_g2958(mul_108_22_n_1061 ,mul_108_22_n_1023 ,mul_108_22_n_1033);
  xnor mul_108_22_g2959(mul_108_22_n_1060 ,mul_108_22_n_1009 ,mul_108_22_n_1021);
  xnor mul_108_22_g2960(mul_108_22_n_1059 ,mul_108_22_n_1010 ,mul_108_22_n_1020);
  xnor mul_108_22_g2961(mul_108_22_n_1070 ,mul_108_22_n_941 ,mul_108_22_n_1011);
  xnor mul_108_22_g2962(mul_108_22_n_1068 ,mul_108_22_n_925 ,mul_108_22_n_4);
  xnor mul_108_22_g2963(mul_108_22_n_1067 ,mul_108_22_n_945 ,mul_108_22_n_1014);
  xnor mul_108_22_g2964(mul_108_22_n_1066 ,mul_108_22_n_942 ,mul_108_22_n_3);
  xnor mul_108_22_g2965(mul_108_22_n_1064 ,mul_108_22_n_912 ,mul_108_22_n_1012);
  xnor mul_108_22_g2966(mul_108_22_n_1063 ,mul_108_22_n_939 ,mul_108_22_n_1013);
  xnor mul_108_22_g2967(mul_108_22_n_1062 ,mul_108_22_n_944 ,mul_108_22_n_1015);
  not mul_108_22_g2968(mul_108_22_n_1057 ,mul_108_22_n_1058);
  not mul_108_22_g2969(mul_108_22_n_1052 ,mul_108_22_n_1053);
  or mul_108_22_g2970(mul_108_22_n_1051 ,mul_108_22_n_1032 ,mul_108_22_n_1022);
  nor mul_108_22_g2971(mul_108_22_n_1050 ,mul_108_22_n_1033 ,mul_108_22_n_1023);
  nor mul_108_22_g2972(mul_108_22_n_1049 ,mul_108_22_n_921 ,mul_108_22_n_1031);
  and mul_108_22_g2973(mul_108_22_n_1058 ,mul_108_22_n_993 ,mul_108_22_n_1024);
  or mul_108_22_g2974(mul_108_22_n_1056 ,mul_108_22_n_1005 ,mul_108_22_n_1030);
  or mul_108_22_g2975(mul_108_22_n_1055 ,mul_108_22_n_997 ,mul_108_22_n_1025);
  and mul_108_22_g2976(mul_108_22_n_1054 ,mul_108_22_n_1007 ,mul_108_22_n_1029);
  and mul_108_22_g2977(mul_108_22_n_1053 ,mul_108_22_n_991 ,mul_108_22_n_1028);
  not mul_108_22_g2978(mul_108_22_n_1047 ,mul_108_22_n_1046);
  or mul_108_22_g2979(mul_108_22_n_1044 ,mul_108_22_n_1010 ,mul_108_22_n_1020);
  and mul_108_22_g2980(mul_108_22_n_1043 ,mul_108_22_n_1010 ,mul_108_22_n_1020);
  or mul_108_22_g2981(mul_108_22_n_1042 ,mul_108_22_n_1009 ,mul_108_22_n_1021);
  and mul_108_22_g2982(mul_108_22_n_1041 ,mul_108_22_n_1009 ,mul_108_22_n_1021);
  xnor mul_108_22_g2983(mul_108_22_n_1040 ,mul_108_22_n_927 ,mul_108_22_n_995);
  xnor mul_108_22_g2984(mul_108_22_n_1048 ,mul_108_22_n_940 ,mul_108_22_n_2);
  xnor mul_108_22_g2985(mul_108_22_n_1046 ,mul_108_22_n_956 ,mul_108_22_n_983);
  xnor mul_108_22_g2986(mul_108_22_n_1045 ,mul_108_22_n_952 ,mul_108_22_n_985);
  not mul_108_22_g2987(mul_108_22_n_1037 ,mul_108_22_n_1036);
  not mul_108_22_g2988(mul_108_22_n_1033 ,mul_108_22_n_1032);
  nor mul_108_22_g2989(mul_108_22_n_1031 ,mul_108_22_n_920 ,mul_108_22_n_1002);
  and mul_108_22_g2990(mul_108_22_n_1030 ,mul_108_22_n_912 ,mul_108_22_n_987);
  or mul_108_22_g2991(mul_108_22_n_1029 ,mul_108_22_n_944 ,mul_108_22_n_1004);
  or mul_108_22_g2992(mul_108_22_n_1028 ,mul_108_22_n_945 ,mul_108_22_n_990);
  or mul_108_22_g2993(mul_108_22_n_1027 ,mul_108_22_n_927 ,mul_108_22_n_995);
  and mul_108_22_g2994(mul_108_22_n_1026 ,mul_108_22_n_927 ,mul_108_22_n_995);
  nor mul_108_22_g2995(mul_108_22_n_1025 ,mul_108_22_n_943 ,mul_108_22_n_1001);
  or mul_108_22_g2996(mul_108_22_n_1024 ,mul_108_22_n_929 ,mul_108_22_n_992);
  and mul_108_22_g2997(mul_108_22_n_1039 ,mul_108_22_n_973 ,mul_108_22_n_994);
  and mul_108_22_g2998(mul_108_22_n_1038 ,mul_108_22_n_969 ,mul_108_22_n_989);
  and mul_108_22_g2999(mul_108_22_n_1036 ,mul_108_22_n_971 ,mul_108_22_n_998);
  or mul_108_22_g3000(mul_108_22_n_1035 ,mul_108_22_n_976 ,mul_108_22_n_986);
  or mul_108_22_g3001(mul_108_22_n_1034 ,mul_108_22_n_978 ,mul_108_22_n_1006);
  or mul_108_22_g3002(mul_108_22_n_1032 ,mul_108_22_n_937 ,mul_108_22_n_1008);
  not mul_108_22_g3003(mul_108_22_n_1022 ,mul_108_22_n_1023);
  not mul_108_22_g3004(mul_108_22_n_1018 ,mul_108_22_n_1017);
  nor mul_108_22_g3006(mul_108_22_n_1016 ,mul_108_22_n_982 ,mul_108_22_n_996);
  xnor mul_108_22_g3007(mul_108_22_n_1015 ,mul_108_22_n_959 ,mul_108_22_n_862);
  xnor mul_108_22_g3008(mul_108_22_n_1014 ,mul_108_22_n_794 ,mul_108_22_n_954);
  xnor mul_108_22_g3009(mul_108_22_n_1013 ,mul_108_22_n_878 ,mul_108_22_n_962);
  xnor mul_108_22_g3010(mul_108_22_n_1012 ,mul_108_22_n_958 ,mul_108_22_n_885);
  xnor mul_108_22_g3011(mul_108_22_n_1011 ,mul_108_22_n_906 ,mul_108_22_n_961);
  xnor mul_108_22_g3014(mul_108_22_n_1023 ,mul_108_22_n_842 ,mul_108_22_n_947);
  xnor mul_108_22_g3015(mul_108_22_n_1021 ,mul_108_22_n_926 ,mul_108_22_n_946);
  xnor mul_108_22_g3016(mul_108_22_n_1020 ,mul_108_22_n_928 ,mul_108_22_n_948);
  or mul_108_22_g3017(mul_108_22_n_1019 ,mul_108_22_n_951 ,mul_108_22_n_988);
  xnor mul_108_22_g3018(mul_108_22_n_1017 ,mul_108_22_n_981 ,mul_108_22_n_949);
  and mul_108_22_g3020(mul_108_22_n_1008 ,mul_108_22_n_981 ,mul_108_22_n_931);
  or mul_108_22_g3021(mul_108_22_n_1007 ,mul_108_22_n_862 ,mul_108_22_n_959);
  and mul_108_22_g3022(mul_108_22_n_1006 ,mul_108_22_n_962 ,mul_108_22_n_977);
  nor mul_108_22_g3023(mul_108_22_n_1005 ,mul_108_22_n_182 ,mul_108_22_n_958);
  and mul_108_22_g3024(mul_108_22_n_1004 ,mul_108_22_n_862 ,mul_108_22_n_959);
  nor mul_108_22_g3025(mul_108_22_n_1003 ,mul_108_22_n_913 ,mul_108_22_n_966);
  nor mul_108_22_g3026(mul_108_22_n_1002 ,mul_108_22_n_935 ,mul_108_22_n_979);
  and mul_108_22_g3027(mul_108_22_n_1001 ,mul_108_22_n_886 ,mul_108_22_n_952);
  nor mul_108_22_g3028(mul_108_22_n_1000 ,mul_108_22_n_848 ,mul_108_22_n_965);
  nor mul_108_22_g3029(mul_108_22_n_999 ,mul_108_22_n_849 ,mul_108_22_n_964);
  or mul_108_22_g3030(mul_108_22_n_998 ,mul_108_22_n_970 ,mul_108_22_n_960);
  nor mul_108_22_g3031(mul_108_22_n_997 ,mul_108_22_n_886 ,mul_108_22_n_952);
  or mul_108_22_g3032(mul_108_22_n_1010 ,mul_108_22_n_923 ,mul_108_22_n_972);
  or mul_108_22_g3033(mul_108_22_n_1009 ,mul_108_22_n_918 ,mul_108_22_n_974);
  or mul_108_22_g3035(mul_108_22_n_994 ,mul_108_22_n_930 ,mul_108_22_n_980);
  or mul_108_22_g3036(mul_108_22_n_993 ,mul_108_22_n_884 ,mul_108_22_n_955);
  nor mul_108_22_g3037(mul_108_22_n_992 ,mul_108_22_n_883 ,mul_108_22_n_956);
  or mul_108_22_g3038(mul_108_22_n_991 ,mul_108_22_n_794 ,mul_108_22_n_953);
  nor mul_108_22_g3039(mul_108_22_n_990 ,mul_108_22_n_793 ,mul_108_22_n_954);
  or mul_108_22_g3040(mul_108_22_n_989 ,mul_108_22_n_968 ,mul_108_22_n_963);
  nor mul_108_22_g3041(mul_108_22_n_988 ,mul_108_22_n_950 ,mul_108_22_n_961);
  or mul_108_22_g3042(mul_108_22_n_987 ,mul_108_22_n_308 ,mul_108_22_n_957);
  nor mul_108_22_g3043(mul_108_22_n_986 ,mul_108_22_n_840 ,mul_108_22_n_975);
  xor mul_108_22_g3044(mul_108_22_n_985 ,mul_108_22_n_943 ,mul_108_22_n_886);
  xnor mul_108_22_g3046(mul_108_22_n_984 ,mul_108_22_n_0 ,mul_108_22_n_916);
  xnor mul_108_22_g3047(mul_108_22_n_996 ,mul_108_22_n_876 ,mul_108_22_n_1);
  xnor mul_108_22_g3048(mul_108_22_n_983 ,mul_108_22_n_929 ,mul_108_22_n_884);
  or mul_108_22_g3049(mul_108_22_n_995 ,mul_108_22_n_933 ,mul_108_22_n_967);
  and mul_108_22_g3051(mul_108_22_n_980 ,mul_108_22_n_890 ,mul_108_22_n_940);
  and mul_108_22_g3052(mul_108_22_n_979 ,mul_108_22_n_802 ,mul_108_22_n_934);
  nor mul_108_22_g3053(mul_108_22_n_978 ,mul_108_22_n_878 ,mul_108_22_n_939);
  or mul_108_22_g3054(mul_108_22_n_977 ,mul_108_22_n_877 ,mul_108_22_n_938);
  nor mul_108_22_g3055(mul_108_22_n_976 ,mul_108_22_n_905 ,mul_108_22_n_926);
  and mul_108_22_g3056(mul_108_22_n_975 ,mul_108_22_n_905 ,mul_108_22_n_926);
  and mul_108_22_g3057(mul_108_22_n_974 ,mul_108_22_n_928 ,mul_108_22_n_917);
  or mul_108_22_g3058(mul_108_22_n_973 ,mul_108_22_n_890 ,mul_108_22_n_940);
  nor mul_108_22_g3059(mul_108_22_n_972 ,mul_108_22_n_847 ,mul_108_22_n_919);
  or mul_108_22_g3060(mul_108_22_n_971 ,mul_108_22_n_889 ,mul_108_22_n_942);
  and mul_108_22_g3061(mul_108_22_n_970 ,mul_108_22_n_889 ,mul_108_22_n_942);
  or mul_108_22_g3062(mul_108_22_n_969 ,mul_108_22_n_882 ,mul_108_22_n_924);
  nor mul_108_22_g3063(mul_108_22_n_968 ,mul_108_22_n_881 ,mul_108_22_n_925);
  and mul_108_22_g3064(mul_108_22_n_967 ,mul_108_22_n_842 ,mul_108_22_n_936);
  or mul_108_22_g3065(mul_108_22_n_982 ,mul_108_22_n_705 ,mul_108_22_n_922);
  or mul_108_22_g3066(mul_108_22_n_981 ,mul_108_22_n_746 ,mul_108_22_n_932);
  not mul_108_22_g3068(mul_108_22_n_965 ,mul_108_22_n_964);
  not mul_108_22_g3071(mul_108_22_n_958 ,mul_108_22_n_957);
  not mul_108_22_g3072(mul_108_22_n_956 ,mul_108_22_n_955);
  not mul_108_22_g3073(mul_108_22_n_953 ,mul_108_22_n_954);
  nor mul_108_22_g3074(mul_108_22_n_951 ,mul_108_22_n_907 ,mul_108_22_n_941);
  and mul_108_22_g3075(mul_108_22_n_950 ,mul_108_22_n_907 ,mul_108_22_n_941);
  xnor mul_108_22_g3076(mul_108_22_n_966 ,mul_108_22_n_910 ,mul_108_22_n_780);
  xnor mul_108_22_g3077(mul_108_22_n_964 ,mul_108_22_n_602 ,mul_108_22_n_875);
  xnor mul_108_22_g3078(mul_108_22_n_949 ,mul_108_22_n_888 ,mul_108_22_n_839);
  xnor mul_108_22_g3079(mul_108_22_n_948 ,mul_108_22_n_880 ,mul_108_22_n_909);
  xnor mul_108_22_g3080(mul_108_22_n_947 ,mul_108_22_n_904 ,mul_108_22_n_649);
  xor mul_108_22_g3081(mul_108_22_n_946 ,mul_108_22_n_905 ,mul_108_22_n_840);
  xnor mul_108_22_g3082(mul_108_22_n_963 ,mul_108_22_n_841 ,mul_108_22_n_868);
  xnor mul_108_22_g3083(mul_108_22_n_962 ,mul_108_22_n_867 ,mul_108_22_n_870);
  xnor mul_108_22_g3084(mul_108_22_n_961 ,mul_108_22_n_866 ,mul_108_22_n_869);
  xnor mul_108_22_g3085(mul_108_22_n_960 ,mul_108_22_n_845 ,mul_108_22_n_874);
  xnor mul_108_22_g3086(mul_108_22_n_959 ,mul_108_22_n_911 ,mul_108_22_n_787);
  xnor mul_108_22_g3087(mul_108_22_n_957 ,mul_108_22_n_865 ,mul_108_22_n_872);
  xnor mul_108_22_g3088(mul_108_22_n_955 ,mul_108_22_n_762 ,mul_108_22_n_871);
  xnor mul_108_22_g3089(mul_108_22_n_954 ,mul_108_22_n_843 ,mul_108_22_n_893);
  xnor mul_108_22_g3090(mul_108_22_n_952 ,mul_108_22_n_864 ,mul_108_22_n_873);
  not mul_108_22_g3091(mul_108_22_n_939 ,mul_108_22_n_938);
  nor mul_108_22_g3092(mul_108_22_n_937 ,mul_108_22_n_839 ,mul_108_22_n_888);
  or mul_108_22_g3093(mul_108_22_n_936 ,mul_108_22_n_204 ,mul_108_22_n_904);
  nor mul_108_22_g3094(mul_108_22_n_935 ,mul_108_22_n_643 ,mul_108_22_n_914);
  or mul_108_22_g3095(mul_108_22_n_934 ,mul_108_22_n_644 ,mul_108_22_n_915);
  and mul_108_22_g3096(mul_108_22_n_933 ,mul_108_22_n_203 ,mul_108_22_n_904);
  and mul_108_22_g3097(mul_108_22_n_932 ,mul_108_22_n_755 ,mul_108_22_n_911);
  or mul_108_22_g3098(mul_108_22_n_931 ,mul_108_22_n_838 ,mul_108_22_n_887);
  and mul_108_22_g3099(mul_108_22_n_945 ,mul_108_22_n_754 ,mul_108_22_n_899);
  and mul_108_22_g3100(mul_108_22_n_944 ,mul_108_22_n_804 ,mul_108_22_n_897);
  and mul_108_22_g3101(mul_108_22_n_943 ,mul_108_22_n_857 ,mul_108_22_n_901);
  and mul_108_22_g3102(mul_108_22_n_942 ,mul_108_22_n_861 ,mul_108_22_n_902);
  and mul_108_22_g3103(mul_108_22_n_941 ,mul_108_22_n_832 ,mul_108_22_n_898);
  and mul_108_22_g3104(mul_108_22_n_940 ,mul_108_22_n_855 ,mul_108_22_n_903);
  or mul_108_22_g3105(mul_108_22_n_938 ,mul_108_22_n_854 ,mul_108_22_n_900);
  not mul_108_22_g3107(mul_108_22_n_924 ,mul_108_22_n_925);
  nor mul_108_22_g3108(mul_108_22_n_923 ,mul_108_22_n_599 ,mul_108_22_n_876);
  and mul_108_22_g3109(mul_108_22_n_922 ,mul_108_22_n_704 ,mul_108_22_n_910);
  nor mul_108_22_g3110(mul_108_22_n_921 ,mul_108_22_n_769 ,mul_108_22_n_891);
  nor mul_108_22_g3111(mul_108_22_n_920 ,mul_108_22_n_768 ,mul_108_22_n_892);
  and mul_108_22_g3112(mul_108_22_n_919 ,mul_108_22_n_599 ,mul_108_22_n_876);
  nor mul_108_22_g3113(mul_108_22_n_918 ,mul_108_22_n_909 ,mul_108_22_n_880);
  or mul_108_22_g3114(mul_108_22_n_917 ,mul_108_22_n_908 ,mul_108_22_n_879);
  or mul_108_22_g3116(mul_108_22_n_916 ,mul_108_22_n_719 ,mul_108_22_n_894);
  xnor mul_108_22_g3117(mul_108_22_n_930 ,mul_108_22_n_844 ,mul_108_22_n_830);
  and mul_108_22_g3118(mul_108_22_n_929 ,mul_108_22_n_851 ,mul_108_22_n_895);
  xnor mul_108_22_g3119(mul_108_22_n_928 ,mul_108_22_n_606 ,mul_108_22_n_831);
  xnor mul_108_22_g3120(mul_108_22_n_927 ,mul_108_22_n_863 ,mul_108_22_n_782);
  xnor mul_108_22_g3121(mul_108_22_n_926 ,mul_108_22_n_846 ,mul_108_22_n_783);
  or mul_108_22_g3122(mul_108_22_n_925 ,mul_108_22_n_835 ,mul_108_22_n_896);
  not mul_108_22_g3123(mul_108_22_n_915 ,mul_108_22_n_914);
  not mul_108_22_g3125(mul_108_22_n_908 ,mul_108_22_n_909);
  not mul_108_22_g3126(mul_108_22_n_907 ,mul_108_22_n_906);
  or mul_108_22_g3127(mul_108_22_n_903 ,mul_108_22_n_858 ,mul_108_22_n_867);
  or mul_108_22_g3128(mul_108_22_n_902 ,mul_108_22_n_860 ,mul_108_22_n_864);
  or mul_108_22_g3129(mul_108_22_n_901 ,mul_108_22_n_856 ,mul_108_22_n_865);
  nor mul_108_22_g3130(mul_108_22_n_900 ,mul_108_22_n_852 ,mul_108_22_n_866);
  or mul_108_22_g3131(mul_108_22_n_899 ,mul_108_22_n_726 ,mul_108_22_n_846);
  or mul_108_22_g3132(mul_108_22_n_898 ,mul_108_22_n_837 ,mul_108_22_n_841);
  or mul_108_22_g3133(mul_108_22_n_897 ,mul_108_22_n_803 ,mul_108_22_n_844);
  nor mul_108_22_g3134(mul_108_22_n_896 ,mul_108_22_n_834 ,mul_108_22_n_845);
  or mul_108_22_g3135(mul_108_22_n_895 ,mul_108_22_n_843 ,mul_108_22_n_850);
  and mul_108_22_g3136(mul_108_22_n_894 ,mul_108_22_n_720 ,mul_108_22_n_863);
  and mul_108_22_g3137(mul_108_22_n_914 ,mul_108_22_n_753 ,mul_108_22_n_859);
  xnor mul_108_22_g3138(mul_108_22_n_893 ,mul_108_22_n_663 ,mul_108_22_n_792);
  xnor mul_108_22_g3139(mul_108_22_n_913 ,mul_108_22_n_731 ,mul_108_22_n_774);
  or mul_108_22_g3140(mul_108_22_n_912 ,mul_108_22_n_816 ,mul_108_22_n_853);
  xnor mul_108_22_g3141(mul_108_22_n_911 ,mul_108_22_n_692 ,mul_108_22_n_800);
  or mul_108_22_g3142(mul_108_22_n_910 ,mul_108_22_n_703 ,mul_108_22_n_833);
  and mul_108_22_g3143(mul_108_22_n_909 ,mul_108_22_n_713 ,mul_108_22_n_836);
  xnor mul_108_22_g3144(mul_108_22_n_906 ,mul_108_22_n_672 ,mul_108_22_n_785);
  xnor mul_108_22_g3145(mul_108_22_n_905 ,mul_108_22_n_661 ,mul_108_22_n_779);
  xnor mul_108_22_g3146(mul_108_22_n_904 ,mul_108_22_n_687 ,mul_108_22_n_777);
  not mul_108_22_g3147(mul_108_22_n_892 ,mul_108_22_n_891);
  not mul_108_22_g3148(mul_108_22_n_888 ,mul_108_22_n_887);
  not mul_108_22_g3150(mul_108_22_n_883 ,mul_108_22_n_884);
  not mul_108_22_g3151(mul_108_22_n_881 ,mul_108_22_n_882);
  not mul_108_22_g3152(mul_108_22_n_879 ,mul_108_22_n_880);
  not mul_108_22_g3153(mul_108_22_n_877 ,mul_108_22_n_878);
  xnor mul_108_22_g3154(mul_108_22_n_875 ,mul_108_22_n_618 ,mul_108_22_n_797);
  xnor mul_108_22_g3155(mul_108_22_n_874 ,mul_108_22_n_758 ,mul_108_22_n_796);
  xnor mul_108_22_g3156(mul_108_22_n_873 ,mul_108_22_n_764 ,mul_108_22_n_829);
  xnor mul_108_22_g3157(mul_108_22_n_872 ,mul_108_22_n_760 ,mul_108_22_n_827);
  xnor mul_108_22_g3158(mul_108_22_n_871 ,mul_108_22_n_767 ,mul_108_22_n_799);
  xnor mul_108_22_g3159(mul_108_22_n_870 ,mul_108_22_n_757 ,mul_108_22_n_825);
  xnor mul_108_22_g3160(mul_108_22_n_869 ,mul_108_22_n_765 ,mul_108_22_n_795);
  xnor mul_108_22_g3161(mul_108_22_n_868 ,mul_108_22_n_730 ,mul_108_22_n_790);
  xnor mul_108_22_g3162(mul_108_22_n_891 ,mul_108_22_n_641 ,mul_108_22_n_775);
  xnor mul_108_22_g3164(mul_108_22_n_890 ,mul_108_22_n_697 ,mul_108_22_n_781);
  xnor mul_108_22_g3165(mul_108_22_n_889 ,mul_108_22_n_608 ,mul_108_22_n_778);
  xnor mul_108_22_g3166(mul_108_22_n_887 ,mul_108_22_n_786 ,mul_108_22_n_204);
  xnor mul_108_22_g3167(mul_108_22_n_886 ,mul_108_22_n_621 ,mul_108_22_n_773);
  xnor mul_108_22_g3168(mul_108_22_n_885 ,mul_108_22_n_632 ,mul_108_22_n_771);
  xnor mul_108_22_g3169(mul_108_22_n_884 ,mul_108_22_n_627 ,mul_108_22_n_770);
  xnor mul_108_22_g3170(mul_108_22_n_882 ,mul_108_22_n_664 ,mul_108_22_n_788);
  xnor mul_108_22_g3171(mul_108_22_n_880 ,mul_108_22_n_631 ,mul_108_22_n_776);
  xnor mul_108_22_g3172(mul_108_22_n_878 ,mul_108_22_n_633 ,mul_108_22_n_772);
  xnor mul_108_22_g3173(mul_108_22_n_876 ,mul_108_22_n_798 ,mul_108_22_n_784);
  or mul_108_22_g3174(mul_108_22_n_861 ,mul_108_22_n_763 ,mul_108_22_n_828);
  nor mul_108_22_g3175(mul_108_22_n_860 ,mul_108_22_n_764 ,mul_108_22_n_829);
  or mul_108_22_g3176(mul_108_22_n_859 ,mul_108_22_n_821 ,mul_108_22_n_751);
  nor mul_108_22_g3177(mul_108_22_n_858 ,mul_108_22_n_757 ,mul_108_22_n_824);
  or mul_108_22_g3178(mul_108_22_n_857 ,mul_108_22_n_760 ,mul_108_22_n_826);
  nor mul_108_22_g3179(mul_108_22_n_856 ,mul_108_22_n_759 ,mul_108_22_n_827);
  or mul_108_22_g3180(mul_108_22_n_855 ,mul_108_22_n_756 ,mul_108_22_n_825);
  and mul_108_22_g3181(mul_108_22_n_854 ,mul_108_22_n_765 ,mul_108_22_n_795);
  and mul_108_22_g3182(mul_108_22_n_853 ,mul_108_22_n_799 ,mul_108_22_n_815);
  nor mul_108_22_g3183(mul_108_22_n_852 ,mul_108_22_n_765 ,mul_108_22_n_795);
  or mul_108_22_g3184(mul_108_22_n_851 ,mul_108_22_n_663 ,mul_108_22_n_791);
  nor mul_108_22_g3185(mul_108_22_n_850 ,mul_108_22_n_662 ,mul_108_22_n_792);
  and mul_108_22_g3186(mul_108_22_n_867 ,mul_108_22_n_715 ,mul_108_22_n_820);
  and mul_108_22_g3187(mul_108_22_n_866 ,mul_108_22_n_736 ,mul_108_22_n_814);
  and mul_108_22_g3188(mul_108_22_n_865 ,mul_108_22_n_743 ,mul_108_22_n_817);
  and mul_108_22_g3189(mul_108_22_n_864 ,mul_108_22_n_752 ,mul_108_22_n_819);
  or mul_108_22_g3190(mul_108_22_n_863 ,mul_108_22_n_741 ,mul_108_22_n_818);
  and mul_108_22_g3191(mul_108_22_n_862 ,mul_108_22_n_737 ,mul_108_22_n_813);
  not mul_108_22_g3192(mul_108_22_n_849 ,mul_108_22_n_848);
  not mul_108_22_g3193(mul_108_22_n_838 ,mul_108_22_n_839);
  nor mul_108_22_g3194(mul_108_22_n_837 ,mul_108_22_n_730 ,mul_108_22_n_790);
  or mul_108_22_g3195(mul_108_22_n_836 ,mul_108_22_n_711 ,mul_108_22_n_798);
  and mul_108_22_g3196(mul_108_22_n_835 ,mul_108_22_n_758 ,mul_108_22_n_796);
  nor mul_108_22_g3197(mul_108_22_n_834 ,mul_108_22_n_758 ,mul_108_22_n_796);
  and mul_108_22_g3198(mul_108_22_n_833 ,mul_108_22_n_750 ,mul_108_22_n_797);
  or mul_108_22_g3199(mul_108_22_n_832 ,mul_108_22_n_729 ,mul_108_22_n_789);
  and mul_108_22_g3200(mul_108_22_n_848 ,mul_108_22_n_747 ,mul_108_22_n_822);
  xnor mul_108_22_g3201(mul_108_22_n_831 ,mul_108_22_n_598 ,mul_108_22_n_733);
  xnor mul_108_22_g3202(mul_108_22_n_830 ,mul_108_22_n_728 ,mul_108_22_n_648);
  and mul_108_22_g3203(mul_108_22_n_847 ,mul_108_22_n_709 ,mul_108_22_n_809);
  and mul_108_22_g3204(mul_108_22_n_846 ,mul_108_22_n_735 ,mul_108_22_n_812);
  and mul_108_22_g3205(mul_108_22_n_845 ,mul_108_22_n_710 ,mul_108_22_n_808);
  and mul_108_22_g3206(mul_108_22_n_844 ,mul_108_22_n_745 ,mul_108_22_n_807);
  and mul_108_22_g3207(mul_108_22_n_843 ,mul_108_22_n_738 ,mul_108_22_n_806);
  or mul_108_22_g3208(mul_108_22_n_842 ,mul_108_22_n_725 ,mul_108_22_n_805);
  and mul_108_22_g3209(mul_108_22_n_841 ,mul_108_22_n_722 ,mul_108_22_n_811);
  and mul_108_22_g3210(mul_108_22_n_840 ,mul_108_22_n_721 ,mul_108_22_n_810);
  and mul_108_22_g3211(mul_108_22_n_839 ,mul_108_22_n_706 ,mul_108_22_n_823);
  not mul_108_22_g3212(mul_108_22_n_828 ,mul_108_22_n_829);
  not mul_108_22_g3213(mul_108_22_n_826 ,mul_108_22_n_827);
  not mul_108_22_g3214(mul_108_22_n_824 ,mul_108_22_n_825);
  or mul_108_22_g3215(mul_108_22_n_823 ,mul_108_22_n_692 ,mul_108_22_n_749);
  or mul_108_22_g3216(mul_108_22_n_822 ,mul_108_22_n_641 ,mul_108_22_n_716);
  or mul_108_22_g3217(mul_108_22_n_821 ,mul_108_22_n_327 ,mul_108_22_n_727);
  or mul_108_22_g3218(mul_108_22_n_820 ,mul_108_22_n_630 ,mul_108_22_n_744);
  or mul_108_22_g3219(mul_108_22_n_819 ,mul_108_22_n_632 ,mul_108_22_n_718);
  and mul_108_22_g3220(mul_108_22_n_818 ,mul_108_22_n_687 ,mul_108_22_n_748);
  or mul_108_22_g3221(mul_108_22_n_817 ,mul_108_22_n_627 ,mul_108_22_n_742);
  nor mul_108_22_g3222(mul_108_22_n_816 ,mul_108_22_n_767 ,mul_108_22_n_761);
  or mul_108_22_g3223(mul_108_22_n_815 ,mul_108_22_n_766 ,mul_108_22_n_762);
  or mul_108_22_g3224(mul_108_22_n_814 ,mul_108_22_n_624 ,mul_108_22_n_739);
  or mul_108_22_g3225(mul_108_22_n_813 ,mul_108_22_n_697 ,mul_108_22_n_723);
  or mul_108_22_g3226(mul_108_22_n_812 ,mul_108_22_n_631 ,mul_108_22_n_724);
  or mul_108_22_g3227(mul_108_22_n_811 ,mul_108_22_n_622 ,mul_108_22_n_714);
  or mul_108_22_g3228(mul_108_22_n_810 ,mul_108_22_n_734 ,mul_108_22_n_717);
  or mul_108_22_g3229(mul_108_22_n_809 ,mul_108_22_n_708 ,mul_108_22_n_732);
  or mul_108_22_g3230(mul_108_22_n_808 ,mul_108_22_n_621 ,mul_108_22_n_707);
  or mul_108_22_g3231(mul_108_22_n_807 ,mul_108_22_n_633 ,mul_108_22_n_702);
  or mul_108_22_g3232(mul_108_22_n_806 ,mul_108_22_n_623 ,mul_108_22_n_740);
  nor mul_108_22_g3233(mul_108_22_n_805 ,mul_108_22_n_203 ,mul_108_22_n_712);
  or mul_108_22_g3234(mul_108_22_n_804 ,mul_108_22_n_156 ,mul_108_22_n_728);
  and mul_108_22_g3235(mul_108_22_n_803 ,mul_108_22_n_157 ,mul_108_22_n_728);
  xnor mul_108_22_g3236(mul_108_22_n_802 ,mul_108_22_n_698 ,mul_108_22_n_547);
  xnor mul_108_22_g3237(mul_108_22_n_801 ,mul_108_22_n_647 ,mul_108_22_n_646);
  xnor mul_108_22_g3238(mul_108_22_n_800 ,mul_108_22_n_604 ,mul_108_22_n_656);
  xnor mul_108_22_g3239(mul_108_22_n_829 ,mul_108_22_n_628 ,mul_108_22_n_636);
  xnor mul_108_22_g3240(mul_108_22_n_827 ,mul_108_22_n_679 ,mul_108_22_n_696);
  xnor mul_108_22_g3241(mul_108_22_n_825 ,mul_108_22_n_645 ,mul_108_22_n_700);
  not mul_108_22_g3242(mul_108_22_n_793 ,mul_108_22_n_794);
  not mul_108_22_g3243(mul_108_22_n_791 ,mul_108_22_n_792);
  not mul_108_22_g3244(mul_108_22_n_789 ,mul_108_22_n_790);
  xnor mul_108_22_g3245(mul_108_22_n_788 ,mul_108_22_n_667 ,mul_108_22_n_624);
  xnor mul_108_22_g3246(mul_108_22_n_787 ,mul_108_22_n_677 ,mul_108_22_n_157);
  xnor mul_108_22_g3247(mul_108_22_n_786 ,mul_108_22_n_670 ,mul_108_22_n_611);
  xor mul_108_22_g3248(mul_108_22_n_785 ,mul_108_22_n_666 ,mul_108_22_n_630);
  xnor mul_108_22_g3249(mul_108_22_n_784 ,mul_108_22_n_609 ,mul_108_22_n_669);
  xnor mul_108_22_g3250(mul_108_22_n_783 ,mul_108_22_n_674 ,mul_108_22_n_654);
  xnor mul_108_22_g3251(mul_108_22_n_782 ,mul_108_22_n_614 ,mul_108_22_n_650);
  xnor mul_108_22_g3252(mul_108_22_n_781 ,mul_108_22_n_657 ,mul_108_22_n_612);
  xnor mul_108_22_g3253(mul_108_22_n_780 ,mul_108_22_n_594 ,mul_108_22_n_596);
  xor mul_108_22_g3254(mul_108_22_n_779 ,mul_108_22_n_659 ,mul_108_22_n_623);
  xnor mul_108_22_g3255(mul_108_22_n_778 ,mul_108_22_n_600 ,mul_108_22_n_622);
  xnor mul_108_22_g3256(mul_108_22_n_777 ,mul_108_22_n_616 ,mul_108_22_n_653);
  xnor mul_108_22_g3257(mul_108_22_n_776 ,mul_108_22_n_449 ,mul_108_22_n_673);
  xnor mul_108_22_g3258(mul_108_22_n_775 ,mul_108_22_n_451 ,mul_108_22_n_651);
  xnor mul_108_22_g3259(mul_108_22_n_774 ,mul_108_22_n_450 ,mul_108_22_n_605);
  xnor mul_108_22_g3260(mul_108_22_n_773 ,mul_108_22_n_592 ,mul_108_22_n_597);
  xnor mul_108_22_g3261(mul_108_22_n_772 ,mul_108_22_n_607 ,mul_108_22_n_665);
  xnor mul_108_22_g3262(mul_108_22_n_771 ,mul_108_22_n_610 ,mul_108_22_n_668);
  xnor mul_108_22_g3263(mul_108_22_n_770 ,mul_108_22_n_678 ,mul_108_22_n_675);
  xnor mul_108_22_g3264(mul_108_22_n_799 ,mul_108_22_n_684 ,mul_108_22_n_682);
  xnor mul_108_22_g3265(mul_108_22_n_798 ,mul_108_22_n_639 ,mul_108_22_n_544);
  xnor mul_108_22_g3266(mul_108_22_n_797 ,mul_108_22_n_546 ,mul_108_22_n_634);
  xnor mul_108_22_g3267(mul_108_22_n_796 ,mul_108_22_n_619 ,mul_108_22_n_629);
  xnor mul_108_22_g3268(mul_108_22_n_795 ,mul_108_22_n_694 ,mul_108_22_n_693);
  xnor mul_108_22_g3269(mul_108_22_n_794 ,mul_108_22_n_690 ,mul_108_22_n_625);
  xnor mul_108_22_g3270(mul_108_22_n_792 ,mul_108_22_n_681 ,mul_108_22_n_685);
  xnor mul_108_22_g3271(mul_108_22_n_790 ,mul_108_22_n_638 ,mul_108_22_n_688);
  not mul_108_22_g3272(mul_108_22_n_769 ,mul_108_22_n_768);
  not mul_108_22_g3273(mul_108_22_n_767 ,mul_108_22_n_766);
  not mul_108_22_g3274(mul_108_22_n_764 ,mul_108_22_n_763);
  not mul_108_22_g3275(mul_108_22_n_761 ,mul_108_22_n_762);
  not mul_108_22_g3276(mul_108_22_n_760 ,mul_108_22_n_759);
  not mul_108_22_g3277(mul_108_22_n_757 ,mul_108_22_n_756);
  or mul_108_22_g3278(mul_108_22_n_755 ,mul_108_22_n_156 ,mul_108_22_n_676);
  or mul_108_22_g3279(mul_108_22_n_754 ,mul_108_22_n_654 ,mul_108_22_n_674);
  or mul_108_22_g3280(mul_108_22_n_753 ,mul_108_22_n_456 ,mul_108_22_n_642);
  or mul_108_22_g3281(mul_108_22_n_752 ,mul_108_22_n_668 ,mul_108_22_n_610);
  and mul_108_22_g3282(mul_108_22_n_751 ,mul_108_22_n_456 ,mul_108_22_n_642);
  or mul_108_22_g3283(mul_108_22_n_750 ,mul_108_22_n_601 ,mul_108_22_n_617);
  nor mul_108_22_g3284(mul_108_22_n_749 ,mul_108_22_n_604 ,mul_108_22_n_655);
  or mul_108_22_g3285(mul_108_22_n_748 ,mul_108_22_n_652 ,mul_108_22_n_615);
  or mul_108_22_g3286(mul_108_22_n_747 ,mul_108_22_n_451 ,mul_108_22_n_651);
  nor mul_108_22_g3287(mul_108_22_n_746 ,mul_108_22_n_306 ,mul_108_22_n_677);
  or mul_108_22_g3288(mul_108_22_n_745 ,mul_108_22_n_665 ,mul_108_22_n_607);
  and mul_108_22_g3289(mul_108_22_n_744 ,mul_108_22_n_672 ,mul_108_22_n_666);
  or mul_108_22_g3290(mul_108_22_n_743 ,mul_108_22_n_675 ,mul_108_22_n_678);
  and mul_108_22_g3291(mul_108_22_n_742 ,mul_108_22_n_675 ,mul_108_22_n_678);
  nor mul_108_22_g3292(mul_108_22_n_741 ,mul_108_22_n_653 ,mul_108_22_n_616);
  nor mul_108_22_g3293(mul_108_22_n_740 ,mul_108_22_n_661 ,mul_108_22_n_658);
  and mul_108_22_g3294(mul_108_22_n_739 ,mul_108_22_n_667 ,mul_108_22_n_664);
  or mul_108_22_g3295(mul_108_22_n_738 ,mul_108_22_n_660 ,mul_108_22_n_659);
  or mul_108_22_g3296(mul_108_22_n_737 ,mul_108_22_n_612 ,mul_108_22_n_657);
  or mul_108_22_g3297(mul_108_22_n_736 ,mul_108_22_n_667 ,mul_108_22_n_664);
  or mul_108_22_g3298(mul_108_22_n_735 ,mul_108_22_n_449 ,mul_108_22_n_673);
  and mul_108_22_g3299(mul_108_22_n_768 ,mul_108_22_n_547 ,mul_108_22_n_699);
  and mul_108_22_g3300(mul_108_22_n_766 ,mul_108_22_n_681 ,mul_108_22_n_686);
  and mul_108_22_g3301(mul_108_22_n_765 ,mul_108_22_n_638 ,mul_108_22_n_689);
  or mul_108_22_g3302(mul_108_22_n_763 ,mul_108_22_n_680 ,mul_108_22_n_696);
  and mul_108_22_g3303(mul_108_22_n_762 ,mul_108_22_n_626 ,mul_108_22_n_691);
  and mul_108_22_g3304(mul_108_22_n_759 ,mul_108_22_n_684 ,mul_108_22_n_683);
  and mul_108_22_g3305(mul_108_22_n_758 ,mul_108_22_n_628 ,mul_108_22_n_637);
  or mul_108_22_g3306(mul_108_22_n_756 ,mul_108_22_n_695 ,mul_108_22_n_693);
  not mul_108_22_g3307(mul_108_22_n_734 ,mul_108_22_n_733);
  not mul_108_22_g3308(mul_108_22_n_732 ,mul_108_22_n_731);
  not mul_108_22_g3309(mul_108_22_n_730 ,mul_108_22_n_729);
  or mul_108_22_g3310(mul_108_22_n_727 ,mul_108_22_n_311 ,mul_108_22_n_591);
  and mul_108_22_g3311(mul_108_22_n_726 ,mul_108_22_n_654 ,mul_108_22_n_674);
  nor mul_108_22_g3312(mul_108_22_n_725 ,mul_108_22_n_671 ,mul_108_22_n_611);
  and mul_108_22_g3313(mul_108_22_n_724 ,mul_108_22_n_449 ,mul_108_22_n_673);
  and mul_108_22_g3314(mul_108_22_n_723 ,mul_108_22_n_612 ,mul_108_22_n_657);
  or mul_108_22_g3315(mul_108_22_n_722 ,mul_108_22_n_600 ,mul_108_22_n_608);
  or mul_108_22_g3316(mul_108_22_n_721 ,mul_108_22_n_598 ,mul_108_22_n_606);
  or mul_108_22_g3317(mul_108_22_n_720 ,mul_108_22_n_307 ,mul_108_22_n_613);
  nor mul_108_22_g3318(mul_108_22_n_719 ,mul_108_22_n_650 ,mul_108_22_n_614);
  and mul_108_22_g3319(mul_108_22_n_718 ,mul_108_22_n_668 ,mul_108_22_n_610);
  and mul_108_22_g3320(mul_108_22_n_717 ,mul_108_22_n_598 ,mul_108_22_n_606);
  and mul_108_22_g3321(mul_108_22_n_716 ,mul_108_22_n_451 ,mul_108_22_n_651);
  or mul_108_22_g3322(mul_108_22_n_715 ,mul_108_22_n_672 ,mul_108_22_n_666);
  and mul_108_22_g3323(mul_108_22_n_714 ,mul_108_22_n_600 ,mul_108_22_n_608);
  or mul_108_22_g3324(mul_108_22_n_713 ,mul_108_22_n_669 ,mul_108_22_n_609);
  and mul_108_22_g3325(mul_108_22_n_712 ,mul_108_22_n_671 ,mul_108_22_n_611);
  and mul_108_22_g3326(mul_108_22_n_711 ,mul_108_22_n_669 ,mul_108_22_n_609);
  or mul_108_22_g3327(mul_108_22_n_710 ,mul_108_22_n_597 ,mul_108_22_n_592);
  or mul_108_22_g3328(mul_108_22_n_709 ,mul_108_22_n_450 ,mul_108_22_n_605);
  and mul_108_22_g3329(mul_108_22_n_708 ,mul_108_22_n_450 ,mul_108_22_n_605);
  and mul_108_22_g3330(mul_108_22_n_707 ,mul_108_22_n_597 ,mul_108_22_n_592);
  or mul_108_22_g3331(mul_108_22_n_706 ,mul_108_22_n_603 ,mul_108_22_n_656);
  nor mul_108_22_g3332(mul_108_22_n_705 ,mul_108_22_n_596 ,mul_108_22_n_594);
  or mul_108_22_g3333(mul_108_22_n_704 ,mul_108_22_n_595 ,mul_108_22_n_593);
  nor mul_108_22_g3334(mul_108_22_n_703 ,mul_108_22_n_602 ,mul_108_22_n_618);
  and mul_108_22_g3335(mul_108_22_n_702 ,mul_108_22_n_665 ,mul_108_22_n_607);
  and mul_108_22_g3336(mul_108_22_n_733 ,mul_108_22_n_545 ,mul_108_22_n_640);
  and mul_108_22_g3337(mul_108_22_n_731 ,mul_108_22_n_546 ,mul_108_22_n_635);
  or mul_108_22_g3338(mul_108_22_n_729 ,mul_108_22_n_620 ,mul_108_22_n_629);
  and mul_108_22_g3339(mul_108_22_n_728 ,mul_108_22_n_645 ,mul_108_22_n_701);
  not mul_108_22_g3340(mul_108_22_n_701 ,mul_108_22_n_700);
  not mul_108_22_g3341(mul_108_22_n_699 ,mul_108_22_n_698);
  not mul_108_22_g3342(mul_108_22_n_695 ,mul_108_22_n_694);
  not mul_108_22_g3343(mul_108_22_n_691 ,mul_108_22_n_690);
  not mul_108_22_g3344(mul_108_22_n_689 ,mul_108_22_n_688);
  not mul_108_22_g3345(mul_108_22_n_686 ,mul_108_22_n_685);
  not mul_108_22_g3346(mul_108_22_n_683 ,mul_108_22_n_682);
  not mul_108_22_g3347(mul_108_22_n_680 ,mul_108_22_n_679);
  not mul_108_22_g3348(mul_108_22_n_676 ,mul_108_22_n_677);
  not mul_108_22_g3349(mul_108_22_n_671 ,mul_108_22_n_670);
  not mul_108_22_g3350(mul_108_22_n_662 ,mul_108_22_n_663);
  not mul_108_22_g3351(mul_108_22_n_660 ,mul_108_22_n_661);
  not mul_108_22_g3352(mul_108_22_n_658 ,mul_108_22_n_659);
  not mul_108_22_g3353(mul_108_22_n_655 ,mul_108_22_n_656);
  not mul_108_22_g3354(mul_108_22_n_652 ,mul_108_22_n_653);
  or mul_108_22_g3358(mul_108_22_n_700 ,mul_108_22_n_502 ,mul_108_22_n_578);
  and mul_108_22_g3359(mul_108_22_n_698 ,mul_108_22_n_422 ,mul_108_22_n_536);
  or mul_108_22_g3360(mul_108_22_n_647 ,mul_108_22_n_457 ,mul_108_22_n_506);
  or mul_108_22_g3361(mul_108_22_n_646 ,mul_108_22_n_497 ,mul_108_22_n_580);
  and mul_108_22_g3362(mul_108_22_n_697 ,mul_108_22_n_429 ,mul_108_22_n_565);
  and mul_108_22_g3363(mul_108_22_n_696 ,mul_108_22_n_460 ,mul_108_22_n_561);
  or mul_108_22_g3364(mul_108_22_n_694 ,mul_108_22_n_500 ,mul_108_22_n_588);
  and mul_108_22_g3365(mul_108_22_n_693 ,mul_108_22_n_466 ,mul_108_22_n_573);
  and mul_108_22_g3366(mul_108_22_n_692 ,mul_108_22_n_461 ,mul_108_22_n_517);
  and mul_108_22_g3367(mul_108_22_n_690 ,mul_108_22_n_470 ,mul_108_22_n_526);
  and mul_108_22_g3368(mul_108_22_n_688 ,mul_108_22_n_472 ,mul_108_22_n_562);
  or mul_108_22_g3369(mul_108_22_n_687 ,mul_108_22_n_495 ,mul_108_22_n_587);
  and mul_108_22_g3370(mul_108_22_n_685 ,mul_108_22_n_412 ,mul_108_22_n_563);
  or mul_108_22_g3371(mul_108_22_n_684 ,mul_108_22_n_499 ,mul_108_22_n_585);
  and mul_108_22_g3372(mul_108_22_n_682 ,mul_108_22_n_441 ,mul_108_22_n_568);
  or mul_108_22_g3373(mul_108_22_n_681 ,mul_108_22_n_491 ,mul_108_22_n_582);
  or mul_108_22_g3374(mul_108_22_n_679 ,mul_108_22_n_501 ,mul_108_22_n_589);
  and mul_108_22_g3375(mul_108_22_n_678 ,mul_108_22_n_471 ,mul_108_22_n_528);
  and mul_108_22_g3376(mul_108_22_n_677 ,mul_108_22_n_440 ,mul_108_22_n_567);
  and mul_108_22_g3377(mul_108_22_n_675 ,mul_108_22_n_464 ,mul_108_22_n_529);
  and mul_108_22_g3378(mul_108_22_n_674 ,mul_108_22_n_467 ,mul_108_22_n_538);
  and mul_108_22_g3379(mul_108_22_n_673 ,mul_108_22_n_443 ,mul_108_22_n_555);
  and mul_108_22_g3380(mul_108_22_n_672 ,mul_108_22_n_459 ,mul_108_22_n_521);
  or mul_108_22_g3381(mul_108_22_n_670 ,mul_108_22_n_492 ,mul_108_22_n_579);
  and mul_108_22_g3382(mul_108_22_n_669 ,mul_108_22_n_434 ,mul_108_22_n_514);
  and mul_108_22_g3383(mul_108_22_n_668 ,mul_108_22_n_462 ,mul_108_22_n_535);
  and mul_108_22_g3384(mul_108_22_n_667 ,mul_108_22_n_473 ,mul_108_22_n_524);
  and mul_108_22_g3385(mul_108_22_n_666 ,mul_108_22_n_436 ,mul_108_22_n_533);
  and mul_108_22_g3386(mul_108_22_n_665 ,mul_108_22_n_432 ,mul_108_22_n_552);
  and mul_108_22_g3387(mul_108_22_n_664 ,mul_108_22_n_423 ,mul_108_22_n_523);
  and mul_108_22_g3388(mul_108_22_n_663 ,mul_108_22_n_426 ,mul_108_22_n_518);
  or mul_108_22_g3389(mul_108_22_n_661 ,mul_108_22_n_494 ,mul_108_22_n_540);
  and mul_108_22_g3390(mul_108_22_n_659 ,mul_108_22_n_433 ,mul_108_22_n_558);
  and mul_108_22_g3391(mul_108_22_n_657 ,mul_108_22_n_431 ,mul_108_22_n_531);
  or mul_108_22_g3392(mul_108_22_n_656 ,mul_108_22_n_454 ,mul_108_22_n_504);
  and mul_108_22_g3393(mul_108_22_n_654 ,mul_108_22_n_418 ,mul_108_22_n_527);
  or mul_108_22_g3394(mul_108_22_n_653 ,mul_108_22_n_452 ,mul_108_22_n_505);
  and mul_108_22_g3395(mul_108_22_n_651 ,mul_108_22_n_413 ,mul_108_22_n_532);
  or mul_108_22_g3396(mul_108_22_n_650 ,mul_108_22_n_493 ,mul_108_22_n_577);
  and mul_108_22_g3397(mul_108_22_n_649 ,mul_108_22_n_425 ,mul_108_22_n_559);
  or mul_108_22_g3398(mul_108_22_n_648 ,mul_108_22_n_498 ,mul_108_22_n_584);
  not mul_108_22_g3399(mul_108_22_n_644 ,mul_108_22_n_643);
  not mul_108_22_g3400(mul_108_22_n_640 ,mul_108_22_n_639);
  not mul_108_22_g3401(mul_108_22_n_637 ,mul_108_22_n_636);
  not mul_108_22_g3402(mul_108_22_n_635 ,mul_108_22_n_634);
  not mul_108_22_g3403(mul_108_22_n_626 ,mul_108_22_n_625);
  not mul_108_22_g3404(mul_108_22_n_620 ,mul_108_22_n_619);
  not mul_108_22_g3405(mul_108_22_n_617 ,mul_108_22_n_618);
  not mul_108_22_g3406(mul_108_22_n_615 ,mul_108_22_n_616);
  not mul_108_22_g3407(mul_108_22_n_613 ,mul_108_22_n_614);
  not mul_108_22_g3408(mul_108_22_n_603 ,mul_108_22_n_604);
  not mul_108_22_g3409(mul_108_22_n_601 ,mul_108_22_n_602);
  not mul_108_22_g3411(mul_108_22_n_595 ,mul_108_22_n_596);
  not mul_108_22_g3412(mul_108_22_n_593 ,mul_108_22_n_594);
  nor mul_108_22_g3413(mul_108_22_n_591 ,mul_108_22_n_486 ,mul_108_22_n_574);
  or mul_108_22_g3414(mul_108_22_n_645 ,mul_108_22_n_324 ,mul_108_22_n_507);
  and mul_108_22_g3415(mul_108_22_n_643 ,mul_108_22_n_488 ,mul_108_22_n_571);
  and mul_108_22_g3416(mul_108_22_n_642 ,mul_108_22_n_478 ,mul_108_22_n_570);
  and mul_108_22_g3417(mul_108_22_n_641 ,mul_108_22_n_481 ,mul_108_22_n_572);
  and mul_108_22_g3418(mul_108_22_n_639 ,mul_108_22_n_421 ,mul_108_22_n_575);
  or mul_108_22_g3419(mul_108_22_n_638 ,mul_108_22_n_490 ,mul_108_22_n_581);
  and mul_108_22_g3420(mul_108_22_n_636 ,mul_108_22_n_428 ,mul_108_22_n_512);
  and mul_108_22_g3421(mul_108_22_n_634 ,mul_108_22_n_468 ,mul_108_22_n_539);
  and mul_108_22_g3422(mul_108_22_n_633 ,mul_108_22_n_430 ,mul_108_22_n_509);
  and mul_108_22_g3423(mul_108_22_n_632 ,mul_108_22_n_484 ,mul_108_22_n_590);
  and mul_108_22_g3424(mul_108_22_n_631 ,mul_108_22_n_437 ,mul_108_22_n_520);
  and mul_108_22_g3425(mul_108_22_n_630 ,mul_108_22_n_325 ,mul_108_22_n_556);
  and mul_108_22_g3426(mul_108_22_n_629 ,mul_108_22_n_427 ,mul_108_22_n_519);
  or mul_108_22_g3427(mul_108_22_n_628 ,mul_108_22_n_496 ,mul_108_22_n_569);
  and mul_108_22_g3428(mul_108_22_n_627 ,mul_108_22_n_482 ,mul_108_22_n_566);
  and mul_108_22_g3429(mul_108_22_n_625 ,mul_108_22_n_479 ,mul_108_22_n_560);
  and mul_108_22_g3430(mul_108_22_n_624 ,mul_108_22_n_477 ,mul_108_22_n_576);
  and mul_108_22_g3431(mul_108_22_n_623 ,mul_108_22_n_475 ,mul_108_22_n_557);
  and mul_108_22_g3432(mul_108_22_n_622 ,mul_108_22_n_474 ,mul_108_22_n_553);
  and mul_108_22_g3433(mul_108_22_n_621 ,mul_108_22_n_487 ,mul_108_22_n_541);
  or mul_108_22_g3434(mul_108_22_n_619 ,mul_108_22_n_503 ,mul_108_22_n_583);
  and mul_108_22_g3435(mul_108_22_n_618 ,mul_108_22_n_416 ,mul_108_22_n_530);
  and mul_108_22_g3436(mul_108_22_n_616 ,mul_108_22_n_420 ,mul_108_22_n_542);
  and mul_108_22_g3437(mul_108_22_n_614 ,mul_108_22_n_458 ,mul_108_22_n_564);
  and mul_108_22_g3438(mul_108_22_n_612 ,mul_108_22_n_455 ,mul_108_22_n_543);
  and mul_108_22_g3439(mul_108_22_n_611 ,mul_108_22_n_453 ,mul_108_22_n_515);
  and mul_108_22_g3440(mul_108_22_n_610 ,mul_108_22_n_438 ,mul_108_22_n_534);
  and mul_108_22_g3441(mul_108_22_n_609 ,mul_108_22_n_469 ,mul_108_22_n_513);
  and mul_108_22_g3442(mul_108_22_n_608 ,mul_108_22_n_442 ,mul_108_22_n_537);
  and mul_108_22_g3443(mul_108_22_n_607 ,mul_108_22_n_419 ,mul_108_22_n_510);
  and mul_108_22_g3444(mul_108_22_n_606 ,mul_108_22_n_463 ,mul_108_22_n_516);
  and mul_108_22_g3445(mul_108_22_n_605 ,mul_108_22_n_465 ,mul_108_22_n_511);
  or mul_108_22_g3446(mul_108_22_n_604 ,mul_108_22_n_489 ,mul_108_22_n_586);
  and mul_108_22_g3447(mul_108_22_n_602 ,mul_108_22_n_485 ,mul_108_22_n_522);
  and mul_108_22_g3448(mul_108_22_n_600 ,mul_108_22_n_435 ,mul_108_22_n_548);
  and mul_108_22_g3449(mul_108_22_n_599 ,mul_108_22_n_483 ,mul_108_22_n_551);
  and mul_108_22_g3450(mul_108_22_n_598 ,mul_108_22_n_476 ,mul_108_22_n_554);
  and mul_108_22_g3451(mul_108_22_n_597 ,mul_108_22_n_417 ,mul_108_22_n_550);
  and mul_108_22_g3452(mul_108_22_n_596 ,mul_108_22_n_480 ,mul_108_22_n_549);
  and mul_108_22_g3453(mul_108_22_n_594 ,mul_108_22_n_411 ,mul_108_22_n_525);
  and mul_108_22_g3454(mul_108_22_n_592 ,mul_108_22_n_414 ,mul_108_22_n_508);
  or mul_108_22_g3455(mul_108_22_n_590 ,mul_108_22_n_353 ,mul_108_22_n_66);
  and mul_108_22_g3456(mul_108_22_n_589 ,mul_108_22_n_140 ,mul_108_22_n_33);
  and mul_108_22_g3457(mul_108_22_n_588 ,mul_108_22_n_90 ,mul_108_22_n_45);
  and mul_108_22_g3458(mul_108_22_n_587 ,mul_108_22_n_132 ,mul_108_22_n_16);
  and mul_108_22_g3459(mul_108_22_n_586 ,mul_108_22_n_128 ,mul_108_22_n_33);
  and mul_108_22_g3460(mul_108_22_n_585 ,mul_108_22_n_110 ,mul_108_22_n_34);
  and mul_108_22_g3461(mul_108_22_n_584 ,mul_108_22_n_92 ,mul_108_22_n_46);
  and mul_108_22_g3462(mul_108_22_n_583 ,mul_108_22_n_142 ,mul_108_22_n_22);
  and mul_108_22_g3463(mul_108_22_n_582 ,mul_108_22_n_144 ,mul_108_22_n_21);
  and mul_108_22_g3464(mul_108_22_n_581 ,mul_108_22_n_134 ,mul_108_22_n_34);
  and mul_108_22_g3465(mul_108_22_n_580 ,mul_108_22_n_138 ,mul_108_22_n_21);
  and mul_108_22_g3466(mul_108_22_n_579 ,mul_108_22_n_120 ,mul_108_22_n_46);
  and mul_108_22_g3467(mul_108_22_n_578 ,mul_108_22_n_94 ,mul_108_22_n_45);
  and mul_108_22_g3468(mul_108_22_n_577 ,mul_108_22_n_126 ,mul_108_22_n_170);
  or mul_108_22_g3469(mul_108_22_n_576 ,mul_108_22_n_351 ,mul_108_22_n_76);
  or mul_108_22_g3470(mul_108_22_n_575 ,mul_108_22_n_328 ,mul_108_22_n_25);
  nor mul_108_22_g3471(mul_108_22_n_574 ,mul_108_22_n_76 ,mul_108_22_n_330);
  or mul_108_22_g3472(mul_108_22_n_573 ,mul_108_22_n_344 ,mul_108_22_n_58);
  or mul_108_22_g3473(mul_108_22_n_572 ,mul_108_22_n_338 ,mul_108_22_n_75);
  or mul_108_22_g3474(mul_108_22_n_571 ,mul_108_22_n_347 ,mul_108_22_n_40);
  or mul_108_22_g3475(mul_108_22_n_570 ,mul_108_22_n_365 ,mul_108_22_n_39);
  and mul_108_22_g3476(mul_108_22_n_569 ,mul_108_22_n_136 ,mul_108_22_n_22);
  or mul_108_22_g3477(mul_108_22_n_568 ,mul_108_22_n_362 ,mul_108_22_n_37);
  or mul_108_22_g3478(mul_108_22_n_567 ,mul_108_22_n_349 ,mul_108_22_n_57);
  or mul_108_22_g3479(mul_108_22_n_566 ,mul_108_22_n_360 ,mul_108_22_n_40);
  or mul_108_22_g3480(mul_108_22_n_565 ,mul_108_22_n_341 ,mul_108_22_n_81);
  or mul_108_22_g3481(mul_108_22_n_564 ,mul_108_22_n_346 ,mul_108_22_n_36);
  or mul_108_22_g3482(mul_108_22_n_563 ,mul_108_22_n_366 ,mul_108_22_n_25);
  or mul_108_22_g3483(mul_108_22_n_562 ,mul_108_22_n_354 ,mul_108_22_n_24);
  or mul_108_22_g3484(mul_108_22_n_561 ,mul_108_22_n_369 ,mul_108_22_n_24);
  or mul_108_22_g3485(mul_108_22_n_560 ,mul_108_22_n_350 ,mul_108_22_n_14);
  or mul_108_22_g3486(mul_108_22_n_559 ,mul_108_22_n_368 ,mul_108_22_n_37);
  or mul_108_22_g3487(mul_108_22_n_558 ,mul_108_22_n_345 ,mul_108_22_n_57);
  or mul_108_22_g3488(mul_108_22_n_557 ,mul_108_22_n_355 ,mul_108_22_n_88);
  or mul_108_22_g3489(mul_108_22_n_556 ,mul_108_22_n_364 ,mul_108_22_n_39);
  or mul_108_22_g3490(mul_108_22_n_555 ,mul_108_22_n_358 ,mul_108_22_n_81);
  or mul_108_22_g3491(mul_108_22_n_554 ,mul_108_22_n_352 ,mul_108_22_n_66);
  or mul_108_22_g3492(mul_108_22_n_553 ,mul_108_22_n_337 ,mul_108_22_n_75);
  or mul_108_22_g3493(mul_108_22_n_552 ,mul_108_22_n_343 ,mul_108_22_n_36);
  or mul_108_22_g3494(mul_108_22_n_551 ,mul_108_22_n_361 ,mul_108_22_n_67);
  or mul_108_22_g3495(mul_108_22_n_550 ,mul_108_22_n_359 ,mul_108_22_n_10);
  or mul_108_22_g3496(mul_108_22_n_549 ,mul_108_22_n_357 ,mul_108_22_n_87);
  or mul_108_22_g3497(mul_108_22_n_548 ,mul_108_22_n_342 ,mul_108_22_n_10);
  not mul_108_22_g3498(mul_108_22_n_545 ,mul_108_22_n_544);
  or mul_108_22_g3499(mul_108_22_n_543 ,mul_108_22_n_392 ,mul_108_22_n_49);
  or mul_108_22_g3500(mul_108_22_n_542 ,mul_108_22_n_356 ,mul_108_22_n_82);
  or mul_108_22_g3501(mul_108_22_n_541 ,mul_108_22_n_340 ,mul_108_22_n_87);
  and mul_108_22_g3502(mul_108_22_n_540 ,mul_108_22_n_165 ,mul_108_22_n_16);
  or mul_108_22_g3503(mul_108_22_n_539 ,mul_108_22_n_377 ,mul_108_22_n_31);
  or mul_108_22_g3504(mul_108_22_n_538 ,mul_108_22_n_388 ,mul_108_22_n_64);
  or mul_108_22_g3505(mul_108_22_n_537 ,mul_108_22_n_407 ,mul_108_22_n_28);
  or mul_108_22_g3506(mul_108_22_n_536 ,mul_108_22_n_370 ,mul_108_22_n_63);
  or mul_108_22_g3507(mul_108_22_n_535 ,mul_108_22_n_405 ,mul_108_22_n_61);
  or mul_108_22_g3508(mul_108_22_n_534 ,mul_108_22_n_404 ,mul_108_22_n_84);
  or mul_108_22_g3509(mul_108_22_n_533 ,mul_108_22_n_386 ,mul_108_22_n_27);
  or mul_108_22_g3510(mul_108_22_n_532 ,mul_108_22_n_399 ,mul_108_22_n_49);
  or mul_108_22_g3511(mul_108_22_n_531 ,mul_108_22_n_390 ,mul_108_22_n_52);
  or mul_108_22_g3512(mul_108_22_n_530 ,mul_108_22_n_339 ,mul_108_22_n_48);
  or mul_108_22_g3513(mul_108_22_n_529 ,mul_108_22_n_410 ,mul_108_22_n_60);
  or mul_108_22_g3514(mul_108_22_n_528 ,mul_108_22_n_385 ,mul_108_22_n_48);
  or mul_108_22_g3515(mul_108_22_n_527 ,mul_108_22_n_389 ,mul_108_22_n_78);
  or mul_108_22_g3516(mul_108_22_n_526 ,mul_108_22_n_408 ,mul_108_22_n_28);
  or mul_108_22_g3517(mul_108_22_n_525 ,mul_108_22_n_397 ,mul_108_22_n_63);
  or mul_108_22_g3518(mul_108_22_n_524 ,mul_108_22_n_395 ,mul_108_22_n_51);
  or mul_108_22_g3519(mul_108_22_n_523 ,mul_108_22_n_403 ,mul_108_22_n_84);
  or mul_108_22_g3520(mul_108_22_n_522 ,mul_108_22_n_348 ,mul_108_22_n_14);
  or mul_108_22_g3521(mul_108_22_n_521 ,mul_108_22_n_406 ,mul_108_22_n_31);
  or mul_108_22_g3522(mul_108_22_n_520 ,mul_108_22_n_396 ,mul_108_22_n_30);
  or mul_108_22_g3523(mul_108_22_n_519 ,mul_108_22_n_363 ,mul_108_22_n_30);
  or mul_108_22_g3524(mul_108_22_n_518 ,mul_108_22_n_391 ,mul_108_22_n_52);
  or mul_108_22_g3525(mul_108_22_n_517 ,mul_108_22_n_394 ,mul_108_22_n_60);
  or mul_108_22_g3526(mul_108_22_n_516 ,mul_108_22_n_400 ,mul_108_22_n_27);
  or mul_108_22_g3527(mul_108_22_n_515 ,mul_108_22_n_387 ,mul_108_22_n_78);
  or mul_108_22_g3528(mul_108_22_n_514 ,mul_108_22_n_384 ,mul_108_22_n_51);
  or mul_108_22_g3529(mul_108_22_n_513 ,mul_108_22_n_409 ,mul_108_22_n_8);
  or mul_108_22_g3530(mul_108_22_n_512 ,mul_108_22_n_393 ,mul_108_22_n_12);
  or mul_108_22_g3531(mul_108_22_n_511 ,mul_108_22_n_401 ,mul_108_22_n_12);
  or mul_108_22_g3532(mul_108_22_n_510 ,mul_108_22_n_367 ,mul_108_22_n_79);
  or mul_108_22_g3533(mul_108_22_n_509 ,mul_108_22_n_402 ,mul_108_22_n_8);
  or mul_108_22_g3534(mul_108_22_n_508 ,mul_108_22_n_398 ,mul_108_22_n_85);
  nor mul_108_22_g3535(mul_108_22_n_507 ,mul_108_22_n_67 ,mul_108_22_n_311);
  nor mul_108_22_g3536(mul_108_22_n_506 ,mul_108_22_n_58 ,mul_108_22_n_310);
  nor mul_108_22_g3537(mul_108_22_n_505 ,mul_108_22_n_61 ,mul_108_22_n_315);
  nor mul_108_22_g3538(mul_108_22_n_504 ,mul_108_22_n_64 ,mul_108_22_n_316);
  and mul_108_22_g3539(mul_108_22_n_547 ,in24[3] ,mul_108_22_n_439);
  and mul_108_22_g3540(mul_108_22_n_546 ,in24[5] ,mul_108_22_n_415);
  or mul_108_22_g3541(mul_108_22_n_544 ,mul_108_22_n_310 ,mul_108_22_n_424);
  and mul_108_22_g3542(mul_108_22_n_503 ,mul_108_22_n_134 ,mul_108_22_n_246);
  and mul_108_22_g3543(mul_108_22_n_502 ,mul_108_22_n_92 ,mul_108_22_n_236);
  and mul_108_22_g3544(mul_108_22_n_501 ,mul_108_22_n_136 ,mul_108_22_n_209);
  and mul_108_22_g3545(mul_108_22_n_500 ,mul_108_22_n_94 ,mul_108_22_n_237);
  and mul_108_22_g3546(mul_108_22_n_499 ,mul_108_22_n_140 ,mul_108_22_n_209);
  and mul_108_22_g3547(mul_108_22_n_498 ,mul_108_22_n_128 ,mul_108_22_n_210);
  and mul_108_22_g3548(mul_108_22_n_497 ,mul_108_22_n_252 ,mul_108_22_n_210);
  and mul_108_22_g3549(mul_108_22_n_496 ,mul_108_22_n_142 ,mul_108_22_n_237);
  and mul_108_22_g3550(mul_108_22_n_495 ,mul_108_22_n_126 ,mul_108_22_n_200);
  and mul_108_22_g3551(mul_108_22_n_494 ,mul_108_22_n_144 ,mul_108_22_n_199);
  and mul_108_22_g3552(mul_108_22_n_493 ,mul_108_22_n_138 ,mul_108_22_n_236);
  and mul_108_22_g3553(mul_108_22_n_492 ,mul_108_22_n_132 ,mul_108_22_n_246);
  and mul_108_22_g3554(mul_108_22_n_491 ,mul_108_22_n_110 ,mul_108_22_n_200);
  and mul_108_22_g3555(mul_108_22_n_490 ,mul_108_22_n_90 ,mul_108_22_n_245);
  and mul_108_22_g3556(mul_108_22_n_489 ,mul_108_22_n_120 ,mul_108_22_n_245);
  or mul_108_22_g3557(mul_108_22_n_488 ,mul_108_22_n_70 ,mul_108_22_n_338);
  or mul_108_22_g3558(mul_108_22_n_487 ,mul_108_22_n_42 ,mul_108_22_n_337);
  nor mul_108_22_g3559(mul_108_22_n_486 ,mul_108_22_n_73 ,mul_108_22_n_365);
  or mul_108_22_g3560(mul_108_22_n_485 ,mul_108_22_n_54 ,mul_108_22_n_357);
  or mul_108_22_g3561(mul_108_22_n_484 ,mul_108_22_n_72 ,mul_108_22_n_340);
  or mul_108_22_g3562(mul_108_22_n_483 ,mul_108_22_n_69 ,mul_108_22_n_352);
  or mul_108_22_g3563(mul_108_22_n_482 ,mul_108_22_n_43 ,mul_108_22_n_353);
  or mul_108_22_g3564(mul_108_22_n_481 ,mul_108_22_n_55 ,mul_108_22_n_348);
  or mul_108_22_g3565(mul_108_22_n_480 ,mul_108_22_n_72 ,mul_108_22_n_361);
  or mul_108_22_g3566(mul_108_22_n_479 ,mul_108_22_n_69 ,mul_108_22_n_360);
  or mul_108_22_g3567(mul_108_22_n_478 ,mul_108_22_n_42 ,mul_108_22_n_347);
  or mul_108_22_g3568(mul_108_22_n_477 ,mul_108_22_n_54 ,mul_108_22_n_364);
  or mul_108_22_g3569(mul_108_22_n_476 ,mul_108_22_n_55 ,mul_108_22_n_355);
  or mul_108_22_g3570(mul_108_22_n_475 ,mul_108_22_n_43 ,mul_108_22_n_350);
  or mul_108_22_g3571(mul_108_22_n_474 ,mul_108_22_n_73 ,mul_108_22_n_351);
  or mul_108_22_g3572(mul_108_22_n_473 ,mul_108_22_n_406 ,mul_108_22_n_224);
  or mul_108_22_g3573(mul_108_22_n_472 ,mul_108_22_n_344 ,mul_108_22_n_215);
  or mul_108_22_g3574(mul_108_22_n_471 ,mul_108_22_n_404 ,mul_108_22_n_239);
  or mul_108_22_g3575(mul_108_22_n_470 ,mul_108_22_n_385 ,mul_108_22_n_206);
  or mul_108_22_g3576(mul_108_22_n_469 ,mul_108_22_n_400 ,mul_108_22_n_206);
  or mul_108_22_g3577(mul_108_22_n_468 ,mul_108_22_n_401 ,mul_108_22_n_233);
  or mul_108_22_g3578(mul_108_22_n_467 ,mul_108_22_n_408 ,mul_108_22_n_240);
  or mul_108_22_g3579(mul_108_22_n_466 ,mul_108_22_n_343 ,mul_108_22_n_218);
  or mul_108_22_g3580(mul_108_22_n_465 ,mul_108_22_n_384 ,mul_108_22_n_233);
  or mul_108_22_g3581(mul_108_22_n_464 ,mul_108_22_n_405 ,mul_108_22_n_225);
  or mul_108_22_g3582(mul_108_22_n_463 ,mul_108_22_n_388 ,mul_108_22_n_243);
  or mul_108_22_g3583(mul_108_22_n_462 ,mul_108_22_n_393 ,mul_108_22_n_228);
  or mul_108_22_g3584(mul_108_22_n_461 ,mul_108_22_n_387 ,mul_108_22_n_224);
  or mul_108_22_g3585(mul_108_22_n_460 ,mul_108_22_n_359 ,mul_108_22_n_218);
  or mul_108_22_g3586(mul_108_22_n_459 ,mul_108_22_n_367 ,mul_108_22_n_227);
  not mul_108_22_g3587(mul_108_22_n_458 ,mul_108_22_n_457);
  not mul_108_22_g3588(mul_108_22_n_455 ,mul_108_22_n_454);
  not mul_108_22_g3589(mul_108_22_n_453 ,mul_108_22_n_452);
  or mul_108_22_g3590(mul_108_22_n_443 ,mul_108_22_n_345 ,mul_108_22_n_216);
  or mul_108_22_g3591(mul_108_22_n_442 ,mul_108_22_n_403 ,mul_108_22_n_239);
  or mul_108_22_g3592(mul_108_22_n_441 ,mul_108_22_n_369 ,mul_108_22_n_249);
  or mul_108_22_g3593(mul_108_22_n_440 ,mul_108_22_n_368 ,mul_108_22_n_215);
  or mul_108_22_g3594(mul_108_22_n_439 ,mul_108_22_n_321 ,mul_108_22_n_376);
  or mul_108_22_g3595(mul_108_22_n_438 ,mul_108_22_n_398 ,mul_108_22_n_242);
  or mul_108_22_g3596(mul_108_22_n_437 ,mul_108_22_n_389 ,mul_108_22_n_230);
  or mul_108_22_g3597(mul_108_22_n_436 ,mul_108_22_n_402 ,mul_108_22_n_212);
  or mul_108_22_g3598(mul_108_22_n_435 ,mul_108_22_n_354 ,mul_108_22_n_248);
  or mul_108_22_g3599(mul_108_22_n_434 ,mul_108_22_n_396 ,mul_108_22_n_230);
  or mul_108_22_g3600(mul_108_22_n_433 ,mul_108_22_n_366 ,mul_108_22_n_221);
  or mul_108_22_g3601(mul_108_22_n_432 ,mul_108_22_n_341 ,mul_108_22_n_221);
  or mul_108_22_g3602(mul_108_22_n_431 ,mul_108_22_n_394 ,mul_108_22_n_227);
  or mul_108_22_g3603(mul_108_22_n_430 ,mul_108_22_n_392 ,mul_108_22_n_212);
  or mul_108_22_g3604(mul_108_22_n_429 ,mul_108_22_n_349 ,mul_108_22_n_248);
  or mul_108_22_g3605(mul_108_22_n_428 ,mul_108_22_n_363 ,mul_108_22_n_234);
  or mul_108_22_g3606(mul_108_22_n_427 ,mul_108_22_n_395 ,mul_108_22_n_228);
  or mul_108_22_g3607(mul_108_22_n_426 ,mul_108_22_n_410 ,mul_108_22_n_231);
  or mul_108_22_g3608(mul_108_22_n_425 ,mul_108_22_n_356 ,mul_108_22_n_219);
  nor mul_108_22_g3609(mul_108_22_n_424 ,mul_108_22_n_320 ,mul_108_22_n_374);
  or mul_108_22_g3610(mul_108_22_n_423 ,mul_108_22_n_386 ,mul_108_22_n_242);
  or mul_108_22_g3611(mul_108_22_n_422 ,mul_108_22_n_399 ,mul_108_22_n_207);
  or mul_108_22_g3612(mul_108_22_n_421 ,mul_108_22_n_358 ,mul_108_22_n_249);
  or mul_108_22_g3613(mul_108_22_n_420 ,mul_108_22_n_346 ,mul_108_22_n_222);
  or mul_108_22_g3614(mul_108_22_n_419 ,mul_108_22_n_390 ,mul_108_22_n_225);
  or mul_108_22_g3615(mul_108_22_n_418 ,mul_108_22_n_391 ,mul_108_22_n_234);
  or mul_108_22_g3616(mul_108_22_n_417 ,mul_108_22_n_342 ,mul_108_22_n_216);
  or mul_108_22_g3617(mul_108_22_n_416 ,mul_108_22_n_397 ,mul_108_22_n_243);
  or mul_108_22_g3618(mul_108_22_n_415 ,mul_108_22_n_326 ,mul_108_22_n_373);
  or mul_108_22_g3619(mul_108_22_n_414 ,mul_108_22_n_407 ,mul_108_22_n_213);
  or mul_108_22_g3620(mul_108_22_n_413 ,mul_108_22_n_339 ,mul_108_22_n_240);
  or mul_108_22_g3621(mul_108_22_n_412 ,mul_108_22_n_362 ,mul_108_22_n_219);
  or mul_108_22_g3622(mul_108_22_n_411 ,mul_108_22_n_409 ,mul_108_22_n_207);
  and mul_108_22_g3623(mul_108_22_n_457 ,in24[7] ,mul_108_22_n_150);
  or mul_108_22_g3624(mul_108_22_n_456 ,mul_108_22_n_159 ,mul_108_22_n_213);
  and mul_108_22_g3625(mul_108_22_n_454 ,in24[3] ,mul_108_22_n_154);
  and mul_108_22_g3626(mul_108_22_n_452 ,in24[5] ,mul_108_22_n_152);
  or mul_108_22_g3627(mul_108_22_n_451 ,mul_108_22_n_163 ,mul_108_22_n_231);
  or mul_108_22_g3628(mul_108_22_n_450 ,mul_108_22_n_162 ,mul_108_22_n_222);
  or mul_108_22_g3629(mul_108_22_n_449 ,mul_108_22_n_162 ,mul_108_22_n_148);
  and mul_108_22_g3630(mul_108_22_n_448 ,in24[8] ,mul_108_22_n_147);
  or mul_108_22_g3631(mul_108_22_n_447 ,mul_108_22_n_371 ,mul_108_22_n_151);
  or mul_108_22_g3632(mul_108_22_n_446 ,in24[0] ,mul_108_22_n_375);
  or mul_108_22_g3633(mul_108_22_n_445 ,mul_108_22_n_329 ,mul_108_22_n_149);
  or mul_108_22_g3634(mul_108_22_n_444 ,mul_108_22_n_372 ,mul_108_22_n_153);
  not mul_108_22_g3635(mul_108_22_n_383 ,mul_108_22_n_152);
  not mul_108_22_g3636(mul_108_22_n_382 ,mul_108_22_n_151);
  not mul_108_22_g3639(mul_108_22_n_380 ,mul_108_22_n_150);
  not mul_108_22_g3640(mul_108_22_n_379 ,mul_108_22_n_149);
  xnor mul_108_22_g3643(mul_108_22_n_377 ,mul_108_22_n_18 ,in24[5]);
  and mul_108_22_g3644(mul_108_22_n_376 ,mul_108_22_n_202 ,mul_108_22_n_322);
  and mul_108_22_g3646(mul_108_22_n_374 ,mul_108_22_n_315 ,mul_108_22_n_319);
  and mul_108_22_g3647(mul_108_22_n_373 ,mul_108_22_n_316 ,mul_108_22_n_323);
  xnor mul_108_22_g3648(mul_108_22_n_372 ,in24[3] ,in24[2]);
  xnor mul_108_22_g3649(mul_108_22_n_371 ,in24[5] ,in24[4]);
  xnor mul_108_22_g3650(mul_108_22_n_370 ,mul_108_22_n_18 ,in24[3]);
  xnor mul_108_22_g3651(mul_108_22_n_410 ,mul_108_22_n_260 ,in24[5]);
  xnor mul_108_22_g3652(mul_108_22_n_409 ,mul_108_22_n_281 ,in24[3]);
  xnor mul_108_22_g3653(mul_108_22_n_408 ,mul_108_22_n_287 ,in24[3]);
  xnor mul_108_22_g3654(mul_108_22_n_407 ,mul_108_22_n_269 ,in24[3]);
  xnor mul_108_22_g3655(mul_108_22_n_406 ,mul_108_22_n_270 ,in24[5]);
  xnor mul_108_22_g3656(mul_108_22_n_405 ,mul_108_22_n_288 ,in24[5]);
  xnor mul_108_22_g3657(mul_108_22_n_404 ,mul_108_22_n_278 ,in24[3]);
  xnor mul_108_22_g3658(mul_108_22_n_403 ,mul_108_22_n_263 ,in24[3]);
  xnor mul_108_22_g3659(mul_108_22_n_402 ,mul_108_22_n_254 ,in24[3]);
  xnor mul_108_22_g3660(mul_108_22_n_401 ,mul_108_22_n_290 ,in24[5]);
  xnor mul_108_22_g3661(mul_108_22_n_400 ,mul_108_22_n_272 ,in24[3]);
  xnor mul_108_22_g3662(mul_108_22_n_399 ,mul_108_22_n_291 ,in24[3]);
  xnor mul_108_22_g3663(mul_108_22_n_398 ,mul_108_22_n_275 ,in24[3]);
  xnor mul_108_22_g3664(mul_108_22_n_397 ,mul_108_22_n_293 ,in24[3]);
  xnor mul_108_22_g3665(mul_108_22_n_396 ,mul_108_22_n_294 ,in24[5]);
  xnor mul_108_22_g3666(mul_108_22_n_395 ,mul_108_22_n_276 ,in24[5]);
  xnor mul_108_22_g3667(mul_108_22_n_394 ,mul_108_22_n_255 ,in24[5]);
  xnor mul_108_22_g3668(mul_108_22_n_393 ,mul_108_22_n_284 ,in24[5]);
  xnor mul_108_22_g3669(mul_108_22_n_392 ,mul_108_22_n_251 ,in24[3]);
  xnor mul_108_22_g3670(mul_108_22_n_391 ,mul_108_22_n_273 ,in24[5]);
  xnor mul_108_22_g3671(mul_108_22_n_390 ,mul_108_22_n_257 ,in24[5]);
  xnor mul_108_22_g3672(mul_108_22_n_389 ,mul_108_22_n_282 ,in24[5]);
  xnor mul_108_22_g3673(mul_108_22_n_388 ,mul_108_22_n_261 ,in24[3]);
  xnor mul_108_22_g3674(mul_108_22_n_387 ,mul_108_22_n_122 ,in24[5]);
  xnor mul_108_22_g3675(mul_108_22_n_386 ,mul_108_22_n_258 ,in24[3]);
  xnor mul_108_22_g3676(mul_108_22_n_385 ,mul_108_22_n_285 ,in24[3]);
  xnor mul_108_22_g3677(mul_108_22_n_384 ,mul_108_22_n_266 ,in24[5]);
  xnor mul_108_22_g3678(mul_108_22_n_381 ,mul_108_22_n_316 ,in24[4]);
  xnor mul_108_22_g3679(mul_108_22_n_378 ,mul_108_22_n_315 ,in24[6]);
  not mul_108_22_g3680(mul_108_22_n_336 ,mul_108_22_n_148);
  not mul_108_22_g3681(mul_108_22_n_335 ,mul_108_22_n_147);
  not mul_108_22_g3684(mul_108_22_n_333 ,mul_108_22_n_154);
  not mul_108_22_g3685(mul_108_22_n_332 ,mul_108_22_n_153);
  xnor mul_108_22_g3689(mul_108_22_n_329 ,in24[7] ,in24[6]);
  xnor mul_108_22_g3690(mul_108_22_n_328 ,mul_108_22_n_168 ,in24[7]);
  xnor mul_108_22_g3691(mul_108_22_n_369 ,mul_108_22_n_98 ,in24[7]);
  xnor mul_108_22_g3692(mul_108_22_n_368 ,mul_108_22_n_100 ,in24[7]);
  xnor mul_108_22_g3693(mul_108_22_n_367 ,mul_108_22_n_264 ,in24[5]);
  xnor mul_108_22_g3694(mul_108_22_n_366 ,mul_108_22_n_112 ,in24[7]);
  xnor mul_108_22_g3695(mul_108_22_n_365 ,mul_108_22_n_114 ,in24[1]);
  xnor mul_108_22_g3696(mul_108_22_n_364 ,mul_108_22_n_251 ,in24[1]);
  xnor mul_108_22_g3697(mul_108_22_n_363 ,mul_108_22_n_279 ,in24[5]);
  xnor mul_108_22_g3698(mul_108_22_n_362 ,mul_108_22_n_146 ,in24[7]);
  xnor mul_108_22_g3699(mul_108_22_n_361 ,mul_108_22_n_124 ,in24[1]);
  xnor mul_108_22_g3700(mul_108_22_n_360 ,mul_108_22_n_102 ,in24[1]);
  xnor mul_108_22_g3701(mul_108_22_n_359 ,mul_108_22_n_124 ,in24[7]);
  xnor mul_108_22_g3702(mul_108_22_n_358 ,mul_108_22_n_114 ,in24[7]);
  xnor mul_108_22_g3703(mul_108_22_n_357 ,mul_108_22_n_98 ,in24[1]);
  xnor mul_108_22_g3704(mul_108_22_n_356 ,mul_108_22_n_118 ,in24[7]);
  xnor mul_108_22_g3705(mul_108_22_n_355 ,mul_108_22_n_108 ,in24[1]);
  xnor mul_108_22_g3706(mul_108_22_n_354 ,mul_108_22_n_108 ,in24[7]);
  xnor mul_108_22_g3707(mul_108_22_n_353 ,mul_108_22_n_106 ,in24[1]);
  xnor mul_108_22_g3708(mul_108_22_n_352 ,mul_108_22_n_96 ,in24[1]);
  xnor mul_108_22_g3709(mul_108_22_n_351 ,mul_108_22_n_118 ,in24[1]);
  xnor mul_108_22_g3710(mul_108_22_n_350 ,mul_108_22_n_104 ,in24[1]);
  xnor mul_108_22_g3711(mul_108_22_n_349 ,mul_108_22_n_116 ,in24[7]);
  xnor mul_108_22_g3712(mul_108_22_n_348 ,mul_108_22_n_146 ,in24[1]);
  xnor mul_108_22_g3713(mul_108_22_n_347 ,mul_108_22_n_267 ,in24[1]);
  xnor mul_108_22_g3714(mul_108_22_n_346 ,mul_108_22_n_122 ,in24[7]);
  xnor mul_108_22_g3715(mul_108_22_n_345 ,mul_108_22_n_130 ,in24[7]);
  xnor mul_108_22_g3716(mul_108_22_n_344 ,mul_108_22_n_104 ,in24[7]);
  xnor mul_108_22_g3717(mul_108_22_n_343 ,mul_108_22_n_102 ,in24[7]);
  xnor mul_108_22_g3718(mul_108_22_n_342 ,mul_108_22_n_96 ,in24[7]);
  xnor mul_108_22_g3719(mul_108_22_n_341 ,mul_108_22_n_106 ,in24[7]);
  xnor mul_108_22_g3720(mul_108_22_n_340 ,mul_108_22_n_116 ,in24[1]);
  xnor mul_108_22_g3721(mul_108_22_n_339 ,mul_108_22_n_130 ,in24[3]);
  xnor mul_108_22_g3722(mul_108_22_n_338 ,mul_108_22_n_112 ,in24[1]);
  xnor mul_108_22_g3723(mul_108_22_n_337 ,mul_108_22_n_100 ,in24[1]);
  xnor mul_108_22_g3724(mul_108_22_n_334 ,in24[8] ,in24[7]);
  xnor mul_108_22_g3725(mul_108_22_n_331 ,mul_108_22_n_202 ,in24[2]);
  nor mul_108_22_g3726(mul_108_22_n_327 ,mul_108_22_n_70 ,mul_108_22_n_163);
  nor mul_108_22_g3727(mul_108_22_n_326 ,mul_108_22_n_166 ,in24[4]);
  not mul_108_22_g3728(mul_108_22_n_325 ,mul_108_22_n_324);
  and mul_108_22_g3729(mul_108_22_n_324 ,in24[1] ,in24[0]);
  or mul_108_22_g3730(mul_108_22_n_323 ,mul_108_22_n_159 ,mul_108_22_n_313);
  or mul_108_22_g3731(mul_108_22_n_322 ,mul_108_22_n_160 ,mul_108_22_n_318);
  nor mul_108_22_g3732(mul_108_22_n_321 ,mul_108_22_n_19 ,in24[2]);
  nor mul_108_22_g3733(mul_108_22_n_320 ,mul_108_22_n_168 ,in24[6]);
  or mul_108_22_g3734(mul_108_22_n_319 ,mul_108_22_n_160 ,mul_108_22_n_314);
  not mul_108_22_g3735(mul_108_22_n_318 ,in24[2]);
  not mul_108_22_g3736(mul_108_22_n_317 ,in24[0]);
  not mul_108_22_g3737(mul_108_22_n_316 ,in24[3]);
  not mul_108_22_g3738(mul_108_22_n_315 ,in24[5]);
  not mul_108_22_g3739(mul_108_22_n_314 ,in24[6]);
  not mul_108_22_g3740(mul_108_22_n_313 ,in24[4]);
  not mul_108_22_g3741(mul_108_22_n_312 ,mul_108_22_n_165);
  not mul_108_22_g3742(mul_108_22_n_311 ,in24[1]);
  not mul_108_22_g3743(mul_108_22_n_310 ,in24[7]);
  not mul_108_22_drc_bufs3784(mul_108_22_n_297 ,mul_108_22_n_295);
  not mul_108_22_drc_bufs3785(mul_108_22_n_296 ,mul_108_22_n_295);
  not mul_108_22_drc_bufs3786(mul_108_22_n_295 ,n_255);
  not mul_108_22_drc_bufs3814(mul_108_22_n_294 ,mul_108_22_n_292);
  not mul_108_22_drc_bufs3815(mul_108_22_n_293 ,mul_108_22_n_292);
  not mul_108_22_drc_bufs3816(mul_108_22_n_292 ,n_258);
  not mul_108_22_drc_bufs3818(mul_108_22_n_291 ,mul_108_22_n_289);
  not mul_108_22_drc_bufs3819(mul_108_22_n_290 ,mul_108_22_n_289);
  not mul_108_22_drc_bufs3820(mul_108_22_n_289 ,n_256);
  not mul_108_22_drc_bufs3822(mul_108_22_n_288 ,mul_108_22_n_286);
  not mul_108_22_drc_bufs3823(mul_108_22_n_287 ,mul_108_22_n_286);
  not mul_108_22_drc_bufs3824(mul_108_22_n_286 ,n_262);
  not mul_108_22_drc_bufs3826(mul_108_22_n_285 ,mul_108_22_n_283);
  not mul_108_22_drc_bufs3827(mul_108_22_n_284 ,mul_108_22_n_283);
  not mul_108_22_drc_bufs3828(mul_108_22_n_283 ,n_263);
  not mul_108_22_drc_bufs3830(mul_108_22_n_282 ,mul_108_22_n_280);
  not mul_108_22_drc_bufs3831(mul_108_22_n_281 ,mul_108_22_n_280);
  not mul_108_22_drc_bufs3832(mul_108_22_n_280 ,n_259);
  not mul_108_22_drc_bufs3834(mul_108_22_n_279 ,mul_108_22_n_277);
  not mul_108_22_drc_bufs3835(mul_108_22_n_278 ,mul_108_22_n_277);
  not mul_108_22_drc_bufs3836(mul_108_22_n_277 ,n_264);
  not mul_108_22_drc_bufs3838(mul_108_22_n_276 ,mul_108_22_n_274);
  not mul_108_22_drc_bufs3839(mul_108_22_n_275 ,mul_108_22_n_274);
  not mul_108_22_drc_bufs3840(mul_108_22_n_274 ,n_265);
  not mul_108_22_drc_bufs3842(mul_108_22_n_273 ,mul_108_22_n_271);
  not mul_108_22_drc_bufs3843(mul_108_22_n_272 ,mul_108_22_n_271);
  not mul_108_22_drc_bufs3844(mul_108_22_n_271 ,n_260);
  not mul_108_22_drc_bufs3846(mul_108_22_n_270 ,mul_108_22_n_268);
  not mul_108_22_drc_bufs3847(mul_108_22_n_269 ,mul_108_22_n_268);
  not mul_108_22_drc_bufs3848(mul_108_22_n_268 ,n_266);
  not mul_108_22_drc_bufs3850(mul_108_22_n_267 ,mul_108_22_n_265);
  not mul_108_22_drc_bufs3851(mul_108_22_n_266 ,mul_108_22_n_265);
  not mul_108_22_drc_bufs3852(mul_108_22_n_265 ,n_257);
  not mul_108_22_drc_bufs3854(mul_108_22_n_264 ,mul_108_22_n_262);
  not mul_108_22_drc_bufs3855(mul_108_22_n_263 ,mul_108_22_n_262);
  not mul_108_22_drc_bufs3856(mul_108_22_n_262 ,n_267);
  not mul_108_22_drc_bufs3858(mul_108_22_n_261 ,mul_108_22_n_259);
  not mul_108_22_drc_bufs3859(mul_108_22_n_260 ,mul_108_22_n_259);
  not mul_108_22_drc_bufs3860(mul_108_22_n_259 ,n_261);
  not mul_108_22_drc_bufs3862(mul_108_22_n_258 ,mul_108_22_n_256);
  not mul_108_22_drc_bufs3863(mul_108_22_n_257 ,mul_108_22_n_256);
  not mul_108_22_drc_bufs3864(mul_108_22_n_256 ,n_268);
  not mul_108_22_drc_bufs3866(mul_108_22_n_255 ,mul_108_22_n_253);
  not mul_108_22_drc_bufs3867(mul_108_22_n_254 ,mul_108_22_n_253);
  not mul_108_22_drc_bufs3868(mul_108_22_n_253 ,n_269);
  not mul_108_22_drc_bufs3870(mul_108_22_n_252 ,mul_108_22_n_250);
  not mul_108_22_drc_bufs3871(mul_108_22_n_251 ,mul_108_22_n_250);
  not mul_108_22_drc_bufs3872(mul_108_22_n_250 ,n_270);
  not mul_108_22_drc_bufs3874(mul_108_22_n_249 ,mul_108_22_n_247);
  not mul_108_22_drc_bufs3875(mul_108_22_n_248 ,mul_108_22_n_247);
  not mul_108_22_drc_bufs3876(mul_108_22_n_247 ,mul_108_22_n_303);
  not mul_108_22_drc_bufs3878(mul_108_22_n_246 ,mul_108_22_n_244);
  not mul_108_22_drc_bufs3879(mul_108_22_n_245 ,mul_108_22_n_244);
  not mul_108_22_drc_bufs3880(mul_108_22_n_244 ,mul_108_22_n_335);
  not mul_108_22_drc_bufs3882(mul_108_22_n_243 ,mul_108_22_n_241);
  not mul_108_22_drc_bufs3883(mul_108_22_n_242 ,mul_108_22_n_241);
  not mul_108_22_drc_bufs3884(mul_108_22_n_241 ,mul_108_22_n_299);
  not mul_108_22_drc_bufs3886(mul_108_22_n_240 ,mul_108_22_n_238);
  not mul_108_22_drc_bufs3887(mul_108_22_n_239 ,mul_108_22_n_238);
  not mul_108_22_drc_bufs3888(mul_108_22_n_238 ,mul_108_22_n_298);
  not mul_108_22_drc_bufs3890(mul_108_22_n_237 ,mul_108_22_n_235);
  not mul_108_22_drc_bufs3891(mul_108_22_n_236 ,mul_108_22_n_235);
  not mul_108_22_drc_bufs3892(mul_108_22_n_235 ,mul_108_22_n_336);
  not mul_108_22_drc_bufs3894(mul_108_22_n_234 ,mul_108_22_n_232);
  not mul_108_22_drc_bufs3895(mul_108_22_n_233 ,mul_108_22_n_232);
  not mul_108_22_drc_bufs3896(mul_108_22_n_232 ,mul_108_22_n_383);
  not mul_108_22_drc_bufs3898(mul_108_22_n_231 ,mul_108_22_n_229);
  not mul_108_22_drc_bufs3899(mul_108_22_n_230 ,mul_108_22_n_229);
  not mul_108_22_drc_bufs3900(mul_108_22_n_229 ,mul_108_22_n_382);
  not mul_108_22_drc_bufs3902(mul_108_22_n_228 ,mul_108_22_n_226);
  not mul_108_22_drc_bufs3903(mul_108_22_n_227 ,mul_108_22_n_226);
  not mul_108_22_drc_bufs3904(mul_108_22_n_226 ,mul_108_22_n_305);
  not mul_108_22_drc_bufs3906(mul_108_22_n_225 ,mul_108_22_n_223);
  not mul_108_22_drc_bufs3907(mul_108_22_n_224 ,mul_108_22_n_223);
  not mul_108_22_drc_bufs3908(mul_108_22_n_223 ,mul_108_22_n_304);
  not mul_108_22_drc_bufs3910(mul_108_22_n_222 ,mul_108_22_n_220);
  not mul_108_22_drc_bufs3911(mul_108_22_n_221 ,mul_108_22_n_220);
  not mul_108_22_drc_bufs3912(mul_108_22_n_220 ,mul_108_22_n_379);
  not mul_108_22_drc_bufs3914(mul_108_22_n_219 ,mul_108_22_n_217);
  not mul_108_22_drc_bufs3915(mul_108_22_n_218 ,mul_108_22_n_217);
  not mul_108_22_drc_bufs3916(mul_108_22_n_217 ,mul_108_22_n_380);
  not mul_108_22_drc_bufs3918(mul_108_22_n_216 ,mul_108_22_n_214);
  not mul_108_22_drc_bufs3919(mul_108_22_n_215 ,mul_108_22_n_214);
  not mul_108_22_drc_bufs3920(mul_108_22_n_214 ,mul_108_22_n_302);
  not mul_108_22_drc_bufs3922(mul_108_22_n_213 ,mul_108_22_n_211);
  not mul_108_22_drc_bufs3923(mul_108_22_n_212 ,mul_108_22_n_211);
  not mul_108_22_drc_bufs3924(mul_108_22_n_211 ,mul_108_22_n_332);
  not mul_108_22_drc_bufs3926(mul_108_22_n_210 ,mul_108_22_n_208);
  not mul_108_22_drc_bufs3927(mul_108_22_n_209 ,mul_108_22_n_208);
  not mul_108_22_drc_bufs3928(mul_108_22_n_208 ,mul_108_22_n_300);
  not mul_108_22_drc_bufs3930(mul_108_22_n_207 ,mul_108_22_n_205);
  not mul_108_22_drc_bufs3931(mul_108_22_n_206 ,mul_108_22_n_205);
  not mul_108_22_drc_bufs3932(mul_108_22_n_205 ,mul_108_22_n_333);
  not mul_108_22_drc_bufs3934(mul_108_22_n_204 ,mul_108_22_n_649);
  not mul_108_22_drc_bufs3935(mul_108_22_n_203 ,mul_108_22_n_649);
  not mul_108_22_drc_bufs3940(mul_108_22_n_307 ,mul_108_22_n_650);
  not mul_108_22_drc_bufs3943(mul_108_22_n_202 ,mul_108_22_n_201);
  not mul_108_22_drc_bufs3944(mul_108_22_n_201 ,mul_108_22_n_311);
  not mul_108_22_drc_bufs3946(mul_108_22_n_200 ,mul_108_22_n_198);
  not mul_108_22_drc_bufs3947(mul_108_22_n_199 ,mul_108_22_n_198);
  not mul_108_22_drc_bufs3948(mul_108_22_n_198 ,mul_108_22_n_301);
  buf mul_108_22_drc_bufs3957(n_248 ,mul_108_22_n_1140);
  buf mul_108_22_drc_bufs3958(n_249 ,mul_108_22_n_1143);
  buf mul_108_22_drc_bufs3959(n_242 ,mul_108_22_n_1121);
  buf mul_108_22_drc_bufs3960(n_244 ,mul_108_22_n_1127);
  buf mul_108_22_drc_bufs3961(n_245 ,mul_108_22_n_1130);
  buf mul_108_22_drc_bufs3962(n_252 ,mul_108_22_n_1153);
  buf mul_108_22_drc_bufs3963(n_247 ,mul_108_22_n_1137);
  buf mul_108_22_drc_bufs3964(n_246 ,mul_108_22_n_1134);
  buf mul_108_22_drc_bufs3965(n_243 ,mul_108_22_n_1124);
  buf mul_108_22_drc_bufs3966(n_253 ,mul_108_22_n_1156);
  buf mul_108_22_drc_bufs3967(n_250 ,mul_108_22_n_1147);
  buf mul_108_22_drc_bufs3968(n_251 ,mul_108_22_n_1150);
  buf mul_108_22_drc_bufs3969(n_239 ,mul_108_22_n_1112);
  buf mul_108_22_drc_bufs3970(n_240 ,mul_108_22_n_1115);
  buf mul_108_22_drc_bufs3971(n_241 ,mul_108_22_n_1118);
  not mul_108_22_drc_bufs3973(mul_108_22_n_182 ,mul_108_22_n_308);
  not mul_108_22_drc_bufs3974(mul_108_22_n_308 ,mul_108_22_n_885);
  not mul_108_22_drc_bufs3996(mul_108_22_n_181 ,mul_108_22_n_180);
  not mul_108_22_drc_bufs3998(mul_108_22_n_180 ,mul_108_22_n_446);
  not mul_108_22_drc_bufs4001(mul_108_22_n_179 ,mul_108_22_n_178);
  not mul_108_22_drc_bufs4003(mul_108_22_n_178 ,mul_108_22_n_444);
  not mul_108_22_drc_bufs4006(mul_108_22_n_177 ,mul_108_22_n_176);
  not mul_108_22_drc_bufs4008(mul_108_22_n_176 ,mul_108_22_n_447);
  not mul_108_22_drc_bufs4011(mul_108_22_n_175 ,mul_108_22_n_174);
  not mul_108_22_drc_bufs4013(mul_108_22_n_174 ,mul_108_22_n_445);
  not mul_108_22_drc_bufs4021(mul_108_22_n_173 ,mul_108_22_n_172);
  not mul_108_22_drc_bufs4023(mul_108_22_n_172 ,mul_108_22_n_317);
  not mul_108_22_drc_bufs4031(mul_108_22_n_171 ,mul_108_22_n_169);
  not mul_108_22_drc_bufs4032(mul_108_22_n_170 ,mul_108_22_n_169);
  not mul_108_22_drc_bufs4033(mul_108_22_n_169 ,mul_108_22_n_448);
  not mul_108_22_drc_bufs4036(mul_108_22_n_168 ,mul_108_22_n_167);
  not mul_108_22_drc_bufs4037(mul_108_22_n_167 ,mul_108_22_n_297);
  not mul_108_22_drc_bufs4039(mul_108_22_n_166 ,mul_108_22_n_164);
  not mul_108_22_drc_bufs4040(mul_108_22_n_165 ,mul_108_22_n_164);
  not mul_108_22_drc_bufs4041(mul_108_22_n_164 ,mul_108_22_n_296);
  not mul_108_22_drc_bufs4043(mul_108_22_n_163 ,mul_108_22_n_161);
  not mul_108_22_drc_bufs4044(mul_108_22_n_162 ,mul_108_22_n_161);
  not mul_108_22_drc_bufs4045(mul_108_22_n_161 ,mul_108_22_n_312);
  not mul_108_22_drc_bufs4047(mul_108_22_n_160 ,mul_108_22_n_158);
  not mul_108_22_drc_bufs4048(mul_108_22_n_159 ,mul_108_22_n_158);
  not mul_108_22_drc_bufs4049(mul_108_22_n_158 ,mul_108_22_n_312);
  not mul_108_22_drc_bufs4051(mul_108_22_n_157 ,mul_108_22_n_306);
  not mul_108_22_drc_bufs4053(mul_108_22_n_306 ,mul_108_22_n_648);
  not mul_108_22_drc_bufs4056(mul_108_22_n_156 ,mul_108_22_n_155);
  not mul_108_22_drc_bufs4057(mul_108_22_n_155 ,mul_108_22_n_648);
  not mul_108_22_drc_bufs4059(mul_108_22_n_154 ,mul_108_22_n_299);
  not mul_108_22_drc_bufs4061(mul_108_22_n_299 ,mul_108_22_n_331);
  not mul_108_22_drc_bufs4063(mul_108_22_n_153 ,mul_108_22_n_298);
  not mul_108_22_drc_bufs4065(mul_108_22_n_298 ,mul_108_22_n_331);
  not mul_108_22_drc_bufs4067(mul_108_22_n_152 ,mul_108_22_n_305);
  not mul_108_22_drc_bufs4069(mul_108_22_n_305 ,mul_108_22_n_381);
  not mul_108_22_drc_bufs4071(mul_108_22_n_151 ,mul_108_22_n_304);
  not mul_108_22_drc_bufs4073(mul_108_22_n_304 ,mul_108_22_n_381);
  not mul_108_22_drc_bufs4075(mul_108_22_n_150 ,mul_108_22_n_303);
  not mul_108_22_drc_bufs4077(mul_108_22_n_303 ,mul_108_22_n_378);
  not mul_108_22_drc_bufs4079(mul_108_22_n_149 ,mul_108_22_n_302);
  not mul_108_22_drc_bufs4081(mul_108_22_n_302 ,mul_108_22_n_378);
  not mul_108_22_drc_bufs4083(mul_108_22_n_148 ,mul_108_22_n_301);
  not mul_108_22_drc_bufs4085(mul_108_22_n_301 ,mul_108_22_n_334);
  not mul_108_22_drc_bufs4087(mul_108_22_n_147 ,mul_108_22_n_300);
  not mul_108_22_drc_bufs4089(mul_108_22_n_300 ,mul_108_22_n_334);
  not mul_108_22_drc_bufs4091(mul_108_22_n_146 ,mul_108_22_n_145);
  not mul_108_22_drc_bufs4093(mul_108_22_n_145 ,mul_108_22_n_281);
  not mul_108_22_drc_bufs4095(mul_108_22_n_144 ,mul_108_22_n_143);
  not mul_108_22_drc_bufs4097(mul_108_22_n_143 ,mul_108_22_n_291);
  not mul_108_22_drc_bufs4099(mul_108_22_n_142 ,mul_108_22_n_141);
  not mul_108_22_drc_bufs4101(mul_108_22_n_141 ,mul_108_22_n_273);
  not mul_108_22_drc_bufs4103(mul_108_22_n_140 ,mul_108_22_n_139);
  not mul_108_22_drc_bufs4105(mul_108_22_n_139 ,mul_108_22_n_294);
  not mul_108_22_drc_bufs4107(mul_108_22_n_138 ,mul_108_22_n_137);
  not mul_108_22_drc_bufs4109(mul_108_22_n_137 ,mul_108_22_n_255);
  not mul_108_22_drc_bufs4111(mul_108_22_n_136 ,mul_108_22_n_135);
  not mul_108_22_drc_bufs4113(mul_108_22_n_135 ,mul_108_22_n_282);
  not mul_108_22_drc_bufs4115(mul_108_22_n_134 ,mul_108_22_n_133);
  not mul_108_22_drc_bufs4117(mul_108_22_n_133 ,mul_108_22_n_261);
  not mul_108_22_drc_bufs4119(mul_108_22_n_132 ,mul_108_22_n_131);
  not mul_108_22_drc_bufs4121(mul_108_22_n_131 ,mul_108_22_n_264);
  not mul_108_22_drc_bufs4123(mul_108_22_n_130 ,mul_108_22_n_129);
  not mul_108_22_drc_bufs4125(mul_108_22_n_129 ,mul_108_22_n_266);
  not mul_108_22_drc_bufs4127(mul_108_22_n_128 ,mul_108_22_n_127);
  not mul_108_22_drc_bufs4129(mul_108_22_n_127 ,mul_108_22_n_276);
  not mul_108_22_drc_bufs4131(mul_108_22_n_126 ,mul_108_22_n_125);
  not mul_108_22_drc_bufs4133(mul_108_22_n_125 ,mul_108_22_n_258);
  not mul_108_22_drc_bufs4135(mul_108_22_n_124 ,mul_108_22_n_123);
  not mul_108_22_drc_bufs4137(mul_108_22_n_123 ,mul_108_22_n_260);
  not mul_108_22_drc_bufs4139(mul_108_22_n_122 ,mul_108_22_n_121);
  not mul_108_22_drc_bufs4141(mul_108_22_n_121 ,mul_108_22_n_252);
  not mul_108_22_drc_bufs4143(mul_108_22_n_120 ,mul_108_22_n_119);
  not mul_108_22_drc_bufs4145(mul_108_22_n_119 ,mul_108_22_n_270);
  not mul_108_22_drc_bufs4147(mul_108_22_n_118 ,mul_108_22_n_117);
  not mul_108_22_drc_bufs4149(mul_108_22_n_117 ,mul_108_22_n_254);
  not mul_108_22_drc_bufs4151(mul_108_22_n_116 ,mul_108_22_n_115);
  not mul_108_22_drc_bufs4153(mul_108_22_n_115 ,mul_108_22_n_263);
  not mul_108_22_drc_bufs4155(mul_108_22_n_114 ,mul_108_22_n_113);
  not mul_108_22_drc_bufs4157(mul_108_22_n_113 ,mul_108_22_n_290);
  not mul_108_22_drc_bufs4159(mul_108_22_n_112 ,mul_108_22_n_111);
  not mul_108_22_drc_bufs4161(mul_108_22_n_111 ,mul_108_22_n_293);
  not mul_108_22_drc_bufs4163(mul_108_22_n_110 ,mul_108_22_n_109);
  not mul_108_22_drc_bufs4165(mul_108_22_n_109 ,mul_108_22_n_267);
  not mul_108_22_drc_bufs4167(mul_108_22_n_108 ,mul_108_22_n_107);
  not mul_108_22_drc_bufs4169(mul_108_22_n_107 ,mul_108_22_n_284);
  not mul_108_22_drc_bufs4171(mul_108_22_n_106 ,mul_108_22_n_105);
  not mul_108_22_drc_bufs4173(mul_108_22_n_105 ,mul_108_22_n_269);
  not mul_108_22_drc_bufs4175(mul_108_22_n_104 ,mul_108_22_n_103);
  not mul_108_22_drc_bufs4177(mul_108_22_n_103 ,mul_108_22_n_278);
  not mul_108_22_drc_bufs4179(mul_108_22_n_102 ,mul_108_22_n_101);
  not mul_108_22_drc_bufs4181(mul_108_22_n_101 ,mul_108_22_n_275);
  not mul_108_22_drc_bufs4183(mul_108_22_n_100 ,mul_108_22_n_99);
  not mul_108_22_drc_bufs4185(mul_108_22_n_99 ,mul_108_22_n_257);
  not mul_108_22_drc_bufs4187(mul_108_22_n_98 ,mul_108_22_n_97);
  not mul_108_22_drc_bufs4189(mul_108_22_n_97 ,mul_108_22_n_272);
  not mul_108_22_drc_bufs4191(mul_108_22_n_96 ,mul_108_22_n_95);
  not mul_108_22_drc_bufs4193(mul_108_22_n_95 ,mul_108_22_n_287);
  not mul_108_22_drc_bufs4195(mul_108_22_n_94 ,mul_108_22_n_93);
  not mul_108_22_drc_bufs4197(mul_108_22_n_93 ,mul_108_22_n_285);
  not mul_108_22_drc_bufs4199(mul_108_22_n_92 ,mul_108_22_n_91);
  not mul_108_22_drc_bufs4201(mul_108_22_n_91 ,mul_108_22_n_279);
  not mul_108_22_drc_bufs4203(mul_108_22_n_90 ,mul_108_22_n_89);
  not mul_108_22_drc_bufs4205(mul_108_22_n_89 ,mul_108_22_n_288);
  not mul_108_22_drc_bufs4207(mul_108_22_n_88 ,mul_108_22_n_86);
  not mul_108_22_drc_bufs4208(mul_108_22_n_87 ,mul_108_22_n_86);
  not mul_108_22_drc_bufs4209(mul_108_22_n_86 ,mul_108_22_n_446);
  not mul_108_22_drc_bufs4211(mul_108_22_n_85 ,mul_108_22_n_83);
  not mul_108_22_drc_bufs4212(mul_108_22_n_84 ,mul_108_22_n_83);
  not mul_108_22_drc_bufs4213(mul_108_22_n_83 ,mul_108_22_n_444);
  not mul_108_22_drc_bufs4215(mul_108_22_n_82 ,mul_108_22_n_80);
  not mul_108_22_drc_bufs4216(mul_108_22_n_81 ,mul_108_22_n_80);
  not mul_108_22_drc_bufs4217(mul_108_22_n_80 ,mul_108_22_n_445);
  not mul_108_22_drc_bufs4219(mul_108_22_n_79 ,mul_108_22_n_77);
  not mul_108_22_drc_bufs4220(mul_108_22_n_78 ,mul_108_22_n_77);
  not mul_108_22_drc_bufs4221(mul_108_22_n_77 ,mul_108_22_n_447);
  not mul_108_22_drc_bufs4223(mul_108_22_n_76 ,mul_108_22_n_74);
  not mul_108_22_drc_bufs4224(mul_108_22_n_75 ,mul_108_22_n_74);
  not mul_108_22_drc_bufs4225(mul_108_22_n_74 ,mul_108_22_n_181);
  not mul_108_22_drc_bufs4227(mul_108_22_n_73 ,mul_108_22_n_71);
  not mul_108_22_drc_bufs4228(mul_108_22_n_72 ,mul_108_22_n_71);
  not mul_108_22_drc_bufs4229(mul_108_22_n_71 ,mul_108_22_n_317);
  not mul_108_22_drc_bufs4231(mul_108_22_n_70 ,mul_108_22_n_68);
  not mul_108_22_drc_bufs4232(mul_108_22_n_69 ,mul_108_22_n_68);
  not mul_108_22_drc_bufs4233(mul_108_22_n_68 ,mul_108_22_n_173);
  not mul_108_22_drc_bufs4235(mul_108_22_n_67 ,mul_108_22_n_65);
  not mul_108_22_drc_bufs4236(mul_108_22_n_66 ,mul_108_22_n_65);
  not mul_108_22_drc_bufs4237(mul_108_22_n_65 ,mul_108_22_n_446);
  not mul_108_22_drc_bufs4239(mul_108_22_n_64 ,mul_108_22_n_62);
  not mul_108_22_drc_bufs4240(mul_108_22_n_63 ,mul_108_22_n_62);
  not mul_108_22_drc_bufs4241(mul_108_22_n_62 ,mul_108_22_n_179);
  not mul_108_22_drc_bufs4243(mul_108_22_n_61 ,mul_108_22_n_59);
  not mul_108_22_drc_bufs4244(mul_108_22_n_60 ,mul_108_22_n_59);
  not mul_108_22_drc_bufs4245(mul_108_22_n_59 ,mul_108_22_n_177);
  not mul_108_22_drc_bufs4247(mul_108_22_n_58 ,mul_108_22_n_56);
  not mul_108_22_drc_bufs4248(mul_108_22_n_57 ,mul_108_22_n_56);
  not mul_108_22_drc_bufs4249(mul_108_22_n_56 ,mul_108_22_n_175);
  not mul_108_22_drc_bufs4251(mul_108_22_n_55 ,mul_108_22_n_53);
  not mul_108_22_drc_bufs4252(mul_108_22_n_54 ,mul_108_22_n_53);
  not mul_108_22_drc_bufs4253(mul_108_22_n_53 ,mul_108_22_n_317);
  not mul_108_22_drc_bufs4255(mul_108_22_n_52 ,mul_108_22_n_50);
  not mul_108_22_drc_bufs4256(mul_108_22_n_51 ,mul_108_22_n_50);
  not mul_108_22_drc_bufs4257(mul_108_22_n_50 ,mul_108_22_n_177);
  not mul_108_22_drc_bufs4259(mul_108_22_n_49 ,mul_108_22_n_47);
  not mul_108_22_drc_bufs4260(mul_108_22_n_48 ,mul_108_22_n_47);
  not mul_108_22_drc_bufs4261(mul_108_22_n_47 ,mul_108_22_n_444);
  not mul_108_22_drc_bufs4263(mul_108_22_n_46 ,mul_108_22_n_44);
  not mul_108_22_drc_bufs4264(mul_108_22_n_45 ,mul_108_22_n_44);
  not mul_108_22_drc_bufs4265(mul_108_22_n_44 ,mul_108_22_n_448);
  not mul_108_22_drc_bufs4267(mul_108_22_n_43 ,mul_108_22_n_41);
  not mul_108_22_drc_bufs4268(mul_108_22_n_42 ,mul_108_22_n_41);
  not mul_108_22_drc_bufs4269(mul_108_22_n_41 ,mul_108_22_n_173);
  not mul_108_22_drc_bufs4271(mul_108_22_n_40 ,mul_108_22_n_38);
  not mul_108_22_drc_bufs4272(mul_108_22_n_39 ,mul_108_22_n_38);
  not mul_108_22_drc_bufs4273(mul_108_22_n_38 ,mul_108_22_n_181);
  not mul_108_22_drc_bufs4275(mul_108_22_n_37 ,mul_108_22_n_35);
  not mul_108_22_drc_bufs4276(mul_108_22_n_36 ,mul_108_22_n_35);
  not mul_108_22_drc_bufs4277(mul_108_22_n_35 ,mul_108_22_n_175);
  not mul_108_22_drc_bufs4279(mul_108_22_n_34 ,mul_108_22_n_32);
  not mul_108_22_drc_bufs4280(mul_108_22_n_33 ,mul_108_22_n_32);
  not mul_108_22_drc_bufs4281(mul_108_22_n_32 ,mul_108_22_n_448);
  not mul_108_22_drc_bufs4283(mul_108_22_n_31 ,mul_108_22_n_29);
  not mul_108_22_drc_bufs4284(mul_108_22_n_30 ,mul_108_22_n_29);
  not mul_108_22_drc_bufs4285(mul_108_22_n_29 ,mul_108_22_n_447);
  not mul_108_22_drc_bufs4287(mul_108_22_n_28 ,mul_108_22_n_26);
  not mul_108_22_drc_bufs4288(mul_108_22_n_27 ,mul_108_22_n_26);
  not mul_108_22_drc_bufs4289(mul_108_22_n_26 ,mul_108_22_n_179);
  not mul_108_22_drc_bufs4291(mul_108_22_n_25 ,mul_108_22_n_23);
  not mul_108_22_drc_bufs4292(mul_108_22_n_24 ,mul_108_22_n_23);
  not mul_108_22_drc_bufs4293(mul_108_22_n_23 ,mul_108_22_n_445);
  not mul_108_22_drc_bufs4295(mul_108_22_n_22 ,mul_108_22_n_20);
  not mul_108_22_drc_bufs4296(mul_108_22_n_21 ,mul_108_22_n_20);
  not mul_108_22_drc_bufs4297(mul_108_22_n_20 ,mul_108_22_n_171);
  not mul_108_22_drc_bufs4299(mul_108_22_n_19 ,mul_108_22_n_17);
  not mul_108_22_drc_bufs4300(mul_108_22_n_18 ,mul_108_22_n_17);
  not mul_108_22_drc_bufs4301(mul_108_22_n_17 ,mul_108_22_n_297);
  not mul_108_22_drc_bufs4303(mul_108_22_n_16 ,mul_108_22_n_15);
  not mul_108_22_drc_bufs4305(mul_108_22_n_15 ,mul_108_22_n_170);
  not mul_108_22_drc_bufs4307(mul_108_22_n_14 ,mul_108_22_n_13);
  not mul_108_22_drc_bufs4309(mul_108_22_n_13 ,mul_108_22_n_88);
  not mul_108_22_drc_bufs4311(mul_108_22_n_12 ,mul_108_22_n_11);
  not mul_108_22_drc_bufs4313(mul_108_22_n_11 ,mul_108_22_n_79);
  not mul_108_22_drc_bufs4315(mul_108_22_n_10 ,mul_108_22_n_9);
  not mul_108_22_drc_bufs4317(mul_108_22_n_9 ,mul_108_22_n_82);
  not mul_108_22_drc_bufs4319(mul_108_22_n_8 ,mul_108_22_n_7);
  not mul_108_22_drc_bufs4321(mul_108_22_n_7 ,mul_108_22_n_85);
  and mul_108_22_g2(mul_108_22_n_6 ,mul_108_22_n_982 ,mul_108_22_n_996);
  and mul_108_22_g4323(mul_108_22_n_5 ,mul_108_22_n_913 ,mul_108_22_n_966);
  xor mul_108_22_g4324(mul_108_22_n_4 ,mul_108_22_n_882 ,mul_108_22_n_963);
  xor mul_108_22_g4325(mul_108_22_n_3 ,mul_108_22_n_889 ,mul_108_22_n_960);
  xor mul_108_22_g4326(mul_108_22_n_2 ,mul_108_22_n_890 ,mul_108_22_n_930);
  xor mul_108_22_g4327(mul_108_22_n_1 ,mul_108_22_n_599 ,mul_108_22_n_847);
  xor mul_108_22_g4328(mul_108_22_n_0 ,mul_108_22_n_801 ,mul_108_22_n_307);
  or mul_113_23_g1494(mul_113_23_n_664 ,mul_113_23_n_476 ,mul_113_23_n_662);
  xnor mul_113_23_g1495(n_338 ,mul_113_23_n_661 ,mul_113_23_n_490);
  and mul_113_23_g1496(mul_113_23_n_662 ,mul_113_23_n_474 ,mul_113_23_n_661);
  and mul_113_23_g1497(mul_113_23_n_661 ,mul_113_23_n_533 ,mul_113_23_n_659);
  xnor mul_113_23_g1498(mul_113_23_n_660 ,mul_113_23_n_657 ,mul_113_23_n_547);
  or mul_113_23_g1499(mul_113_23_n_659 ,mul_113_23_n_541 ,mul_113_23_n_658);
  not mul_113_23_g1500(mul_113_23_n_658 ,mul_113_23_n_657);
  or mul_113_23_g1501(mul_113_23_n_657 ,mul_113_23_n_560 ,mul_113_23_n_655);
  xnor mul_113_23_g1502(mul_113_23_n_656 ,mul_113_23_n_654 ,mul_113_23_n_572);
  and mul_113_23_g1503(mul_113_23_n_655 ,mul_113_23_n_548 ,mul_113_23_n_654);
  or mul_113_23_g1504(mul_113_23_n_654 ,mul_113_23_n_586 ,mul_113_23_n_652);
  xnor mul_113_23_g1505(mul_113_23_n_653 ,mul_113_23_n_651 ,mul_113_23_n_595);
  and mul_113_23_g1506(mul_113_23_n_652 ,mul_113_23_n_589 ,mul_113_23_n_651);
  or mul_113_23_g1507(mul_113_23_n_651 ,mul_113_23_n_585 ,mul_113_23_n_649);
  xnor mul_113_23_g1508(mul_113_23_n_650 ,mul_113_23_n_648 ,mul_113_23_n_594);
  nor mul_113_23_g1509(mul_113_23_n_649 ,mul_113_23_n_588 ,mul_113_23_n_648);
  and mul_113_23_g1510(mul_113_23_n_648 ,mul_113_23_n_605 ,mul_113_23_n_646);
  xnor mul_113_23_g1511(mul_113_23_n_647 ,mul_113_23_n_645 ,mul_113_23_n_619);
  or mul_113_23_g1512(mul_113_23_n_646 ,mul_113_23_n_600 ,mul_113_23_n_645);
  and mul_113_23_g1513(mul_113_23_n_645 ,mul_113_23_n_599 ,mul_113_23_n_643);
  xnor mul_113_23_g1514(mul_113_23_n_644 ,mul_113_23_n_642 ,mul_113_23_n_618);
  or mul_113_23_g1515(mul_113_23_n_643 ,mul_113_23_n_604 ,mul_113_23_n_642);
  and mul_113_23_g1516(mul_113_23_n_642 ,mul_113_23_n_611 ,mul_113_23_n_640);
  xnor mul_113_23_g1517(mul_113_23_n_641 ,mul_113_23_n_639 ,mul_113_23_n_617);
  or mul_113_23_g1518(mul_113_23_n_640 ,mul_113_23_n_609 ,mul_113_23_n_639);
  and mul_113_23_g1519(mul_113_23_n_639 ,mul_113_23_n_608 ,mul_113_23_n_637);
  xnor mul_113_23_g1520(mul_113_23_n_638 ,mul_113_23_n_636 ,mul_113_23_n_616);
  or mul_113_23_g1521(mul_113_23_n_637 ,mul_113_23_n_607 ,mul_113_23_n_636);
  and mul_113_23_g1522(mul_113_23_n_636 ,mul_113_23_n_606 ,mul_113_23_n_634);
  xnor mul_113_23_g1523(mul_113_23_n_635 ,mul_113_23_n_633 ,mul_113_23_n_615);
  or mul_113_23_g1524(mul_113_23_n_634 ,mul_113_23_n_612 ,mul_113_23_n_633);
  and mul_113_23_g1525(mul_113_23_n_633 ,mul_113_23_n_603 ,mul_113_23_n_631);
  xnor mul_113_23_g1526(mul_113_23_n_632 ,mul_113_23_n_630 ,mul_113_23_n_614);
  or mul_113_23_g1527(mul_113_23_n_631 ,mul_113_23_n_602 ,mul_113_23_n_630);
  and mul_113_23_g1528(mul_113_23_n_630 ,mul_113_23_n_601 ,mul_113_23_n_628);
  xnor mul_113_23_g1529(mul_113_23_n_629 ,mul_113_23_n_627 ,mul_113_23_n_620);
  or mul_113_23_g1530(mul_113_23_n_628 ,mul_113_23_n_598 ,mul_113_23_n_627);
  and mul_113_23_g1531(mul_113_23_n_627 ,mul_113_23_n_597 ,mul_113_23_n_625);
  xor mul_113_23_g1532(n_326 ,mul_113_23_n_624 ,mul_113_23_n_613);
  or mul_113_23_g1533(mul_113_23_n_625 ,mul_113_23_n_596 ,mul_113_23_n_624);
  and mul_113_23_g1534(mul_113_23_n_624 ,mul_113_23_n_550 ,mul_113_23_n_623);
  or mul_113_23_g1535(mul_113_23_n_623 ,mul_113_23_n_561 ,mul_113_23_n_622);
  nor mul_113_23_g1536(mul_113_23_n_622 ,mul_113_23_n_6 ,mul_113_23_n_621);
  nor mul_113_23_g1537(mul_113_23_n_621 ,mul_113_23_n_549 ,mul_113_23_n_610);
  xnor mul_113_23_g1538(mul_113_23_n_620 ,mul_113_23_n_552 ,mul_113_23_n_580);
  xnor mul_113_23_g1539(mul_113_23_n_619 ,mul_113_23_n_564 ,mul_113_23_n_581);
  xnor mul_113_23_g1540(mul_113_23_n_618 ,mul_113_23_n_558 ,mul_113_23_n_593);
  xnor mul_113_23_g1541(mul_113_23_n_617 ,mul_113_23_n_563 ,mul_113_23_n_591);
  xnor mul_113_23_g1542(mul_113_23_n_616 ,mul_113_23_n_568 ,mul_113_23_n_576);
  xnor mul_113_23_g1543(mul_113_23_n_615 ,mul_113_23_n_566 ,mul_113_23_n_574);
  xnor mul_113_23_g1544(mul_113_23_n_614 ,mul_113_23_n_571 ,mul_113_23_n_584);
  xnor mul_113_23_g1545(mul_113_23_n_613 ,mul_113_23_n_528 ,mul_113_23_n_578);
  nor mul_113_23_g1546(mul_113_23_n_612 ,mul_113_23_n_565 ,mul_113_23_n_574);
  or mul_113_23_g1547(mul_113_23_n_611 ,mul_113_23_n_563 ,mul_113_23_n_590);
  nor mul_113_23_g1548(mul_113_23_n_610 ,mul_113_23_n_515 ,mul_113_23_n_587);
  nor mul_113_23_g1549(mul_113_23_n_609 ,mul_113_23_n_562 ,mul_113_23_n_591);
  or mul_113_23_g1550(mul_113_23_n_608 ,mul_113_23_n_568 ,mul_113_23_n_575);
  nor mul_113_23_g1551(mul_113_23_n_607 ,mul_113_23_n_567 ,mul_113_23_n_576);
  or mul_113_23_g1552(mul_113_23_n_606 ,mul_113_23_n_566 ,mul_113_23_n_573);
  or mul_113_23_g1553(mul_113_23_n_605 ,mul_113_23_n_564 ,mul_113_23_n_582);
  nor mul_113_23_g1554(mul_113_23_n_604 ,mul_113_23_n_557 ,mul_113_23_n_593);
  or mul_113_23_g1555(mul_113_23_n_603 ,mul_113_23_n_571 ,mul_113_23_n_583);
  nor mul_113_23_g1556(mul_113_23_n_602 ,mul_113_23_n_570 ,mul_113_23_n_584);
  or mul_113_23_g1557(mul_113_23_n_601 ,mul_113_23_n_552 ,mul_113_23_n_579);
  and mul_113_23_g1558(mul_113_23_n_600 ,mul_113_23_n_564 ,mul_113_23_n_582);
  or mul_113_23_g1559(mul_113_23_n_599 ,mul_113_23_n_558 ,mul_113_23_n_592);
  nor mul_113_23_g1560(mul_113_23_n_598 ,mul_113_23_n_551 ,mul_113_23_n_580);
  or mul_113_23_g1561(mul_113_23_n_597 ,mul_113_23_n_527 ,mul_113_23_n_577);
  nor mul_113_23_g1562(mul_113_23_n_596 ,mul_113_23_n_528 ,mul_113_23_n_578);
  xnor mul_113_23_g1563(mul_113_23_n_595 ,mul_113_23_n_556 ,mul_113_23_n_546);
  xnor mul_113_23_g1564(mul_113_23_n_594 ,mul_113_23_n_569 ,mul_113_23_n_553);
  not mul_113_23_g1565(mul_113_23_n_592 ,mul_113_23_n_593);
  not mul_113_23_g1566(mul_113_23_n_590 ,mul_113_23_n_591);
  or mul_113_23_g1567(mul_113_23_n_589 ,mul_113_23_n_545 ,mul_113_23_n_555);
  and mul_113_23_g1568(mul_113_23_n_588 ,mul_113_23_n_569 ,mul_113_23_n_554);
  nor mul_113_23_g1569(mul_113_23_n_587 ,mul_113_23_n_514 ,mul_113_23_n_559);
  nor mul_113_23_g1570(mul_113_23_n_586 ,mul_113_23_n_546 ,mul_113_23_n_556);
  nor mul_113_23_g1571(mul_113_23_n_585 ,mul_113_23_n_569 ,mul_113_23_n_554);
  xnor mul_113_23_g1572(mul_113_23_n_593 ,mul_113_23_n_484 ,mul_113_23_n_525);
  xnor mul_113_23_g1573(mul_113_23_n_591 ,mul_113_23_n_467 ,mul_113_23_n_524);
  not mul_113_23_g1574(mul_113_23_n_583 ,mul_113_23_n_584);
  not mul_113_23_g1575(mul_113_23_n_582 ,mul_113_23_n_581);
  not mul_113_23_g1576(mul_113_23_n_579 ,mul_113_23_n_580);
  not mul_113_23_g1577(mul_113_23_n_577 ,mul_113_23_n_578);
  not mul_113_23_g1578(mul_113_23_n_575 ,mul_113_23_n_576);
  not mul_113_23_g1579(mul_113_23_n_573 ,mul_113_23_n_574);
  xnor mul_113_23_g1580(mul_113_23_n_572 ,mul_113_23_n_530 ,mul_113_23_n_544);
  xnor mul_113_23_g1581(mul_113_23_n_584 ,mul_113_23_n_486 ,mul_113_23_n_521);
  xnor mul_113_23_g1582(mul_113_23_n_581 ,mul_113_23_n_487 ,mul_113_23_n_520);
  xnor mul_113_23_g1583(mul_113_23_n_580 ,mul_113_23_n_485 ,mul_113_23_n_519);
  xnor mul_113_23_g1584(mul_113_23_n_578 ,mul_113_23_n_481 ,mul_113_23_n_518);
  xnor mul_113_23_g1585(mul_113_23_n_576 ,mul_113_23_n_482 ,mul_113_23_n_523);
  xnor mul_113_23_g1586(mul_113_23_n_574 ,mul_113_23_n_483 ,mul_113_23_n_522);
  not mul_113_23_g1587(mul_113_23_n_570 ,mul_113_23_n_571);
  not mul_113_23_g1588(mul_113_23_n_567 ,mul_113_23_n_568);
  not mul_113_23_g1589(mul_113_23_n_565 ,mul_113_23_n_566);
  not mul_113_23_g1590(mul_113_23_n_562 ,mul_113_23_n_563);
  and mul_113_23_g1591(mul_113_23_n_561 ,mul_113_23_n_503 ,mul_113_23_n_531);
  nor mul_113_23_g1592(mul_113_23_n_560 ,mul_113_23_n_544 ,mul_113_23_n_530);
  nor mul_113_23_g1593(mul_113_23_n_559 ,mul_113_23_n_513 ,mul_113_23_n_539);
  and mul_113_23_g1594(mul_113_23_n_571 ,mul_113_23_n_492 ,mul_113_23_n_534);
  and mul_113_23_g1595(mul_113_23_n_569 ,mul_113_23_n_511 ,mul_113_23_n_542);
  and mul_113_23_g1596(mul_113_23_n_568 ,mul_113_23_n_500 ,mul_113_23_n_538);
  and mul_113_23_g1597(mul_113_23_n_566 ,mul_113_23_n_507 ,mul_113_23_n_537);
  and mul_113_23_g1598(mul_113_23_n_564 ,mul_113_23_n_517 ,mul_113_23_n_535);
  and mul_113_23_g1599(mul_113_23_n_563 ,mul_113_23_n_516 ,mul_113_23_n_536);
  not mul_113_23_g1600(mul_113_23_n_557 ,mul_113_23_n_558);
  not mul_113_23_g1601(mul_113_23_n_556 ,mul_113_23_n_555);
  not mul_113_23_g1602(mul_113_23_n_554 ,mul_113_23_n_553);
  not mul_113_23_g1603(mul_113_23_n_551 ,mul_113_23_n_552);
  or mul_113_23_g1604(mul_113_23_n_550 ,mul_113_23_n_503 ,mul_113_23_n_531);
  nor mul_113_23_g1605(mul_113_23_n_549 ,mul_113_23_n_488 ,mul_113_23_n_532);
  or mul_113_23_g1606(mul_113_23_n_548 ,mul_113_23_n_543 ,mul_113_23_n_529);
  xnor mul_113_23_g1608(mul_113_23_n_547 ,mul_113_23_n_430 ,mul_113_23_n_502);
  and mul_113_23_g1609(mul_113_23_n_558 ,mul_113_23_n_494 ,mul_113_23_n_526);
  xnor mul_113_23_g1610(mul_113_23_n_555 ,mul_113_23_n_431 ,mul_113_23_n_491);
  xnor mul_113_23_g1611(mul_113_23_n_553 ,mul_113_23_n_468 ,mul_113_23_n_489);
  and mul_113_23_g1612(mul_113_23_n_552 ,mul_113_23_n_498 ,mul_113_23_n_540);
  not mul_113_23_g1613(mul_113_23_n_545 ,mul_113_23_n_546);
  not mul_113_23_g1614(mul_113_23_n_543 ,mul_113_23_n_544);
  or mul_113_23_g1615(mul_113_23_n_542 ,mul_113_23_n_487 ,mul_113_23_n_506);
  nor mul_113_23_g1616(mul_113_23_n_541 ,mul_113_23_n_430 ,mul_113_23_n_502);
  or mul_113_23_g1617(mul_113_23_n_540 ,mul_113_23_n_481 ,mul_113_23_n_495);
  nor mul_113_23_g1618(mul_113_23_n_539 ,mul_113_23_n_438 ,mul_113_23_n_510);
  or mul_113_23_g1619(mul_113_23_n_538 ,mul_113_23_n_483 ,mul_113_23_n_508);
  or mul_113_23_g1620(mul_113_23_n_537 ,mul_113_23_n_486 ,mul_113_23_n_505);
  or mul_113_23_g1621(mul_113_23_n_536 ,mul_113_23_n_482 ,mul_113_23_n_512);
  or mul_113_23_g1622(mul_113_23_n_535 ,mul_113_23_n_484 ,mul_113_23_n_497);
  or mul_113_23_g1623(mul_113_23_n_534 ,mul_113_23_n_485 ,mul_113_23_n_499);
  or mul_113_23_g1624(mul_113_23_n_533 ,mul_113_23_n_429 ,mul_113_23_n_501);
  and mul_113_23_g1625(mul_113_23_n_546 ,mul_113_23_n_479 ,mul_113_23_n_496);
  and mul_113_23_g1626(mul_113_23_n_544 ,mul_113_23_n_477 ,mul_113_23_n_509);
  not mul_113_23_g1628(mul_113_23_n_530 ,mul_113_23_n_529);
  not mul_113_23_g1629(mul_113_23_n_527 ,mul_113_23_n_528);
  or mul_113_23_g1630(mul_113_23_n_526 ,mul_113_23_n_467 ,mul_113_23_n_504);
  xnor mul_113_23_g1631(mul_113_23_n_525 ,mul_113_23_n_375 ,mul_113_23_n_461);
  xnor mul_113_23_g1632(mul_113_23_n_524 ,mul_113_23_n_374 ,mul_113_23_n_460);
  xnor mul_113_23_g1633(mul_113_23_n_523 ,mul_113_23_n_391 ,mul_113_23_n_456);
  xnor mul_113_23_g1634(mul_113_23_n_522 ,mul_113_23_n_393 ,mul_113_23_n_464);
  xnor mul_113_23_g1635(mul_113_23_n_521 ,mul_113_23_n_385 ,mul_113_23_n_452);
  xnor mul_113_23_g1636(mul_113_23_n_520 ,mul_113_23_n_389 ,mul_113_23_n_458);
  xnor mul_113_23_g1637(mul_113_23_n_519 ,mul_113_23_n_372 ,mul_113_23_n_454);
  xnor mul_113_23_g1638(mul_113_23_n_518 ,mul_113_23_n_364 ,mul_113_23_n_466);
  xnor mul_113_23_g1639(mul_113_23_n_532 ,mul_113_23_n_404 ,mul_113_23_n_449);
  xnor mul_113_23_g1640(mul_113_23_n_531 ,mul_113_23_n_469 ,mul_113_23_n_423);
  xnor mul_113_23_g1641(mul_113_23_n_529 ,mul_113_23_n_435 ,mul_113_23_n_448);
  or mul_113_23_g1642(mul_113_23_n_528 ,mul_113_23_n_409 ,mul_113_23_n_493);
  or mul_113_23_g1643(mul_113_23_n_517 ,mul_113_23_n_375 ,mul_113_23_n_462);
  or mul_113_23_g1644(mul_113_23_n_516 ,mul_113_23_n_391 ,mul_113_23_n_455);
  nor mul_113_23_g1645(mul_113_23_n_515 ,mul_113_23_n_422 ,mul_113_23_n_472);
  nor mul_113_23_g1646(mul_113_23_n_514 ,mul_113_23_n_421 ,mul_113_23_n_473);
  nor mul_113_23_g1647(mul_113_23_n_513 ,mul_113_23_n_291 ,mul_113_23_n_470);
  nor mul_113_23_g1648(mul_113_23_n_512 ,mul_113_23_n_390 ,mul_113_23_n_456);
  or mul_113_23_g1649(mul_113_23_n_511 ,mul_113_23_n_389 ,mul_113_23_n_457);
  nor mul_113_23_g1650(mul_113_23_n_510 ,mul_113_23_n_290 ,mul_113_23_n_471);
  or mul_113_23_g1651(mul_113_23_n_509 ,mul_113_23_n_434 ,mul_113_23_n_475);
  nor mul_113_23_g1652(mul_113_23_n_508 ,mul_113_23_n_392 ,mul_113_23_n_464);
  or mul_113_23_g1653(mul_113_23_n_507 ,mul_113_23_n_385 ,mul_113_23_n_451);
  nor mul_113_23_g1654(mul_113_23_n_506 ,mul_113_23_n_388 ,mul_113_23_n_458);
  nor mul_113_23_g1655(mul_113_23_n_505 ,mul_113_23_n_384 ,mul_113_23_n_452);
  nor mul_113_23_g1656(mul_113_23_n_504 ,mul_113_23_n_373 ,mul_113_23_n_460);
  not mul_113_23_g1657(mul_113_23_n_502 ,mul_113_23_n_501);
  or mul_113_23_g1658(mul_113_23_n_500 ,mul_113_23_n_393 ,mul_113_23_n_463);
  nor mul_113_23_g1659(mul_113_23_n_499 ,mul_113_23_n_371 ,mul_113_23_n_454);
  or mul_113_23_g1660(mul_113_23_n_498 ,mul_113_23_n_364 ,mul_113_23_n_465);
  and mul_113_23_g1661(mul_113_23_n_497 ,mul_113_23_n_375 ,mul_113_23_n_462);
  or mul_113_23_g1662(mul_113_23_n_496 ,mul_113_23_n_468 ,mul_113_23_n_478);
  nor mul_113_23_g1663(mul_113_23_n_495 ,mul_113_23_n_363 ,mul_113_23_n_466);
  or mul_113_23_g1664(mul_113_23_n_494 ,mul_113_23_n_374 ,mul_113_23_n_459);
  and mul_113_23_g1665(mul_113_23_n_493 ,mul_113_23_n_408 ,mul_113_23_n_469);
  or mul_113_23_g1666(mul_113_23_n_492 ,mul_113_23_n_372 ,mul_113_23_n_453);
  and mul_113_23_g1667(mul_113_23_n_503 ,mul_113_23_n_428 ,mul_113_23_n_480);
  xnor mul_113_23_g1668(mul_113_23_n_491 ,mul_113_23_n_399 ,mul_113_23_n_434);
  xnor mul_113_23_g1669(mul_113_23_n_490 ,mul_113_23_n_166 ,mul_113_23_n_447);
  xnor mul_113_23_g1670(mul_113_23_n_489 ,mul_113_23_n_417 ,mul_113_23_n_433);
  and mul_113_23_g1671(mul_113_23_n_501 ,mul_113_23_n_440 ,mul_113_23_n_450);
  or mul_113_23_g1673(mul_113_23_n_480 ,mul_113_23_n_404 ,mul_113_23_n_442);
  or mul_113_23_g1674(mul_113_23_n_479 ,mul_113_23_n_416 ,mul_113_23_n_433);
  nor mul_113_23_g1675(mul_113_23_n_478 ,mul_113_23_n_417 ,mul_113_23_n_432);
  or mul_113_23_g1676(mul_113_23_n_477 ,mul_113_23_n_399 ,mul_113_23_n_5);
  nor mul_113_23_g1677(mul_113_23_n_476 ,mul_113_23_n_165 ,mul_113_23_n_447);
  nor mul_113_23_g1678(mul_113_23_n_475 ,mul_113_23_n_398 ,mul_113_23_n_431);
  or mul_113_23_g1679(mul_113_23_n_474 ,mul_113_23_n_166 ,mul_113_23_n_446);
  or mul_113_23_g1680(mul_113_23_n_488 ,mul_113_23_n_381 ,mul_113_23_n_441);
  and mul_113_23_g1681(mul_113_23_n_487 ,mul_113_23_n_286 ,mul_113_23_n_439);
  and mul_113_23_g1682(mul_113_23_n_486 ,mul_113_23_n_268 ,mul_113_23_n_436);
  and mul_113_23_g1683(mul_113_23_n_485 ,mul_113_23_n_266 ,mul_113_23_n_426);
  and mul_113_23_g1684(mul_113_23_n_484 ,mul_113_23_n_318 ,mul_113_23_n_427);
  and mul_113_23_g1685(mul_113_23_n_483 ,mul_113_23_n_320 ,mul_113_23_n_437);
  and mul_113_23_g1686(mul_113_23_n_482 ,mul_113_23_n_310 ,mul_113_23_n_445);
  and mul_113_23_g1687(mul_113_23_n_481 ,mul_113_23_n_288 ,mul_113_23_n_425);
  not mul_113_23_g1688(mul_113_23_n_473 ,mul_113_23_n_472);
  not mul_113_23_g1689(mul_113_23_n_471 ,mul_113_23_n_470);
  not mul_113_23_g1690(mul_113_23_n_465 ,mul_113_23_n_466);
  not mul_113_23_g1691(mul_113_23_n_463 ,mul_113_23_n_464);
  not mul_113_23_g1692(mul_113_23_n_462 ,mul_113_23_n_461);
  not mul_113_23_g1693(mul_113_23_n_459 ,mul_113_23_n_460);
  not mul_113_23_g1694(mul_113_23_n_457 ,mul_113_23_n_458);
  not mul_113_23_g1695(mul_113_23_n_455 ,mul_113_23_n_456);
  not mul_113_23_g1696(mul_113_23_n_453 ,mul_113_23_n_454);
  not mul_113_23_g1697(mul_113_23_n_451 ,mul_113_23_n_452);
  or mul_113_23_g1698(mul_113_23_n_450 ,mul_113_23_n_435 ,mul_113_23_n_443);
  xnor mul_113_23_g1699(mul_113_23_n_472 ,mul_113_23_n_418 ,mul_113_23_n_394);
  xnor mul_113_23_g1700(mul_113_23_n_470 ,mul_113_23_n_246 ,mul_113_23_n_395);
  xnor mul_113_23_g1701(mul_113_23_n_449 ,mul_113_23_n_366 ,mul_113_23_n_415);
  xnor mul_113_23_g1702(mul_113_23_n_448 ,mul_113_23_n_387 ,mul_113_23_n_397);
  xnor mul_113_23_g1703(mul_113_23_n_469 ,mul_113_23_n_401 ,mul_113_23_n_335);
  and mul_113_23_g1704(mul_113_23_n_468 ,mul_113_23_n_309 ,mul_113_23_n_444);
  and mul_113_23_g1705(mul_113_23_n_467 ,mul_113_23_n_303 ,mul_113_23_n_424);
  xnor mul_113_23_g1706(mul_113_23_n_466 ,mul_113_23_n_403 ,mul_113_23_n_337);
  xnor mul_113_23_g1707(mul_113_23_n_464 ,mul_113_23_n_420 ,mul_113_23_n_338);
  xnor mul_113_23_g1708(mul_113_23_n_461 ,mul_113_23_n_407 ,mul_113_23_n_340);
  xnor mul_113_23_g1709(mul_113_23_n_460 ,mul_113_23_n_402 ,mul_113_23_n_336);
  xnor mul_113_23_g1710(mul_113_23_n_458 ,mul_113_23_n_419 ,mul_113_23_n_346);
  xnor mul_113_23_g1711(mul_113_23_n_456 ,mul_113_23_n_406 ,mul_113_23_n_344);
  xnor mul_113_23_g1712(mul_113_23_n_454 ,mul_113_23_n_405 ,mul_113_23_n_339);
  xnor mul_113_23_g1713(mul_113_23_n_452 ,mul_113_23_n_400 ,mul_113_23_n_324);
  not mul_113_23_g1714(mul_113_23_n_446 ,mul_113_23_n_447);
  or mul_113_23_g1715(mul_113_23_n_445 ,mul_113_23_n_278 ,mul_113_23_n_420);
  or mul_113_23_g1716(mul_113_23_n_444 ,mul_113_23_n_311 ,mul_113_23_n_419);
  nor mul_113_23_g1717(mul_113_23_n_443 ,mul_113_23_n_387 ,mul_113_23_n_396);
  nor mul_113_23_g1718(mul_113_23_n_442 ,mul_113_23_n_366 ,mul_113_23_n_414);
  nor mul_113_23_g1719(mul_113_23_n_441 ,mul_113_23_n_382 ,mul_113_23_n_418);
  or mul_113_23_g1720(mul_113_23_n_440 ,mul_113_23_n_386 ,mul_113_23_n_397);
  or mul_113_23_g1721(mul_113_23_n_439 ,mul_113_23_n_292 ,mul_113_23_n_407);
  nor mul_113_23_g1722(mul_113_23_n_438 ,mul_113_23_n_379 ,mul_113_23_n_412);
  or mul_113_23_g1723(mul_113_23_n_437 ,mul_113_23_n_314 ,mul_113_23_n_400);
  or mul_113_23_g1724(mul_113_23_n_436 ,mul_113_23_n_281 ,mul_113_23_n_405);
  or mul_113_23_g1725(mul_113_23_n_447 ,mul_113_23_n_264 ,mul_113_23_n_410);
  not mul_113_23_g1726(mul_113_23_n_432 ,mul_113_23_n_433);
  not mul_113_23_g1727(mul_113_23_n_431 ,mul_113_23_n_5);
  not mul_113_23_g1728(mul_113_23_n_429 ,mul_113_23_n_430);
  or mul_113_23_g1729(mul_113_23_n_428 ,mul_113_23_n_365 ,mul_113_23_n_415);
  or mul_113_23_g1730(mul_113_23_n_427 ,mul_113_23_n_317 ,mul_113_23_n_402);
  or mul_113_23_g1731(mul_113_23_n_426 ,mul_113_23_n_287 ,mul_113_23_n_403);
  or mul_113_23_g1732(mul_113_23_n_425 ,mul_113_23_n_285 ,mul_113_23_n_401);
  or mul_113_23_g1733(mul_113_23_n_424 ,mul_113_23_n_313 ,mul_113_23_n_406);
  xnor mul_113_23_g1734(mul_113_23_n_423 ,mul_113_23_n_370 ,mul_113_23_n_368);
  and mul_113_23_g1735(mul_113_23_n_435 ,mul_113_23_n_269 ,mul_113_23_n_413);
  and mul_113_23_g1736(mul_113_23_n_434 ,mul_113_23_n_302 ,mul_113_23_n_411);
  xnor mul_113_23_g1737(mul_113_23_n_433 ,mul_113_23_n_378 ,mul_113_23_n_0);
  xnor mul_113_23_g1739(mul_113_23_n_430 ,mul_113_23_n_376 ,mul_113_23_n_326);
  not mul_113_23_g1740(mul_113_23_n_422 ,mul_113_23_n_421);
  not mul_113_23_g1741(mul_113_23_n_416 ,mul_113_23_n_417);
  not mul_113_23_g1742(mul_113_23_n_414 ,mul_113_23_n_415);
  or mul_113_23_g1743(mul_113_23_n_413 ,mul_113_23_n_295 ,mul_113_23_n_377);
  nor mul_113_23_g1744(mul_113_23_n_412 ,mul_113_23_n_380 ,mul_113_23_n_3);
  or mul_113_23_g1745(mul_113_23_n_411 ,mul_113_23_n_282 ,mul_113_23_n_378);
  and mul_113_23_g1746(mul_113_23_n_410 ,mul_113_23_n_299 ,mul_113_23_n_376);
  nor mul_113_23_g1747(mul_113_23_n_409 ,mul_113_23_n_370 ,mul_113_23_n_367);
  or mul_113_23_g1748(mul_113_23_n_408 ,mul_113_23_n_369 ,mul_113_23_n_368);
  xnor mul_113_23_g1749(mul_113_23_n_421 ,mul_113_23_n_234 ,mul_113_23_n_2);
  xnor mul_113_23_g1750(mul_113_23_n_420 ,mul_113_23_n_198 ,mul_113_23_n_329);
  xnor mul_113_23_g1751(mul_113_23_n_419 ,mul_113_23_n_200 ,mul_113_23_n_342);
  and mul_113_23_g1752(mul_113_23_n_418 ,mul_113_23_n_294 ,mul_113_23_n_383);
  xnor mul_113_23_g1753(mul_113_23_n_417 ,mul_113_23_n_250 ,mul_113_23_n_322);
  xnor mul_113_23_g1754(mul_113_23_n_415 ,mul_113_23_n_196 ,mul_113_23_n_332);
  not mul_113_23_g1755(mul_113_23_n_398 ,mul_113_23_n_399);
  not mul_113_23_g1756(mul_113_23_n_396 ,mul_113_23_n_397);
  xnor mul_113_23_g1757(mul_113_23_n_395 ,mul_113_23_n_1 ,mul_113_23_n_158);
  xnor mul_113_23_g1758(mul_113_23_n_394 ,mul_113_23_n_289 ,mul_113_23_n_4);
  xnor mul_113_23_g1759(mul_113_23_n_407 ,mul_113_23_n_249 ,mul_113_23_n_333);
  xnor mul_113_23_g1760(mul_113_23_n_406 ,mul_113_23_n_253 ,mul_113_23_n_330);
  xnor mul_113_23_g1761(mul_113_23_n_405 ,mul_113_23_n_252 ,mul_113_23_n_327);
  xnor mul_113_23_g1762(mul_113_23_n_404 ,mul_113_23_n_321 ,mul_113_23_n_345);
  xnor mul_113_23_g1763(mul_113_23_n_403 ,mul_113_23_n_201 ,mul_113_23_n_325);
  xnor mul_113_23_g1764(mul_113_23_n_402 ,mul_113_23_n_256 ,mul_113_23_n_328);
  xnor mul_113_23_g1765(mul_113_23_n_401 ,mul_113_23_n_202 ,mul_113_23_n_323);
  xnor mul_113_23_g1766(mul_113_23_n_400 ,mul_113_23_n_257 ,mul_113_23_n_331);
  xnor mul_113_23_g1767(mul_113_23_n_399 ,mul_113_23_n_203 ,mul_113_23_n_343);
  xnor mul_113_23_g1768(mul_113_23_n_397 ,mul_113_23_n_197 ,mul_113_23_n_341);
  not mul_113_23_g1769(mul_113_23_n_392 ,mul_113_23_n_393);
  not mul_113_23_g1770(mul_113_23_n_390 ,mul_113_23_n_391);
  not mul_113_23_g1771(mul_113_23_n_388 ,mul_113_23_n_389);
  not mul_113_23_g1772(mul_113_23_n_386 ,mul_113_23_n_387);
  not mul_113_23_g1773(mul_113_23_n_384 ,mul_113_23_n_385);
  or mul_113_23_g1774(mul_113_23_n_383 ,mul_113_23_n_280 ,mul_113_23_n_1);
  nor mul_113_23_g1775(mul_113_23_n_382 ,mul_113_23_n_289 ,mul_113_23_n_4);
  and mul_113_23_g1776(mul_113_23_n_381 ,mul_113_23_n_289 ,mul_113_23_n_4);
  and mul_113_23_g1777(mul_113_23_n_380 ,mul_113_23_n_258 ,mul_113_23_n_362);
  nor mul_113_23_g1778(mul_113_23_n_379 ,mul_113_23_n_258 ,mul_113_23_n_362);
  and mul_113_23_g1779(mul_113_23_n_393 ,mul_113_23_n_261 ,mul_113_23_n_359);
  and mul_113_23_g1780(mul_113_23_n_391 ,mul_113_23_n_262 ,mul_113_23_n_361);
  and mul_113_23_g1781(mul_113_23_n_389 ,mul_113_23_n_296 ,mul_113_23_n_360);
  or mul_113_23_g1782(mul_113_23_n_387 ,mul_113_23_n_297 ,mul_113_23_n_353);
  and mul_113_23_g1783(mul_113_23_n_385 ,mul_113_23_n_270 ,mul_113_23_n_358);
  not mul_113_23_g1785(mul_113_23_n_373 ,mul_113_23_n_374);
  not mul_113_23_g1786(mul_113_23_n_371 ,mul_113_23_n_372);
  not mul_113_23_g1787(mul_113_23_n_369 ,mul_113_23_n_370);
  not mul_113_23_g1788(mul_113_23_n_367 ,mul_113_23_n_368);
  not mul_113_23_g1789(mul_113_23_n_366 ,mul_113_23_n_365);
  not mul_113_23_g1790(mul_113_23_n_363 ,mul_113_23_n_364);
  and mul_113_23_g1791(mul_113_23_n_378 ,mul_113_23_n_273 ,mul_113_23_n_357);
  and mul_113_23_g1792(mul_113_23_n_377 ,mul_113_23_n_304 ,mul_113_23_n_355);
  or mul_113_23_g1793(mul_113_23_n_376 ,mul_113_23_n_307 ,mul_113_23_n_347);
  and mul_113_23_g1794(mul_113_23_n_375 ,mul_113_23_n_279 ,mul_113_23_n_356);
  and mul_113_23_g1795(mul_113_23_n_374 ,mul_113_23_n_301 ,mul_113_23_n_351);
  and mul_113_23_g1796(mul_113_23_n_372 ,mul_113_23_n_308 ,mul_113_23_n_354);
  and mul_113_23_g1797(mul_113_23_n_370 ,mul_113_23_n_265 ,mul_113_23_n_350);
  or mul_113_23_g1798(mul_113_23_n_368 ,mul_113_23_n_305 ,mul_113_23_n_349);
  and mul_113_23_g1799(mul_113_23_n_365 ,mul_113_23_n_271 ,mul_113_23_n_348);
  and mul_113_23_g1800(mul_113_23_n_364 ,mul_113_23_n_284 ,mul_113_23_n_352);
  or mul_113_23_g1802(mul_113_23_n_361 ,mul_113_23_n_198 ,mul_113_23_n_263);
  or mul_113_23_g1803(mul_113_23_n_360 ,mul_113_23_n_249 ,mul_113_23_n_277);
  or mul_113_23_g1804(mul_113_23_n_359 ,mul_113_23_n_257 ,mul_113_23_n_283);
  or mul_113_23_g1805(mul_113_23_n_358 ,mul_113_23_n_252 ,mul_113_23_n_272);
  or mul_113_23_g1806(mul_113_23_n_357 ,mul_113_23_n_200 ,mul_113_23_n_276);
  or mul_113_23_g1807(mul_113_23_n_356 ,mul_113_23_n_256 ,mul_113_23_n_275);
  or mul_113_23_g1808(mul_113_23_n_355 ,mul_113_23_n_251 ,mul_113_23_n_312);
  or mul_113_23_g1809(mul_113_23_n_354 ,mul_113_23_n_201 ,mul_113_23_n_274);
  and mul_113_23_g1810(mul_113_23_n_353 ,mul_113_23_n_203 ,mul_113_23_n_293);
  or mul_113_23_g1811(mul_113_23_n_352 ,mul_113_23_n_202 ,mul_113_23_n_319);
  or mul_113_23_g1812(mul_113_23_n_351 ,mul_113_23_n_253 ,mul_113_23_n_267);
  or mul_113_23_g1813(mul_113_23_n_350 ,mul_113_23_n_196 ,mul_113_23_n_298);
  and mul_113_23_g1814(mul_113_23_n_349 ,mul_113_23_n_321 ,mul_113_23_n_316);
  or mul_113_23_g1815(mul_113_23_n_348 ,mul_113_23_n_204 ,mul_113_23_n_315);
  and mul_113_23_g1816(mul_113_23_n_347 ,mul_113_23_n_197 ,mul_113_23_n_300);
  or mul_113_23_g1817(mul_113_23_n_362 ,mul_113_23_n_147 ,mul_113_23_n_306);
  xnor mul_113_23_g1818(mul_113_23_n_346 ,mul_113_23_n_231 ,mul_113_23_n_229);
  xnor mul_113_23_g1819(mul_113_23_n_345 ,mul_113_23_n_242 ,mul_113_23_n_191);
  xnor mul_113_23_g1820(mul_113_23_n_344 ,mul_113_23_n_174 ,mul_113_23_n_248);
  xnor mul_113_23_g1821(mul_113_23_n_343 ,mul_113_23_n_170 ,mul_113_23_n_221);
  xnor mul_113_23_g1824(mul_113_23_n_342 ,mul_113_23_n_218 ,mul_113_23_n_164);
  xnor mul_113_23_g1825(mul_113_23_n_341 ,mul_113_23_n_210 ,mul_113_23_n_176);
  xnor mul_113_23_g1826(mul_113_23_n_340 ,mul_113_23_n_225 ,mul_113_23_n_168);
  xnor mul_113_23_g1827(mul_113_23_n_339 ,mul_113_23_n_233 ,mul_113_23_n_178);
  xnor mul_113_23_g1828(mul_113_23_n_338 ,mul_113_23_n_213 ,mul_113_23_n_237);
  xnor mul_113_23_g1829(mul_113_23_n_337 ,mul_113_23_n_212 ,mul_113_23_n_180);
  xnor mul_113_23_g1830(mul_113_23_n_336 ,mul_113_23_n_217 ,mul_113_23_n_182);
  xnor mul_113_23_g1831(mul_113_23_n_335 ,mul_113_23_n_185 ,mul_113_23_n_157);
  xnor mul_113_23_g1832(mul_113_23_n_334 ,mul_113_23_n_163 ,mul_113_23_n_207);
  xnor mul_113_23_g1834(mul_113_23_n_333 ,mul_113_23_n_159 ,mul_113_23_n_186);
  xnor mul_113_23_g1835(mul_113_23_n_332 ,mul_113_23_n_160 ,mul_113_23_n_236);
  xnor mul_113_23_g1836(mul_113_23_n_331 ,mul_113_23_n_193 ,mul_113_23_n_243);
  xnor mul_113_23_g1837(mul_113_23_n_330 ,mul_113_23_n_222 ,mul_113_23_n_235);
  xnor mul_113_23_g1838(mul_113_23_n_329 ,mul_113_23_n_171 ,mul_113_23_n_227);
  xnor mul_113_23_g1839(mul_113_23_n_328 ,mul_113_23_n_183 ,mul_113_23_n_194);
  xnor mul_113_23_g1840(mul_113_23_n_327 ,mul_113_23_n_245 ,mul_113_23_n_172);
  xnor mul_113_23_g1841(mul_113_23_n_326 ,mul_113_23_n_215 ,mul_113_23_n_219);
  xnor mul_113_23_g1842(mul_113_23_n_325 ,mul_113_23_n_244 ,mul_113_23_n_187);
  xnor mul_113_23_g1843(mul_113_23_n_324 ,mul_113_23_n_162 ,mul_113_23_n_239);
  xnor mul_113_23_g1844(mul_113_23_n_323 ,mul_113_23_n_226 ,mul_113_23_n_189);
  xnor mul_113_23_g1845(mul_113_23_n_322 ,mul_113_23_n_240 ,mul_113_23_n_192);
  or mul_113_23_g1847(mul_113_23_n_320 ,mul_113_23_n_161 ,mul_113_23_n_239);
  and mul_113_23_g1848(mul_113_23_n_319 ,mul_113_23_n_226 ,mul_113_23_n_189);
  or mul_113_23_g1849(mul_113_23_n_318 ,mul_113_23_n_216 ,mul_113_23_n_182);
  nor mul_113_23_g1850(mul_113_23_n_317 ,mul_113_23_n_181 ,mul_113_23_n_217);
  or mul_113_23_g1851(mul_113_23_n_316 ,mul_113_23_n_190 ,mul_113_23_n_242);
  and mul_113_23_g1852(mul_113_23_n_315 ,mul_113_23_n_234 ,mul_113_23_n_223);
  nor mul_113_23_g1853(mul_113_23_n_314 ,mul_113_23_n_238 ,mul_113_23_n_162);
  nor mul_113_23_g1854(mul_113_23_n_313 ,mul_113_23_n_247 ,mul_113_23_n_174);
  and mul_113_23_g1855(mul_113_23_n_312 ,mul_113_23_n_240 ,mul_113_23_n_192);
  nor mul_113_23_g1856(mul_113_23_n_311 ,mul_113_23_n_228 ,mul_113_23_n_231);
  or mul_113_23_g1857(mul_113_23_n_310 ,mul_113_23_n_214 ,mul_113_23_n_237);
  or mul_113_23_g1858(mul_113_23_n_309 ,mul_113_23_n_230 ,mul_113_23_n_229);
  or mul_113_23_g1859(mul_113_23_n_308 ,mul_113_23_n_244 ,mul_113_23_n_187);
  nor mul_113_23_g1860(mul_113_23_n_307 ,mul_113_23_n_175 ,mul_113_23_n_210);
  or mul_113_23_g1861(mul_113_23_n_306 ,mul_113_23_n_33 ,mul_113_23_n_255);
  nor mul_113_23_g1862(mul_113_23_n_305 ,mul_113_23_n_241 ,mul_113_23_n_191);
  or mul_113_23_g1863(mul_113_23_n_304 ,mul_113_23_n_240 ,mul_113_23_n_192);
  or mul_113_23_g1864(mul_113_23_n_303 ,mul_113_23_n_173 ,mul_113_23_n_248);
  or mul_113_23_g1865(mul_113_23_n_302 ,mul_113_23_n_188 ,mul_113_23_n_70);
  or mul_113_23_g1866(mul_113_23_n_301 ,mul_113_23_n_222 ,mul_113_23_n_235);
  or mul_113_23_g1867(mul_113_23_n_300 ,mul_113_23_n_209 ,mul_113_23_n_176);
  or mul_113_23_g1868(mul_113_23_n_299 ,mul_113_23_n_215 ,mul_113_23_n_219);
  and mul_113_23_g1869(mul_113_23_n_298 ,mul_113_23_n_160 ,mul_113_23_n_236);
  nor mul_113_23_g1870(mul_113_23_n_297 ,mul_113_23_n_220 ,mul_113_23_n_170);
  or mul_113_23_g1871(mul_113_23_n_296 ,mul_113_23_n_159 ,mul_113_23_n_186);
  and mul_113_23_g1872(mul_113_23_n_295 ,mul_113_23_n_163 ,mul_113_23_n_208);
  or mul_113_23_g1873(mul_113_23_n_294 ,mul_113_23_n_246 ,mul_113_23_n_158);
  or mul_113_23_g1874(mul_113_23_n_293 ,mul_113_23_n_169 ,mul_113_23_n_221);
  nor mul_113_23_g1875(mul_113_23_n_292 ,mul_113_23_n_167 ,mul_113_23_n_225);
  or mul_113_23_g1876(mul_113_23_n_321 ,mul_113_23_n_260 ,mul_113_23_n_206);
  not mul_113_23_g1877(mul_113_23_n_291 ,mul_113_23_n_290);
  or mul_113_23_g1878(mul_113_23_n_288 ,mul_113_23_n_184 ,mul_113_23_n_157);
  nor mul_113_23_g1879(mul_113_23_n_287 ,mul_113_23_n_179 ,mul_113_23_n_212);
  or mul_113_23_g1880(mul_113_23_n_286 ,mul_113_23_n_224 ,mul_113_23_n_168);
  nor mul_113_23_g1881(mul_113_23_n_285 ,mul_113_23_n_156 ,mul_113_23_n_185);
  or mul_113_23_g1882(mul_113_23_n_284 ,mul_113_23_n_226 ,mul_113_23_n_189);
  and mul_113_23_g1883(mul_113_23_n_283 ,mul_113_23_n_193 ,mul_113_23_n_243);
  and mul_113_23_g1884(mul_113_23_n_282 ,mul_113_23_n_188 ,mul_113_23_n_70);
  nor mul_113_23_g1885(mul_113_23_n_281 ,mul_113_23_n_177 ,mul_113_23_n_233);
  and mul_113_23_g1886(mul_113_23_n_280 ,mul_113_23_n_246 ,mul_113_23_n_158);
  or mul_113_23_g1887(mul_113_23_n_279 ,mul_113_23_n_183 ,mul_113_23_n_194);
  and mul_113_23_g1888(mul_113_23_n_278 ,mul_113_23_n_237 ,mul_113_23_n_214);
  and mul_113_23_g1889(mul_113_23_n_277 ,mul_113_23_n_159 ,mul_113_23_n_186);
  and mul_113_23_g1890(mul_113_23_n_276 ,mul_113_23_n_218 ,mul_113_23_n_164);
  and mul_113_23_g1891(mul_113_23_n_275 ,mul_113_23_n_183 ,mul_113_23_n_194);
  and mul_113_23_g1892(mul_113_23_n_274 ,mul_113_23_n_244 ,mul_113_23_n_187);
  or mul_113_23_g1893(mul_113_23_n_273 ,mul_113_23_n_218 ,mul_113_23_n_164);
  and mul_113_23_g1894(mul_113_23_n_272 ,mul_113_23_n_245 ,mul_113_23_n_172);
  or mul_113_23_g1895(mul_113_23_n_271 ,mul_113_23_n_234 ,mul_113_23_n_223);
  or mul_113_23_g1896(mul_113_23_n_270 ,mul_113_23_n_245 ,mul_113_23_n_172);
  or mul_113_23_g1897(mul_113_23_n_269 ,mul_113_23_n_208 ,mul_113_23_n_163);
  or mul_113_23_g1898(mul_113_23_n_268 ,mul_113_23_n_232 ,mul_113_23_n_178);
  and mul_113_23_g1899(mul_113_23_n_267 ,mul_113_23_n_222 ,mul_113_23_n_235);
  or mul_113_23_g1900(mul_113_23_n_266 ,mul_113_23_n_211 ,mul_113_23_n_180);
  or mul_113_23_g1901(mul_113_23_n_265 ,mul_113_23_n_160 ,mul_113_23_n_236);
  and mul_113_23_g1902(mul_113_23_n_264 ,mul_113_23_n_215 ,mul_113_23_n_219);
  and mul_113_23_g1903(mul_113_23_n_263 ,mul_113_23_n_171 ,mul_113_23_n_227);
  or mul_113_23_g1904(mul_113_23_n_262 ,mul_113_23_n_171 ,mul_113_23_n_227);
  or mul_113_23_g1905(mul_113_23_n_261 ,mul_113_23_n_193 ,mul_113_23_n_243);
  and mul_113_23_g1906(mul_113_23_n_290 ,mul_113_23_n_254 ,mul_113_23_n_205);
  and mul_113_23_g1907(mul_113_23_n_289 ,mul_113_23_n_195 ,mul_113_23_n_199);
  not mul_113_23_g1908(mul_113_23_n_260 ,mul_113_23_n_259);
  not mul_113_23_g1909(mul_113_23_n_254 ,mul_113_23_n_255);
  not mul_113_23_g1910(mul_113_23_n_251 ,mul_113_23_n_250);
  not mul_113_23_g1911(mul_113_23_n_247 ,mul_113_23_n_248);
  not mul_113_23_g1912(mul_113_23_n_241 ,mul_113_23_n_242);
  not mul_113_23_g1913(mul_113_23_n_238 ,mul_113_23_n_239);
  not mul_113_23_g1914(mul_113_23_n_232 ,mul_113_23_n_233);
  not mul_113_23_g1915(mul_113_23_n_230 ,mul_113_23_n_231);
  not mul_113_23_g1916(mul_113_23_n_228 ,mul_113_23_n_229);
  not mul_113_23_g1917(mul_113_23_n_224 ,mul_113_23_n_225);
  not mul_113_23_g1918(mul_113_23_n_220 ,mul_113_23_n_221);
  not mul_113_23_g1919(mul_113_23_n_216 ,mul_113_23_n_217);
  not mul_113_23_g1920(mul_113_23_n_214 ,mul_113_23_n_213);
  not mul_113_23_g1921(mul_113_23_n_211 ,mul_113_23_n_212);
  not mul_113_23_g1922(mul_113_23_n_209 ,mul_113_23_n_210);
  not mul_113_23_g1923(mul_113_23_n_208 ,mul_113_23_n_207);
  or mul_113_23_g1924(mul_113_23_n_259 ,mul_113_23_n_141 ,mul_113_23_n_40);
  or mul_113_23_g1925(mul_113_23_n_258 ,mul_113_23_n_147 ,mul_113_23_n_49);
  or mul_113_23_g1926(mul_113_23_n_257 ,mul_113_23_n_117 ,mul_113_23_n_48);
  or mul_113_23_g1927(mul_113_23_n_256 ,mul_113_23_n_111 ,mul_113_23_n_37);
  or mul_113_23_g1928(mul_113_23_n_255 ,mul_113_23_n_119 ,mul_113_23_n_39);
  or mul_113_23_g1929(mul_113_23_n_253 ,mul_113_23_n_115 ,mul_113_23_n_35);
  or mul_113_23_g1930(mul_113_23_n_252 ,mul_113_23_n_52 ,mul_113_23_n_46);
  or mul_113_23_g1931(mul_113_23_n_250 ,mul_113_23_n_61 ,mul_113_23_n_11);
  or mul_113_23_g1932(mul_113_23_n_249 ,mul_113_23_n_151 ,mul_113_23_n_49);
  or mul_113_23_g1933(mul_113_23_n_248 ,mul_113_23_n_55 ,mul_113_23_n_14);
  or mul_113_23_g1934(mul_113_23_n_246 ,mul_113_23_n_147 ,mul_113_23_n_21);
  or mul_113_23_g1935(mul_113_23_n_245 ,mul_113_23_n_117 ,mul_113_23_n_18);
  or mul_113_23_g1936(mul_113_23_n_244 ,mul_113_23_n_150 ,mul_113_23_n_23);
  or mul_113_23_g1937(mul_113_23_n_243 ,mul_113_23_n_115 ,mul_113_23_n_16);
  or mul_113_23_g1938(mul_113_23_n_242 ,mul_113_23_n_119 ,mul_113_23_n_29);
  or mul_113_23_g1939(mul_113_23_n_240 ,mul_113_23_n_58 ,mul_113_23_n_93);
  or mul_113_23_g1940(mul_113_23_n_239 ,mul_113_23_n_52 ,mul_113_23_n_75);
  or mul_113_23_g1941(mul_113_23_n_237 ,mul_113_23_n_149 ,mul_113_23_n_77);
  or mul_113_23_g1942(mul_113_23_n_236 ,mul_113_23_n_154 ,mul_113_23_n_8);
  or mul_113_23_g1943(mul_113_23_n_235 ,mul_113_23_n_61 ,mul_113_23_n_31);
  or mul_113_23_g1944(mul_113_23_n_234 ,mul_113_23_n_155 ,mul_113_23_n_21);
  or mul_113_23_g1945(mul_113_23_n_233 ,mul_113_23_n_144 ,mul_113_23_n_26);
  or mul_113_23_g1946(mul_113_23_n_231 ,mul_113_23_n_111 ,mul_113_23_n_79);
  or mul_113_23_g1947(mul_113_23_n_229 ,mul_113_23_n_151 ,mul_113_23_n_14);
  or mul_113_23_g1948(mul_113_23_n_227 ,mul_113_23_n_140 ,mul_113_23_n_81);
  or mul_113_23_g1949(mul_113_23_n_226 ,mul_113_23_n_154 ,mul_113_23_n_43);
  or mul_113_23_g1950(mul_113_23_n_225 ,mul_113_23_n_145 ,mul_113_23_n_28);
  or mul_113_23_g1951(mul_113_23_n_223 ,mul_113_23_n_153 ,mul_113_23_n_96);
  or mul_113_23_g1952(mul_113_23_n_222 ,mul_113_23_n_140 ,mul_113_23_n_40);
  or mul_113_23_g1953(mul_113_23_n_221 ,mul_113_23_n_142 ,mul_113_23_n_90);
  or mul_113_23_g1954(mul_113_23_n_219 ,mul_113_23_n_142 ,mul_113_23_n_75);
  or mul_113_23_g1955(mul_113_23_n_218 ,mul_113_23_n_152 ,mul_113_23_n_87);
  or mul_113_23_g1956(mul_113_23_n_217 ,mul_113_23_n_143 ,mul_113_23_n_26);
  or mul_113_23_g1957(mul_113_23_n_215 ,mul_113_23_n_113 ,mul_113_23_n_25);
  or mul_113_23_g1958(mul_113_23_n_213 ,mul_113_23_n_150 ,mul_113_23_n_79);
  or mul_113_23_g1959(mul_113_23_n_212 ,mul_113_23_n_141 ,mul_113_23_n_29);
  or mul_113_23_g1960(mul_113_23_n_210 ,mul_113_23_n_113 ,mul_113_23_n_77);
  or mul_113_23_g1961(mul_113_23_n_207 ,mul_113_23_n_142 ,mul_113_23_n_31);
  not mul_113_23_g1967(mul_113_23_n_191 ,mul_113_23_n_190);
  not mul_113_23_g1968(mul_113_23_n_185 ,mul_113_23_n_184);
  not mul_113_23_g1969(mul_113_23_n_182 ,mul_113_23_n_181);
  not mul_113_23_g1970(mul_113_23_n_180 ,mul_113_23_n_179);
  not mul_113_23_g1971(mul_113_23_n_178 ,mul_113_23_n_177);
  not mul_113_23_g1972(mul_113_23_n_176 ,mul_113_23_n_175);
  not mul_113_23_g1973(mul_113_23_n_174 ,mul_113_23_n_173);
  not mul_113_23_g1974(mul_113_23_n_170 ,mul_113_23_n_169);
  not mul_113_23_g1975(mul_113_23_n_168 ,mul_113_23_n_167);
  not mul_113_23_g1976(mul_113_23_n_166 ,mul_113_23_n_165);
  not mul_113_23_g1977(mul_113_23_n_162 ,mul_113_23_n_161);
  not mul_113_23_g1978(mul_113_23_n_157 ,mul_113_23_n_156);
  and mul_113_23_g1979(mul_113_23_n_206 ,in31[4] ,mul_113_23_n_121);
  and mul_113_23_g1980(mul_113_23_n_205 ,in31[2] ,mul_113_23_n_121);
  and mul_113_23_g1981(mul_113_23_n_204 ,in31[0] ,mul_113_23_n_67);
  or mul_113_23_g1982(mul_113_23_n_203 ,mul_113_23_n_64 ,mul_113_23_n_10);
  or mul_113_23_g1983(mul_113_23_n_202 ,mul_113_23_n_144 ,mul_113_23_n_45);
  or mul_113_23_g1984(mul_113_23_n_201 ,mul_113_23_n_154 ,mul_113_23_n_48);
  or mul_113_23_g1985(mul_113_23_n_200 ,mul_113_23_n_146 ,mul_113_23_n_37);
  and mul_113_23_g1986(mul_113_23_n_199 ,in31[3] ,mul_113_23_n_122);
  or mul_113_23_g1987(mul_113_23_n_198 ,mul_113_23_n_55 ,mul_113_23_n_35);
  or mul_113_23_g1988(mul_113_23_n_197 ,mul_113_23_n_58 ,mul_113_23_n_11);
  or mul_113_23_g1989(mul_113_23_n_196 ,mul_113_23_n_141 ,mul_113_23_n_45);
  and mul_113_23_g1990(mul_113_23_n_195 ,in31[2] ,n_341);
  or mul_113_23_g1991(mul_113_23_n_194 ,mul_113_23_n_64 ,mul_113_23_n_82);
  or mul_113_23_g1992(mul_113_23_n_193 ,mul_113_23_n_143 ,mul_113_23_n_42);
  or mul_113_23_g1993(mul_113_23_n_192 ,mul_113_23_n_139 ,mul_113_23_n_39);
  and mul_113_23_g1994(mul_113_23_n_190 ,in31[2] ,mul_113_23_n_72);
  or mul_113_23_g1995(mul_113_23_n_189 ,mul_113_23_n_51 ,mul_113_23_n_85);
  or mul_113_23_g1996(mul_113_23_n_188 ,mul_113_23_n_146 ,mul_113_23_n_20);
  or mul_113_23_g1997(mul_113_23_n_187 ,mul_113_23_n_149 ,mul_113_23_n_16);
  or mul_113_23_g1998(mul_113_23_n_186 ,mul_113_23_n_152 ,mul_113_23_n_33);
  and mul_113_23_g1999(mul_113_23_n_184 ,in31[2] ,mul_113_23_n_67);
  or mul_113_23_g2000(mul_113_23_n_183 ,mul_113_23_n_60 ,mul_113_23_n_18);
  and mul_113_23_g2001(mul_113_23_n_181 ,in31[9] ,mul_113_23_n_73);
  and mul_113_23_g2002(mul_113_23_n_179 ,in31[4] ,mul_113_23_n_68);
  and mul_113_23_g2003(mul_113_23_n_177 ,in31[5] ,mul_113_23_n_73);
  and mul_113_23_g2004(mul_113_23_n_175 ,in31[15] ,n_342);
  and mul_113_23_g2005(mul_113_23_n_173 ,in31[7] ,mul_113_23_n_124);
  or mul_113_23_g2006(mul_113_23_n_172 ,mul_113_23_n_54 ,mul_113_23_n_8);
  or mul_113_23_g2007(mul_113_23_n_171 ,mul_113_23_n_145 ,mul_113_23_n_23);
  and mul_113_23_g2008(mul_113_23_n_169 ,in31[14] ,n_342);
  and mul_113_23_g2009(mul_113_23_n_167 ,in31[10] ,mul_113_23_n_68);
  and mul_113_23_g2010(mul_113_23_n_165 ,in31[15] ,mul_113_23_n_66);
  or mul_113_23_g2011(mul_113_23_n_164 ,mul_113_23_n_139 ,mul_113_23_n_84);
  or mul_113_23_g2012(mul_113_23_n_163 ,mul_113_23_n_57 ,mul_113_23_n_13);
  and mul_113_23_g2013(mul_113_23_n_161 ,in31[5] ,mul_113_23_n_66);
  or mul_113_23_g2014(mul_113_23_n_160 ,mul_113_23_n_144 ,mul_113_23_n_42);
  or mul_113_23_g2015(mul_113_23_n_159 ,mul_113_23_n_63 ,mul_113_23_n_43);
  or mul_113_23_g2016(mul_113_23_n_158 ,mul_113_23_n_155 ,mul_113_23_n_46);
  and mul_113_23_g2017(mul_113_23_n_156 ,in31[3] ,mul_113_23_n_72);
  not mul_113_23_g2018(mul_113_23_n_155 ,in31[1]);
  not mul_113_23_g2019(mul_113_23_n_154 ,in31[5]);
  not mul_113_23_g2020(mul_113_23_n_153 ,in31[2]);
  not mul_113_23_g2021(mul_113_23_n_152 ,in31[13]);
  not mul_113_23_g2022(mul_113_23_n_151 ,in31[11]);
  not mul_113_23_g2023(mul_113_23_n_150 ,in31[6]);
  not mul_113_23_g2024(mul_113_23_n_149 ,in31[7]);
  not mul_113_23_g2025(mul_113_23_n_148 ,n_341);
  not mul_113_23_g2028(mul_113_23_n_147 ,in31[0]);
  not mul_113_23_g2029(mul_113_23_n_146 ,in31[12]);
  not mul_113_23_g2030(mul_113_23_n_145 ,in31[9]);
  not mul_113_23_g2031(mul_113_23_n_144 ,in31[4]);
  not mul_113_23_g2032(mul_113_23_n_143 ,in31[8]);
  not mul_113_23_g2033(mul_113_23_n_142 ,in31[15]);
  not mul_113_23_g2034(mul_113_23_n_141 ,in31[3]);
  not mul_113_23_g2035(mul_113_23_n_140 ,in31[10]);
  not mul_113_23_g2036(mul_113_23_n_139 ,in31[14]);
  not mul_113_23_g2037(mul_113_23_n_138 ,mul_113_23_n_122);
  not mul_113_23_g2038(mul_113_23_n_137 ,n_342);
  not mul_113_23_drc_bufs2056(mul_113_23_n_133 ,mul_113_23_n_131);
  not mul_113_23_drc_bufs2057(mul_113_23_n_132 ,mul_113_23_n_131);
  not mul_113_23_drc_bufs2058(mul_113_23_n_131 ,mul_113_23_n_135);
  not mul_113_23_drc_bufs2061(mul_113_23_n_130 ,mul_113_23_n_128);
  not mul_113_23_drc_bufs2062(mul_113_23_n_129 ,mul_113_23_n_128);
  not mul_113_23_drc_bufs2063(mul_113_23_n_128 ,mul_113_23_n_134);
  not mul_113_23_drc_bufs2066(mul_113_23_n_127 ,mul_113_23_n_126);
  not mul_113_23_drc_bufs2068(mul_113_23_n_126 ,n_343);
  not mul_113_23_drc_bufs2070(mul_113_23_n_125 ,mul_113_23_n_123);
  not mul_113_23_drc_bufs2071(mul_113_23_n_124 ,mul_113_23_n_123);
  not mul_113_23_drc_bufs2072(mul_113_23_n_123 ,n_344);
  not mul_113_23_drc_bufs2098(mul_113_23_n_122 ,mul_113_23_n_120);
  not mul_113_23_drc_bufs2099(mul_113_23_n_121 ,mul_113_23_n_120);
  not mul_113_23_drc_bufs2100(mul_113_23_n_120 ,n_340);
  not mul_113_23_drc_bufs2103(mul_113_23_n_119 ,mul_113_23_n_118);
  not mul_113_23_drc_bufs2104(mul_113_23_n_118 ,mul_113_23_n_155);
  not mul_113_23_drc_bufs2107(mul_113_23_n_117 ,mul_113_23_n_116);
  not mul_113_23_drc_bufs2108(mul_113_23_n_116 ,mul_113_23_n_149);
  not mul_113_23_drc_bufs2111(mul_113_23_n_115 ,mul_113_23_n_114);
  not mul_113_23_drc_bufs2112(mul_113_23_n_114 ,mul_113_23_n_145);
  not mul_113_23_drc_bufs2115(mul_113_23_n_113 ,mul_113_23_n_112);
  not mul_113_23_drc_bufs2116(mul_113_23_n_112 ,mul_113_23_n_139);
  not mul_113_23_drc_bufs2119(mul_113_23_n_111 ,mul_113_23_n_110);
  not mul_113_23_drc_bufs2120(mul_113_23_n_110 ,mul_113_23_n_140);
  buf mul_113_23_drc_bufs2122(n_339 ,mul_113_23_n_664);
  buf mul_113_23_drc_bufs2123(n_334 ,mul_113_23_n_650);
  buf mul_113_23_drc_bufs2124(n_333 ,mul_113_23_n_647);
  buf mul_113_23_drc_bufs2125(n_331 ,mul_113_23_n_641);
  buf mul_113_23_drc_bufs2126(n_332 ,mul_113_23_n_644);
  buf mul_113_23_drc_bufs2127(n_337 ,mul_113_23_n_660);
  buf mul_113_23_drc_bufs2128(n_335 ,mul_113_23_n_653);
  buf mul_113_23_drc_bufs2129(n_336 ,mul_113_23_n_656);
  buf mul_113_23_drc_bufs2130(n_327 ,mul_113_23_n_629);
  buf mul_113_23_drc_bufs2131(n_329 ,mul_113_23_n_635);
  buf mul_113_23_drc_bufs2132(n_328 ,mul_113_23_n_632);
  buf mul_113_23_drc_bufs2133(n_330 ,mul_113_23_n_638);
  not mul_113_23_drc_bufs2134(mul_113_23_n_97 ,mul_113_23_n_95);
  not mul_113_23_drc_bufs2135(mul_113_23_n_96 ,mul_113_23_n_95);
  not mul_113_23_drc_bufs2136(mul_113_23_n_95 ,mul_113_23_n_137);
  not mul_113_23_drc_bufs2138(mul_113_23_n_94 ,mul_113_23_n_92);
  not mul_113_23_drc_bufs2139(mul_113_23_n_93 ,mul_113_23_n_92);
  not mul_113_23_drc_bufs2140(mul_113_23_n_92 ,mul_113_23_n_137);
  not mul_113_23_drc_bufs2142(mul_113_23_n_91 ,mul_113_23_n_89);
  not mul_113_23_drc_bufs2143(mul_113_23_n_90 ,mul_113_23_n_89);
  not mul_113_23_drc_bufs2144(mul_113_23_n_89 ,mul_113_23_n_148);
  not mul_113_23_drc_bufs2146(mul_113_23_n_88 ,mul_113_23_n_86);
  not mul_113_23_drc_bufs2147(mul_113_23_n_87 ,mul_113_23_n_86);
  not mul_113_23_drc_bufs2148(mul_113_23_n_86 ,mul_113_23_n_148);
  not mul_113_23_drc_bufs2154(mul_113_23_n_85 ,mul_113_23_n_83);
  not mul_113_23_drc_bufs2155(mul_113_23_n_84 ,mul_113_23_n_83);
  not mul_113_23_drc_bufs2156(mul_113_23_n_83 ,mul_113_23_n_138);
  not mul_113_23_drc_bufs2158(mul_113_23_n_82 ,mul_113_23_n_80);
  not mul_113_23_drc_bufs2159(mul_113_23_n_81 ,mul_113_23_n_80);
  not mul_113_23_drc_bufs2160(mul_113_23_n_80 ,mul_113_23_n_138);
  not mul_113_23_drc_bufs2163(mul_113_23_n_79 ,mul_113_23_n_78);
  not mul_113_23_drc_bufs2164(mul_113_23_n_78 ,mul_113_23_n_132);
  not mul_113_23_drc_bufs2167(mul_113_23_n_77 ,mul_113_23_n_76);
  not mul_113_23_drc_bufs2168(mul_113_23_n_76 ,mul_113_23_n_130);
  not mul_113_23_drc_bufs2171(mul_113_23_n_75 ,mul_113_23_n_74);
  not mul_113_23_drc_bufs2172(mul_113_23_n_74 ,mul_113_23_n_129);
  not mul_113_23_drc_bufs2174(mul_113_23_n_73 ,mul_113_23_n_71);
  not mul_113_23_drc_bufs2175(mul_113_23_n_72 ,mul_113_23_n_71);
  not mul_113_23_drc_bufs2176(mul_113_23_n_71 ,mul_113_23_n_127);
  not mul_113_23_drc_bufs2179(mul_113_23_n_70 ,mul_113_23_n_69);
  not mul_113_23_drc_bufs2180(mul_113_23_n_69 ,mul_113_23_n_207);
  not mul_113_23_drc_bufs2183(mul_113_23_n_68 ,mul_113_23_n_134);
  not mul_113_23_drc_bufs2184(mul_113_23_n_134 ,mul_113_23_n_127);
  not mul_113_23_drc_bufs2187(mul_113_23_n_67 ,mul_113_23_n_135);
  not mul_113_23_drc_bufs2188(mul_113_23_n_135 ,mul_113_23_n_125);
  not mul_113_23_drc_bufs2190(mul_113_23_n_66 ,mul_113_23_n_65);
  not mul_113_23_drc_bufs2192(mul_113_23_n_65 ,mul_113_23_n_124);
  not mul_113_23_drc_bufs2194(mul_113_23_n_64 ,mul_113_23_n_62);
  not mul_113_23_drc_bufs2195(mul_113_23_n_63 ,mul_113_23_n_62);
  not mul_113_23_drc_bufs2196(mul_113_23_n_62 ,mul_113_23_n_146);
  not mul_113_23_drc_bufs2198(mul_113_23_n_61 ,mul_113_23_n_59);
  not mul_113_23_drc_bufs2199(mul_113_23_n_60 ,mul_113_23_n_59);
  not mul_113_23_drc_bufs2200(mul_113_23_n_59 ,mul_113_23_n_151);
  not mul_113_23_drc_bufs2202(mul_113_23_n_58 ,mul_113_23_n_56);
  not mul_113_23_drc_bufs2203(mul_113_23_n_57 ,mul_113_23_n_56);
  not mul_113_23_drc_bufs2204(mul_113_23_n_56 ,mul_113_23_n_152);
  not mul_113_23_drc_bufs2206(mul_113_23_n_55 ,mul_113_23_n_53);
  not mul_113_23_drc_bufs2207(mul_113_23_n_54 ,mul_113_23_n_53);
  not mul_113_23_drc_bufs2208(mul_113_23_n_53 ,mul_113_23_n_143);
  not mul_113_23_drc_bufs2210(mul_113_23_n_52 ,mul_113_23_n_50);
  not mul_113_23_drc_bufs2211(mul_113_23_n_51 ,mul_113_23_n_50);
  not mul_113_23_drc_bufs2212(mul_113_23_n_50 ,mul_113_23_n_150);
  not mul_113_23_drc_bufs2214(mul_113_23_n_49 ,mul_113_23_n_47);
  not mul_113_23_drc_bufs2215(mul_113_23_n_48 ,mul_113_23_n_47);
  not mul_113_23_drc_bufs2216(mul_113_23_n_47 ,mul_113_23_n_97);
  not mul_113_23_drc_bufs2218(mul_113_23_n_46 ,mul_113_23_n_44);
  not mul_113_23_drc_bufs2219(mul_113_23_n_45 ,mul_113_23_n_44);
  not mul_113_23_drc_bufs2220(mul_113_23_n_44 ,mul_113_23_n_94);
  not mul_113_23_drc_bufs2222(mul_113_23_n_43 ,mul_113_23_n_41);
  not mul_113_23_drc_bufs2223(mul_113_23_n_42 ,mul_113_23_n_41);
  not mul_113_23_drc_bufs2224(mul_113_23_n_41 ,mul_113_23_n_91);
  not mul_113_23_drc_bufs2226(mul_113_23_n_40 ,mul_113_23_n_38);
  not mul_113_23_drc_bufs2227(mul_113_23_n_39 ,mul_113_23_n_38);
  not mul_113_23_drc_bufs2228(mul_113_23_n_38 ,mul_113_23_n_88);
  not mul_113_23_drc_bufs2230(mul_113_23_n_37 ,mul_113_23_n_36);
  not mul_113_23_drc_bufs2232(mul_113_23_n_36 ,mul_113_23_n_93);
  not mul_113_23_drc_bufs2234(mul_113_23_n_35 ,mul_113_23_n_34);
  not mul_113_23_drc_bufs2236(mul_113_23_n_34 ,mul_113_23_n_96);
  not mul_113_23_drc_bufs2238(mul_113_23_n_33 ,mul_113_23_n_32);
  not mul_113_23_drc_bufs2240(mul_113_23_n_32 ,mul_113_23_n_84);
  not mul_113_23_drc_bufs2242(mul_113_23_n_31 ,mul_113_23_n_30);
  not mul_113_23_drc_bufs2244(mul_113_23_n_30 ,mul_113_23_n_85);
  not mul_113_23_drc_bufs2246(mul_113_23_n_29 ,mul_113_23_n_27);
  not mul_113_23_drc_bufs2247(mul_113_23_n_28 ,mul_113_23_n_27);
  not mul_113_23_drc_bufs2248(mul_113_23_n_27 ,mul_113_23_n_133);
  not mul_113_23_drc_bufs2250(mul_113_23_n_26 ,mul_113_23_n_24);
  not mul_113_23_drc_bufs2251(mul_113_23_n_25 ,mul_113_23_n_24);
  not mul_113_23_drc_bufs2252(mul_113_23_n_24 ,mul_113_23_n_133);
  not mul_113_23_drc_bufs2254(mul_113_23_n_23 ,mul_113_23_n_22);
  not mul_113_23_drc_bufs2256(mul_113_23_n_22 ,mul_113_23_n_87);
  not mul_113_23_drc_bufs2258(mul_113_23_n_21 ,mul_113_23_n_19);
  not mul_113_23_drc_bufs2259(mul_113_23_n_20 ,mul_113_23_n_19);
  not mul_113_23_drc_bufs2260(mul_113_23_n_19 ,mul_113_23_n_129);
  not mul_113_23_drc_bufs2262(mul_113_23_n_18 ,mul_113_23_n_17);
  not mul_113_23_drc_bufs2264(mul_113_23_n_17 ,mul_113_23_n_90);
  not mul_113_23_drc_bufs2266(mul_113_23_n_16 ,mul_113_23_n_15);
  not mul_113_23_drc_bufs2268(mul_113_23_n_15 ,mul_113_23_n_81);
  not mul_113_23_drc_bufs2270(mul_113_23_n_14 ,mul_113_23_n_12);
  not mul_113_23_drc_bufs2271(mul_113_23_n_13 ,mul_113_23_n_12);
  not mul_113_23_drc_bufs2272(mul_113_23_n_12 ,mul_113_23_n_130);
  not mul_113_23_drc_bufs2274(mul_113_23_n_11 ,mul_113_23_n_9);
  not mul_113_23_drc_bufs2275(mul_113_23_n_10 ,mul_113_23_n_9);
  not mul_113_23_drc_bufs2276(mul_113_23_n_9 ,mul_113_23_n_132);
  not mul_113_23_drc_bufs2278(mul_113_23_n_8 ,mul_113_23_n_7);
  not mul_113_23_drc_bufs2280(mul_113_23_n_7 ,mul_113_23_n_82);
  and mul_113_23_g2(mul_113_23_n_6 ,mul_113_23_n_488 ,mul_113_23_n_532);
  xor mul_113_23_g2282(mul_113_23_n_5 ,mul_113_23_n_377 ,mul_113_23_n_334);
  xor mul_113_23_g2283(mul_113_23_n_4 ,mul_113_23_n_259 ,mul_113_23_n_206);
  xor mul_113_23_g2284(mul_113_23_n_3 ,mul_113_23_n_255 ,mul_113_23_n_205);
  xor mul_113_23_g2285(mul_113_23_n_2 ,mul_113_23_n_204 ,mul_113_23_n_223);
  xnor mul_113_23_g2286(mul_113_23_n_1 ,mul_113_23_n_195 ,mul_113_23_n_199);
  xor mul_113_23_g2287(mul_113_23_n_0 ,mul_113_23_n_188 ,mul_113_23_n_69);
  or sub_112_23_g97(n_344 ,sub_112_23_n_9 ,sub_112_23_n_23);
  xnor sub_112_23_g98(n_343 ,sub_112_23_n_22 ,sub_112_23_n_14);
  and sub_112_23_g99(sub_112_23_n_23 ,sub_112_23_n_10 ,sub_112_23_n_22);
  and sub_112_23_g100(sub_112_23_n_22 ,sub_112_23_n_12 ,sub_112_23_n_20);
  xnor sub_112_23_g101(sub_112_23_n_21 ,sub_112_23_n_18 ,sub_112_23_n_13);
  or sub_112_23_g102(sub_112_23_n_20 ,sub_112_23_n_7 ,sub_112_23_n_18);
  xnor sub_112_23_g103(n_341 ,sub_112_23_n_8 ,sub_112_23_n_15);
  and sub_112_23_g104(sub_112_23_n_18 ,sub_112_23_n_6 ,sub_112_23_n_17);
  or sub_112_23_g105(sub_112_23_n_17 ,sub_112_23_n_11 ,sub_112_23_n_8);
  xor sub_112_23_g106(n_340 ,in32[0] ,in33[0]);
  xnor sub_112_23_g107(sub_112_23_n_15 ,in32[1] ,in33[1]);
  xnor sub_112_23_g108(sub_112_23_n_14 ,in32[3] ,in33[3]);
  xnor sub_112_23_g109(sub_112_23_n_13 ,in32[2] ,in33[2]);
  or sub_112_23_g110(sub_112_23_n_12 ,sub_112_23_n_4 ,in33[2]);
  nor sub_112_23_g111(sub_112_23_n_11 ,sub_112_23_n_5 ,in32[1]);
  or sub_112_23_g112(sub_112_23_n_10 ,sub_112_23_n_3 ,in33[3]);
  and sub_112_23_g113(sub_112_23_n_9 ,in33[3] ,sub_112_23_n_3);
  and sub_112_23_g114(sub_112_23_n_8 ,in33[0] ,sub_112_23_n_2);
  and sub_112_23_g115(sub_112_23_n_7 ,in33[2] ,sub_112_23_n_4);
  or sub_112_23_g116(sub_112_23_n_6 ,sub_112_23_n_1 ,in33[1]);
  not sub_112_23_g117(sub_112_23_n_5 ,in33[1]);
  not sub_112_23_g118(sub_112_23_n_4 ,in32[2]);
  not sub_112_23_g119(sub_112_23_n_3 ,in32[3]);
  not sub_112_23_g120(sub_112_23_n_2 ,in32[0]);
  not sub_112_23_g121(sub_112_23_n_1 ,in32[1]);
  buf sub_112_23_drc_bufs(n_342 ,sub_112_23_n_21);
  not g6124(csa_tree_add_110_49_pad_groupi_n_421 ,in16[1]);
  not g6125(mul_90_22_n_375 ,in12[1]);
  not g6126(mul_108_22_n_375 ,in24[1]);
  not g6127(mul_102_22_n_375 ,in20[1]);
  not g6128(mul_84_22_n_375 ,in7[1]);
  not g6134(csa_tree_add_117_21_pad_groupi_n_352 ,in4[1]);
  not g6135(csa_tree_add_117_21_pad_groupi_n_354 ,in4[1]);
  buf g6136(csa_tree_add_95_22_pad_groupi_n_708 ,in9[0]);
  buf g6137(csa_tree_add_107_22_pad_groupi_n_708 ,in9[0]);
  buf g6138(csa_tree_add_101_22_pad_groupi_n_708 ,in9[0]);
  buf g6139(csa_tree_add_83_21_pad_groupi_n_708 ,in9[0]);
  not g6140(csa_tree_add_101_22_pad_groupi_n_584 ,in9[15]);
  not g6141(csa_tree_add_95_22_pad_groupi_n_584 ,in9[15]);
  not g6142(csa_tree_add_107_22_pad_groupi_n_584 ,in9[15]);
  not g6143(csa_tree_add_83_21_pad_groupi_n_584 ,in9[15]);
  not g6144(csa_tree_add_89_22_pad_groupi_n_584 ,in9[15]);
  buf g6145(csa_tree_add_95_22_pad_groupi_n_412 ,n_556);
  buf g6146(csa_tree_add_89_22_pad_groupi_n_412 ,n_724);
  buf g6147(csa_tree_add_107_22_pad_groupi_n_412 ,n_586);
  buf g6148(csa_tree_add_101_22_pad_groupi_n_412 ,n_632);
  buf g6149(csa_tree_add_83_21_pad_groupi_n_412 ,n_678);
  buf g6150(csa_tree_add_101_22_pad_groupi_n_978 ,in21[12]);
  buf g6151(csa_tree_add_95_22_pad_groupi_n_978 ,in17[12]);
  buf g6152(csa_tree_add_107_22_pad_groupi_n_978 ,in25[12]);
  buf g6153(csa_tree_add_83_21_pad_groupi_n_978 ,in8[12]);
  buf g6154(csa_tree_add_89_22_pad_groupi_n_978 ,in13[12]);
  buf g6155(csa_tree_add_117_21_pad_groupi_n_269 ,n_469);
  buf g6158(csa_tree_add_95_22_pad_groupi_n_559 ,csa_tree_add_95_22_pad_groupi_n_200);
  buf g6159(csa_tree_add_95_22_pad_groupi_n_567 ,csa_tree_add_95_22_pad_groupi_n_245);
  buf g6160(csa_tree_add_95_22_pad_groupi_n_561 ,csa_tree_add_95_22_pad_groupi_n_62);
  buf g6161(csa_tree_add_95_22_pad_groupi_n_565 ,csa_tree_add_95_22_pad_groupi_n_182);
  buf g6162(csa_tree_add_95_22_pad_groupi_n_569 ,csa_tree_add_95_22_pad_groupi_n_205);
  buf g6165(csa_tree_add_89_22_pad_groupi_n_559 ,csa_tree_add_89_22_pad_groupi_n_200);
  buf g6166(csa_tree_add_89_22_pad_groupi_n_567 ,csa_tree_add_89_22_pad_groupi_n_245);
  buf g6167(csa_tree_add_89_22_pad_groupi_n_561 ,csa_tree_add_89_22_pad_groupi_n_62);
  buf g6168(csa_tree_add_89_22_pad_groupi_n_708 ,in9[0]);
  buf g6169(csa_tree_add_89_22_pad_groupi_n_565 ,csa_tree_add_89_22_pad_groupi_n_182);
  buf g6170(csa_tree_add_89_22_pad_groupi_n_569 ,csa_tree_add_89_22_pad_groupi_n_205);
  buf g6171(csa_tree_add_89_22_pad_groupi_n_570 ,csa_tree_add_89_22_pad_groupi_n_234);
  buf g6174(csa_tree_add_107_22_pad_groupi_n_559 ,csa_tree_add_107_22_pad_groupi_n_200);
  buf g6175(csa_tree_add_107_22_pad_groupi_n_567 ,csa_tree_add_107_22_pad_groupi_n_245);
  buf g6176(csa_tree_add_107_22_pad_groupi_n_561 ,csa_tree_add_107_22_pad_groupi_n_62);
  buf g6177(csa_tree_add_107_22_pad_groupi_n_565 ,csa_tree_add_107_22_pad_groupi_n_182);
  buf g6178(csa_tree_add_107_22_pad_groupi_n_569 ,csa_tree_add_107_22_pad_groupi_n_205);
  buf g6179(csa_tree_add_107_22_pad_groupi_n_570 ,csa_tree_add_107_22_pad_groupi_n_234);
  buf g6182(csa_tree_add_101_22_pad_groupi_n_559 ,csa_tree_add_101_22_pad_groupi_n_200);
  buf g6183(csa_tree_add_101_22_pad_groupi_n_567 ,csa_tree_add_101_22_pad_groupi_n_245);
  buf g6184(csa_tree_add_101_22_pad_groupi_n_561 ,csa_tree_add_101_22_pad_groupi_n_62);
  buf g6185(csa_tree_add_101_22_pad_groupi_n_565 ,csa_tree_add_101_22_pad_groupi_n_182);
  buf g6186(csa_tree_add_101_22_pad_groupi_n_569 ,csa_tree_add_101_22_pad_groupi_n_205);
  buf g6187(csa_tree_add_101_22_pad_groupi_n_570 ,csa_tree_add_101_22_pad_groupi_n_234);
  buf g6190(csa_tree_add_83_21_pad_groupi_n_559 ,csa_tree_add_83_21_pad_groupi_n_200);
  buf g6191(csa_tree_add_83_21_pad_groupi_n_567 ,csa_tree_add_83_21_pad_groupi_n_245);
  buf g6192(csa_tree_add_83_21_pad_groupi_n_561 ,csa_tree_add_83_21_pad_groupi_n_62);
  buf g6193(csa_tree_add_83_21_pad_groupi_n_565 ,csa_tree_add_83_21_pad_groupi_n_182);
  buf g6194(csa_tree_add_83_21_pad_groupi_n_569 ,csa_tree_add_83_21_pad_groupi_n_205);
  buf g6195(csa_tree_add_83_21_pad_groupi_n_570 ,csa_tree_add_83_21_pad_groupi_n_234);
  buf g6196(csa_tree_add_95_22_pad_groupi_n_570 ,csa_tree_add_95_22_pad_groupi_n_234);
  buf g6197(csa_tree_add_101_22_pad_groupi_n_1075 ,csa_tree_add_101_22_pad_groupi_n_978);
  buf g6198(csa_tree_add_101_22_pad_groupi_n_563 ,csa_tree_add_101_22_pad_groupi_n_198);
  not g6200(csa_tree_add_101_22_pad_groupi_n_578 ,csa_tree_add_101_22_pad_groupi_n_161);
  buf g6201(csa_tree_add_101_22_pad_groupi_n_568 ,csa_tree_add_101_22_pad_groupi_n_228);
  buf g6202(csa_tree_add_101_22_pad_groupi_n_572 ,csa_tree_add_101_22_pad_groupi_n_80);
  buf g6203(csa_tree_add_101_22_pad_groupi_n_562 ,csa_tree_add_101_22_pad_groupi_n_224);
  buf g6204(csa_tree_add_95_22_pad_groupi_n_562 ,csa_tree_add_95_22_pad_groupi_n_224);
  buf g6205(csa_tree_add_95_22_pad_groupi_n_572 ,csa_tree_add_95_22_pad_groupi_n_80);
  buf g6206(csa_tree_add_95_22_pad_groupi_n_1075 ,csa_tree_add_95_22_pad_groupi_n_978);
  buf g6207(csa_tree_add_95_22_pad_groupi_n_563 ,csa_tree_add_95_22_pad_groupi_n_198);
  not g6209(csa_tree_add_95_22_pad_groupi_n_578 ,csa_tree_add_95_22_pad_groupi_n_161);
  buf g6210(csa_tree_add_95_22_pad_groupi_n_568 ,csa_tree_add_95_22_pad_groupi_n_228);
  buf g6211(csa_tree_add_107_22_pad_groupi_n_1075 ,csa_tree_add_107_22_pad_groupi_n_978);
  buf g6212(csa_tree_add_107_22_pad_groupi_n_563 ,csa_tree_add_107_22_pad_groupi_n_198);
  not g6214(csa_tree_add_107_22_pad_groupi_n_578 ,csa_tree_add_107_22_pad_groupi_n_161);
  buf g6215(csa_tree_add_107_22_pad_groupi_n_568 ,csa_tree_add_107_22_pad_groupi_n_228);
  buf g6216(csa_tree_add_107_22_pad_groupi_n_572 ,csa_tree_add_107_22_pad_groupi_n_80);
  buf g6217(csa_tree_add_107_22_pad_groupi_n_562 ,csa_tree_add_107_22_pad_groupi_n_224);
  buf g6218(csa_tree_add_83_21_pad_groupi_n_1075 ,csa_tree_add_83_21_pad_groupi_n_978);
  buf g6219(csa_tree_add_83_21_pad_groupi_n_563 ,csa_tree_add_83_21_pad_groupi_n_198);
  not g6221(csa_tree_add_83_21_pad_groupi_n_578 ,csa_tree_add_83_21_pad_groupi_n_161);
  buf g6222(csa_tree_add_83_21_pad_groupi_n_568 ,csa_tree_add_83_21_pad_groupi_n_228);
  buf g6223(csa_tree_add_83_21_pad_groupi_n_572 ,csa_tree_add_83_21_pad_groupi_n_80);
  buf g6224(csa_tree_add_83_21_pad_groupi_n_562 ,csa_tree_add_83_21_pad_groupi_n_224);
  not g6225(csa_tree_add_89_22_pad_groupi_n_578 ,csa_tree_add_89_22_pad_groupi_n_161);
  buf g6226(csa_tree_add_89_22_pad_groupi_n_563 ,csa_tree_add_89_22_pad_groupi_n_198);
  buf g6228(csa_tree_add_89_22_pad_groupi_n_568 ,csa_tree_add_89_22_pad_groupi_n_228);
  buf g6229(csa_tree_add_89_22_pad_groupi_n_572 ,csa_tree_add_89_22_pad_groupi_n_80);
  buf g6230(csa_tree_add_89_22_pad_groupi_n_562 ,csa_tree_add_89_22_pad_groupi_n_224);
  buf g6231(csa_tree_add_117_21_pad_groupi_n_257 ,n_464);
  buf g6234(csa_tree_add_95_22_pad_groupi_n_592 ,csa_tree_add_95_22_pad_groupi_n_559);
  buf g6235(csa_tree_add_95_22_pad_groupi_n_668 ,csa_tree_add_95_22_pad_groupi_n_567);
  buf g6236(csa_tree_add_95_22_pad_groupi_n_664 ,csa_tree_add_95_22_pad_groupi_n_561);
  buf g6237(csa_tree_add_95_22_pad_groupi_n_686 ,csa_tree_add_95_22_pad_groupi_n_565);
  buf g6238(csa_tree_add_95_22_pad_groupi_n_684 ,csa_tree_add_95_22_pad_groupi_n_569);
  buf g6241(csa_tree_add_89_22_pad_groupi_n_592 ,csa_tree_add_89_22_pad_groupi_n_559);
  buf g6242(csa_tree_add_89_22_pad_groupi_n_668 ,csa_tree_add_89_22_pad_groupi_n_567);
  buf g6243(csa_tree_add_89_22_pad_groupi_n_664 ,csa_tree_add_89_22_pad_groupi_n_561);
  buf g6244(csa_tree_add_89_22_pad_groupi_n_686 ,csa_tree_add_89_22_pad_groupi_n_565);
  buf g6245(csa_tree_add_89_22_pad_groupi_n_684 ,csa_tree_add_89_22_pad_groupi_n_569);
  buf g6246(csa_tree_add_89_22_pad_groupi_n_641 ,csa_tree_add_89_22_pad_groupi_n_570);
  buf g6249(csa_tree_add_107_22_pad_groupi_n_592 ,csa_tree_add_107_22_pad_groupi_n_559);
  buf g6250(csa_tree_add_107_22_pad_groupi_n_668 ,csa_tree_add_107_22_pad_groupi_n_567);
  buf g6251(csa_tree_add_107_22_pad_groupi_n_664 ,csa_tree_add_107_22_pad_groupi_n_561);
  buf g6252(csa_tree_add_107_22_pad_groupi_n_686 ,csa_tree_add_107_22_pad_groupi_n_565);
  buf g6253(csa_tree_add_107_22_pad_groupi_n_684 ,csa_tree_add_107_22_pad_groupi_n_569);
  buf g6254(csa_tree_add_107_22_pad_groupi_n_641 ,csa_tree_add_107_22_pad_groupi_n_570);
  buf g6257(csa_tree_add_101_22_pad_groupi_n_592 ,csa_tree_add_101_22_pad_groupi_n_559);
  buf g6258(csa_tree_add_101_22_pad_groupi_n_668 ,csa_tree_add_101_22_pad_groupi_n_567);
  buf g6259(csa_tree_add_101_22_pad_groupi_n_664 ,csa_tree_add_101_22_pad_groupi_n_561);
  buf g6260(csa_tree_add_101_22_pad_groupi_n_686 ,csa_tree_add_101_22_pad_groupi_n_565);
  buf g6261(csa_tree_add_101_22_pad_groupi_n_684 ,csa_tree_add_101_22_pad_groupi_n_569);
  buf g6262(csa_tree_add_101_22_pad_groupi_n_641 ,csa_tree_add_101_22_pad_groupi_n_570);
  buf g6265(csa_tree_add_83_21_pad_groupi_n_592 ,csa_tree_add_83_21_pad_groupi_n_559);
  buf g6266(csa_tree_add_83_21_pad_groupi_n_668 ,csa_tree_add_83_21_pad_groupi_n_567);
  buf g6267(csa_tree_add_83_21_pad_groupi_n_664 ,csa_tree_add_83_21_pad_groupi_n_561);
  buf g6268(csa_tree_add_83_21_pad_groupi_n_686 ,csa_tree_add_83_21_pad_groupi_n_565);
  buf g6269(csa_tree_add_83_21_pad_groupi_n_684 ,csa_tree_add_83_21_pad_groupi_n_569);
  buf g6270(csa_tree_add_83_21_pad_groupi_n_641 ,csa_tree_add_83_21_pad_groupi_n_570);
  buf g6271(csa_tree_add_95_22_pad_groupi_n_641 ,csa_tree_add_95_22_pad_groupi_n_570);
  buf g6272(csa_tree_add_101_22_pad_groupi_n_615 ,csa_tree_add_101_22_pad_groupi_n_563);
  not g6273(csa_tree_add_101_22_pad_groupi_n_829 ,csa_tree_add_101_22_pad_groupi_n_584);
  buf g6274(csa_tree_add_101_22_pad_groupi_n_601 ,csa_tree_add_101_22_pad_groupi_n_568);
  buf g6275(csa_tree_add_101_22_pad_groupi_n_614 ,csa_tree_add_101_22_pad_groupi_n_572);
  buf g6276(csa_tree_add_101_22_pad_groupi_n_678 ,csa_tree_add_101_22_pad_groupi_n_562);
  buf g6277(csa_tree_add_95_22_pad_groupi_n_678 ,csa_tree_add_95_22_pad_groupi_n_562);
  buf g6278(csa_tree_add_95_22_pad_groupi_n_614 ,csa_tree_add_95_22_pad_groupi_n_572);
  buf g6279(csa_tree_add_95_22_pad_groupi_n_615 ,csa_tree_add_95_22_pad_groupi_n_563);
  not g6280(csa_tree_add_95_22_pad_groupi_n_829 ,csa_tree_add_95_22_pad_groupi_n_584);
  buf g6281(csa_tree_add_95_22_pad_groupi_n_601 ,csa_tree_add_95_22_pad_groupi_n_568);
  buf g6282(csa_tree_add_107_22_pad_groupi_n_615 ,csa_tree_add_107_22_pad_groupi_n_563);
  not g6283(csa_tree_add_107_22_pad_groupi_n_829 ,csa_tree_add_107_22_pad_groupi_n_584);
  buf g6284(csa_tree_add_107_22_pad_groupi_n_601 ,csa_tree_add_107_22_pad_groupi_n_568);
  buf g6285(csa_tree_add_107_22_pad_groupi_n_614 ,csa_tree_add_107_22_pad_groupi_n_572);
  buf g6286(csa_tree_add_107_22_pad_groupi_n_678 ,csa_tree_add_107_22_pad_groupi_n_562);
  buf g6287(csa_tree_add_83_21_pad_groupi_n_615 ,csa_tree_add_83_21_pad_groupi_n_563);
  not g6288(csa_tree_add_83_21_pad_groupi_n_829 ,csa_tree_add_83_21_pad_groupi_n_584);
  buf g6289(csa_tree_add_83_21_pad_groupi_n_601 ,csa_tree_add_83_21_pad_groupi_n_568);
  buf g6290(csa_tree_add_83_21_pad_groupi_n_614 ,csa_tree_add_83_21_pad_groupi_n_572);
  buf g6291(csa_tree_add_83_21_pad_groupi_n_678 ,csa_tree_add_83_21_pad_groupi_n_562);
  buf g6292(csa_tree_add_89_22_pad_groupi_n_615 ,csa_tree_add_89_22_pad_groupi_n_563);
  not g6293(csa_tree_add_89_22_pad_groupi_n_829 ,csa_tree_add_89_22_pad_groupi_n_584);
  buf g6294(csa_tree_add_89_22_pad_groupi_n_601 ,csa_tree_add_89_22_pad_groupi_n_568);
  buf g6295(csa_tree_add_89_22_pad_groupi_n_614 ,csa_tree_add_89_22_pad_groupi_n_572);
  buf g6296(csa_tree_add_89_22_pad_groupi_n_678 ,csa_tree_add_89_22_pad_groupi_n_562);
  not g6297(csa_tree_add_95_22_pad_groupi_n_780 ,csa_tree_add_95_22_pad_groupi_n_188);
  not g6298(csa_tree_add_95_22_pad_groupi_n_497 ,csa_tree_add_95_22_pad_groupi_n_349);
  not g6299(csa_tree_add_95_22_pad_groupi_n_830 ,csa_tree_add_95_22_pad_groupi_n_51);
  buf g6300(csa_tree_add_95_22_pad_groupi_n_774 ,csa_tree_add_95_22_pad_groupi_n_592);
  buf g6301(csa_tree_add_95_22_pad_groupi_n_740 ,csa_tree_add_95_22_pad_groupi_n_668);
  buf g6303(csa_tree_add_95_22_pad_groupi_n_835 ,csa_tree_add_95_22_pad_groupi_n_686);
  buf g6304(csa_tree_add_95_22_pad_groupi_n_838 ,csa_tree_add_95_22_pad_groupi_n_684);
  not g6305(csa_tree_add_89_22_pad_groupi_n_780 ,csa_tree_add_89_22_pad_groupi_n_188);
  not g6306(csa_tree_add_89_22_pad_groupi_n_497 ,csa_tree_add_89_22_pad_groupi_n_349);
  not g6307(csa_tree_add_89_22_pad_groupi_n_830 ,csa_tree_add_89_22_pad_groupi_n_51);
  buf g6308(csa_tree_add_89_22_pad_groupi_n_774 ,csa_tree_add_89_22_pad_groupi_n_592);
  buf g6309(csa_tree_add_89_22_pad_groupi_n_740 ,csa_tree_add_89_22_pad_groupi_n_668);
  buf g6311(csa_tree_add_89_22_pad_groupi_n_835 ,csa_tree_add_89_22_pad_groupi_n_686);
  buf g6312(csa_tree_add_89_22_pad_groupi_n_838 ,csa_tree_add_89_22_pad_groupi_n_684);
  buf g6313(csa_tree_add_89_22_pad_groupi_n_782 ,csa_tree_add_89_22_pad_groupi_n_641);
  not g6314(csa_tree_add_107_22_pad_groupi_n_780 ,csa_tree_add_107_22_pad_groupi_n_188);
  not g6315(csa_tree_add_107_22_pad_groupi_n_497 ,csa_tree_add_107_22_pad_groupi_n_349);
  not g6316(csa_tree_add_107_22_pad_groupi_n_830 ,csa_tree_add_107_22_pad_groupi_n_51);
  buf g6317(csa_tree_add_107_22_pad_groupi_n_774 ,csa_tree_add_107_22_pad_groupi_n_592);
  buf g6318(csa_tree_add_107_22_pad_groupi_n_740 ,csa_tree_add_107_22_pad_groupi_n_668);
  buf g6320(csa_tree_add_107_22_pad_groupi_n_835 ,csa_tree_add_107_22_pad_groupi_n_686);
  buf g6321(csa_tree_add_107_22_pad_groupi_n_838 ,csa_tree_add_107_22_pad_groupi_n_684);
  buf g6322(csa_tree_add_107_22_pad_groupi_n_782 ,csa_tree_add_107_22_pad_groupi_n_641);
  not g6323(csa_tree_add_101_22_pad_groupi_n_780 ,csa_tree_add_101_22_pad_groupi_n_188);
  not g6324(csa_tree_add_101_22_pad_groupi_n_497 ,csa_tree_add_101_22_pad_groupi_n_349);
  not g6325(csa_tree_add_101_22_pad_groupi_n_830 ,csa_tree_add_101_22_pad_groupi_n_51);
  buf g6326(csa_tree_add_101_22_pad_groupi_n_774 ,csa_tree_add_101_22_pad_groupi_n_592);
  buf g6327(csa_tree_add_101_22_pad_groupi_n_740 ,csa_tree_add_101_22_pad_groupi_n_668);
  buf g6329(csa_tree_add_101_22_pad_groupi_n_835 ,csa_tree_add_101_22_pad_groupi_n_686);
  buf g6330(csa_tree_add_101_22_pad_groupi_n_838 ,csa_tree_add_101_22_pad_groupi_n_684);
  buf g6331(csa_tree_add_101_22_pad_groupi_n_782 ,csa_tree_add_101_22_pad_groupi_n_641);
  not g6332(csa_tree_add_83_21_pad_groupi_n_780 ,csa_tree_add_83_21_pad_groupi_n_188);
  not g6333(csa_tree_add_83_21_pad_groupi_n_497 ,csa_tree_add_83_21_pad_groupi_n_349);
  not g6334(csa_tree_add_83_21_pad_groupi_n_830 ,csa_tree_add_83_21_pad_groupi_n_51);
  buf g6335(csa_tree_add_83_21_pad_groupi_n_774 ,csa_tree_add_83_21_pad_groupi_n_592);
  buf g6336(csa_tree_add_83_21_pad_groupi_n_740 ,csa_tree_add_83_21_pad_groupi_n_668);
  buf g6338(csa_tree_add_83_21_pad_groupi_n_835 ,csa_tree_add_83_21_pad_groupi_n_686);
  buf g6339(csa_tree_add_83_21_pad_groupi_n_838 ,csa_tree_add_83_21_pad_groupi_n_684);
  buf g6340(csa_tree_add_83_21_pad_groupi_n_782 ,csa_tree_add_83_21_pad_groupi_n_641);
  buf g6341(csa_tree_add_95_22_pad_groupi_n_782 ,csa_tree_add_95_22_pad_groupi_n_641);
  buf g6342(csa_tree_add_101_22_pad_groupi_n_828 ,csa_tree_add_101_22_pad_groupi_n_615);
  buf g6343(csa_tree_add_101_22_pad_groupi_n_822 ,csa_tree_add_101_22_pad_groupi_n_601);
  buf g6344(csa_tree_add_101_22_pad_groupi_n_566 ,csa_tree_add_101_22_pad_groupi_n_68);
  buf g6345(csa_tree_add_101_22_pad_groupi_n_766 ,csa_tree_add_101_22_pad_groupi_n_614);
  buf g6346(csa_tree_add_101_22_pad_groupi_n_831 ,csa_tree_add_101_22_pad_groupi_n_678);
  buf g6347(csa_tree_add_95_22_pad_groupi_n_831 ,csa_tree_add_95_22_pad_groupi_n_678);
  buf g6348(csa_tree_add_95_22_pad_groupi_n_766 ,csa_tree_add_95_22_pad_groupi_n_614);
  buf g6349(csa_tree_add_95_22_pad_groupi_n_828 ,csa_tree_add_95_22_pad_groupi_n_615);
  buf g6350(csa_tree_add_95_22_pad_groupi_n_822 ,csa_tree_add_95_22_pad_groupi_n_601);
  buf g6351(csa_tree_add_95_22_pad_groupi_n_566 ,csa_tree_add_95_22_pad_groupi_n_68);
  buf g6352(csa_tree_add_107_22_pad_groupi_n_828 ,csa_tree_add_107_22_pad_groupi_n_615);
  buf g6353(csa_tree_add_107_22_pad_groupi_n_822 ,csa_tree_add_107_22_pad_groupi_n_601);
  buf g6354(csa_tree_add_107_22_pad_groupi_n_566 ,csa_tree_add_107_22_pad_groupi_n_68);
  buf g6355(csa_tree_add_107_22_pad_groupi_n_766 ,csa_tree_add_107_22_pad_groupi_n_614);
  buf g6356(csa_tree_add_107_22_pad_groupi_n_831 ,csa_tree_add_107_22_pad_groupi_n_678);
  buf g6357(csa_tree_add_83_21_pad_groupi_n_828 ,csa_tree_add_83_21_pad_groupi_n_615);
  buf g6358(csa_tree_add_83_21_pad_groupi_n_822 ,csa_tree_add_83_21_pad_groupi_n_601);
  buf g6359(csa_tree_add_83_21_pad_groupi_n_566 ,csa_tree_add_83_21_pad_groupi_n_68);
  buf g6360(csa_tree_add_83_21_pad_groupi_n_766 ,csa_tree_add_83_21_pad_groupi_n_614);
  buf g6361(csa_tree_add_83_21_pad_groupi_n_831 ,csa_tree_add_83_21_pad_groupi_n_678);
  buf g6362(csa_tree_add_89_22_pad_groupi_n_828 ,csa_tree_add_89_22_pad_groupi_n_615);
  buf g6363(csa_tree_add_89_22_pad_groupi_n_822 ,csa_tree_add_89_22_pad_groupi_n_601);
  buf g6364(csa_tree_add_89_22_pad_groupi_n_566 ,csa_tree_add_89_22_pad_groupi_n_68);
  buf g6365(csa_tree_add_89_22_pad_groupi_n_766 ,csa_tree_add_89_22_pad_groupi_n_614);
  buf g6366(csa_tree_add_89_22_pad_groupi_n_831 ,csa_tree_add_89_22_pad_groupi_n_678);
  buf g6368(csa_tree_add_95_22_pad_groupi_n_802 ,csa_tree_add_95_22_pad_groupi_n_664);
  buf g6370(csa_tree_add_89_22_pad_groupi_n_802 ,csa_tree_add_89_22_pad_groupi_n_664);
  buf g6372(csa_tree_add_107_22_pad_groupi_n_802 ,csa_tree_add_107_22_pad_groupi_n_664);
  buf g6374(csa_tree_add_101_22_pad_groupi_n_802 ,csa_tree_add_101_22_pad_groupi_n_664);
  buf g6376(csa_tree_add_83_21_pad_groupi_n_802 ,csa_tree_add_83_21_pad_groupi_n_664);
  buf g6377(csa_tree_add_101_22_pad_groupi_n_630 ,csa_tree_add_101_22_pad_groupi_n_566);
  buf g6378(csa_tree_add_95_22_pad_groupi_n_630 ,csa_tree_add_95_22_pad_groupi_n_566);
  buf g6379(csa_tree_add_107_22_pad_groupi_n_630 ,csa_tree_add_107_22_pad_groupi_n_566);
  buf g6380(csa_tree_add_83_21_pad_groupi_n_630 ,csa_tree_add_83_21_pad_groupi_n_566);
  buf g6381(csa_tree_add_89_22_pad_groupi_n_630 ,csa_tree_add_89_22_pad_groupi_n_566);
  not g6382(csa_tree_add_95_22_pad_groupi_n_770 ,csa_tree_add_95_22_pad_groupi_n_58);
  not g6383(csa_tree_add_89_22_pad_groupi_n_770 ,csa_tree_add_89_22_pad_groupi_n_58);
  not g6384(csa_tree_add_107_22_pad_groupi_n_770 ,csa_tree_add_107_22_pad_groupi_n_58);
  not g6385(csa_tree_add_101_22_pad_groupi_n_770 ,csa_tree_add_101_22_pad_groupi_n_58);
  not g6386(csa_tree_add_83_21_pad_groupi_n_770 ,csa_tree_add_83_21_pad_groupi_n_58);
  buf g6387(csa_tree_add_101_22_pad_groupi_n_836 ,csa_tree_add_101_22_pad_groupi_n_630);
  buf g6388(csa_tree_add_95_22_pad_groupi_n_836 ,csa_tree_add_95_22_pad_groupi_n_630);
  buf g6389(csa_tree_add_107_22_pad_groupi_n_836 ,csa_tree_add_107_22_pad_groupi_n_630);
  buf g6390(csa_tree_add_83_21_pad_groupi_n_836 ,csa_tree_add_83_21_pad_groupi_n_630);
  buf g6391(csa_tree_add_89_22_pad_groupi_n_836 ,csa_tree_add_89_22_pad_groupi_n_630);
  not g6392(csa_tree_add_95_22_pad_groupi_n_459 ,csa_tree_add_95_22_pad_groupi_n_259);
  not g6393(csa_tree_add_89_22_pad_groupi_n_459 ,csa_tree_add_89_22_pad_groupi_n_259);
  not g6394(csa_tree_add_107_22_pad_groupi_n_459 ,csa_tree_add_107_22_pad_groupi_n_259);
  not g6395(csa_tree_add_101_22_pad_groupi_n_459 ,csa_tree_add_101_22_pad_groupi_n_259);
  not g6396(csa_tree_add_83_21_pad_groupi_n_459 ,csa_tree_add_83_21_pad_groupi_n_259);
  buf g6397(csa_tree_add_117_21_pad_groupi_n_341 ,csa_tree_add_117_21_pad_groupi_n_314);
  buf g6398(csa_tree_add_117_21_pad_groupi_n_550 ,csa_tree_add_117_21_pad_groupi_n_396);
  buf g6399(csa_tree_add_117_21_pad_groupi_n_710 ,csa_tree_add_117_21_pad_groupi_n_600);
  buf g6400(csa_tree_add_117_21_pad_groupi_n_554 ,csa_tree_add_117_21_pad_groupi_n_378);
  buf g6401(csa_tree_add_117_21_pad_groupi_n_558 ,csa_tree_add_117_21_pad_groupi_n_400);
  buf g6402(csa_tree_add_117_21_pad_groupi_n_556 ,csa_tree_add_117_21_pad_groupi_n_398);
  buf g6403(csa_tree_add_117_21_pad_groupi_n_526 ,csa_tree_add_117_21_pad_groupi_n_355);
  buf g6404(csa_tree_add_117_21_pad_groupi_n_522 ,csa_tree_add_117_21_pad_groupi_n_388);
  buf g6405(csa_tree_add_117_21_pad_groupi_n_564 ,csa_tree_add_117_21_pad_groupi_n_401);
  buf g6406(csa_tree_add_117_21_pad_groupi_n_542 ,csa_tree_add_117_21_pad_groupi_n_403);
  buf g6407(csa_tree_add_117_21_pad_groupi_n_561 ,csa_tree_add_117_21_pad_groupi_n_387);
  buf g6408(csa_tree_add_117_21_pad_groupi_n_567 ,csa_tree_add_117_21_pad_groupi_n_399);
  buf g6409(csa_tree_add_117_21_pad_groupi_n_579 ,csa_tree_add_117_21_pad_groupi_n_423);
  buf g6410(csa_tree_add_117_21_pad_groupi_n_565 ,csa_tree_add_117_21_pad_groupi_n_404);
  buf g6411(csa_tree_add_117_21_pad_groupi_n_537 ,csa_tree_add_117_21_pad_groupi_n_434);
  buf g6412(csa_tree_add_117_21_pad_groupi_n_525 ,csa_tree_add_117_21_pad_groupi_n_402);
  buf g6413(csa_tree_add_117_21_pad_groupi_n_515 ,csa_tree_add_117_21_pad_groupi_n_386);
  not g6414(csa_tree_add_117_21_pad_groupi_n_667 ,csa_tree_add_117_21_pad_groupi_n_554);
  not g6415(csa_tree_add_117_21_pad_groupi_n_709 ,csa_tree_add_117_21_pad_groupi_n_558);
  not g6416(csa_tree_add_117_21_pad_groupi_n_697 ,csa_tree_add_117_21_pad_groupi_n_556);
  not g6417(csa_tree_add_117_21_pad_groupi_n_703 ,csa_tree_add_117_21_pad_groupi_n_526);
  not g6418(csa_tree_add_117_21_pad_groupi_n_698 ,csa_tree_add_117_21_pad_groupi_n_522);
  not g6419(csa_tree_add_117_21_pad_groupi_n_706 ,csa_tree_add_117_21_pad_groupi_n_564);
  not g6420(csa_tree_add_117_21_pad_groupi_n_702 ,csa_tree_add_117_21_pad_groupi_n_542);
  not g6421(csa_tree_add_117_21_pad_groupi_n_699 ,csa_tree_add_117_21_pad_groupi_n_561);
  not g6422(csa_tree_add_117_21_pad_groupi_n_713 ,csa_tree_add_117_21_pad_groupi_n_567);
  not g6423(csa_tree_add_117_21_pad_groupi_n_708 ,csa_tree_add_117_21_pad_groupi_n_579);
  not g6424(csa_tree_add_117_21_pad_groupi_n_707 ,csa_tree_add_117_21_pad_groupi_n_565);
  not g6425(csa_tree_add_117_21_pad_groupi_n_705 ,csa_tree_add_117_21_pad_groupi_n_537);
  not g6426(csa_tree_add_117_21_pad_groupi_n_701 ,csa_tree_add_117_21_pad_groupi_n_525);
  not g6427(csa_tree_add_117_21_pad_groupi_n_688 ,csa_tree_add_117_21_pad_groupi_n_515);
  not g6428(csa_tree_add_110_49_pad_groupi_n_467 ,csa_tree_add_110_49_pad_groupi_n_234);
  not g6429(csa_tree_add_110_49_pad_groupi_n_420 ,csa_tree_add_110_49_pad_groupi_n_171);
  not g6430(mul_90_22_n_330 ,mul_90_22_n_164);
  not g6431(mul_108_22_n_330 ,mul_108_22_n_164);
  not g6432(mul_102_22_n_330 ,mul_102_22_n_164);
  not g6433(mul_84_22_n_330 ,mul_84_22_n_164);
  not g6434(add_115_23_pad_n_96 ,add_115_23_pad_n_94);
endmodule
