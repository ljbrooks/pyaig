module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, out1, out2);
  input [15:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61;
  input in62;
  output [28:0] out1;
  output [16:0] out2;
  wire [15:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61;
  wire in62;
  wire [28:0] out1;
  wire [16:0] out2;
  wire add_128_19_n_0, add_128_19_n_1, add_128_19_n_2, add_128_19_n_3, add_128_19_n_4, add_128_19_n_5, add_128_19_n_6, add_128_19_n_7;
  wire add_128_19_n_8, add_128_19_n_9, add_128_19_n_10, add_128_19_n_11, add_128_19_n_12, add_128_19_n_13, add_128_19_n_14, add_128_19_n_15;
  wire add_128_19_n_16, add_128_19_n_17, add_128_19_n_18, add_128_19_n_19, add_128_19_n_20, add_128_19_n_21, add_128_19_n_22, add_128_19_n_23;
  wire add_128_19_n_24, add_128_19_n_25, add_128_19_n_26, add_128_19_n_27, add_128_19_n_28, add_128_19_n_29, add_128_19_n_30, add_128_19_n_31;
  wire add_128_19_n_32, add_128_19_n_33, add_128_19_n_34, add_128_19_n_35, add_128_19_n_36, add_128_19_n_37, add_128_19_n_38, add_128_19_n_39;
  wire add_128_19_n_40, add_128_19_n_41, add_128_19_n_42, add_128_19_n_43, add_128_19_n_44, add_128_19_n_45, add_128_19_n_46, add_128_19_n_47;
  wire add_128_19_n_48, add_128_19_n_49, add_128_19_n_51, add_128_19_n_53, add_128_19_n_55, add_128_19_n_56, add_128_19_n_58, add_128_19_n_59;
  wire add_128_19_n_61, add_128_19_n_62, add_128_19_n_64, add_128_19_n_65, add_128_19_n_67, add_128_19_n_68, add_128_19_n_70, add_128_19_n_71;
  wire add_128_19_n_73, add_128_19_n_74, add_128_19_n_76, add_128_19_n_77, add_128_19_n_79, add_128_19_n_80, add_128_19_n_82, add_128_19_n_83;
  wire add_128_19_n_85, add_128_19_n_86, add_128_19_n_88, add_128_19_n_89, add_128_19_n_91, add_128_19_n_92, add_130_19_n_0, add_130_19_n_1;
  wire add_130_19_n_2, add_130_19_n_3, add_130_19_n_4, add_130_19_n_5, add_130_19_n_6, add_130_19_n_7, add_130_19_n_8, add_130_19_n_9;
  wire add_130_19_n_10, add_130_19_n_11, add_130_19_n_12, add_130_19_n_13, add_130_19_n_14, add_130_19_n_15, add_130_19_n_16, add_130_19_n_17;
  wire add_130_19_n_18, add_130_19_n_19, add_130_19_n_20, add_130_19_n_21, add_130_19_n_22, add_130_19_n_23, add_130_19_n_24, add_130_19_n_25;
  wire add_130_19_n_26, add_130_19_n_27, add_130_19_n_28, add_130_19_n_29, add_130_19_n_30, add_130_19_n_31, add_130_19_n_32, add_130_19_n_33;
  wire add_130_19_n_34, add_130_19_n_35, add_130_19_n_36, add_130_19_n_37, add_130_19_n_38, add_130_19_n_39, add_130_19_n_40, add_130_19_n_41;
  wire add_130_19_n_42, add_130_19_n_43, add_130_19_n_44, add_130_19_n_45, add_130_19_n_46, add_130_19_n_47, add_130_19_n_48, add_130_19_n_49;
  wire add_130_19_n_51, add_130_19_n_53, add_130_19_n_55, add_130_19_n_56, add_130_19_n_58, add_130_19_n_59, add_130_19_n_61, add_130_19_n_62;
  wire add_130_19_n_64, add_130_19_n_65, add_130_19_n_67, add_130_19_n_68, add_130_19_n_70, add_130_19_n_71, add_130_19_n_73, add_130_19_n_74;
  wire add_130_19_n_76, add_130_19_n_77, add_130_19_n_79, add_130_19_n_80, add_130_19_n_82, add_130_19_n_83, add_130_19_n_85, add_130_19_n_86;
  wire add_130_19_n_88, add_130_19_n_89, add_130_19_n_91, add_130_19_n_92, add_132_19_n_0, add_132_19_n_1, add_132_19_n_2, add_132_19_n_3;
  wire add_132_19_n_4, add_132_19_n_5, add_132_19_n_6, add_132_19_n_7, add_132_19_n_8, add_132_19_n_9, add_132_19_n_10, add_132_19_n_11;
  wire add_132_19_n_12, add_132_19_n_13, add_132_19_n_14, add_132_19_n_15, add_132_19_n_16, add_132_19_n_17, add_132_19_n_18, add_132_19_n_19;
  wire add_132_19_n_20, add_132_19_n_21, add_132_19_n_22, add_132_19_n_23, add_132_19_n_24, add_132_19_n_25, add_132_19_n_26, add_132_19_n_27;
  wire add_132_19_n_28, add_132_19_n_29, add_132_19_n_30, add_132_19_n_31, add_132_19_n_32, add_132_19_n_33, add_132_19_n_34, add_132_19_n_35;
  wire add_132_19_n_36, add_132_19_n_37, add_132_19_n_38, add_132_19_n_39, add_132_19_n_40, add_132_19_n_41, add_132_19_n_42, add_132_19_n_43;
  wire add_132_19_n_44, add_132_19_n_45, add_132_19_n_46, add_132_19_n_47, add_132_19_n_48, add_132_19_n_49, add_132_19_n_51, add_132_19_n_53;
  wire add_132_19_n_55, add_132_19_n_56, add_132_19_n_58, add_132_19_n_59, add_132_19_n_61, add_132_19_n_62, add_132_19_n_64, add_132_19_n_65;
  wire add_132_19_n_67, add_132_19_n_68, add_132_19_n_70, add_132_19_n_71, add_132_19_n_73, add_132_19_n_74, add_132_19_n_76, add_132_19_n_77;
  wire add_132_19_n_79, add_132_19_n_80, add_132_19_n_82, add_132_19_n_83, add_132_19_n_85, add_132_19_n_86, add_132_19_n_88, add_132_19_n_89;
  wire add_132_19_n_91, add_132_19_n_92, add_134_19_n_0, add_134_19_n_1, add_134_19_n_2, add_134_19_n_3, add_134_19_n_4, add_134_19_n_5;
  wire add_134_19_n_6, add_134_19_n_7, add_134_19_n_8, add_134_19_n_9, add_134_19_n_10, add_134_19_n_11, add_134_19_n_12, add_134_19_n_13;
  wire add_134_19_n_14, add_134_19_n_15, add_134_19_n_16, add_134_19_n_17, add_134_19_n_18, add_134_19_n_19, add_134_19_n_20, add_134_19_n_21;
  wire add_134_19_n_22, add_134_19_n_23, add_134_19_n_24, add_134_19_n_25, add_134_19_n_26, add_134_19_n_27, add_134_19_n_28, add_134_19_n_29;
  wire add_134_19_n_30, add_134_19_n_31, add_134_19_n_32, add_134_19_n_33, add_134_19_n_34, add_134_19_n_35, add_134_19_n_36, add_134_19_n_37;
  wire add_134_19_n_38, add_134_19_n_39, add_134_19_n_40, add_134_19_n_41, add_134_19_n_42, add_134_19_n_43, add_134_19_n_44, add_134_19_n_45;
  wire add_134_19_n_46, add_134_19_n_47, add_134_19_n_48, add_134_19_n_49, add_134_19_n_51, add_134_19_n_53, add_134_19_n_55, add_134_19_n_56;
  wire add_134_19_n_58, add_134_19_n_59, add_134_19_n_61, add_134_19_n_62, add_134_19_n_64, add_134_19_n_65, add_134_19_n_67, add_134_19_n_68;
  wire add_134_19_n_70, add_134_19_n_71, add_134_19_n_73, add_134_19_n_74, add_134_19_n_76, add_134_19_n_77, add_134_19_n_79, add_134_19_n_80;
  wire add_134_19_n_82, add_134_19_n_83, add_134_19_n_85, add_134_19_n_86, add_134_19_n_88, add_134_19_n_89, add_134_19_n_91, add_134_19_n_92;
  wire add_136_19_n_0, add_136_19_n_1, add_136_19_n_2, add_136_19_n_3, add_136_19_n_4, add_136_19_n_5, add_136_19_n_6, add_136_19_n_7;
  wire add_136_19_n_8, add_136_19_n_9, add_136_19_n_10, add_136_19_n_11, add_136_19_n_12, add_136_19_n_13, add_136_19_n_14, add_136_19_n_15;
  wire add_136_19_n_16, add_136_19_n_17, add_136_19_n_18, add_136_19_n_19, add_136_19_n_20, add_136_19_n_21, add_136_19_n_22, add_136_19_n_23;
  wire add_136_19_n_24, add_136_19_n_25, add_136_19_n_26, add_136_19_n_27, add_136_19_n_28, add_136_19_n_29, add_136_19_n_30, add_136_19_n_31;
  wire add_136_19_n_32, add_136_19_n_33, add_136_19_n_34, add_136_19_n_35, add_136_19_n_36, add_136_19_n_37, add_136_19_n_38, add_136_19_n_39;
  wire add_136_19_n_40, add_136_19_n_41, add_136_19_n_42, add_136_19_n_43, add_136_19_n_44, add_136_19_n_45, add_136_19_n_46, add_136_19_n_47;
  wire add_136_19_n_48, add_136_19_n_49, add_136_19_n_51, add_136_19_n_53, add_136_19_n_55, add_136_19_n_56, add_136_19_n_58, add_136_19_n_59;
  wire add_136_19_n_61, add_136_19_n_62, add_136_19_n_64, add_136_19_n_65, add_136_19_n_67, add_136_19_n_68, add_136_19_n_70, add_136_19_n_71;
  wire add_136_19_n_73, add_136_19_n_74, add_136_19_n_76, add_136_19_n_77, add_136_19_n_79, add_136_19_n_80, add_136_19_n_82, add_136_19_n_83;
  wire add_136_19_n_85, add_136_19_n_86, add_136_19_n_88, add_136_19_n_89, add_136_19_n_91, add_136_19_n_92, add_138_20_n_0, add_138_20_n_1;
  wire add_138_20_n_2, add_138_20_n_3, add_138_20_n_4, add_138_20_n_5, add_138_20_n_6, add_138_20_n_7, add_138_20_n_8, add_138_20_n_9;
  wire add_138_20_n_10, add_138_20_n_11, add_138_20_n_12, add_138_20_n_13, add_138_20_n_14, add_138_20_n_15, add_138_20_n_16, add_138_20_n_17;
  wire add_138_20_n_18, add_138_20_n_19, add_138_20_n_20, add_138_20_n_21, add_138_20_n_22, add_138_20_n_23, add_138_20_n_24, add_138_20_n_25;
  wire add_138_20_n_26, add_138_20_n_27, add_138_20_n_28, add_138_20_n_29, add_138_20_n_30, add_138_20_n_31, add_138_20_n_32, add_138_20_n_33;
  wire add_138_20_n_34, add_138_20_n_35, add_138_20_n_36, add_138_20_n_37, add_138_20_n_38, add_138_20_n_39, add_138_20_n_40, add_138_20_n_41;
  wire add_138_20_n_42, add_138_20_n_43, add_138_20_n_44, add_138_20_n_45, add_138_20_n_46, add_138_20_n_47, add_138_20_n_48, add_138_20_n_49;
  wire add_138_20_n_51, add_138_20_n_53, add_138_20_n_55, add_138_20_n_56, add_138_20_n_58, add_138_20_n_59, add_138_20_n_61, add_138_20_n_62;
  wire add_138_20_n_64, add_138_20_n_65, add_138_20_n_67, add_138_20_n_68, add_138_20_n_70, add_138_20_n_71, add_138_20_n_73, add_138_20_n_74;
  wire add_138_20_n_76, add_138_20_n_77, add_138_20_n_79, add_138_20_n_80, add_138_20_n_82, add_138_20_n_83, add_138_20_n_85, add_138_20_n_86;
  wire add_138_20_n_88, add_138_20_n_89, add_138_20_n_91, add_138_20_n_92, add_140_21_n_0, add_140_21_n_1, add_140_21_n_2, add_140_21_n_3;
  wire add_140_21_n_4, add_140_21_n_5, add_140_21_n_6, add_140_21_n_7, add_140_21_n_8, add_140_21_n_9, add_140_21_n_10, add_140_21_n_11;
  wire add_140_21_n_12, add_140_21_n_13, add_140_21_n_14, add_140_21_n_15, add_140_21_n_16, add_140_21_n_17, add_140_21_n_18, add_140_21_n_19;
  wire add_140_21_n_20, add_140_21_n_21, add_140_21_n_22, add_140_21_n_23, add_140_21_n_24, add_140_21_n_25, add_140_21_n_26, add_140_21_n_27;
  wire add_140_21_n_28, add_140_21_n_29, add_140_21_n_30, add_140_21_n_31, add_140_21_n_32, add_140_21_n_33, add_140_21_n_34, add_140_21_n_35;
  wire add_140_21_n_36, add_140_21_n_37, add_140_21_n_38, add_140_21_n_39, add_140_21_n_40, add_140_21_n_41, add_140_21_n_42, add_140_21_n_43;
  wire add_140_21_n_44, add_140_21_n_45, add_140_21_n_46, add_140_21_n_47, add_140_21_n_48, add_140_21_n_49, add_140_21_n_51, add_140_21_n_53;
  wire add_140_21_n_55, add_140_21_n_56, add_140_21_n_58, add_140_21_n_59, add_140_21_n_61, add_140_21_n_62, add_140_21_n_64, add_140_21_n_65;
  wire add_140_21_n_67, add_140_21_n_68, add_140_21_n_70, add_140_21_n_71, add_140_21_n_73, add_140_21_n_74, add_140_21_n_76, add_140_21_n_77;
  wire add_140_21_n_79, add_140_21_n_80, add_140_21_n_82, add_140_21_n_83, add_140_21_n_85, add_140_21_n_86, add_140_21_n_88, add_140_21_n_89;
  wire add_140_21_n_91, add_140_21_n_92, add_142_21_n_0, add_142_21_n_1, add_142_21_n_2, add_142_21_n_3, add_142_21_n_4, add_142_21_n_5;
  wire add_142_21_n_6, add_142_21_n_7, add_142_21_n_8, add_142_21_n_9, add_142_21_n_10, add_142_21_n_11, add_142_21_n_12, add_142_21_n_13;
  wire add_142_21_n_14, add_142_21_n_15, add_142_21_n_16, add_142_21_n_17, add_142_21_n_18, add_142_21_n_19, add_142_21_n_20, add_142_21_n_21;
  wire add_142_21_n_22, add_142_21_n_23, add_142_21_n_24, add_142_21_n_25, add_142_21_n_26, add_142_21_n_27, add_142_21_n_28, add_142_21_n_29;
  wire add_142_21_n_30, add_142_21_n_31, add_142_21_n_32, add_142_21_n_33, add_142_21_n_34, add_142_21_n_35, add_142_21_n_36, add_142_21_n_37;
  wire add_142_21_n_38, add_142_21_n_39, add_142_21_n_40, add_142_21_n_41, add_142_21_n_42, add_142_21_n_43, add_142_21_n_44, add_142_21_n_45;
  wire add_142_21_n_46, add_142_21_n_47, add_142_21_n_48, add_142_21_n_49, add_142_21_n_51, add_142_21_n_53, add_142_21_n_55, add_142_21_n_56;
  wire add_142_21_n_58, add_142_21_n_59, add_142_21_n_61, add_142_21_n_62, add_142_21_n_64, add_142_21_n_65, add_142_21_n_67, add_142_21_n_68;
  wire add_142_21_n_70, add_142_21_n_71, add_142_21_n_73, add_142_21_n_74, add_142_21_n_76, add_142_21_n_77, add_142_21_n_79, add_142_21_n_80;
  wire add_142_21_n_82, add_142_21_n_83, add_142_21_n_85, add_142_21_n_86, add_142_21_n_88, add_142_21_n_89, add_142_21_n_91, add_142_21_n_92;
  wire add_144_21_n_0, add_144_21_n_1, add_144_21_n_2, add_144_21_n_3, add_144_21_n_4, add_144_21_n_5, add_144_21_n_6, add_144_21_n_7;
  wire add_144_21_n_8, add_144_21_n_9, add_144_21_n_10, add_144_21_n_11, add_144_21_n_12, add_144_21_n_13, add_144_21_n_14, add_144_21_n_15;
  wire add_144_21_n_16, add_144_21_n_17, add_144_21_n_18, add_144_21_n_19, add_144_21_n_20, add_144_21_n_21, add_144_21_n_22, add_144_21_n_23;
  wire add_144_21_n_24, add_144_21_n_25, add_144_21_n_26, add_144_21_n_27, add_144_21_n_28, add_144_21_n_29, add_144_21_n_30, add_144_21_n_31;
  wire add_144_21_n_32, add_144_21_n_33, add_144_21_n_34, add_144_21_n_35, add_144_21_n_36, add_144_21_n_37, add_144_21_n_38, add_144_21_n_39;
  wire add_144_21_n_40, add_144_21_n_41, add_144_21_n_42, add_144_21_n_43, add_144_21_n_44, add_144_21_n_45, add_144_21_n_46, add_144_21_n_47;
  wire add_144_21_n_48, add_144_21_n_49, add_144_21_n_51, add_144_21_n_53, add_144_21_n_55, add_144_21_n_56, add_144_21_n_58, add_144_21_n_59;
  wire add_144_21_n_61, add_144_21_n_62, add_144_21_n_64, add_144_21_n_65, add_144_21_n_67, add_144_21_n_68, add_144_21_n_70, add_144_21_n_71;
  wire add_144_21_n_73, add_144_21_n_74, add_144_21_n_76, add_144_21_n_77, add_144_21_n_79, add_144_21_n_80, add_144_21_n_82, add_144_21_n_83;
  wire add_144_21_n_85, add_144_21_n_86, add_144_21_n_88, add_144_21_n_89, add_144_21_n_91, add_144_21_n_92, add_146_21_n_0, add_146_21_n_1;
  wire add_146_21_n_2, add_146_21_n_3, add_146_21_n_4, add_146_21_n_5, add_146_21_n_6, add_146_21_n_7, add_146_21_n_8, add_146_21_n_9;
  wire add_146_21_n_10, add_146_21_n_11, add_146_21_n_12, add_146_21_n_13, add_146_21_n_14, add_146_21_n_15, add_146_21_n_16, add_146_21_n_17;
  wire add_146_21_n_18, add_146_21_n_19, add_146_21_n_20, add_146_21_n_21, add_146_21_n_22, add_146_21_n_23, add_146_21_n_24, add_146_21_n_25;
  wire add_146_21_n_26, add_146_21_n_27, add_146_21_n_28, add_146_21_n_29, add_146_21_n_30, add_146_21_n_31, add_146_21_n_32, add_146_21_n_33;
  wire add_146_21_n_34, add_146_21_n_35, add_146_21_n_36, add_146_21_n_37, add_146_21_n_38, add_146_21_n_39, add_146_21_n_40, add_146_21_n_41;
  wire add_146_21_n_42, add_146_21_n_43, add_146_21_n_44, add_146_21_n_45, add_146_21_n_46, add_146_21_n_47, add_146_21_n_48, add_146_21_n_49;
  wire add_146_21_n_51, add_146_21_n_53, add_146_21_n_55, add_146_21_n_56, add_146_21_n_58, add_146_21_n_59, add_146_21_n_61, add_146_21_n_62;
  wire add_146_21_n_64, add_146_21_n_65, add_146_21_n_67, add_146_21_n_68, add_146_21_n_70, add_146_21_n_71, add_146_21_n_73, add_146_21_n_74;
  wire add_146_21_n_76, add_146_21_n_77, add_146_21_n_79, add_146_21_n_80, add_146_21_n_82, add_146_21_n_83, add_146_21_n_85, add_146_21_n_86;
  wire add_146_21_n_88, add_146_21_n_89, add_146_21_n_91, add_146_21_n_92, add_148_21_n_0, add_148_21_n_1, add_148_21_n_2, add_148_21_n_3;
  wire add_148_21_n_4, add_148_21_n_5, add_148_21_n_6, add_148_21_n_7, add_148_21_n_8, add_148_21_n_9, add_148_21_n_10, add_148_21_n_11;
  wire add_148_21_n_12, add_148_21_n_13, add_148_21_n_14, add_148_21_n_15, add_148_21_n_16, add_148_21_n_17, add_148_21_n_18, add_148_21_n_19;
  wire add_148_21_n_20, add_148_21_n_21, add_148_21_n_22, add_148_21_n_23, add_148_21_n_24, add_148_21_n_25, add_148_21_n_26, add_148_21_n_27;
  wire add_148_21_n_28, add_148_21_n_29, add_148_21_n_30, add_148_21_n_31, add_148_21_n_32, add_148_21_n_33, add_148_21_n_34, add_148_21_n_35;
  wire add_148_21_n_36, add_148_21_n_37, add_148_21_n_38, add_148_21_n_39, add_148_21_n_40, add_148_21_n_41, add_148_21_n_42, add_148_21_n_43;
  wire add_148_21_n_44, add_148_21_n_45, add_148_21_n_46, add_148_21_n_47, add_148_21_n_48, add_148_21_n_49, add_148_21_n_51, add_148_21_n_53;
  wire add_148_21_n_55, add_148_21_n_56, add_148_21_n_58, add_148_21_n_59, add_148_21_n_61, add_148_21_n_62, add_148_21_n_64, add_148_21_n_65;
  wire add_148_21_n_67, add_148_21_n_68, add_148_21_n_70, add_148_21_n_71, add_148_21_n_73, add_148_21_n_74, add_148_21_n_76, add_148_21_n_77;
  wire add_148_21_n_79, add_148_21_n_80, add_148_21_n_82, add_148_21_n_83, add_148_21_n_85, add_148_21_n_86, add_148_21_n_88, add_148_21_n_89;
  wire add_148_21_n_91, add_148_21_n_92, add_150_21_n_0, add_150_21_n_1, add_150_21_n_2, add_150_21_n_3, add_150_21_n_4, add_150_21_n_5;
  wire add_150_21_n_6, add_150_21_n_7, add_150_21_n_8, add_150_21_n_9, add_150_21_n_10, add_150_21_n_11, add_150_21_n_12, add_150_21_n_13;
  wire add_150_21_n_14, add_150_21_n_15, add_150_21_n_16, add_150_21_n_17, add_150_21_n_18, add_150_21_n_19, add_150_21_n_20, add_150_21_n_21;
  wire add_150_21_n_22, add_150_21_n_23, add_150_21_n_24, add_150_21_n_25, add_150_21_n_26, add_150_21_n_27, add_150_21_n_28, add_150_21_n_29;
  wire add_150_21_n_30, add_150_21_n_31, add_150_21_n_32, add_150_21_n_33, add_150_21_n_34, add_150_21_n_35, add_150_21_n_36, add_150_21_n_37;
  wire add_150_21_n_38, add_150_21_n_39, add_150_21_n_40, add_150_21_n_41, add_150_21_n_42, add_150_21_n_43, add_150_21_n_44, add_150_21_n_45;
  wire add_150_21_n_46, add_150_21_n_47, add_150_21_n_48, add_150_21_n_49, add_150_21_n_51, add_150_21_n_53, add_150_21_n_55, add_150_21_n_56;
  wire add_150_21_n_58, add_150_21_n_59, add_150_21_n_61, add_150_21_n_62, add_150_21_n_64, add_150_21_n_65, add_150_21_n_67, add_150_21_n_68;
  wire add_150_21_n_70, add_150_21_n_71, add_150_21_n_73, add_150_21_n_74, add_150_21_n_76, add_150_21_n_77, add_150_21_n_79, add_150_21_n_80;
  wire add_150_21_n_82, add_150_21_n_83, add_150_21_n_85, add_150_21_n_86, add_150_21_n_88, add_150_21_n_89, add_150_21_n_91, add_150_21_n_92;
  wire add_152_21_n_0, add_152_21_n_1, add_152_21_n_2, add_152_21_n_3, add_152_21_n_4, add_152_21_n_5, add_152_21_n_6, add_152_21_n_7;
  wire add_152_21_n_8, add_152_21_n_9, add_152_21_n_10, add_152_21_n_11, add_152_21_n_12, add_152_21_n_13, add_152_21_n_14, add_152_21_n_15;
  wire add_152_21_n_16, add_152_21_n_17, add_152_21_n_18, add_152_21_n_19, add_152_21_n_20, add_152_21_n_21, add_152_21_n_22, add_152_21_n_23;
  wire add_152_21_n_24, add_152_21_n_25, add_152_21_n_26, add_152_21_n_27, add_152_21_n_28, add_152_21_n_29, add_152_21_n_30, add_152_21_n_31;
  wire add_152_21_n_32, add_152_21_n_33, add_152_21_n_34, add_152_21_n_35, add_152_21_n_36, add_152_21_n_37, add_152_21_n_38, add_152_21_n_39;
  wire add_152_21_n_40, add_152_21_n_41, add_152_21_n_42, add_152_21_n_43, add_152_21_n_44, add_152_21_n_45, add_152_21_n_46, add_152_21_n_47;
  wire add_152_21_n_48, add_152_21_n_49, add_152_21_n_51, add_152_21_n_53, add_152_21_n_55, add_152_21_n_56, add_152_21_n_58, add_152_21_n_59;
  wire add_152_21_n_61, add_152_21_n_62, add_152_21_n_64, add_152_21_n_65, add_152_21_n_67, add_152_21_n_68, add_152_21_n_70, add_152_21_n_71;
  wire add_152_21_n_73, add_152_21_n_74, add_152_21_n_76, add_152_21_n_77, add_152_21_n_79, add_152_21_n_80, add_152_21_n_82, add_152_21_n_83;
  wire add_152_21_n_85, add_152_21_n_86, add_152_21_n_88, add_152_21_n_89, add_152_21_n_91, add_152_21_n_92, add_154_21_n_0, add_154_21_n_1;
  wire add_154_21_n_2, add_154_21_n_3, add_154_21_n_4, add_154_21_n_5, add_154_21_n_6, add_154_21_n_7, add_154_21_n_8, add_154_21_n_9;
  wire add_154_21_n_10, add_154_21_n_11, add_154_21_n_12, add_154_21_n_13, add_154_21_n_14, add_154_21_n_15, add_154_21_n_16, add_154_21_n_17;
  wire add_154_21_n_18, add_154_21_n_19, add_154_21_n_20, add_154_21_n_21, add_154_21_n_22, add_154_21_n_23, add_154_21_n_24, add_154_21_n_25;
  wire add_154_21_n_26, add_154_21_n_27, add_154_21_n_28, add_154_21_n_29, add_154_21_n_30, add_154_21_n_31, add_154_21_n_32, add_154_21_n_33;
  wire add_154_21_n_34, add_154_21_n_35, add_154_21_n_36, add_154_21_n_37, add_154_21_n_38, add_154_21_n_39, add_154_21_n_40, add_154_21_n_41;
  wire add_154_21_n_42, add_154_21_n_43, add_154_21_n_44, add_154_21_n_45, add_154_21_n_46, add_154_21_n_47, add_154_21_n_48, add_154_21_n_49;
  wire add_154_21_n_51, add_154_21_n_53, add_154_21_n_55, add_154_21_n_56, add_154_21_n_58, add_154_21_n_59, add_154_21_n_61, add_154_21_n_62;
  wire add_154_21_n_64, add_154_21_n_65, add_154_21_n_67, add_154_21_n_68, add_154_21_n_70, add_154_21_n_71, add_154_21_n_73, add_154_21_n_74;
  wire add_154_21_n_76, add_154_21_n_77, add_154_21_n_79, add_154_21_n_80, add_154_21_n_82, add_154_21_n_83, add_154_21_n_85, add_154_21_n_86;
  wire add_154_21_n_88, add_154_21_n_89, add_154_21_n_91, add_154_21_n_92, add_156_21_n_0, add_156_21_n_1, add_156_21_n_2, add_156_21_n_3;
  wire add_156_21_n_4, add_156_21_n_5, add_156_21_n_6, add_156_21_n_7, add_156_21_n_8, add_156_21_n_9, add_156_21_n_10, add_156_21_n_11;
  wire add_156_21_n_12, add_156_21_n_13, add_156_21_n_14, add_156_21_n_15, add_156_21_n_16, add_156_21_n_17, add_156_21_n_18, add_156_21_n_19;
  wire add_156_21_n_20, add_156_21_n_21, add_156_21_n_22, add_156_21_n_23, add_156_21_n_24, add_156_21_n_25, add_156_21_n_26, add_156_21_n_27;
  wire add_156_21_n_28, add_156_21_n_29, add_156_21_n_30, add_156_21_n_31, add_156_21_n_32, add_156_21_n_33, add_156_21_n_34, add_156_21_n_35;
  wire add_156_21_n_36, add_156_21_n_37, add_156_21_n_38, add_156_21_n_39, add_156_21_n_40, add_156_21_n_41, add_156_21_n_42, add_156_21_n_43;
  wire add_156_21_n_44, add_156_21_n_45, add_156_21_n_46, add_156_21_n_47, add_156_21_n_48, add_156_21_n_49, add_156_21_n_51, add_156_21_n_53;
  wire add_156_21_n_55, add_156_21_n_56, add_156_21_n_58, add_156_21_n_59, add_156_21_n_61, add_156_21_n_62, add_156_21_n_64, add_156_21_n_65;
  wire add_156_21_n_67, add_156_21_n_68, add_156_21_n_70, add_156_21_n_71, add_156_21_n_73, add_156_21_n_74, add_156_21_n_76, add_156_21_n_77;
  wire add_156_21_n_79, add_156_21_n_80, add_156_21_n_82, add_156_21_n_83, add_156_21_n_85, add_156_21_n_86, add_156_21_n_88, add_156_21_n_89;
  wire add_156_21_n_91, add_156_21_n_92, add_158_21_n_0, add_158_21_n_1, add_158_21_n_2, add_158_21_n_3, add_158_21_n_4, add_158_21_n_5;
  wire add_158_21_n_6, add_158_21_n_7, add_158_21_n_8, add_158_21_n_9, add_158_21_n_10, add_158_21_n_11, add_158_21_n_12, add_158_21_n_13;
  wire add_158_21_n_14, add_158_21_n_15, add_158_21_n_16, add_158_21_n_17, add_158_21_n_18, add_158_21_n_19, add_158_21_n_20, add_158_21_n_21;
  wire add_158_21_n_22, add_158_21_n_23, add_158_21_n_24, add_158_21_n_25, add_158_21_n_26, add_158_21_n_27, add_158_21_n_28, add_158_21_n_29;
  wire add_158_21_n_30, add_158_21_n_31, add_158_21_n_32, add_158_21_n_33, add_158_21_n_34, add_158_21_n_35, add_158_21_n_36, add_158_21_n_37;
  wire add_158_21_n_38, add_158_21_n_39, add_158_21_n_40, add_158_21_n_41, add_158_21_n_42, add_158_21_n_43, add_158_21_n_44, add_158_21_n_45;
  wire add_158_21_n_46, add_158_21_n_47, add_158_21_n_48, add_158_21_n_49, add_158_21_n_51, add_158_21_n_53, add_158_21_n_55, add_158_21_n_56;
  wire add_158_21_n_58, add_158_21_n_59, add_158_21_n_61, add_158_21_n_62, add_158_21_n_64, add_158_21_n_65, add_158_21_n_67, add_158_21_n_68;
  wire add_158_21_n_70, add_158_21_n_71, add_158_21_n_73, add_158_21_n_74, add_158_21_n_76, add_158_21_n_77, add_158_21_n_79, add_158_21_n_80;
  wire add_158_21_n_82, add_158_21_n_83, add_158_21_n_85, add_158_21_n_86, add_158_21_n_88, add_158_21_n_89, add_158_21_n_91, add_158_21_n_92;
  wire add_160_21_n_0, add_160_21_n_1, add_160_21_n_2, add_160_21_n_3, add_160_21_n_4, add_160_21_n_5, add_160_21_n_6, add_160_21_n_7;
  wire add_160_21_n_8, add_160_21_n_9, add_160_21_n_10, add_160_21_n_11, add_160_21_n_12, add_160_21_n_13, add_160_21_n_14, add_160_21_n_15;
  wire add_160_21_n_16, add_160_21_n_17, add_160_21_n_18, add_160_21_n_19, add_160_21_n_20, add_160_21_n_21, add_160_21_n_22, add_160_21_n_23;
  wire add_160_21_n_24, add_160_21_n_25, add_160_21_n_26, add_160_21_n_27, add_160_21_n_28, add_160_21_n_29, add_160_21_n_30, add_160_21_n_31;
  wire add_160_21_n_32, add_160_21_n_33, add_160_21_n_34, add_160_21_n_35, add_160_21_n_36, add_160_21_n_37, add_160_21_n_38, add_160_21_n_39;
  wire add_160_21_n_40, add_160_21_n_41, add_160_21_n_42, add_160_21_n_43, add_160_21_n_44, add_160_21_n_45, add_160_21_n_46, add_160_21_n_47;
  wire add_160_21_n_48, add_160_21_n_49, add_160_21_n_51, add_160_21_n_53, add_160_21_n_55, add_160_21_n_56, add_160_21_n_58, add_160_21_n_59;
  wire add_160_21_n_61, add_160_21_n_62, add_160_21_n_64, add_160_21_n_65, add_160_21_n_67, add_160_21_n_68, add_160_21_n_70, add_160_21_n_71;
  wire add_160_21_n_73, add_160_21_n_74, add_160_21_n_76, add_160_21_n_77, add_160_21_n_79, add_160_21_n_80, add_160_21_n_82, add_160_21_n_83;
  wire add_160_21_n_85, add_160_21_n_86, add_160_21_n_88, add_160_21_n_89, add_160_21_n_91, add_160_21_n_92, add_162_21_n_0, add_162_21_n_1;
  wire add_162_21_n_2, add_162_21_n_3, add_162_21_n_4, add_162_21_n_5, add_162_21_n_6, add_162_21_n_7, add_162_21_n_8, add_162_21_n_9;
  wire add_162_21_n_10, add_162_21_n_11, add_162_21_n_12, add_162_21_n_13, add_162_21_n_14, add_162_21_n_15, add_162_21_n_16, add_162_21_n_17;
  wire add_162_21_n_18, add_162_21_n_19, add_162_21_n_20, add_162_21_n_21, add_162_21_n_22, add_162_21_n_23, add_162_21_n_24, add_162_21_n_25;
  wire add_162_21_n_26, add_162_21_n_27, add_162_21_n_28, add_162_21_n_29, add_162_21_n_30, add_162_21_n_31, add_162_21_n_32, add_162_21_n_33;
  wire add_162_21_n_34, add_162_21_n_35, add_162_21_n_36, add_162_21_n_37, add_162_21_n_38, add_162_21_n_39, add_162_21_n_40, add_162_21_n_41;
  wire add_162_21_n_42, add_162_21_n_43, add_162_21_n_44, add_162_21_n_45, add_162_21_n_46, add_162_21_n_47, add_162_21_n_48, add_162_21_n_49;
  wire add_162_21_n_51, add_162_21_n_53, add_162_21_n_55, add_162_21_n_56, add_162_21_n_58, add_162_21_n_59, add_162_21_n_61, add_162_21_n_62;
  wire add_162_21_n_64, add_162_21_n_65, add_162_21_n_67, add_162_21_n_68, add_162_21_n_70, add_162_21_n_71, add_162_21_n_73, add_162_21_n_74;
  wire add_162_21_n_76, add_162_21_n_77, add_162_21_n_79, add_162_21_n_80, add_162_21_n_82, add_162_21_n_83, add_162_21_n_85, add_162_21_n_86;
  wire add_162_21_n_88, add_162_21_n_89, add_162_21_n_91, add_162_21_n_92, add_164_21_n_0, add_164_21_n_1, add_164_21_n_2, add_164_21_n_3;
  wire add_164_21_n_4, add_164_21_n_5, add_164_21_n_6, add_164_21_n_7, add_164_21_n_8, add_164_21_n_9, add_164_21_n_10, add_164_21_n_11;
  wire add_164_21_n_12, add_164_21_n_13, add_164_21_n_14, add_164_21_n_15, add_164_21_n_16, add_164_21_n_17, add_164_21_n_18, add_164_21_n_19;
  wire add_164_21_n_20, add_164_21_n_21, add_164_21_n_22, add_164_21_n_23, add_164_21_n_24, add_164_21_n_25, add_164_21_n_26, add_164_21_n_27;
  wire add_164_21_n_28, add_164_21_n_29, add_164_21_n_30, add_164_21_n_31, add_164_21_n_32, add_164_21_n_33, add_164_21_n_34, add_164_21_n_35;
  wire add_164_21_n_36, add_164_21_n_37, add_164_21_n_38, add_164_21_n_39, add_164_21_n_40, add_164_21_n_41, add_164_21_n_42, add_164_21_n_43;
  wire add_164_21_n_44, add_164_21_n_45, add_164_21_n_46, add_164_21_n_47, add_164_21_n_48, add_164_21_n_49, add_164_21_n_51, add_164_21_n_53;
  wire add_164_21_n_55, add_164_21_n_56, add_164_21_n_58, add_164_21_n_59, add_164_21_n_61, add_164_21_n_62, add_164_21_n_64, add_164_21_n_65;
  wire add_164_21_n_67, add_164_21_n_68, add_164_21_n_70, add_164_21_n_71, add_164_21_n_73, add_164_21_n_74, add_164_21_n_76, add_164_21_n_77;
  wire add_164_21_n_79, add_164_21_n_80, add_164_21_n_82, add_164_21_n_83, add_164_21_n_85, add_164_21_n_86, add_164_21_n_88, add_164_21_n_89;
  wire add_164_21_n_91, add_164_21_n_92, add_166_21_n_0, add_166_21_n_1, add_166_21_n_2, add_166_21_n_3, add_166_21_n_4, add_166_21_n_5;
  wire add_166_21_n_6, add_166_21_n_7, add_166_21_n_8, add_166_21_n_9, add_166_21_n_10, add_166_21_n_11, add_166_21_n_12, add_166_21_n_13;
  wire add_166_21_n_14, add_166_21_n_15, add_166_21_n_16, add_166_21_n_17, add_166_21_n_18, add_166_21_n_19, add_166_21_n_20, add_166_21_n_21;
  wire add_166_21_n_22, add_166_21_n_23, add_166_21_n_24, add_166_21_n_25, add_166_21_n_26, add_166_21_n_27, add_166_21_n_28, add_166_21_n_29;
  wire add_166_21_n_30, add_166_21_n_31, add_166_21_n_32, add_166_21_n_33, add_166_21_n_34, add_166_21_n_35, add_166_21_n_36, add_166_21_n_37;
  wire add_166_21_n_38, add_166_21_n_39, add_166_21_n_40, add_166_21_n_41, add_166_21_n_42, add_166_21_n_43, add_166_21_n_44, add_166_21_n_45;
  wire add_166_21_n_46, add_166_21_n_47, add_166_21_n_48, add_166_21_n_49, add_166_21_n_51, add_166_21_n_53, add_166_21_n_55, add_166_21_n_56;
  wire add_166_21_n_58, add_166_21_n_59, add_166_21_n_61, add_166_21_n_62, add_166_21_n_64, add_166_21_n_65, add_166_21_n_67, add_166_21_n_68;
  wire add_166_21_n_70, add_166_21_n_71, add_166_21_n_73, add_166_21_n_74, add_166_21_n_76, add_166_21_n_77, add_166_21_n_79, add_166_21_n_80;
  wire add_166_21_n_82, add_166_21_n_83, add_166_21_n_85, add_166_21_n_86, add_166_21_n_88, add_166_21_n_89, add_166_21_n_91, add_166_21_n_92;
  wire add_168_21_n_0, add_168_21_n_1, add_168_21_n_2, add_168_21_n_3, add_168_21_n_4, add_168_21_n_5, add_168_21_n_6, add_168_21_n_7;
  wire add_168_21_n_8, add_168_21_n_9, add_168_21_n_10, add_168_21_n_11, add_168_21_n_12, add_168_21_n_13, add_168_21_n_14, add_168_21_n_15;
  wire add_168_21_n_16, add_168_21_n_17, add_168_21_n_18, add_168_21_n_19, add_168_21_n_20, add_168_21_n_21, add_168_21_n_22, add_168_21_n_23;
  wire add_168_21_n_24, add_168_21_n_25, add_168_21_n_26, add_168_21_n_27, add_168_21_n_28, add_168_21_n_29, add_168_21_n_30, add_168_21_n_31;
  wire add_168_21_n_32, add_168_21_n_33, add_168_21_n_34, add_168_21_n_35, add_168_21_n_36, add_168_21_n_37, add_168_21_n_38, add_168_21_n_39;
  wire add_168_21_n_40, add_168_21_n_41, add_168_21_n_42, add_168_21_n_43, add_168_21_n_44, add_168_21_n_45, add_168_21_n_46, add_168_21_n_47;
  wire add_168_21_n_48, add_168_21_n_49, add_168_21_n_51, add_168_21_n_53, add_168_21_n_55, add_168_21_n_56, add_168_21_n_58, add_168_21_n_59;
  wire add_168_21_n_61, add_168_21_n_62, add_168_21_n_64, add_168_21_n_65, add_168_21_n_67, add_168_21_n_68, add_168_21_n_70, add_168_21_n_71;
  wire add_168_21_n_73, add_168_21_n_74, add_168_21_n_76, add_168_21_n_77, add_168_21_n_79, add_168_21_n_80, add_168_21_n_82, add_168_21_n_83;
  wire add_168_21_n_85, add_168_21_n_86, add_168_21_n_88, add_168_21_n_89, add_168_21_n_91, add_168_21_n_92, add_170_21_n_0, add_170_21_n_1;
  wire add_170_21_n_2, add_170_21_n_3, add_170_21_n_4, add_170_21_n_5, add_170_21_n_6, add_170_21_n_7, add_170_21_n_8, add_170_21_n_9;
  wire add_170_21_n_10, add_170_21_n_11, add_170_21_n_12, add_170_21_n_13, add_170_21_n_14, add_170_21_n_15, add_170_21_n_16, add_170_21_n_17;
  wire add_170_21_n_18, add_170_21_n_19, add_170_21_n_20, add_170_21_n_21, add_170_21_n_22, add_170_21_n_23, add_170_21_n_24, add_170_21_n_25;
  wire add_170_21_n_26, add_170_21_n_27, add_170_21_n_28, add_170_21_n_29, add_170_21_n_30, add_170_21_n_31, add_170_21_n_32, add_170_21_n_33;
  wire add_170_21_n_34, add_170_21_n_35, add_170_21_n_36, add_170_21_n_37, add_170_21_n_38, add_170_21_n_39, add_170_21_n_40, add_170_21_n_41;
  wire add_170_21_n_42, add_170_21_n_43, add_170_21_n_44, add_170_21_n_45, add_170_21_n_46, add_170_21_n_47, add_170_21_n_48, add_170_21_n_49;
  wire add_170_21_n_51, add_170_21_n_53, add_170_21_n_55, add_170_21_n_56, add_170_21_n_58, add_170_21_n_59, add_170_21_n_61, add_170_21_n_62;
  wire add_170_21_n_64, add_170_21_n_65, add_170_21_n_67, add_170_21_n_68, add_170_21_n_70, add_170_21_n_71, add_170_21_n_73, add_170_21_n_74;
  wire add_170_21_n_76, add_170_21_n_77, add_170_21_n_79, add_170_21_n_80, add_170_21_n_82, add_170_21_n_83, add_170_21_n_85, add_170_21_n_86;
  wire add_170_21_n_88, add_170_21_n_89, add_170_21_n_91, add_170_21_n_92, add_172_21_n_0, add_172_21_n_1, add_172_21_n_2, add_172_21_n_3;
  wire add_172_21_n_4, add_172_21_n_5, add_172_21_n_6, add_172_21_n_7, add_172_21_n_8, add_172_21_n_9, add_172_21_n_10, add_172_21_n_11;
  wire add_172_21_n_12, add_172_21_n_13, add_172_21_n_14, add_172_21_n_15, add_172_21_n_16, add_172_21_n_17, add_172_21_n_18, add_172_21_n_19;
  wire add_172_21_n_20, add_172_21_n_21, add_172_21_n_22, add_172_21_n_23, add_172_21_n_24, add_172_21_n_25, add_172_21_n_26, add_172_21_n_27;
  wire add_172_21_n_28, add_172_21_n_29, add_172_21_n_30, add_172_21_n_31, add_172_21_n_32, add_172_21_n_33, add_172_21_n_34, add_172_21_n_35;
  wire add_172_21_n_36, add_172_21_n_37, add_172_21_n_38, add_172_21_n_39, add_172_21_n_40, add_172_21_n_41, add_172_21_n_42, add_172_21_n_43;
  wire add_172_21_n_44, add_172_21_n_45, add_172_21_n_46, add_172_21_n_47, add_172_21_n_48, add_172_21_n_49, add_172_21_n_51, add_172_21_n_53;
  wire add_172_21_n_55, add_172_21_n_56, add_172_21_n_58, add_172_21_n_59, add_172_21_n_61, add_172_21_n_62, add_172_21_n_64, add_172_21_n_65;
  wire add_172_21_n_67, add_172_21_n_68, add_172_21_n_70, add_172_21_n_71, add_172_21_n_73, add_172_21_n_74, add_172_21_n_76, add_172_21_n_77;
  wire add_172_21_n_79, add_172_21_n_80, add_172_21_n_82, add_172_21_n_83, add_172_21_n_85, add_172_21_n_86, add_172_21_n_88, add_172_21_n_89;
  wire add_172_21_n_91, add_172_21_n_92, add_174_21_n_0, add_174_21_n_1, add_174_21_n_2, add_174_21_n_3, add_174_21_n_4, add_174_21_n_5;
  wire add_174_21_n_6, add_174_21_n_7, add_174_21_n_8, add_174_21_n_9, add_174_21_n_10, add_174_21_n_11, add_174_21_n_12, add_174_21_n_13;
  wire add_174_21_n_14, add_174_21_n_15, add_174_21_n_16, add_174_21_n_17, add_174_21_n_18, add_174_21_n_19, add_174_21_n_20, add_174_21_n_21;
  wire add_174_21_n_22, add_174_21_n_23, add_174_21_n_24, add_174_21_n_25, add_174_21_n_26, add_174_21_n_27, add_174_21_n_28, add_174_21_n_29;
  wire add_174_21_n_30, add_174_21_n_31, add_174_21_n_32, add_174_21_n_33, add_174_21_n_34, add_174_21_n_35, add_174_21_n_36, add_174_21_n_37;
  wire add_174_21_n_38, add_174_21_n_39, add_174_21_n_40, add_174_21_n_41, add_174_21_n_42, add_174_21_n_43, add_174_21_n_44, add_174_21_n_45;
  wire add_174_21_n_46, add_174_21_n_47, add_174_21_n_48, add_174_21_n_49, add_174_21_n_51, add_174_21_n_53, add_174_21_n_55, add_174_21_n_56;
  wire add_174_21_n_58, add_174_21_n_59, add_174_21_n_61, add_174_21_n_62, add_174_21_n_64, add_174_21_n_65, add_174_21_n_67, add_174_21_n_68;
  wire add_174_21_n_70, add_174_21_n_71, add_174_21_n_73, add_174_21_n_74, add_174_21_n_76, add_174_21_n_77, add_174_21_n_79, add_174_21_n_80;
  wire add_174_21_n_82, add_174_21_n_83, add_174_21_n_85, add_174_21_n_86, add_174_21_n_88, add_174_21_n_89, add_174_21_n_91, add_174_21_n_92;
  wire add_176_21_n_0, add_176_21_n_1, add_176_21_n_2, add_176_21_n_3, add_176_21_n_4, add_176_21_n_5, add_176_21_n_6, add_176_21_n_7;
  wire add_176_21_n_8, add_176_21_n_9, add_176_21_n_10, add_176_21_n_11, add_176_21_n_12, add_176_21_n_13, add_176_21_n_14, add_176_21_n_15;
  wire add_176_21_n_16, add_176_21_n_17, add_176_21_n_18, add_176_21_n_19, add_176_21_n_20, add_176_21_n_21, add_176_21_n_22, add_176_21_n_23;
  wire add_176_21_n_24, add_176_21_n_25, add_176_21_n_26, add_176_21_n_27, add_176_21_n_28, add_176_21_n_29, add_176_21_n_30, add_176_21_n_31;
  wire add_176_21_n_32, add_176_21_n_33, add_176_21_n_34, add_176_21_n_35, add_176_21_n_36, add_176_21_n_37, add_176_21_n_38, add_176_21_n_39;
  wire add_176_21_n_40, add_176_21_n_41, add_176_21_n_42, add_176_21_n_43, add_176_21_n_44, add_176_21_n_45, add_176_21_n_46, add_176_21_n_47;
  wire add_176_21_n_48, add_176_21_n_49, add_176_21_n_51, add_176_21_n_53, add_176_21_n_55, add_176_21_n_56, add_176_21_n_58, add_176_21_n_59;
  wire add_176_21_n_61, add_176_21_n_62, add_176_21_n_64, add_176_21_n_65, add_176_21_n_67, add_176_21_n_68, add_176_21_n_70, add_176_21_n_71;
  wire add_176_21_n_73, add_176_21_n_74, add_176_21_n_76, add_176_21_n_77, add_176_21_n_79, add_176_21_n_80, add_176_21_n_82, add_176_21_n_83;
  wire add_176_21_n_85, add_176_21_n_86, add_176_21_n_88, add_176_21_n_89, add_176_21_n_91, add_176_21_n_92, add_178_21_n_0, add_178_21_n_1;
  wire add_178_21_n_2, add_178_21_n_3, add_178_21_n_4, add_178_21_n_5, add_178_21_n_6, add_178_21_n_7, add_178_21_n_8, add_178_21_n_9;
  wire add_178_21_n_10, add_178_21_n_11, add_178_21_n_12, add_178_21_n_13, add_178_21_n_14, add_178_21_n_15, add_178_21_n_16, add_178_21_n_17;
  wire add_178_21_n_18, add_178_21_n_19, add_178_21_n_20, add_178_21_n_21, add_178_21_n_22, add_178_21_n_23, add_178_21_n_24, add_178_21_n_25;
  wire add_178_21_n_26, add_178_21_n_27, add_178_21_n_28, add_178_21_n_29, add_178_21_n_30, add_178_21_n_31, add_178_21_n_32, add_178_21_n_33;
  wire add_178_21_n_34, add_178_21_n_35, add_178_21_n_36, add_178_21_n_37, add_178_21_n_38, add_178_21_n_39, add_178_21_n_40, add_178_21_n_41;
  wire add_178_21_n_42, add_178_21_n_43, add_178_21_n_44, add_178_21_n_45, add_178_21_n_46, add_178_21_n_47, add_178_21_n_48, add_178_21_n_49;
  wire add_178_21_n_51, add_178_21_n_53, add_178_21_n_55, add_178_21_n_56, add_178_21_n_58, add_178_21_n_59, add_178_21_n_61, add_178_21_n_62;
  wire add_178_21_n_64, add_178_21_n_65, add_178_21_n_67, add_178_21_n_68, add_178_21_n_70, add_178_21_n_71, add_178_21_n_73, add_178_21_n_74;
  wire add_178_21_n_76, add_178_21_n_77, add_178_21_n_79, add_178_21_n_80, add_178_21_n_82, add_178_21_n_83, add_178_21_n_85, add_178_21_n_86;
  wire add_178_21_n_88, add_178_21_n_89, add_178_21_n_91, add_178_21_n_92, add_180_21_n_0, add_180_21_n_1, add_180_21_n_2, add_180_21_n_3;
  wire add_180_21_n_4, add_180_21_n_5, add_180_21_n_6, add_180_21_n_7, add_180_21_n_8, add_180_21_n_9, add_180_21_n_10, add_180_21_n_11;
  wire add_180_21_n_12, add_180_21_n_13, add_180_21_n_14, add_180_21_n_15, add_180_21_n_16, add_180_21_n_17, add_180_21_n_18, add_180_21_n_19;
  wire add_180_21_n_20, add_180_21_n_21, add_180_21_n_22, add_180_21_n_23, add_180_21_n_24, add_180_21_n_25, add_180_21_n_26, add_180_21_n_27;
  wire add_180_21_n_28, add_180_21_n_29, add_180_21_n_30, add_180_21_n_31, add_180_21_n_32, add_180_21_n_33, add_180_21_n_34, add_180_21_n_35;
  wire add_180_21_n_36, add_180_21_n_37, add_180_21_n_38, add_180_21_n_39, add_180_21_n_40, add_180_21_n_41, add_180_21_n_42, add_180_21_n_43;
  wire add_180_21_n_44, add_180_21_n_45, add_180_21_n_46, add_180_21_n_47, add_180_21_n_48, add_180_21_n_49, add_180_21_n_51, add_180_21_n_53;
  wire add_180_21_n_55, add_180_21_n_56, add_180_21_n_58, add_180_21_n_59, add_180_21_n_61, add_180_21_n_62, add_180_21_n_64, add_180_21_n_65;
  wire add_180_21_n_67, add_180_21_n_68, add_180_21_n_70, add_180_21_n_71, add_180_21_n_73, add_180_21_n_74, add_180_21_n_76, add_180_21_n_77;
  wire add_180_21_n_79, add_180_21_n_80, add_180_21_n_82, add_180_21_n_83, add_180_21_n_85, add_180_21_n_86, add_180_21_n_88, add_180_21_n_89;
  wire add_180_21_n_91, add_180_21_n_92, csa_tree_add_190_195_groupi_n_0, csa_tree_add_190_195_groupi_n_1, csa_tree_add_190_195_groupi_n_2, csa_tree_add_190_195_groupi_n_3, csa_tree_add_190_195_groupi_n_4, csa_tree_add_190_195_groupi_n_5;
  wire csa_tree_add_190_195_groupi_n_6, csa_tree_add_190_195_groupi_n_7, csa_tree_add_190_195_groupi_n_8, csa_tree_add_190_195_groupi_n_9, csa_tree_add_190_195_groupi_n_10, csa_tree_add_190_195_groupi_n_11, csa_tree_add_190_195_groupi_n_12, csa_tree_add_190_195_groupi_n_13;
  wire csa_tree_add_190_195_groupi_n_14, csa_tree_add_190_195_groupi_n_15, csa_tree_add_190_195_groupi_n_16, csa_tree_add_190_195_groupi_n_17, csa_tree_add_190_195_groupi_n_18, csa_tree_add_190_195_groupi_n_19, csa_tree_add_190_195_groupi_n_20, csa_tree_add_190_195_groupi_n_21;
  wire csa_tree_add_190_195_groupi_n_22, csa_tree_add_190_195_groupi_n_23, csa_tree_add_190_195_groupi_n_24, csa_tree_add_190_195_groupi_n_25, csa_tree_add_190_195_groupi_n_26, csa_tree_add_190_195_groupi_n_27, csa_tree_add_190_195_groupi_n_28, csa_tree_add_190_195_groupi_n_29;
  wire csa_tree_add_190_195_groupi_n_30, csa_tree_add_190_195_groupi_n_31, csa_tree_add_190_195_groupi_n_32, csa_tree_add_190_195_groupi_n_33, csa_tree_add_190_195_groupi_n_34, csa_tree_add_190_195_groupi_n_35, csa_tree_add_190_195_groupi_n_36, csa_tree_add_190_195_groupi_n_37;
  wire csa_tree_add_190_195_groupi_n_38, csa_tree_add_190_195_groupi_n_39, csa_tree_add_190_195_groupi_n_40, csa_tree_add_190_195_groupi_n_41, csa_tree_add_190_195_groupi_n_42, csa_tree_add_190_195_groupi_n_43, csa_tree_add_190_195_groupi_n_44, csa_tree_add_190_195_groupi_n_45;
  wire csa_tree_add_190_195_groupi_n_46, csa_tree_add_190_195_groupi_n_47, csa_tree_add_190_195_groupi_n_48, csa_tree_add_190_195_groupi_n_49, csa_tree_add_190_195_groupi_n_50, csa_tree_add_190_195_groupi_n_51, csa_tree_add_190_195_groupi_n_52, csa_tree_add_190_195_groupi_n_53;
  wire csa_tree_add_190_195_groupi_n_54, csa_tree_add_190_195_groupi_n_55, csa_tree_add_190_195_groupi_n_56, csa_tree_add_190_195_groupi_n_57, csa_tree_add_190_195_groupi_n_58, csa_tree_add_190_195_groupi_n_59, csa_tree_add_190_195_groupi_n_60, csa_tree_add_190_195_groupi_n_61;
  wire csa_tree_add_190_195_groupi_n_62, csa_tree_add_190_195_groupi_n_63, csa_tree_add_190_195_groupi_n_64, csa_tree_add_190_195_groupi_n_65, csa_tree_add_190_195_groupi_n_66, csa_tree_add_190_195_groupi_n_67, csa_tree_add_190_195_groupi_n_68, csa_tree_add_190_195_groupi_n_69;
  wire csa_tree_add_190_195_groupi_n_70, csa_tree_add_190_195_groupi_n_71, csa_tree_add_190_195_groupi_n_72, csa_tree_add_190_195_groupi_n_73, csa_tree_add_190_195_groupi_n_74, csa_tree_add_190_195_groupi_n_75, csa_tree_add_190_195_groupi_n_76, csa_tree_add_190_195_groupi_n_77;
  wire csa_tree_add_190_195_groupi_n_78, csa_tree_add_190_195_groupi_n_79, csa_tree_add_190_195_groupi_n_80, csa_tree_add_190_195_groupi_n_81, csa_tree_add_190_195_groupi_n_82, csa_tree_add_190_195_groupi_n_83, csa_tree_add_190_195_groupi_n_84, csa_tree_add_190_195_groupi_n_85;
  wire csa_tree_add_190_195_groupi_n_86, csa_tree_add_190_195_groupi_n_87, csa_tree_add_190_195_groupi_n_88, csa_tree_add_190_195_groupi_n_89, csa_tree_add_190_195_groupi_n_90, csa_tree_add_190_195_groupi_n_91, csa_tree_add_190_195_groupi_n_92, csa_tree_add_190_195_groupi_n_93;
  wire csa_tree_add_190_195_groupi_n_94, csa_tree_add_190_195_groupi_n_95, csa_tree_add_190_195_groupi_n_96, csa_tree_add_190_195_groupi_n_97, csa_tree_add_190_195_groupi_n_98, csa_tree_add_190_195_groupi_n_99, csa_tree_add_190_195_groupi_n_100, csa_tree_add_190_195_groupi_n_101;
  wire csa_tree_add_190_195_groupi_n_102, csa_tree_add_190_195_groupi_n_103, csa_tree_add_190_195_groupi_n_104, csa_tree_add_190_195_groupi_n_105, csa_tree_add_190_195_groupi_n_106, csa_tree_add_190_195_groupi_n_107, csa_tree_add_190_195_groupi_n_108, csa_tree_add_190_195_groupi_n_109;
  wire csa_tree_add_190_195_groupi_n_110, csa_tree_add_190_195_groupi_n_111, csa_tree_add_190_195_groupi_n_112, csa_tree_add_190_195_groupi_n_113, csa_tree_add_190_195_groupi_n_114, csa_tree_add_190_195_groupi_n_115, csa_tree_add_190_195_groupi_n_116, csa_tree_add_190_195_groupi_n_117;
  wire csa_tree_add_190_195_groupi_n_118, csa_tree_add_190_195_groupi_n_119, csa_tree_add_190_195_groupi_n_120, csa_tree_add_190_195_groupi_n_121, csa_tree_add_190_195_groupi_n_122, csa_tree_add_190_195_groupi_n_123, csa_tree_add_190_195_groupi_n_124, csa_tree_add_190_195_groupi_n_125;
  wire csa_tree_add_190_195_groupi_n_126, csa_tree_add_190_195_groupi_n_127, csa_tree_add_190_195_groupi_n_128, csa_tree_add_190_195_groupi_n_129, csa_tree_add_190_195_groupi_n_130, csa_tree_add_190_195_groupi_n_131, csa_tree_add_190_195_groupi_n_132, csa_tree_add_190_195_groupi_n_133;
  wire csa_tree_add_190_195_groupi_n_134, csa_tree_add_190_195_groupi_n_135, csa_tree_add_190_195_groupi_n_136, csa_tree_add_190_195_groupi_n_137, csa_tree_add_190_195_groupi_n_138, csa_tree_add_190_195_groupi_n_139, csa_tree_add_190_195_groupi_n_140, csa_tree_add_190_195_groupi_n_141;
  wire csa_tree_add_190_195_groupi_n_142, csa_tree_add_190_195_groupi_n_143, csa_tree_add_190_195_groupi_n_144, csa_tree_add_190_195_groupi_n_145, csa_tree_add_190_195_groupi_n_146, csa_tree_add_190_195_groupi_n_147, csa_tree_add_190_195_groupi_n_148, csa_tree_add_190_195_groupi_n_149;
  wire csa_tree_add_190_195_groupi_n_150, csa_tree_add_190_195_groupi_n_151, csa_tree_add_190_195_groupi_n_152, csa_tree_add_190_195_groupi_n_153, csa_tree_add_190_195_groupi_n_154, csa_tree_add_190_195_groupi_n_155, csa_tree_add_190_195_groupi_n_156, csa_tree_add_190_195_groupi_n_157;
  wire csa_tree_add_190_195_groupi_n_158, csa_tree_add_190_195_groupi_n_159, csa_tree_add_190_195_groupi_n_160, csa_tree_add_190_195_groupi_n_161, csa_tree_add_190_195_groupi_n_162, csa_tree_add_190_195_groupi_n_163, csa_tree_add_190_195_groupi_n_164, csa_tree_add_190_195_groupi_n_165;
  wire csa_tree_add_190_195_groupi_n_166, csa_tree_add_190_195_groupi_n_167, csa_tree_add_190_195_groupi_n_168, csa_tree_add_190_195_groupi_n_169, csa_tree_add_190_195_groupi_n_170, csa_tree_add_190_195_groupi_n_171, csa_tree_add_190_195_groupi_n_172, csa_tree_add_190_195_groupi_n_173;
  wire csa_tree_add_190_195_groupi_n_174, csa_tree_add_190_195_groupi_n_175, csa_tree_add_190_195_groupi_n_176, csa_tree_add_190_195_groupi_n_177, csa_tree_add_190_195_groupi_n_180, csa_tree_add_190_195_groupi_n_182, csa_tree_add_190_195_groupi_n_183, csa_tree_add_190_195_groupi_n_184;
  wire csa_tree_add_190_195_groupi_n_185, csa_tree_add_190_195_groupi_n_186, csa_tree_add_190_195_groupi_n_187, csa_tree_add_190_195_groupi_n_188, csa_tree_add_190_195_groupi_n_189, csa_tree_add_190_195_groupi_n_190, csa_tree_add_190_195_groupi_n_191, csa_tree_add_190_195_groupi_n_192;
  wire csa_tree_add_190_195_groupi_n_193, csa_tree_add_190_195_groupi_n_194, csa_tree_add_190_195_groupi_n_195, csa_tree_add_190_195_groupi_n_196, csa_tree_add_190_195_groupi_n_197, csa_tree_add_190_195_groupi_n_198, csa_tree_add_190_195_groupi_n_199, csa_tree_add_190_195_groupi_n_200;
  wire csa_tree_add_190_195_groupi_n_201, csa_tree_add_190_195_groupi_n_202, csa_tree_add_190_195_groupi_n_203, csa_tree_add_190_195_groupi_n_204, csa_tree_add_190_195_groupi_n_205, csa_tree_add_190_195_groupi_n_206, csa_tree_add_190_195_groupi_n_207, csa_tree_add_190_195_groupi_n_208;
  wire csa_tree_add_190_195_groupi_n_209, csa_tree_add_190_195_groupi_n_210, csa_tree_add_190_195_groupi_n_211, csa_tree_add_190_195_groupi_n_212, csa_tree_add_190_195_groupi_n_213, csa_tree_add_190_195_groupi_n_214, csa_tree_add_190_195_groupi_n_215, csa_tree_add_190_195_groupi_n_216;
  wire csa_tree_add_190_195_groupi_n_217, csa_tree_add_190_195_groupi_n_218, csa_tree_add_190_195_groupi_n_219, csa_tree_add_190_195_groupi_n_220, csa_tree_add_190_195_groupi_n_221, csa_tree_add_190_195_groupi_n_222, csa_tree_add_190_195_groupi_n_223, csa_tree_add_190_195_groupi_n_224;
  wire csa_tree_add_190_195_groupi_n_225, csa_tree_add_190_195_groupi_n_226, csa_tree_add_190_195_groupi_n_227, csa_tree_add_190_195_groupi_n_228, csa_tree_add_190_195_groupi_n_229, csa_tree_add_190_195_groupi_n_230, csa_tree_add_190_195_groupi_n_231, csa_tree_add_190_195_groupi_n_232;
  wire csa_tree_add_190_195_groupi_n_233, csa_tree_add_190_195_groupi_n_234, csa_tree_add_190_195_groupi_n_235, csa_tree_add_190_195_groupi_n_236, csa_tree_add_190_195_groupi_n_237, csa_tree_add_190_195_groupi_n_238, csa_tree_add_190_195_groupi_n_239, csa_tree_add_190_195_groupi_n_240;
  wire csa_tree_add_190_195_groupi_n_241, csa_tree_add_190_195_groupi_n_242, csa_tree_add_190_195_groupi_n_243, csa_tree_add_190_195_groupi_n_244, csa_tree_add_190_195_groupi_n_245, csa_tree_add_190_195_groupi_n_246, csa_tree_add_190_195_groupi_n_247, csa_tree_add_190_195_groupi_n_248;
  wire csa_tree_add_190_195_groupi_n_249, csa_tree_add_190_195_groupi_n_250, csa_tree_add_190_195_groupi_n_251, csa_tree_add_190_195_groupi_n_252, csa_tree_add_190_195_groupi_n_253, csa_tree_add_190_195_groupi_n_254, csa_tree_add_190_195_groupi_n_255, csa_tree_add_190_195_groupi_n_256;
  wire csa_tree_add_190_195_groupi_n_257, csa_tree_add_190_195_groupi_n_258, csa_tree_add_190_195_groupi_n_259, csa_tree_add_190_195_groupi_n_260, csa_tree_add_190_195_groupi_n_261, csa_tree_add_190_195_groupi_n_262, csa_tree_add_190_195_groupi_n_263, csa_tree_add_190_195_groupi_n_264;
  wire csa_tree_add_190_195_groupi_n_265, csa_tree_add_190_195_groupi_n_266, csa_tree_add_190_195_groupi_n_267, csa_tree_add_190_195_groupi_n_268, csa_tree_add_190_195_groupi_n_269, csa_tree_add_190_195_groupi_n_270, csa_tree_add_190_195_groupi_n_271, csa_tree_add_190_195_groupi_n_272;
  wire csa_tree_add_190_195_groupi_n_273, csa_tree_add_190_195_groupi_n_274, csa_tree_add_190_195_groupi_n_275, csa_tree_add_190_195_groupi_n_276, csa_tree_add_190_195_groupi_n_277, csa_tree_add_190_195_groupi_n_278, csa_tree_add_190_195_groupi_n_279, csa_tree_add_190_195_groupi_n_280;
  wire csa_tree_add_190_195_groupi_n_281, csa_tree_add_190_195_groupi_n_282, csa_tree_add_190_195_groupi_n_283, csa_tree_add_190_195_groupi_n_284, csa_tree_add_190_195_groupi_n_285, csa_tree_add_190_195_groupi_n_286, csa_tree_add_190_195_groupi_n_287, csa_tree_add_190_195_groupi_n_288;
  wire csa_tree_add_190_195_groupi_n_289, csa_tree_add_190_195_groupi_n_290, csa_tree_add_190_195_groupi_n_291, csa_tree_add_190_195_groupi_n_292, csa_tree_add_190_195_groupi_n_293, csa_tree_add_190_195_groupi_n_294, csa_tree_add_190_195_groupi_n_295, csa_tree_add_190_195_groupi_n_296;
  wire csa_tree_add_190_195_groupi_n_297, csa_tree_add_190_195_groupi_n_298, csa_tree_add_190_195_groupi_n_299, csa_tree_add_190_195_groupi_n_300, csa_tree_add_190_195_groupi_n_301, csa_tree_add_190_195_groupi_n_302, csa_tree_add_190_195_groupi_n_303, csa_tree_add_190_195_groupi_n_304;
  wire csa_tree_add_190_195_groupi_n_305, csa_tree_add_190_195_groupi_n_306, csa_tree_add_190_195_groupi_n_307, csa_tree_add_190_195_groupi_n_308, csa_tree_add_190_195_groupi_n_309, csa_tree_add_190_195_groupi_n_310, csa_tree_add_190_195_groupi_n_311, csa_tree_add_190_195_groupi_n_312;
  wire csa_tree_add_190_195_groupi_n_313, csa_tree_add_190_195_groupi_n_314, csa_tree_add_190_195_groupi_n_315, csa_tree_add_190_195_groupi_n_316, csa_tree_add_190_195_groupi_n_317, csa_tree_add_190_195_groupi_n_318, csa_tree_add_190_195_groupi_n_319, csa_tree_add_190_195_groupi_n_320;
  wire csa_tree_add_190_195_groupi_n_321, csa_tree_add_190_195_groupi_n_322, csa_tree_add_190_195_groupi_n_323, csa_tree_add_190_195_groupi_n_324, csa_tree_add_190_195_groupi_n_325, csa_tree_add_190_195_groupi_n_326, csa_tree_add_190_195_groupi_n_327, csa_tree_add_190_195_groupi_n_328;
  wire csa_tree_add_190_195_groupi_n_329, csa_tree_add_190_195_groupi_n_330, csa_tree_add_190_195_groupi_n_331, csa_tree_add_190_195_groupi_n_332, csa_tree_add_190_195_groupi_n_333, csa_tree_add_190_195_groupi_n_334, csa_tree_add_190_195_groupi_n_335, csa_tree_add_190_195_groupi_n_336;
  wire csa_tree_add_190_195_groupi_n_337, csa_tree_add_190_195_groupi_n_338, csa_tree_add_190_195_groupi_n_339, csa_tree_add_190_195_groupi_n_340, csa_tree_add_190_195_groupi_n_341, csa_tree_add_190_195_groupi_n_342, csa_tree_add_190_195_groupi_n_343, csa_tree_add_190_195_groupi_n_344;
  wire csa_tree_add_190_195_groupi_n_345, csa_tree_add_190_195_groupi_n_346, csa_tree_add_190_195_groupi_n_347, csa_tree_add_190_195_groupi_n_348, csa_tree_add_190_195_groupi_n_349, csa_tree_add_190_195_groupi_n_350, csa_tree_add_190_195_groupi_n_351, csa_tree_add_190_195_groupi_n_352;
  wire csa_tree_add_190_195_groupi_n_353, csa_tree_add_190_195_groupi_n_354, csa_tree_add_190_195_groupi_n_355, csa_tree_add_190_195_groupi_n_356, csa_tree_add_190_195_groupi_n_357, csa_tree_add_190_195_groupi_n_358, csa_tree_add_190_195_groupi_n_359, csa_tree_add_190_195_groupi_n_360;
  wire csa_tree_add_190_195_groupi_n_361, csa_tree_add_190_195_groupi_n_362, csa_tree_add_190_195_groupi_n_363, csa_tree_add_190_195_groupi_n_364, csa_tree_add_190_195_groupi_n_365, csa_tree_add_190_195_groupi_n_366, csa_tree_add_190_195_groupi_n_367, csa_tree_add_190_195_groupi_n_368;
  wire csa_tree_add_190_195_groupi_n_369, csa_tree_add_190_195_groupi_n_370, csa_tree_add_190_195_groupi_n_371, csa_tree_add_190_195_groupi_n_372, csa_tree_add_190_195_groupi_n_373, csa_tree_add_190_195_groupi_n_374, csa_tree_add_190_195_groupi_n_375, csa_tree_add_190_195_groupi_n_376;
  wire csa_tree_add_190_195_groupi_n_377, csa_tree_add_190_195_groupi_n_378, csa_tree_add_190_195_groupi_n_379, csa_tree_add_190_195_groupi_n_380, csa_tree_add_190_195_groupi_n_381, csa_tree_add_190_195_groupi_n_382, csa_tree_add_190_195_groupi_n_383, csa_tree_add_190_195_groupi_n_384;
  wire csa_tree_add_190_195_groupi_n_385, csa_tree_add_190_195_groupi_n_386, csa_tree_add_190_195_groupi_n_387, csa_tree_add_190_195_groupi_n_388, csa_tree_add_190_195_groupi_n_389, csa_tree_add_190_195_groupi_n_390, csa_tree_add_190_195_groupi_n_391, csa_tree_add_190_195_groupi_n_392;
  wire csa_tree_add_190_195_groupi_n_393, csa_tree_add_190_195_groupi_n_394, csa_tree_add_190_195_groupi_n_395, csa_tree_add_190_195_groupi_n_396, csa_tree_add_190_195_groupi_n_397, csa_tree_add_190_195_groupi_n_398, csa_tree_add_190_195_groupi_n_399, csa_tree_add_190_195_groupi_n_400;
  wire csa_tree_add_190_195_groupi_n_401, csa_tree_add_190_195_groupi_n_402, csa_tree_add_190_195_groupi_n_403, csa_tree_add_190_195_groupi_n_404, csa_tree_add_190_195_groupi_n_405, csa_tree_add_190_195_groupi_n_406, csa_tree_add_190_195_groupi_n_407, csa_tree_add_190_195_groupi_n_408;
  wire csa_tree_add_190_195_groupi_n_409, csa_tree_add_190_195_groupi_n_410, csa_tree_add_190_195_groupi_n_411, csa_tree_add_190_195_groupi_n_412, csa_tree_add_190_195_groupi_n_413, csa_tree_add_190_195_groupi_n_414, csa_tree_add_190_195_groupi_n_415, csa_tree_add_190_195_groupi_n_416;
  wire csa_tree_add_190_195_groupi_n_417, csa_tree_add_190_195_groupi_n_418, csa_tree_add_190_195_groupi_n_419, csa_tree_add_190_195_groupi_n_420, csa_tree_add_190_195_groupi_n_421, csa_tree_add_190_195_groupi_n_422, csa_tree_add_190_195_groupi_n_423, csa_tree_add_190_195_groupi_n_424;
  wire csa_tree_add_190_195_groupi_n_425, csa_tree_add_190_195_groupi_n_426, csa_tree_add_190_195_groupi_n_427, csa_tree_add_190_195_groupi_n_428, csa_tree_add_190_195_groupi_n_429, csa_tree_add_190_195_groupi_n_430, csa_tree_add_190_195_groupi_n_431, csa_tree_add_190_195_groupi_n_432;
  wire csa_tree_add_190_195_groupi_n_433, csa_tree_add_190_195_groupi_n_434, csa_tree_add_190_195_groupi_n_435, csa_tree_add_190_195_groupi_n_436, csa_tree_add_190_195_groupi_n_437, csa_tree_add_190_195_groupi_n_438, csa_tree_add_190_195_groupi_n_439, csa_tree_add_190_195_groupi_n_440;
  wire csa_tree_add_190_195_groupi_n_441, csa_tree_add_190_195_groupi_n_442, csa_tree_add_190_195_groupi_n_443, csa_tree_add_190_195_groupi_n_444, csa_tree_add_190_195_groupi_n_445, csa_tree_add_190_195_groupi_n_446, csa_tree_add_190_195_groupi_n_447, csa_tree_add_190_195_groupi_n_448;
  wire csa_tree_add_190_195_groupi_n_449, csa_tree_add_190_195_groupi_n_450, csa_tree_add_190_195_groupi_n_451, csa_tree_add_190_195_groupi_n_452, csa_tree_add_190_195_groupi_n_453, csa_tree_add_190_195_groupi_n_454, csa_tree_add_190_195_groupi_n_455, csa_tree_add_190_195_groupi_n_456;
  wire csa_tree_add_190_195_groupi_n_457, csa_tree_add_190_195_groupi_n_458, csa_tree_add_190_195_groupi_n_459, csa_tree_add_190_195_groupi_n_460, csa_tree_add_190_195_groupi_n_461, csa_tree_add_190_195_groupi_n_462, csa_tree_add_190_195_groupi_n_463, csa_tree_add_190_195_groupi_n_464;
  wire csa_tree_add_190_195_groupi_n_465, csa_tree_add_190_195_groupi_n_466, csa_tree_add_190_195_groupi_n_467, csa_tree_add_190_195_groupi_n_468, csa_tree_add_190_195_groupi_n_469, csa_tree_add_190_195_groupi_n_470, csa_tree_add_190_195_groupi_n_471, csa_tree_add_190_195_groupi_n_472;
  wire csa_tree_add_190_195_groupi_n_473, csa_tree_add_190_195_groupi_n_474, csa_tree_add_190_195_groupi_n_475, csa_tree_add_190_195_groupi_n_476, csa_tree_add_190_195_groupi_n_477, csa_tree_add_190_195_groupi_n_478, csa_tree_add_190_195_groupi_n_479, csa_tree_add_190_195_groupi_n_480;
  wire csa_tree_add_190_195_groupi_n_481, csa_tree_add_190_195_groupi_n_482, csa_tree_add_190_195_groupi_n_483, csa_tree_add_190_195_groupi_n_484, csa_tree_add_190_195_groupi_n_485, csa_tree_add_190_195_groupi_n_486, csa_tree_add_190_195_groupi_n_487, csa_tree_add_190_195_groupi_n_488;
  wire csa_tree_add_190_195_groupi_n_489, csa_tree_add_190_195_groupi_n_490, csa_tree_add_190_195_groupi_n_491, csa_tree_add_190_195_groupi_n_492, csa_tree_add_190_195_groupi_n_493, csa_tree_add_190_195_groupi_n_494, csa_tree_add_190_195_groupi_n_495, csa_tree_add_190_195_groupi_n_496;
  wire csa_tree_add_190_195_groupi_n_497, csa_tree_add_190_195_groupi_n_498, csa_tree_add_190_195_groupi_n_499, csa_tree_add_190_195_groupi_n_500, csa_tree_add_190_195_groupi_n_501, csa_tree_add_190_195_groupi_n_502, csa_tree_add_190_195_groupi_n_503, csa_tree_add_190_195_groupi_n_504;
  wire csa_tree_add_190_195_groupi_n_505, csa_tree_add_190_195_groupi_n_506, csa_tree_add_190_195_groupi_n_507, csa_tree_add_190_195_groupi_n_508, csa_tree_add_190_195_groupi_n_509, csa_tree_add_190_195_groupi_n_510, csa_tree_add_190_195_groupi_n_511, csa_tree_add_190_195_groupi_n_512;
  wire csa_tree_add_190_195_groupi_n_513, csa_tree_add_190_195_groupi_n_514, csa_tree_add_190_195_groupi_n_515, csa_tree_add_190_195_groupi_n_516, csa_tree_add_190_195_groupi_n_517, csa_tree_add_190_195_groupi_n_518, csa_tree_add_190_195_groupi_n_519, csa_tree_add_190_195_groupi_n_520;
  wire csa_tree_add_190_195_groupi_n_521, csa_tree_add_190_195_groupi_n_522, csa_tree_add_190_195_groupi_n_523, csa_tree_add_190_195_groupi_n_524, csa_tree_add_190_195_groupi_n_525, csa_tree_add_190_195_groupi_n_526, csa_tree_add_190_195_groupi_n_527, csa_tree_add_190_195_groupi_n_528;
  wire csa_tree_add_190_195_groupi_n_529, csa_tree_add_190_195_groupi_n_530, csa_tree_add_190_195_groupi_n_531, csa_tree_add_190_195_groupi_n_532, csa_tree_add_190_195_groupi_n_533, csa_tree_add_190_195_groupi_n_534, csa_tree_add_190_195_groupi_n_535, csa_tree_add_190_195_groupi_n_536;
  wire csa_tree_add_190_195_groupi_n_537, csa_tree_add_190_195_groupi_n_538, csa_tree_add_190_195_groupi_n_539, csa_tree_add_190_195_groupi_n_540, csa_tree_add_190_195_groupi_n_541, csa_tree_add_190_195_groupi_n_542, csa_tree_add_190_195_groupi_n_543, csa_tree_add_190_195_groupi_n_544;
  wire csa_tree_add_190_195_groupi_n_545, csa_tree_add_190_195_groupi_n_546, csa_tree_add_190_195_groupi_n_547, csa_tree_add_190_195_groupi_n_548, csa_tree_add_190_195_groupi_n_549, csa_tree_add_190_195_groupi_n_550, csa_tree_add_190_195_groupi_n_551, csa_tree_add_190_195_groupi_n_552;
  wire csa_tree_add_190_195_groupi_n_553, csa_tree_add_190_195_groupi_n_554, csa_tree_add_190_195_groupi_n_555, csa_tree_add_190_195_groupi_n_556, csa_tree_add_190_195_groupi_n_557, csa_tree_add_190_195_groupi_n_558, csa_tree_add_190_195_groupi_n_559, csa_tree_add_190_195_groupi_n_560;
  wire csa_tree_add_190_195_groupi_n_561, csa_tree_add_190_195_groupi_n_562, csa_tree_add_190_195_groupi_n_563, csa_tree_add_190_195_groupi_n_564, csa_tree_add_190_195_groupi_n_565, csa_tree_add_190_195_groupi_n_566, csa_tree_add_190_195_groupi_n_567, csa_tree_add_190_195_groupi_n_568;
  wire csa_tree_add_190_195_groupi_n_569, csa_tree_add_190_195_groupi_n_570, csa_tree_add_190_195_groupi_n_571, csa_tree_add_190_195_groupi_n_572, csa_tree_add_190_195_groupi_n_573, csa_tree_add_190_195_groupi_n_574, csa_tree_add_190_195_groupi_n_575, csa_tree_add_190_195_groupi_n_576;
  wire csa_tree_add_190_195_groupi_n_577, csa_tree_add_190_195_groupi_n_578, csa_tree_add_190_195_groupi_n_579, csa_tree_add_190_195_groupi_n_580, csa_tree_add_190_195_groupi_n_581, csa_tree_add_190_195_groupi_n_582, csa_tree_add_190_195_groupi_n_583, csa_tree_add_190_195_groupi_n_584;
  wire csa_tree_add_190_195_groupi_n_585, csa_tree_add_190_195_groupi_n_586, csa_tree_add_190_195_groupi_n_587, csa_tree_add_190_195_groupi_n_588, csa_tree_add_190_195_groupi_n_589, csa_tree_add_190_195_groupi_n_590, csa_tree_add_190_195_groupi_n_591, csa_tree_add_190_195_groupi_n_592;
  wire csa_tree_add_190_195_groupi_n_593, csa_tree_add_190_195_groupi_n_594, csa_tree_add_190_195_groupi_n_595, csa_tree_add_190_195_groupi_n_596, csa_tree_add_190_195_groupi_n_597, csa_tree_add_190_195_groupi_n_598, csa_tree_add_190_195_groupi_n_599, csa_tree_add_190_195_groupi_n_600;
  wire csa_tree_add_190_195_groupi_n_601, csa_tree_add_190_195_groupi_n_602, csa_tree_add_190_195_groupi_n_603, csa_tree_add_190_195_groupi_n_604, csa_tree_add_190_195_groupi_n_605, csa_tree_add_190_195_groupi_n_606, csa_tree_add_190_195_groupi_n_607, csa_tree_add_190_195_groupi_n_608;
  wire csa_tree_add_190_195_groupi_n_609, csa_tree_add_190_195_groupi_n_610, csa_tree_add_190_195_groupi_n_611, csa_tree_add_190_195_groupi_n_612, csa_tree_add_190_195_groupi_n_613, csa_tree_add_190_195_groupi_n_614, csa_tree_add_190_195_groupi_n_615, csa_tree_add_190_195_groupi_n_616;
  wire csa_tree_add_190_195_groupi_n_617, csa_tree_add_190_195_groupi_n_618, csa_tree_add_190_195_groupi_n_619, csa_tree_add_190_195_groupi_n_620, csa_tree_add_190_195_groupi_n_621, csa_tree_add_190_195_groupi_n_622, csa_tree_add_190_195_groupi_n_623, csa_tree_add_190_195_groupi_n_624;
  wire csa_tree_add_190_195_groupi_n_625, csa_tree_add_190_195_groupi_n_626, csa_tree_add_190_195_groupi_n_627, csa_tree_add_190_195_groupi_n_628, csa_tree_add_190_195_groupi_n_629, csa_tree_add_190_195_groupi_n_630, csa_tree_add_190_195_groupi_n_631, csa_tree_add_190_195_groupi_n_632;
  wire csa_tree_add_190_195_groupi_n_633, csa_tree_add_190_195_groupi_n_634, csa_tree_add_190_195_groupi_n_635, csa_tree_add_190_195_groupi_n_636, csa_tree_add_190_195_groupi_n_637, csa_tree_add_190_195_groupi_n_638, csa_tree_add_190_195_groupi_n_639, csa_tree_add_190_195_groupi_n_640;
  wire csa_tree_add_190_195_groupi_n_641, csa_tree_add_190_195_groupi_n_642, csa_tree_add_190_195_groupi_n_643, csa_tree_add_190_195_groupi_n_644, csa_tree_add_190_195_groupi_n_645, csa_tree_add_190_195_groupi_n_646, csa_tree_add_190_195_groupi_n_647, csa_tree_add_190_195_groupi_n_648;
  wire csa_tree_add_190_195_groupi_n_649, csa_tree_add_190_195_groupi_n_650, csa_tree_add_190_195_groupi_n_651, csa_tree_add_190_195_groupi_n_652, csa_tree_add_190_195_groupi_n_653, csa_tree_add_190_195_groupi_n_654, csa_tree_add_190_195_groupi_n_655, csa_tree_add_190_195_groupi_n_656;
  wire csa_tree_add_190_195_groupi_n_657, csa_tree_add_190_195_groupi_n_658, csa_tree_add_190_195_groupi_n_659, csa_tree_add_190_195_groupi_n_660, csa_tree_add_190_195_groupi_n_661, csa_tree_add_190_195_groupi_n_662, csa_tree_add_190_195_groupi_n_663, csa_tree_add_190_195_groupi_n_664;
  wire csa_tree_add_190_195_groupi_n_665, csa_tree_add_190_195_groupi_n_666, csa_tree_add_190_195_groupi_n_667, csa_tree_add_190_195_groupi_n_668, csa_tree_add_190_195_groupi_n_669, csa_tree_add_190_195_groupi_n_670, csa_tree_add_190_195_groupi_n_671, csa_tree_add_190_195_groupi_n_672;
  wire csa_tree_add_190_195_groupi_n_673, csa_tree_add_190_195_groupi_n_674, csa_tree_add_190_195_groupi_n_675, csa_tree_add_190_195_groupi_n_676, csa_tree_add_190_195_groupi_n_677, csa_tree_add_190_195_groupi_n_678, csa_tree_add_190_195_groupi_n_679, csa_tree_add_190_195_groupi_n_680;
  wire csa_tree_add_190_195_groupi_n_681, csa_tree_add_190_195_groupi_n_682, csa_tree_add_190_195_groupi_n_683, csa_tree_add_190_195_groupi_n_684, csa_tree_add_190_195_groupi_n_685, csa_tree_add_190_195_groupi_n_686, csa_tree_add_190_195_groupi_n_687, csa_tree_add_190_195_groupi_n_688;
  wire csa_tree_add_190_195_groupi_n_689, csa_tree_add_190_195_groupi_n_690, csa_tree_add_190_195_groupi_n_691, csa_tree_add_190_195_groupi_n_692, csa_tree_add_190_195_groupi_n_693, csa_tree_add_190_195_groupi_n_694, csa_tree_add_190_195_groupi_n_695, csa_tree_add_190_195_groupi_n_696;
  wire csa_tree_add_190_195_groupi_n_697, csa_tree_add_190_195_groupi_n_698, csa_tree_add_190_195_groupi_n_699, csa_tree_add_190_195_groupi_n_700, csa_tree_add_190_195_groupi_n_701, csa_tree_add_190_195_groupi_n_702, csa_tree_add_190_195_groupi_n_703, csa_tree_add_190_195_groupi_n_704;
  wire csa_tree_add_190_195_groupi_n_705, csa_tree_add_190_195_groupi_n_706, csa_tree_add_190_195_groupi_n_707, csa_tree_add_190_195_groupi_n_708, csa_tree_add_190_195_groupi_n_709, csa_tree_add_190_195_groupi_n_710, csa_tree_add_190_195_groupi_n_711, csa_tree_add_190_195_groupi_n_712;
  wire csa_tree_add_190_195_groupi_n_713, csa_tree_add_190_195_groupi_n_714, csa_tree_add_190_195_groupi_n_715, csa_tree_add_190_195_groupi_n_716, csa_tree_add_190_195_groupi_n_717, csa_tree_add_190_195_groupi_n_718, csa_tree_add_190_195_groupi_n_719, csa_tree_add_190_195_groupi_n_720;
  wire csa_tree_add_190_195_groupi_n_721, csa_tree_add_190_195_groupi_n_722, csa_tree_add_190_195_groupi_n_723, csa_tree_add_190_195_groupi_n_724, csa_tree_add_190_195_groupi_n_725, csa_tree_add_190_195_groupi_n_726, csa_tree_add_190_195_groupi_n_727, csa_tree_add_190_195_groupi_n_728;
  wire csa_tree_add_190_195_groupi_n_729, csa_tree_add_190_195_groupi_n_730, csa_tree_add_190_195_groupi_n_731, csa_tree_add_190_195_groupi_n_732, csa_tree_add_190_195_groupi_n_733, csa_tree_add_190_195_groupi_n_734, csa_tree_add_190_195_groupi_n_735, csa_tree_add_190_195_groupi_n_736;
  wire csa_tree_add_190_195_groupi_n_737, csa_tree_add_190_195_groupi_n_738, csa_tree_add_190_195_groupi_n_739, csa_tree_add_190_195_groupi_n_740, csa_tree_add_190_195_groupi_n_741, csa_tree_add_190_195_groupi_n_742, csa_tree_add_190_195_groupi_n_743, csa_tree_add_190_195_groupi_n_744;
  wire csa_tree_add_190_195_groupi_n_745, csa_tree_add_190_195_groupi_n_746, csa_tree_add_190_195_groupi_n_747, csa_tree_add_190_195_groupi_n_748, csa_tree_add_190_195_groupi_n_749, csa_tree_add_190_195_groupi_n_750, csa_tree_add_190_195_groupi_n_751, csa_tree_add_190_195_groupi_n_752;
  wire csa_tree_add_190_195_groupi_n_753, csa_tree_add_190_195_groupi_n_754, csa_tree_add_190_195_groupi_n_755, csa_tree_add_190_195_groupi_n_756, csa_tree_add_190_195_groupi_n_757, csa_tree_add_190_195_groupi_n_758, csa_tree_add_190_195_groupi_n_759, csa_tree_add_190_195_groupi_n_760;
  wire csa_tree_add_190_195_groupi_n_761, csa_tree_add_190_195_groupi_n_762, csa_tree_add_190_195_groupi_n_763, csa_tree_add_190_195_groupi_n_764, csa_tree_add_190_195_groupi_n_765, csa_tree_add_190_195_groupi_n_766, csa_tree_add_190_195_groupi_n_767, csa_tree_add_190_195_groupi_n_768;
  wire csa_tree_add_190_195_groupi_n_769, csa_tree_add_190_195_groupi_n_770, csa_tree_add_190_195_groupi_n_771, csa_tree_add_190_195_groupi_n_772, csa_tree_add_190_195_groupi_n_773, csa_tree_add_190_195_groupi_n_774, csa_tree_add_190_195_groupi_n_775, csa_tree_add_190_195_groupi_n_776;
  wire csa_tree_add_190_195_groupi_n_777, csa_tree_add_190_195_groupi_n_778, csa_tree_add_190_195_groupi_n_779, csa_tree_add_190_195_groupi_n_780, csa_tree_add_190_195_groupi_n_781, csa_tree_add_190_195_groupi_n_782, csa_tree_add_190_195_groupi_n_783, csa_tree_add_190_195_groupi_n_784;
  wire csa_tree_add_190_195_groupi_n_785, csa_tree_add_190_195_groupi_n_786, csa_tree_add_190_195_groupi_n_787, csa_tree_add_190_195_groupi_n_788, csa_tree_add_190_195_groupi_n_789, csa_tree_add_190_195_groupi_n_790, csa_tree_add_190_195_groupi_n_791, csa_tree_add_190_195_groupi_n_792;
  wire csa_tree_add_190_195_groupi_n_793, csa_tree_add_190_195_groupi_n_794, csa_tree_add_190_195_groupi_n_795, csa_tree_add_190_195_groupi_n_796, csa_tree_add_190_195_groupi_n_797, csa_tree_add_190_195_groupi_n_798, csa_tree_add_190_195_groupi_n_799, csa_tree_add_190_195_groupi_n_800;
  wire csa_tree_add_190_195_groupi_n_801, csa_tree_add_190_195_groupi_n_802, csa_tree_add_190_195_groupi_n_803, csa_tree_add_190_195_groupi_n_804, csa_tree_add_190_195_groupi_n_805, csa_tree_add_190_195_groupi_n_806, csa_tree_add_190_195_groupi_n_807, csa_tree_add_190_195_groupi_n_808;
  wire csa_tree_add_190_195_groupi_n_809, csa_tree_add_190_195_groupi_n_810, csa_tree_add_190_195_groupi_n_811, csa_tree_add_190_195_groupi_n_812, csa_tree_add_190_195_groupi_n_813, csa_tree_add_190_195_groupi_n_814, csa_tree_add_190_195_groupi_n_815, csa_tree_add_190_195_groupi_n_816;
  wire csa_tree_add_190_195_groupi_n_817, csa_tree_add_190_195_groupi_n_818, csa_tree_add_190_195_groupi_n_819, csa_tree_add_190_195_groupi_n_820, csa_tree_add_190_195_groupi_n_821, csa_tree_add_190_195_groupi_n_822, csa_tree_add_190_195_groupi_n_823, csa_tree_add_190_195_groupi_n_824;
  wire csa_tree_add_190_195_groupi_n_825, csa_tree_add_190_195_groupi_n_826, csa_tree_add_190_195_groupi_n_827, csa_tree_add_190_195_groupi_n_828, csa_tree_add_190_195_groupi_n_829, csa_tree_add_190_195_groupi_n_830, csa_tree_add_190_195_groupi_n_831, csa_tree_add_190_195_groupi_n_832;
  wire csa_tree_add_190_195_groupi_n_833, csa_tree_add_190_195_groupi_n_834, csa_tree_add_190_195_groupi_n_835, csa_tree_add_190_195_groupi_n_836, csa_tree_add_190_195_groupi_n_837, csa_tree_add_190_195_groupi_n_838, csa_tree_add_190_195_groupi_n_839, csa_tree_add_190_195_groupi_n_840;
  wire csa_tree_add_190_195_groupi_n_841, csa_tree_add_190_195_groupi_n_842, csa_tree_add_190_195_groupi_n_843, csa_tree_add_190_195_groupi_n_844, csa_tree_add_190_195_groupi_n_845, csa_tree_add_190_195_groupi_n_846, csa_tree_add_190_195_groupi_n_847, csa_tree_add_190_195_groupi_n_848;
  wire csa_tree_add_190_195_groupi_n_849, csa_tree_add_190_195_groupi_n_850, csa_tree_add_190_195_groupi_n_851, csa_tree_add_190_195_groupi_n_852, csa_tree_add_190_195_groupi_n_853, csa_tree_add_190_195_groupi_n_854, csa_tree_add_190_195_groupi_n_855, csa_tree_add_190_195_groupi_n_856;
  wire csa_tree_add_190_195_groupi_n_857, csa_tree_add_190_195_groupi_n_858, csa_tree_add_190_195_groupi_n_859, csa_tree_add_190_195_groupi_n_860, csa_tree_add_190_195_groupi_n_861, csa_tree_add_190_195_groupi_n_862, csa_tree_add_190_195_groupi_n_863, csa_tree_add_190_195_groupi_n_864;
  wire csa_tree_add_190_195_groupi_n_865, csa_tree_add_190_195_groupi_n_866, csa_tree_add_190_195_groupi_n_867, csa_tree_add_190_195_groupi_n_868, csa_tree_add_190_195_groupi_n_869, csa_tree_add_190_195_groupi_n_870, csa_tree_add_190_195_groupi_n_871, csa_tree_add_190_195_groupi_n_872;
  wire csa_tree_add_190_195_groupi_n_873, csa_tree_add_190_195_groupi_n_874, csa_tree_add_190_195_groupi_n_875, csa_tree_add_190_195_groupi_n_876, csa_tree_add_190_195_groupi_n_877, csa_tree_add_190_195_groupi_n_878, csa_tree_add_190_195_groupi_n_879, csa_tree_add_190_195_groupi_n_880;
  wire csa_tree_add_190_195_groupi_n_881, csa_tree_add_190_195_groupi_n_882, csa_tree_add_190_195_groupi_n_883, csa_tree_add_190_195_groupi_n_884, csa_tree_add_190_195_groupi_n_885, csa_tree_add_190_195_groupi_n_886, csa_tree_add_190_195_groupi_n_887, csa_tree_add_190_195_groupi_n_888;
  wire csa_tree_add_190_195_groupi_n_889, csa_tree_add_190_195_groupi_n_890, csa_tree_add_190_195_groupi_n_891, csa_tree_add_190_195_groupi_n_892, csa_tree_add_190_195_groupi_n_893, csa_tree_add_190_195_groupi_n_894, csa_tree_add_190_195_groupi_n_895, csa_tree_add_190_195_groupi_n_896;
  wire csa_tree_add_190_195_groupi_n_897, csa_tree_add_190_195_groupi_n_898, csa_tree_add_190_195_groupi_n_899, csa_tree_add_190_195_groupi_n_900, csa_tree_add_190_195_groupi_n_901, csa_tree_add_190_195_groupi_n_902, csa_tree_add_190_195_groupi_n_903, csa_tree_add_190_195_groupi_n_904;
  wire csa_tree_add_190_195_groupi_n_905, csa_tree_add_190_195_groupi_n_906, csa_tree_add_190_195_groupi_n_907, csa_tree_add_190_195_groupi_n_908, csa_tree_add_190_195_groupi_n_909, csa_tree_add_190_195_groupi_n_910, csa_tree_add_190_195_groupi_n_911, csa_tree_add_190_195_groupi_n_912;
  wire csa_tree_add_190_195_groupi_n_913, csa_tree_add_190_195_groupi_n_914, csa_tree_add_190_195_groupi_n_915, csa_tree_add_190_195_groupi_n_916, csa_tree_add_190_195_groupi_n_917, csa_tree_add_190_195_groupi_n_918, csa_tree_add_190_195_groupi_n_919, csa_tree_add_190_195_groupi_n_920;
  wire csa_tree_add_190_195_groupi_n_921, csa_tree_add_190_195_groupi_n_922, csa_tree_add_190_195_groupi_n_923, csa_tree_add_190_195_groupi_n_924, csa_tree_add_190_195_groupi_n_925, csa_tree_add_190_195_groupi_n_926, csa_tree_add_190_195_groupi_n_927, csa_tree_add_190_195_groupi_n_928;
  wire csa_tree_add_190_195_groupi_n_929, csa_tree_add_190_195_groupi_n_930, csa_tree_add_190_195_groupi_n_931, csa_tree_add_190_195_groupi_n_932, csa_tree_add_190_195_groupi_n_933, csa_tree_add_190_195_groupi_n_934, csa_tree_add_190_195_groupi_n_935, csa_tree_add_190_195_groupi_n_936;
  wire csa_tree_add_190_195_groupi_n_937, csa_tree_add_190_195_groupi_n_938, csa_tree_add_190_195_groupi_n_939, csa_tree_add_190_195_groupi_n_940, csa_tree_add_190_195_groupi_n_941, csa_tree_add_190_195_groupi_n_942, csa_tree_add_190_195_groupi_n_943, csa_tree_add_190_195_groupi_n_944;
  wire csa_tree_add_190_195_groupi_n_945, csa_tree_add_190_195_groupi_n_946, csa_tree_add_190_195_groupi_n_947, csa_tree_add_190_195_groupi_n_948, csa_tree_add_190_195_groupi_n_949, csa_tree_add_190_195_groupi_n_950, csa_tree_add_190_195_groupi_n_951, csa_tree_add_190_195_groupi_n_952;
  wire csa_tree_add_190_195_groupi_n_953, csa_tree_add_190_195_groupi_n_954, csa_tree_add_190_195_groupi_n_955, csa_tree_add_190_195_groupi_n_956, csa_tree_add_190_195_groupi_n_957, csa_tree_add_190_195_groupi_n_958, csa_tree_add_190_195_groupi_n_959, csa_tree_add_190_195_groupi_n_960;
  wire csa_tree_add_190_195_groupi_n_961, csa_tree_add_190_195_groupi_n_962, csa_tree_add_190_195_groupi_n_963, csa_tree_add_190_195_groupi_n_964, csa_tree_add_190_195_groupi_n_965, csa_tree_add_190_195_groupi_n_966, csa_tree_add_190_195_groupi_n_967, csa_tree_add_190_195_groupi_n_968;
  wire csa_tree_add_190_195_groupi_n_969, csa_tree_add_190_195_groupi_n_970, csa_tree_add_190_195_groupi_n_971, csa_tree_add_190_195_groupi_n_972, csa_tree_add_190_195_groupi_n_973, csa_tree_add_190_195_groupi_n_974, csa_tree_add_190_195_groupi_n_975, csa_tree_add_190_195_groupi_n_976;
  wire csa_tree_add_190_195_groupi_n_977, csa_tree_add_190_195_groupi_n_978, csa_tree_add_190_195_groupi_n_979, csa_tree_add_190_195_groupi_n_980, csa_tree_add_190_195_groupi_n_981, csa_tree_add_190_195_groupi_n_982, csa_tree_add_190_195_groupi_n_983, csa_tree_add_190_195_groupi_n_984;
  wire csa_tree_add_190_195_groupi_n_985, csa_tree_add_190_195_groupi_n_986, csa_tree_add_190_195_groupi_n_987, csa_tree_add_190_195_groupi_n_988, csa_tree_add_190_195_groupi_n_989, csa_tree_add_190_195_groupi_n_990, csa_tree_add_190_195_groupi_n_991, csa_tree_add_190_195_groupi_n_992;
  wire csa_tree_add_190_195_groupi_n_993, csa_tree_add_190_195_groupi_n_994, csa_tree_add_190_195_groupi_n_995, csa_tree_add_190_195_groupi_n_996, csa_tree_add_190_195_groupi_n_997, csa_tree_add_190_195_groupi_n_998, csa_tree_add_190_195_groupi_n_999, csa_tree_add_190_195_groupi_n_1000;
  wire csa_tree_add_190_195_groupi_n_1001, csa_tree_add_190_195_groupi_n_1002, csa_tree_add_190_195_groupi_n_1003, csa_tree_add_190_195_groupi_n_1004, csa_tree_add_190_195_groupi_n_1005, csa_tree_add_190_195_groupi_n_1006, csa_tree_add_190_195_groupi_n_1007, csa_tree_add_190_195_groupi_n_1008;
  wire csa_tree_add_190_195_groupi_n_1009, csa_tree_add_190_195_groupi_n_1010, csa_tree_add_190_195_groupi_n_1011, csa_tree_add_190_195_groupi_n_1012, csa_tree_add_190_195_groupi_n_1013, csa_tree_add_190_195_groupi_n_1014, csa_tree_add_190_195_groupi_n_1015, csa_tree_add_190_195_groupi_n_1016;
  wire csa_tree_add_190_195_groupi_n_1017, csa_tree_add_190_195_groupi_n_1018, csa_tree_add_190_195_groupi_n_1019, csa_tree_add_190_195_groupi_n_1020, csa_tree_add_190_195_groupi_n_1021, csa_tree_add_190_195_groupi_n_1022, csa_tree_add_190_195_groupi_n_1023, csa_tree_add_190_195_groupi_n_1024;
  wire csa_tree_add_190_195_groupi_n_1025, csa_tree_add_190_195_groupi_n_1026, csa_tree_add_190_195_groupi_n_1027, csa_tree_add_190_195_groupi_n_1028, csa_tree_add_190_195_groupi_n_1029, csa_tree_add_190_195_groupi_n_1030, csa_tree_add_190_195_groupi_n_1031, csa_tree_add_190_195_groupi_n_1032;
  wire csa_tree_add_190_195_groupi_n_1033, csa_tree_add_190_195_groupi_n_1034, csa_tree_add_190_195_groupi_n_1035, csa_tree_add_190_195_groupi_n_1036, csa_tree_add_190_195_groupi_n_1037, csa_tree_add_190_195_groupi_n_1038, csa_tree_add_190_195_groupi_n_1039, csa_tree_add_190_195_groupi_n_1040;
  wire csa_tree_add_190_195_groupi_n_1041, csa_tree_add_190_195_groupi_n_1042, csa_tree_add_190_195_groupi_n_1043, csa_tree_add_190_195_groupi_n_1044, csa_tree_add_190_195_groupi_n_1045, csa_tree_add_190_195_groupi_n_1046, csa_tree_add_190_195_groupi_n_1047, csa_tree_add_190_195_groupi_n_1048;
  wire csa_tree_add_190_195_groupi_n_1049, csa_tree_add_190_195_groupi_n_1050, csa_tree_add_190_195_groupi_n_1051, csa_tree_add_190_195_groupi_n_1052, csa_tree_add_190_195_groupi_n_1053, csa_tree_add_190_195_groupi_n_1054, csa_tree_add_190_195_groupi_n_1055, csa_tree_add_190_195_groupi_n_1056;
  wire csa_tree_add_190_195_groupi_n_1057, csa_tree_add_190_195_groupi_n_1058, csa_tree_add_190_195_groupi_n_1059, csa_tree_add_190_195_groupi_n_1060, csa_tree_add_190_195_groupi_n_1061, csa_tree_add_190_195_groupi_n_1062, csa_tree_add_190_195_groupi_n_1063, csa_tree_add_190_195_groupi_n_1064;
  wire csa_tree_add_190_195_groupi_n_1065, csa_tree_add_190_195_groupi_n_1066, csa_tree_add_190_195_groupi_n_1067, csa_tree_add_190_195_groupi_n_1068, csa_tree_add_190_195_groupi_n_1069, csa_tree_add_190_195_groupi_n_1070, csa_tree_add_190_195_groupi_n_1071, csa_tree_add_190_195_groupi_n_1072;
  wire csa_tree_add_190_195_groupi_n_1073, csa_tree_add_190_195_groupi_n_1074, csa_tree_add_190_195_groupi_n_1075, csa_tree_add_190_195_groupi_n_1076, csa_tree_add_190_195_groupi_n_1077, csa_tree_add_190_195_groupi_n_1078, csa_tree_add_190_195_groupi_n_1079, csa_tree_add_190_195_groupi_n_1080;
  wire csa_tree_add_190_195_groupi_n_1081, csa_tree_add_190_195_groupi_n_1082, csa_tree_add_190_195_groupi_n_1083, csa_tree_add_190_195_groupi_n_1084, csa_tree_add_190_195_groupi_n_1085, csa_tree_add_190_195_groupi_n_1086, csa_tree_add_190_195_groupi_n_1087, csa_tree_add_190_195_groupi_n_1088;
  wire csa_tree_add_190_195_groupi_n_1089, csa_tree_add_190_195_groupi_n_1090, csa_tree_add_190_195_groupi_n_1091, csa_tree_add_190_195_groupi_n_1092, csa_tree_add_190_195_groupi_n_1093, csa_tree_add_190_195_groupi_n_1094, csa_tree_add_190_195_groupi_n_1095, csa_tree_add_190_195_groupi_n_1096;
  wire csa_tree_add_190_195_groupi_n_1097, csa_tree_add_190_195_groupi_n_1098, csa_tree_add_190_195_groupi_n_1099, csa_tree_add_190_195_groupi_n_1100, csa_tree_add_190_195_groupi_n_1101, csa_tree_add_190_195_groupi_n_1102, csa_tree_add_190_195_groupi_n_1103, csa_tree_add_190_195_groupi_n_1104;
  wire csa_tree_add_190_195_groupi_n_1105, csa_tree_add_190_195_groupi_n_1106, csa_tree_add_190_195_groupi_n_1107, csa_tree_add_190_195_groupi_n_1108, csa_tree_add_190_195_groupi_n_1109, csa_tree_add_190_195_groupi_n_1110, csa_tree_add_190_195_groupi_n_1111, csa_tree_add_190_195_groupi_n_1112;
  wire csa_tree_add_190_195_groupi_n_1113, csa_tree_add_190_195_groupi_n_1114, csa_tree_add_190_195_groupi_n_1115, csa_tree_add_190_195_groupi_n_1116, csa_tree_add_190_195_groupi_n_1117, csa_tree_add_190_195_groupi_n_1118, csa_tree_add_190_195_groupi_n_1119, csa_tree_add_190_195_groupi_n_1120;
  wire csa_tree_add_190_195_groupi_n_1121, csa_tree_add_190_195_groupi_n_1122, csa_tree_add_190_195_groupi_n_1123, csa_tree_add_190_195_groupi_n_1124, csa_tree_add_190_195_groupi_n_1125, csa_tree_add_190_195_groupi_n_1126, csa_tree_add_190_195_groupi_n_1127, csa_tree_add_190_195_groupi_n_1128;
  wire csa_tree_add_190_195_groupi_n_1129, csa_tree_add_190_195_groupi_n_1130, csa_tree_add_190_195_groupi_n_1131, csa_tree_add_190_195_groupi_n_1132, csa_tree_add_190_195_groupi_n_1133, csa_tree_add_190_195_groupi_n_1134, csa_tree_add_190_195_groupi_n_1135, csa_tree_add_190_195_groupi_n_1136;
  wire csa_tree_add_190_195_groupi_n_1137, csa_tree_add_190_195_groupi_n_1138, csa_tree_add_190_195_groupi_n_1139, csa_tree_add_190_195_groupi_n_1140, csa_tree_add_190_195_groupi_n_1141, csa_tree_add_190_195_groupi_n_1142, csa_tree_add_190_195_groupi_n_1143, csa_tree_add_190_195_groupi_n_1144;
  wire csa_tree_add_190_195_groupi_n_1145, csa_tree_add_190_195_groupi_n_1146, csa_tree_add_190_195_groupi_n_1147, csa_tree_add_190_195_groupi_n_1148, csa_tree_add_190_195_groupi_n_1149, csa_tree_add_190_195_groupi_n_1150, csa_tree_add_190_195_groupi_n_1151, csa_tree_add_190_195_groupi_n_1152;
  wire csa_tree_add_190_195_groupi_n_1153, csa_tree_add_190_195_groupi_n_1154, csa_tree_add_190_195_groupi_n_1155, csa_tree_add_190_195_groupi_n_1156, csa_tree_add_190_195_groupi_n_1157, csa_tree_add_190_195_groupi_n_1158, csa_tree_add_190_195_groupi_n_1159, csa_tree_add_190_195_groupi_n_1160;
  wire csa_tree_add_190_195_groupi_n_1161, csa_tree_add_190_195_groupi_n_1162, csa_tree_add_190_195_groupi_n_1163, csa_tree_add_190_195_groupi_n_1164, csa_tree_add_190_195_groupi_n_1165, csa_tree_add_190_195_groupi_n_1166, csa_tree_add_190_195_groupi_n_1167, csa_tree_add_190_195_groupi_n_1168;
  wire csa_tree_add_190_195_groupi_n_1169, csa_tree_add_190_195_groupi_n_1170, csa_tree_add_190_195_groupi_n_1171, csa_tree_add_190_195_groupi_n_1172, csa_tree_add_190_195_groupi_n_1173, csa_tree_add_190_195_groupi_n_1174, csa_tree_add_190_195_groupi_n_1175, csa_tree_add_190_195_groupi_n_1176;
  wire csa_tree_add_190_195_groupi_n_1177, csa_tree_add_190_195_groupi_n_1178, csa_tree_add_190_195_groupi_n_1179, csa_tree_add_190_195_groupi_n_1180, csa_tree_add_190_195_groupi_n_1181, csa_tree_add_190_195_groupi_n_1182, csa_tree_add_190_195_groupi_n_1183, csa_tree_add_190_195_groupi_n_1184;
  wire csa_tree_add_190_195_groupi_n_1185, csa_tree_add_190_195_groupi_n_1186, csa_tree_add_190_195_groupi_n_1187, csa_tree_add_190_195_groupi_n_1188, csa_tree_add_190_195_groupi_n_1189, csa_tree_add_190_195_groupi_n_1190, csa_tree_add_190_195_groupi_n_1191, csa_tree_add_190_195_groupi_n_1192;
  wire csa_tree_add_190_195_groupi_n_1193, csa_tree_add_190_195_groupi_n_1194, csa_tree_add_190_195_groupi_n_1195, csa_tree_add_190_195_groupi_n_1196, csa_tree_add_190_195_groupi_n_1197, csa_tree_add_190_195_groupi_n_1198, csa_tree_add_190_195_groupi_n_1199, csa_tree_add_190_195_groupi_n_1200;
  wire csa_tree_add_190_195_groupi_n_1201, csa_tree_add_190_195_groupi_n_1202, csa_tree_add_190_195_groupi_n_1203, csa_tree_add_190_195_groupi_n_1204, csa_tree_add_190_195_groupi_n_1205, csa_tree_add_190_195_groupi_n_1206, csa_tree_add_190_195_groupi_n_1207, csa_tree_add_190_195_groupi_n_1208;
  wire csa_tree_add_190_195_groupi_n_1209, csa_tree_add_190_195_groupi_n_1210, csa_tree_add_190_195_groupi_n_1211, csa_tree_add_190_195_groupi_n_1212, csa_tree_add_190_195_groupi_n_1213, csa_tree_add_190_195_groupi_n_1214, csa_tree_add_190_195_groupi_n_1215, csa_tree_add_190_195_groupi_n_1216;
  wire csa_tree_add_190_195_groupi_n_1217, csa_tree_add_190_195_groupi_n_1218, csa_tree_add_190_195_groupi_n_1219, csa_tree_add_190_195_groupi_n_1220, csa_tree_add_190_195_groupi_n_1221, csa_tree_add_190_195_groupi_n_1222, csa_tree_add_190_195_groupi_n_1223, csa_tree_add_190_195_groupi_n_1224;
  wire csa_tree_add_190_195_groupi_n_1225, csa_tree_add_190_195_groupi_n_1226, csa_tree_add_190_195_groupi_n_1227, csa_tree_add_190_195_groupi_n_1228, csa_tree_add_190_195_groupi_n_1229, csa_tree_add_190_195_groupi_n_1230, csa_tree_add_190_195_groupi_n_1231, csa_tree_add_190_195_groupi_n_1232;
  wire csa_tree_add_190_195_groupi_n_1233, csa_tree_add_190_195_groupi_n_1234, csa_tree_add_190_195_groupi_n_1235, csa_tree_add_190_195_groupi_n_1236, csa_tree_add_190_195_groupi_n_1237, csa_tree_add_190_195_groupi_n_1238, csa_tree_add_190_195_groupi_n_1239, csa_tree_add_190_195_groupi_n_1240;
  wire csa_tree_add_190_195_groupi_n_1241, csa_tree_add_190_195_groupi_n_1242, csa_tree_add_190_195_groupi_n_1243, csa_tree_add_190_195_groupi_n_1244, csa_tree_add_190_195_groupi_n_1245, csa_tree_add_190_195_groupi_n_1246, csa_tree_add_190_195_groupi_n_1247, csa_tree_add_190_195_groupi_n_1248;
  wire csa_tree_add_190_195_groupi_n_1249, csa_tree_add_190_195_groupi_n_1250, csa_tree_add_190_195_groupi_n_1251, csa_tree_add_190_195_groupi_n_1252, csa_tree_add_190_195_groupi_n_1253, csa_tree_add_190_195_groupi_n_1254, csa_tree_add_190_195_groupi_n_1255, csa_tree_add_190_195_groupi_n_1256;
  wire csa_tree_add_190_195_groupi_n_1257, csa_tree_add_190_195_groupi_n_1258, csa_tree_add_190_195_groupi_n_1259, csa_tree_add_190_195_groupi_n_1260, csa_tree_add_190_195_groupi_n_1261, csa_tree_add_190_195_groupi_n_1262, csa_tree_add_190_195_groupi_n_1263, csa_tree_add_190_195_groupi_n_1264;
  wire csa_tree_add_190_195_groupi_n_1265, csa_tree_add_190_195_groupi_n_1266, csa_tree_add_190_195_groupi_n_1267, csa_tree_add_190_195_groupi_n_1268, csa_tree_add_190_195_groupi_n_1269, csa_tree_add_190_195_groupi_n_1270, csa_tree_add_190_195_groupi_n_1271, csa_tree_add_190_195_groupi_n_1272;
  wire csa_tree_add_190_195_groupi_n_1273, csa_tree_add_190_195_groupi_n_1274, csa_tree_add_190_195_groupi_n_1275, csa_tree_add_190_195_groupi_n_1276, csa_tree_add_190_195_groupi_n_1277, csa_tree_add_190_195_groupi_n_1278, csa_tree_add_190_195_groupi_n_1279, csa_tree_add_190_195_groupi_n_1280;
  wire csa_tree_add_190_195_groupi_n_1281, csa_tree_add_190_195_groupi_n_1282, csa_tree_add_190_195_groupi_n_1283, csa_tree_add_190_195_groupi_n_1284, csa_tree_add_190_195_groupi_n_1285, csa_tree_add_190_195_groupi_n_1286, csa_tree_add_190_195_groupi_n_1287, csa_tree_add_190_195_groupi_n_1288;
  wire csa_tree_add_190_195_groupi_n_1289, csa_tree_add_190_195_groupi_n_1290, csa_tree_add_190_195_groupi_n_1291, csa_tree_add_190_195_groupi_n_1292, csa_tree_add_190_195_groupi_n_1293, csa_tree_add_190_195_groupi_n_1294, csa_tree_add_190_195_groupi_n_1295, csa_tree_add_190_195_groupi_n_1296;
  wire csa_tree_add_190_195_groupi_n_1297, csa_tree_add_190_195_groupi_n_1298, csa_tree_add_190_195_groupi_n_1299, csa_tree_add_190_195_groupi_n_1300, csa_tree_add_190_195_groupi_n_1301, csa_tree_add_190_195_groupi_n_1302, csa_tree_add_190_195_groupi_n_1303, csa_tree_add_190_195_groupi_n_1304;
  wire csa_tree_add_190_195_groupi_n_1305, csa_tree_add_190_195_groupi_n_1306, csa_tree_add_190_195_groupi_n_1307, csa_tree_add_190_195_groupi_n_1308, csa_tree_add_190_195_groupi_n_1309, csa_tree_add_190_195_groupi_n_1310, csa_tree_add_190_195_groupi_n_1311, csa_tree_add_190_195_groupi_n_1312;
  wire csa_tree_add_190_195_groupi_n_1313, csa_tree_add_190_195_groupi_n_1314, csa_tree_add_190_195_groupi_n_1329, csa_tree_add_190_195_groupi_n_1330, csa_tree_add_190_195_groupi_n_1331, csa_tree_add_190_195_groupi_n_1332, csa_tree_add_190_195_groupi_n_1333, csa_tree_add_190_195_groupi_n_1334;
  wire csa_tree_add_190_195_groupi_n_1335, csa_tree_add_190_195_groupi_n_1336, csa_tree_add_190_195_groupi_n_1337, csa_tree_add_190_195_groupi_n_1338, csa_tree_add_190_195_groupi_n_1339, csa_tree_add_190_195_groupi_n_1340, csa_tree_add_190_195_groupi_n_1341, csa_tree_add_190_195_groupi_n_1342;
  wire csa_tree_add_190_195_groupi_n_1343, csa_tree_add_190_195_groupi_n_1344, csa_tree_add_190_195_groupi_n_1345, csa_tree_add_190_195_groupi_n_1346, csa_tree_add_190_195_groupi_n_1347, csa_tree_add_190_195_groupi_n_1348, csa_tree_add_190_195_groupi_n_1349, csa_tree_add_190_195_groupi_n_1350;
  wire csa_tree_add_190_195_groupi_n_1351, csa_tree_add_190_195_groupi_n_1352, csa_tree_add_190_195_groupi_n_1353, csa_tree_add_190_195_groupi_n_1354, csa_tree_add_190_195_groupi_n_1355, csa_tree_add_190_195_groupi_n_1356, csa_tree_add_190_195_groupi_n_1357, csa_tree_add_190_195_groupi_n_1358;
  wire csa_tree_add_190_195_groupi_n_1359, csa_tree_add_190_195_groupi_n_1360, csa_tree_add_190_195_groupi_n_1361, csa_tree_add_190_195_groupi_n_1362, csa_tree_add_190_195_groupi_n_1363, csa_tree_add_190_195_groupi_n_1364, csa_tree_add_190_195_groupi_n_1365, csa_tree_add_190_195_groupi_n_1366;
  wire csa_tree_add_190_195_groupi_n_1367, csa_tree_add_190_195_groupi_n_1368, csa_tree_add_190_195_groupi_n_1369, csa_tree_add_190_195_groupi_n_1370, csa_tree_add_190_195_groupi_n_1371, csa_tree_add_190_195_groupi_n_1372, csa_tree_add_190_195_groupi_n_1373, csa_tree_add_190_195_groupi_n_1374;
  wire csa_tree_add_190_195_groupi_n_1375, csa_tree_add_190_195_groupi_n_1376, csa_tree_add_190_195_groupi_n_1377, csa_tree_add_190_195_groupi_n_1378, csa_tree_add_190_195_groupi_n_1379, csa_tree_add_190_195_groupi_n_1380, csa_tree_add_190_195_groupi_n_1381, csa_tree_add_190_195_groupi_n_1382;
  wire csa_tree_add_190_195_groupi_n_1383, csa_tree_add_190_195_groupi_n_1384, csa_tree_add_190_195_groupi_n_1385, csa_tree_add_190_195_groupi_n_1386, csa_tree_add_190_195_groupi_n_1387, csa_tree_add_190_195_groupi_n_1388, csa_tree_add_190_195_groupi_n_1389, csa_tree_add_190_195_groupi_n_1390;
  wire csa_tree_add_190_195_groupi_n_1391, csa_tree_add_190_195_groupi_n_1392, csa_tree_add_190_195_groupi_n_1393, csa_tree_add_190_195_groupi_n_1394, csa_tree_add_190_195_groupi_n_1395, csa_tree_add_190_195_groupi_n_1396, csa_tree_add_190_195_groupi_n_1397, csa_tree_add_190_195_groupi_n_1398;
  wire csa_tree_add_190_195_groupi_n_1399, csa_tree_add_190_195_groupi_n_1400, csa_tree_add_190_195_groupi_n_1401, csa_tree_add_190_195_groupi_n_1402, csa_tree_add_190_195_groupi_n_1403, csa_tree_add_190_195_groupi_n_1404, csa_tree_add_190_195_groupi_n_1405, csa_tree_add_190_195_groupi_n_1406;
  wire csa_tree_add_190_195_groupi_n_1407, csa_tree_add_190_195_groupi_n_1408, csa_tree_add_190_195_groupi_n_1409, csa_tree_add_190_195_groupi_n_1410, csa_tree_add_190_195_groupi_n_1411, csa_tree_add_190_195_groupi_n_1412, csa_tree_add_190_195_groupi_n_1413, csa_tree_add_190_195_groupi_n_1414;
  wire csa_tree_add_190_195_groupi_n_1415, csa_tree_add_190_195_groupi_n_1416, csa_tree_add_190_195_groupi_n_1417, csa_tree_add_190_195_groupi_n_1418, csa_tree_add_190_195_groupi_n_1419, csa_tree_add_190_195_groupi_n_1420, csa_tree_add_190_195_groupi_n_1421, csa_tree_add_190_195_groupi_n_1422;
  wire csa_tree_add_190_195_groupi_n_1423, csa_tree_add_190_195_groupi_n_1424, csa_tree_add_190_195_groupi_n_1425, csa_tree_add_190_195_groupi_n_1426, csa_tree_add_190_195_groupi_n_1427, csa_tree_add_190_195_groupi_n_1428, csa_tree_add_190_195_groupi_n_1429, csa_tree_add_190_195_groupi_n_1430;
  wire csa_tree_add_190_195_groupi_n_1431, csa_tree_add_190_195_groupi_n_1432, csa_tree_add_190_195_groupi_n_1433, csa_tree_add_190_195_groupi_n_1434, csa_tree_add_190_195_groupi_n_1435, csa_tree_add_190_195_groupi_n_1436, csa_tree_add_190_195_groupi_n_1437, csa_tree_add_190_195_groupi_n_1438;
  wire csa_tree_add_190_195_groupi_n_1439, csa_tree_add_190_195_groupi_n_1440, csa_tree_add_190_195_groupi_n_1441, csa_tree_add_190_195_groupi_n_1442, csa_tree_add_190_195_groupi_n_1443, csa_tree_add_190_195_groupi_n_1444, csa_tree_add_190_195_groupi_n_1445, csa_tree_add_190_195_groupi_n_1446;
  wire csa_tree_add_190_195_groupi_n_1447, csa_tree_add_190_195_groupi_n_1448, csa_tree_add_190_195_groupi_n_1449, csa_tree_add_190_195_groupi_n_1450, csa_tree_add_190_195_groupi_n_1451, csa_tree_add_190_195_groupi_n_1452, csa_tree_add_190_195_groupi_n_1453, csa_tree_add_190_195_groupi_n_1454;
  wire csa_tree_add_190_195_groupi_n_1455, csa_tree_add_190_195_groupi_n_1456, csa_tree_add_190_195_groupi_n_1457, csa_tree_add_190_195_groupi_n_1458, csa_tree_add_190_195_groupi_n_1459, csa_tree_add_190_195_groupi_n_1460, csa_tree_add_190_195_groupi_n_1461, csa_tree_add_190_195_groupi_n_1462;
  wire csa_tree_add_190_195_groupi_n_1463, csa_tree_add_190_195_groupi_n_1464, csa_tree_add_190_195_groupi_n_1465, csa_tree_add_190_195_groupi_n_1466, csa_tree_add_190_195_groupi_n_1467, csa_tree_add_190_195_groupi_n_1468, csa_tree_add_190_195_groupi_n_1469, csa_tree_add_190_195_groupi_n_1470;
  wire csa_tree_add_190_195_groupi_n_1471, csa_tree_add_190_195_groupi_n_1472, csa_tree_add_190_195_groupi_n_1473, csa_tree_add_190_195_groupi_n_1474, csa_tree_add_190_195_groupi_n_1475, csa_tree_add_190_195_groupi_n_1476, csa_tree_add_190_195_groupi_n_1477, csa_tree_add_190_195_groupi_n_1478;
  wire csa_tree_add_190_195_groupi_n_1479, csa_tree_add_190_195_groupi_n_1480, csa_tree_add_190_195_groupi_n_1481, csa_tree_add_190_195_groupi_n_1482, csa_tree_add_190_195_groupi_n_1483, csa_tree_add_190_195_groupi_n_1484, csa_tree_add_190_195_groupi_n_1485, csa_tree_add_190_195_groupi_n_1486;
  wire csa_tree_add_190_195_groupi_n_1487, csa_tree_add_190_195_groupi_n_1488, csa_tree_add_190_195_groupi_n_1489, csa_tree_add_190_195_groupi_n_1490, csa_tree_add_190_195_groupi_n_1491, csa_tree_add_190_195_groupi_n_1492, csa_tree_add_190_195_groupi_n_1493, csa_tree_add_190_195_groupi_n_1494;
  wire csa_tree_add_190_195_groupi_n_1495, csa_tree_add_190_195_groupi_n_1496, csa_tree_add_190_195_groupi_n_1497, csa_tree_add_190_195_groupi_n_1498, csa_tree_add_190_195_groupi_n_1499, csa_tree_add_190_195_groupi_n_1500, csa_tree_add_190_195_groupi_n_1501, csa_tree_add_190_195_groupi_n_1502;
  wire csa_tree_add_190_195_groupi_n_1503, csa_tree_add_190_195_groupi_n_1504, csa_tree_add_190_195_groupi_n_1505, csa_tree_add_190_195_groupi_n_1506, csa_tree_add_190_195_groupi_n_1507, csa_tree_add_190_195_groupi_n_1508, csa_tree_add_190_195_groupi_n_1509, csa_tree_add_190_195_groupi_n_1510;
  wire csa_tree_add_190_195_groupi_n_1511, csa_tree_add_190_195_groupi_n_1512, csa_tree_add_190_195_groupi_n_1513, csa_tree_add_190_195_groupi_n_1514, csa_tree_add_190_195_groupi_n_1515, csa_tree_add_190_195_groupi_n_1516, csa_tree_add_190_195_groupi_n_1517, csa_tree_add_190_195_groupi_n_1518;
  wire csa_tree_add_190_195_groupi_n_1519, csa_tree_add_190_195_groupi_n_1520, csa_tree_add_190_195_groupi_n_1521, csa_tree_add_190_195_groupi_n_1522, csa_tree_add_190_195_groupi_n_1523, csa_tree_add_190_195_groupi_n_1524, csa_tree_add_190_195_groupi_n_1525, csa_tree_add_190_195_groupi_n_1526;
  wire csa_tree_add_190_195_groupi_n_1527, csa_tree_add_190_195_groupi_n_1528, csa_tree_add_190_195_groupi_n_1529, csa_tree_add_190_195_groupi_n_1530, csa_tree_add_190_195_groupi_n_1531, csa_tree_add_190_195_groupi_n_1532, csa_tree_add_190_195_groupi_n_1533, csa_tree_add_190_195_groupi_n_1534;
  wire csa_tree_add_190_195_groupi_n_1535, csa_tree_add_190_195_groupi_n_1536, csa_tree_add_190_195_groupi_n_1537, csa_tree_add_190_195_groupi_n_1538, csa_tree_add_190_195_groupi_n_1539, csa_tree_add_190_195_groupi_n_1540, csa_tree_add_190_195_groupi_n_1541, csa_tree_add_190_195_groupi_n_1542;
  wire csa_tree_add_190_195_groupi_n_1543, csa_tree_add_190_195_groupi_n_1544, csa_tree_add_190_195_groupi_n_1545, csa_tree_add_190_195_groupi_n_1546, csa_tree_add_190_195_groupi_n_1547, csa_tree_add_190_195_groupi_n_1548, csa_tree_add_190_195_groupi_n_1549, csa_tree_add_190_195_groupi_n_1550;
  wire csa_tree_add_190_195_groupi_n_1551, csa_tree_add_190_195_groupi_n_1552, csa_tree_add_190_195_groupi_n_1553, csa_tree_add_190_195_groupi_n_1554, csa_tree_add_190_195_groupi_n_1555, csa_tree_add_190_195_groupi_n_1556, csa_tree_add_190_195_groupi_n_1557, csa_tree_add_190_195_groupi_n_1558;
  wire csa_tree_add_190_195_groupi_n_1559, csa_tree_add_190_195_groupi_n_1560, csa_tree_add_190_195_groupi_n_1561, csa_tree_add_190_195_groupi_n_1562, csa_tree_add_190_195_groupi_n_1563, csa_tree_add_190_195_groupi_n_1564, csa_tree_add_190_195_groupi_n_1565, csa_tree_add_190_195_groupi_n_1566;
  wire csa_tree_add_190_195_groupi_n_1567, csa_tree_add_190_195_groupi_n_1568, csa_tree_add_190_195_groupi_n_1569, csa_tree_add_190_195_groupi_n_1570, csa_tree_add_190_195_groupi_n_1571, csa_tree_add_190_195_groupi_n_1572, csa_tree_add_190_195_groupi_n_1573, csa_tree_add_190_195_groupi_n_1574;
  wire csa_tree_add_190_195_groupi_n_1575, csa_tree_add_190_195_groupi_n_1576, csa_tree_add_190_195_groupi_n_1577, csa_tree_add_190_195_groupi_n_1578, csa_tree_add_190_195_groupi_n_1579, csa_tree_add_190_195_groupi_n_1580, csa_tree_add_190_195_groupi_n_1581, csa_tree_add_190_195_groupi_n_1582;
  wire csa_tree_add_190_195_groupi_n_1583, csa_tree_add_190_195_groupi_n_1584, csa_tree_add_190_195_groupi_n_1585, csa_tree_add_190_195_groupi_n_1586, csa_tree_add_190_195_groupi_n_1587, csa_tree_add_190_195_groupi_n_1588, csa_tree_add_190_195_groupi_n_1589, csa_tree_add_190_195_groupi_n_1590;
  wire csa_tree_add_190_195_groupi_n_1591, csa_tree_add_190_195_groupi_n_1592, csa_tree_add_190_195_groupi_n_1593, csa_tree_add_190_195_groupi_n_1594, csa_tree_add_190_195_groupi_n_1595, csa_tree_add_190_195_groupi_n_1596, csa_tree_add_190_195_groupi_n_1597, csa_tree_add_190_195_groupi_n_1598;
  wire csa_tree_add_190_195_groupi_n_1599, csa_tree_add_190_195_groupi_n_1600, csa_tree_add_190_195_groupi_n_1601, csa_tree_add_190_195_groupi_n_1602, csa_tree_add_190_195_groupi_n_1603, csa_tree_add_190_195_groupi_n_1604, csa_tree_add_190_195_groupi_n_1605, csa_tree_add_190_195_groupi_n_1606;
  wire csa_tree_add_190_195_groupi_n_1607, csa_tree_add_190_195_groupi_n_1608, csa_tree_add_190_195_groupi_n_1609, csa_tree_add_190_195_groupi_n_1610, csa_tree_add_190_195_groupi_n_1611, csa_tree_add_190_195_groupi_n_1612, csa_tree_add_190_195_groupi_n_1613, csa_tree_add_190_195_groupi_n_1614;
  wire csa_tree_add_190_195_groupi_n_1615, csa_tree_add_190_195_groupi_n_1616, csa_tree_add_190_195_groupi_n_1617, csa_tree_add_190_195_groupi_n_1618, csa_tree_add_190_195_groupi_n_1619, csa_tree_add_190_195_groupi_n_1620, csa_tree_add_190_195_groupi_n_1621, csa_tree_add_190_195_groupi_n_1622;
  wire csa_tree_add_190_195_groupi_n_1623, csa_tree_add_190_195_groupi_n_1624, csa_tree_add_190_195_groupi_n_1625, csa_tree_add_190_195_groupi_n_1626, csa_tree_add_190_195_groupi_n_1627, csa_tree_add_190_195_groupi_n_1628, csa_tree_add_190_195_groupi_n_1629, csa_tree_add_190_195_groupi_n_1630;
  wire csa_tree_add_190_195_groupi_n_1631, csa_tree_add_190_195_groupi_n_1632, csa_tree_add_190_195_groupi_n_1633, csa_tree_add_190_195_groupi_n_1634, csa_tree_add_190_195_groupi_n_1635, csa_tree_add_190_195_groupi_n_1636, csa_tree_add_190_195_groupi_n_1637, csa_tree_add_190_195_groupi_n_1638;
  wire csa_tree_add_190_195_groupi_n_1639, csa_tree_add_190_195_groupi_n_1640, csa_tree_add_190_195_groupi_n_1641, csa_tree_add_190_195_groupi_n_1642, csa_tree_add_190_195_groupi_n_1643, csa_tree_add_190_195_groupi_n_1644, csa_tree_add_190_195_groupi_n_1645, csa_tree_add_190_195_groupi_n_1646;
  wire csa_tree_add_190_195_groupi_n_1647, csa_tree_add_190_195_groupi_n_1648, csa_tree_add_190_195_groupi_n_1649, csa_tree_add_190_195_groupi_n_1650, csa_tree_add_190_195_groupi_n_1651, csa_tree_add_190_195_groupi_n_1652, csa_tree_add_190_195_groupi_n_1653, csa_tree_add_190_195_groupi_n_1654;
  wire csa_tree_add_190_195_groupi_n_1655, csa_tree_add_190_195_groupi_n_1656, csa_tree_add_190_195_groupi_n_1657, csa_tree_add_190_195_groupi_n_1658, csa_tree_add_190_195_groupi_n_1659, csa_tree_add_190_195_groupi_n_1660, csa_tree_add_190_195_groupi_n_1661, csa_tree_add_190_195_groupi_n_1662;
  wire csa_tree_add_190_195_groupi_n_1663, csa_tree_add_190_195_groupi_n_1664, csa_tree_add_190_195_groupi_n_1665, csa_tree_add_190_195_groupi_n_1666, csa_tree_add_190_195_groupi_n_1667, csa_tree_add_190_195_groupi_n_1668, csa_tree_add_190_195_groupi_n_1669, csa_tree_add_190_195_groupi_n_1670;
  wire csa_tree_add_190_195_groupi_n_1671, csa_tree_add_190_195_groupi_n_1672, csa_tree_add_190_195_groupi_n_1673, csa_tree_add_190_195_groupi_n_1674, csa_tree_add_190_195_groupi_n_1675, csa_tree_add_190_195_groupi_n_1676, csa_tree_add_190_195_groupi_n_1677, csa_tree_add_190_195_groupi_n_1678;
  wire csa_tree_add_190_195_groupi_n_1679, csa_tree_add_190_195_groupi_n_1680, csa_tree_add_190_195_groupi_n_1681, csa_tree_add_190_195_groupi_n_1682, csa_tree_add_190_195_groupi_n_1683, csa_tree_add_190_195_groupi_n_1684, csa_tree_add_190_195_groupi_n_1685, csa_tree_add_190_195_groupi_n_1686;
  wire csa_tree_add_190_195_groupi_n_1687, csa_tree_add_190_195_groupi_n_1688, csa_tree_add_190_195_groupi_n_1689, csa_tree_add_190_195_groupi_n_1690, csa_tree_add_190_195_groupi_n_1691, csa_tree_add_190_195_groupi_n_1692, csa_tree_add_190_195_groupi_n_1693, csa_tree_add_190_195_groupi_n_1694;
  wire csa_tree_add_190_195_groupi_n_1695, csa_tree_add_190_195_groupi_n_1696, csa_tree_add_190_195_groupi_n_1697, csa_tree_add_190_195_groupi_n_1698, csa_tree_add_190_195_groupi_n_1699, csa_tree_add_190_195_groupi_n_1700, csa_tree_add_190_195_groupi_n_1701, csa_tree_add_190_195_groupi_n_1702;
  wire csa_tree_add_190_195_groupi_n_1703, csa_tree_add_190_195_groupi_n_1704, csa_tree_add_190_195_groupi_n_1705, csa_tree_add_190_195_groupi_n_1706, csa_tree_add_190_195_groupi_n_1707, csa_tree_add_190_195_groupi_n_1708, csa_tree_add_190_195_groupi_n_1709, csa_tree_add_190_195_groupi_n_1710;
  wire csa_tree_add_190_195_groupi_n_1711, csa_tree_add_190_195_groupi_n_1712, csa_tree_add_190_195_groupi_n_1713, csa_tree_add_190_195_groupi_n_1714, csa_tree_add_190_195_groupi_n_1715, csa_tree_add_190_195_groupi_n_1716, csa_tree_add_190_195_groupi_n_1717, csa_tree_add_190_195_groupi_n_1718;
  wire csa_tree_add_190_195_groupi_n_1719, csa_tree_add_190_195_groupi_n_1720, csa_tree_add_190_195_groupi_n_1721, csa_tree_add_190_195_groupi_n_1722, csa_tree_add_190_195_groupi_n_1723, csa_tree_add_190_195_groupi_n_1724, csa_tree_add_190_195_groupi_n_1725, csa_tree_add_190_195_groupi_n_1726;
  wire csa_tree_add_190_195_groupi_n_1727, csa_tree_add_190_195_groupi_n_1728, csa_tree_add_190_195_groupi_n_1729, csa_tree_add_190_195_groupi_n_1730, csa_tree_add_190_195_groupi_n_1731, csa_tree_add_190_195_groupi_n_1732, csa_tree_add_190_195_groupi_n_1733, csa_tree_add_190_195_groupi_n_1734;
  wire csa_tree_add_190_195_groupi_n_1735, csa_tree_add_190_195_groupi_n_1736, csa_tree_add_190_195_groupi_n_1737, csa_tree_add_190_195_groupi_n_1738, csa_tree_add_190_195_groupi_n_1739, csa_tree_add_190_195_groupi_n_1740, csa_tree_add_190_195_groupi_n_1741, csa_tree_add_190_195_groupi_n_1742;
  wire csa_tree_add_190_195_groupi_n_1743, csa_tree_add_190_195_groupi_n_1744, csa_tree_add_190_195_groupi_n_1745, csa_tree_add_190_195_groupi_n_1746, csa_tree_add_190_195_groupi_n_1747, csa_tree_add_190_195_groupi_n_1748, csa_tree_add_190_195_groupi_n_1749, csa_tree_add_190_195_groupi_n_1750;
  wire csa_tree_add_190_195_groupi_n_1751, csa_tree_add_190_195_groupi_n_1752, csa_tree_add_190_195_groupi_n_1753, csa_tree_add_190_195_groupi_n_1754, csa_tree_add_190_195_groupi_n_1755, csa_tree_add_190_195_groupi_n_1756, csa_tree_add_190_195_groupi_n_1757, csa_tree_add_190_195_groupi_n_1758;
  wire csa_tree_add_190_195_groupi_n_1759, csa_tree_add_190_195_groupi_n_1760, csa_tree_add_190_195_groupi_n_1761, csa_tree_add_190_195_groupi_n_1762, csa_tree_add_190_195_groupi_n_1763, csa_tree_add_190_195_groupi_n_1764, csa_tree_add_190_195_groupi_n_1765, csa_tree_add_190_195_groupi_n_1766;
  wire csa_tree_add_190_195_groupi_n_1767, csa_tree_add_190_195_groupi_n_1768, csa_tree_add_190_195_groupi_n_1769, csa_tree_add_190_195_groupi_n_1770, csa_tree_add_190_195_groupi_n_1771, csa_tree_add_190_195_groupi_n_1772, csa_tree_add_190_195_groupi_n_1773, csa_tree_add_190_195_groupi_n_1774;
  wire csa_tree_add_190_195_groupi_n_1775, csa_tree_add_190_195_groupi_n_1776, csa_tree_add_190_195_groupi_n_1777, csa_tree_add_190_195_groupi_n_1778, csa_tree_add_190_195_groupi_n_1779, csa_tree_add_190_195_groupi_n_1780, csa_tree_add_190_195_groupi_n_1781, csa_tree_add_190_195_groupi_n_1782;
  wire csa_tree_add_190_195_groupi_n_1783, csa_tree_add_190_195_groupi_n_1784, csa_tree_add_190_195_groupi_n_1785, csa_tree_add_190_195_groupi_n_1786, csa_tree_add_190_195_groupi_n_1787, csa_tree_add_190_195_groupi_n_1788, csa_tree_add_190_195_groupi_n_1789, csa_tree_add_190_195_groupi_n_1790;
  wire csa_tree_add_190_195_groupi_n_1791, csa_tree_add_190_195_groupi_n_1792, csa_tree_add_190_195_groupi_n_1793, csa_tree_add_190_195_groupi_n_1794, csa_tree_add_190_195_groupi_n_1795, csa_tree_add_190_195_groupi_n_1796, csa_tree_add_190_195_groupi_n_1797, csa_tree_add_190_195_groupi_n_1798;
  wire csa_tree_add_190_195_groupi_n_1799, csa_tree_add_190_195_groupi_n_1800, csa_tree_add_190_195_groupi_n_1801, csa_tree_add_190_195_groupi_n_1802, csa_tree_add_190_195_groupi_n_1803, csa_tree_add_190_195_groupi_n_1804, csa_tree_add_190_195_groupi_n_1805, csa_tree_add_190_195_groupi_n_1806;
  wire csa_tree_add_190_195_groupi_n_1807, csa_tree_add_190_195_groupi_n_1808, csa_tree_add_190_195_groupi_n_1809, csa_tree_add_190_195_groupi_n_1810, csa_tree_add_190_195_groupi_n_1811, csa_tree_add_190_195_groupi_n_1812, csa_tree_add_190_195_groupi_n_1813, csa_tree_add_190_195_groupi_n_1814;
  wire csa_tree_add_190_195_groupi_n_1815, csa_tree_add_190_195_groupi_n_1816, csa_tree_add_190_195_groupi_n_1817, csa_tree_add_190_195_groupi_n_1818, csa_tree_add_190_195_groupi_n_1819, csa_tree_add_190_195_groupi_n_1820, csa_tree_add_190_195_groupi_n_1821, csa_tree_add_190_195_groupi_n_1822;
  wire csa_tree_add_190_195_groupi_n_1823, csa_tree_add_190_195_groupi_n_1824, csa_tree_add_190_195_groupi_n_1825, csa_tree_add_190_195_groupi_n_1826, csa_tree_add_190_195_groupi_n_1827, csa_tree_add_190_195_groupi_n_1828, csa_tree_add_190_195_groupi_n_1829, csa_tree_add_190_195_groupi_n_1830;
  wire csa_tree_add_190_195_groupi_n_1831, csa_tree_add_190_195_groupi_n_1832, csa_tree_add_190_195_groupi_n_1833, csa_tree_add_190_195_groupi_n_1834, csa_tree_add_190_195_groupi_n_1835, csa_tree_add_190_195_groupi_n_1836, csa_tree_add_190_195_groupi_n_1837, csa_tree_add_190_195_groupi_n_1838;
  wire csa_tree_add_190_195_groupi_n_1839, csa_tree_add_190_195_groupi_n_1840, csa_tree_add_190_195_groupi_n_1841, csa_tree_add_190_195_groupi_n_1842, csa_tree_add_190_195_groupi_n_1843, csa_tree_add_190_195_groupi_n_1844, csa_tree_add_190_195_groupi_n_1845, csa_tree_add_190_195_groupi_n_1846;
  wire csa_tree_add_190_195_groupi_n_1847, csa_tree_add_190_195_groupi_n_1848, csa_tree_add_190_195_groupi_n_1849, csa_tree_add_190_195_groupi_n_1850, csa_tree_add_190_195_groupi_n_1851, csa_tree_add_190_195_groupi_n_1852, csa_tree_add_190_195_groupi_n_1853, csa_tree_add_190_195_groupi_n_1854;
  wire csa_tree_add_190_195_groupi_n_1855, csa_tree_add_190_195_groupi_n_1856, csa_tree_add_190_195_groupi_n_1857, csa_tree_add_190_195_groupi_n_1858, csa_tree_add_190_195_groupi_n_1859, csa_tree_add_190_195_groupi_n_1860, csa_tree_add_190_195_groupi_n_1861, csa_tree_add_190_195_groupi_n_1862;
  wire csa_tree_add_190_195_groupi_n_1863, csa_tree_add_190_195_groupi_n_1864, csa_tree_add_190_195_groupi_n_1865, csa_tree_add_190_195_groupi_n_1866, csa_tree_add_190_195_groupi_n_1867, csa_tree_add_190_195_groupi_n_1868, csa_tree_add_190_195_groupi_n_1869, csa_tree_add_190_195_groupi_n_1870;
  wire csa_tree_add_190_195_groupi_n_1871, csa_tree_add_190_195_groupi_n_1872, csa_tree_add_190_195_groupi_n_1873, csa_tree_add_190_195_groupi_n_1874, csa_tree_add_190_195_groupi_n_1875, csa_tree_add_190_195_groupi_n_1876, csa_tree_add_190_195_groupi_n_1877, csa_tree_add_190_195_groupi_n_1878;
  wire csa_tree_add_190_195_groupi_n_1879, csa_tree_add_190_195_groupi_n_1880, csa_tree_add_190_195_groupi_n_1881, csa_tree_add_190_195_groupi_n_1882, csa_tree_add_190_195_groupi_n_1883, csa_tree_add_190_195_groupi_n_1884, csa_tree_add_190_195_groupi_n_1885, csa_tree_add_190_195_groupi_n_1886;
  wire csa_tree_add_190_195_groupi_n_1887, csa_tree_add_190_195_groupi_n_1888, csa_tree_add_190_195_groupi_n_1889, csa_tree_add_190_195_groupi_n_1890, csa_tree_add_190_195_groupi_n_1891, csa_tree_add_190_195_groupi_n_1892, csa_tree_add_190_195_groupi_n_1893, csa_tree_add_190_195_groupi_n_1894;
  wire csa_tree_add_190_195_groupi_n_1895, csa_tree_add_190_195_groupi_n_1896, csa_tree_add_190_195_groupi_n_1897, csa_tree_add_190_195_groupi_n_1898, csa_tree_add_190_195_groupi_n_1899, csa_tree_add_190_195_groupi_n_1900, csa_tree_add_190_195_groupi_n_1901, csa_tree_add_190_195_groupi_n_1902;
  wire csa_tree_add_190_195_groupi_n_1903, csa_tree_add_190_195_groupi_n_1904, csa_tree_add_190_195_groupi_n_1905, csa_tree_add_190_195_groupi_n_1906, csa_tree_add_190_195_groupi_n_1907, csa_tree_add_190_195_groupi_n_1908, csa_tree_add_190_195_groupi_n_1909, csa_tree_add_190_195_groupi_n_1910;
  wire csa_tree_add_190_195_groupi_n_1911, csa_tree_add_190_195_groupi_n_1912, csa_tree_add_190_195_groupi_n_1913, csa_tree_add_190_195_groupi_n_1914, csa_tree_add_190_195_groupi_n_1915, csa_tree_add_190_195_groupi_n_1916, csa_tree_add_190_195_groupi_n_1917, csa_tree_add_190_195_groupi_n_1918;
  wire csa_tree_add_190_195_groupi_n_1919, csa_tree_add_190_195_groupi_n_1920, csa_tree_add_190_195_groupi_n_1921, csa_tree_add_190_195_groupi_n_1922, csa_tree_add_190_195_groupi_n_1923, csa_tree_add_190_195_groupi_n_1924, csa_tree_add_190_195_groupi_n_1925, csa_tree_add_190_195_groupi_n_1926;
  wire csa_tree_add_190_195_groupi_n_1927, csa_tree_add_190_195_groupi_n_1928, csa_tree_add_190_195_groupi_n_1929, csa_tree_add_190_195_groupi_n_1930, csa_tree_add_190_195_groupi_n_1931, csa_tree_add_190_195_groupi_n_1932, csa_tree_add_190_195_groupi_n_1933, csa_tree_add_190_195_groupi_n_1934;
  wire csa_tree_add_190_195_groupi_n_1935, csa_tree_add_190_195_groupi_n_1936, csa_tree_add_190_195_groupi_n_1937, csa_tree_add_190_195_groupi_n_1938, csa_tree_add_190_195_groupi_n_1939, csa_tree_add_190_195_groupi_n_1940, csa_tree_add_190_195_groupi_n_1941, csa_tree_add_190_195_groupi_n_1942;
  wire csa_tree_add_190_195_groupi_n_1943, csa_tree_add_190_195_groupi_n_1944, csa_tree_add_190_195_groupi_n_1945, csa_tree_add_190_195_groupi_n_1946, csa_tree_add_190_195_groupi_n_1947, csa_tree_add_190_195_groupi_n_1948, csa_tree_add_190_195_groupi_n_1949, csa_tree_add_190_195_groupi_n_1950;
  wire csa_tree_add_190_195_groupi_n_1951, csa_tree_add_190_195_groupi_n_1952, csa_tree_add_190_195_groupi_n_1953, csa_tree_add_190_195_groupi_n_1954, csa_tree_add_190_195_groupi_n_1955, csa_tree_add_190_195_groupi_n_1956, csa_tree_add_190_195_groupi_n_1957, csa_tree_add_190_195_groupi_n_1958;
  wire csa_tree_add_190_195_groupi_n_1959, csa_tree_add_190_195_groupi_n_1960, csa_tree_add_190_195_groupi_n_1961, csa_tree_add_190_195_groupi_n_1962, csa_tree_add_190_195_groupi_n_1963, csa_tree_add_190_195_groupi_n_1964, csa_tree_add_190_195_groupi_n_1965, csa_tree_add_190_195_groupi_n_1966;
  wire csa_tree_add_190_195_groupi_n_1967, csa_tree_add_190_195_groupi_n_1968, csa_tree_add_190_195_groupi_n_1969, csa_tree_add_190_195_groupi_n_1970, csa_tree_add_190_195_groupi_n_1971, csa_tree_add_190_195_groupi_n_1972, csa_tree_add_190_195_groupi_n_1973, csa_tree_add_190_195_groupi_n_1974;
  wire csa_tree_add_190_195_groupi_n_1975, csa_tree_add_190_195_groupi_n_1976, csa_tree_add_190_195_groupi_n_1977, csa_tree_add_190_195_groupi_n_1978, csa_tree_add_190_195_groupi_n_1979, csa_tree_add_190_195_groupi_n_1980, csa_tree_add_190_195_groupi_n_1981, csa_tree_add_190_195_groupi_n_1982;
  wire csa_tree_add_190_195_groupi_n_1983, csa_tree_add_190_195_groupi_n_1984, csa_tree_add_190_195_groupi_n_1985, csa_tree_add_190_195_groupi_n_1986, csa_tree_add_190_195_groupi_n_1987, csa_tree_add_190_195_groupi_n_1988, csa_tree_add_190_195_groupi_n_1989, csa_tree_add_190_195_groupi_n_1990;
  wire csa_tree_add_190_195_groupi_n_1991, csa_tree_add_190_195_groupi_n_1992, csa_tree_add_190_195_groupi_n_1993, csa_tree_add_190_195_groupi_n_1994, csa_tree_add_190_195_groupi_n_1995, csa_tree_add_190_195_groupi_n_1996, csa_tree_add_190_195_groupi_n_1997, csa_tree_add_190_195_groupi_n_1998;
  wire csa_tree_add_190_195_groupi_n_1999, csa_tree_add_190_195_groupi_n_2000, csa_tree_add_190_195_groupi_n_2001, csa_tree_add_190_195_groupi_n_2002, csa_tree_add_190_195_groupi_n_2003, csa_tree_add_190_195_groupi_n_2004, csa_tree_add_190_195_groupi_n_2005, csa_tree_add_190_195_groupi_n_2006;
  wire csa_tree_add_190_195_groupi_n_2007, csa_tree_add_190_195_groupi_n_2008, csa_tree_add_190_195_groupi_n_2009, csa_tree_add_190_195_groupi_n_2010, csa_tree_add_190_195_groupi_n_2011, csa_tree_add_190_195_groupi_n_2012, csa_tree_add_190_195_groupi_n_2013, csa_tree_add_190_195_groupi_n_2014;
  wire csa_tree_add_190_195_groupi_n_2015, csa_tree_add_190_195_groupi_n_2016, csa_tree_add_190_195_groupi_n_2017, csa_tree_add_190_195_groupi_n_2018, csa_tree_add_190_195_groupi_n_2019, csa_tree_add_190_195_groupi_n_2020, csa_tree_add_190_195_groupi_n_2021, csa_tree_add_190_195_groupi_n_2022;
  wire csa_tree_add_190_195_groupi_n_2023, csa_tree_add_190_195_groupi_n_2024, csa_tree_add_190_195_groupi_n_2025, csa_tree_add_190_195_groupi_n_2026, csa_tree_add_190_195_groupi_n_2027, csa_tree_add_190_195_groupi_n_2028, csa_tree_add_190_195_groupi_n_2029, csa_tree_add_190_195_groupi_n_2030;
  wire csa_tree_add_190_195_groupi_n_2031, csa_tree_add_190_195_groupi_n_2032, csa_tree_add_190_195_groupi_n_2033, csa_tree_add_190_195_groupi_n_2034, csa_tree_add_190_195_groupi_n_2035, csa_tree_add_190_195_groupi_n_2036, csa_tree_add_190_195_groupi_n_2037, csa_tree_add_190_195_groupi_n_2038;
  wire csa_tree_add_190_195_groupi_n_2039, csa_tree_add_190_195_groupi_n_2040, csa_tree_add_190_195_groupi_n_2041, csa_tree_add_190_195_groupi_n_2042, csa_tree_add_190_195_groupi_n_2043, csa_tree_add_190_195_groupi_n_2044, csa_tree_add_190_195_groupi_n_2045, csa_tree_add_190_195_groupi_n_2046;
  wire csa_tree_add_190_195_groupi_n_2047, csa_tree_add_190_195_groupi_n_2048, csa_tree_add_190_195_groupi_n_2049, csa_tree_add_190_195_groupi_n_2050, csa_tree_add_190_195_groupi_n_2051, csa_tree_add_190_195_groupi_n_2052, csa_tree_add_190_195_groupi_n_2053, csa_tree_add_190_195_groupi_n_2054;
  wire csa_tree_add_190_195_groupi_n_2055, csa_tree_add_190_195_groupi_n_2056, csa_tree_add_190_195_groupi_n_2057, csa_tree_add_190_195_groupi_n_2058, csa_tree_add_190_195_groupi_n_2059, csa_tree_add_190_195_groupi_n_2060, csa_tree_add_190_195_groupi_n_2061, csa_tree_add_190_195_groupi_n_2062;
  wire csa_tree_add_190_195_groupi_n_2063, csa_tree_add_190_195_groupi_n_2064, csa_tree_add_190_195_groupi_n_2065, csa_tree_add_190_195_groupi_n_2066, csa_tree_add_190_195_groupi_n_2067, csa_tree_add_190_195_groupi_n_2068, csa_tree_add_190_195_groupi_n_2069, csa_tree_add_190_195_groupi_n_2070;
  wire csa_tree_add_190_195_groupi_n_2071, csa_tree_add_190_195_groupi_n_2072, csa_tree_add_190_195_groupi_n_2073, csa_tree_add_190_195_groupi_n_2074, csa_tree_add_190_195_groupi_n_2075, csa_tree_add_190_195_groupi_n_2076, csa_tree_add_190_195_groupi_n_2077, csa_tree_add_190_195_groupi_n_2078;
  wire csa_tree_add_190_195_groupi_n_2079, csa_tree_add_190_195_groupi_n_2080, csa_tree_add_190_195_groupi_n_2081, csa_tree_add_190_195_groupi_n_2082, csa_tree_add_190_195_groupi_n_2083, csa_tree_add_190_195_groupi_n_2084, csa_tree_add_190_195_groupi_n_2085, csa_tree_add_190_195_groupi_n_2086;
  wire csa_tree_add_190_195_groupi_n_2087, csa_tree_add_190_195_groupi_n_2088, csa_tree_add_190_195_groupi_n_2089, csa_tree_add_190_195_groupi_n_2090, csa_tree_add_190_195_groupi_n_2091, csa_tree_add_190_195_groupi_n_2092, csa_tree_add_190_195_groupi_n_2093, csa_tree_add_190_195_groupi_n_2094;
  wire csa_tree_add_190_195_groupi_n_2095, csa_tree_add_190_195_groupi_n_2096, csa_tree_add_190_195_groupi_n_2097, csa_tree_add_190_195_groupi_n_2098, csa_tree_add_190_195_groupi_n_2099, csa_tree_add_190_195_groupi_n_2100, csa_tree_add_190_195_groupi_n_2101, csa_tree_add_190_195_groupi_n_2102;
  wire csa_tree_add_190_195_groupi_n_2103, csa_tree_add_190_195_groupi_n_2104, csa_tree_add_190_195_groupi_n_2105, csa_tree_add_190_195_groupi_n_2106, csa_tree_add_190_195_groupi_n_2107, csa_tree_add_190_195_groupi_n_2108, csa_tree_add_190_195_groupi_n_2109, csa_tree_add_190_195_groupi_n_2110;
  wire csa_tree_add_190_195_groupi_n_2111, csa_tree_add_190_195_groupi_n_2112, csa_tree_add_190_195_groupi_n_2113, csa_tree_add_190_195_groupi_n_2114, csa_tree_add_190_195_groupi_n_2115, csa_tree_add_190_195_groupi_n_2116, csa_tree_add_190_195_groupi_n_2117, csa_tree_add_190_195_groupi_n_2118;
  wire csa_tree_add_190_195_groupi_n_2119, csa_tree_add_190_195_groupi_n_2120, csa_tree_add_190_195_groupi_n_2121, csa_tree_add_190_195_groupi_n_2122, csa_tree_add_190_195_groupi_n_2123, csa_tree_add_190_195_groupi_n_2124, csa_tree_add_190_195_groupi_n_2125, csa_tree_add_190_195_groupi_n_2126;
  wire csa_tree_add_190_195_groupi_n_2127, csa_tree_add_190_195_groupi_n_2128, csa_tree_add_190_195_groupi_n_2129, csa_tree_add_190_195_groupi_n_2130, csa_tree_add_190_195_groupi_n_2131, csa_tree_add_190_195_groupi_n_2132, csa_tree_add_190_195_groupi_n_2133, csa_tree_add_190_195_groupi_n_2134;
  wire csa_tree_add_190_195_groupi_n_2135, csa_tree_add_190_195_groupi_n_2136, csa_tree_add_190_195_groupi_n_2137, csa_tree_add_190_195_groupi_n_2138, csa_tree_add_190_195_groupi_n_2139, csa_tree_add_190_195_groupi_n_2140, csa_tree_add_190_195_groupi_n_2141, csa_tree_add_190_195_groupi_n_2142;
  wire csa_tree_add_190_195_groupi_n_2143, csa_tree_add_190_195_groupi_n_2144, csa_tree_add_190_195_groupi_n_2145, csa_tree_add_190_195_groupi_n_2146, csa_tree_add_190_195_groupi_n_2147, csa_tree_add_190_195_groupi_n_2148, csa_tree_add_190_195_groupi_n_2149, csa_tree_add_190_195_groupi_n_2150;
  wire csa_tree_add_190_195_groupi_n_2151, csa_tree_add_190_195_groupi_n_2152, csa_tree_add_190_195_groupi_n_2153, csa_tree_add_190_195_groupi_n_2154, csa_tree_add_190_195_groupi_n_2155, csa_tree_add_190_195_groupi_n_2156, csa_tree_add_190_195_groupi_n_2157, csa_tree_add_190_195_groupi_n_2158;
  wire csa_tree_add_190_195_groupi_n_2159, csa_tree_add_190_195_groupi_n_2160, csa_tree_add_190_195_groupi_n_2161, csa_tree_add_190_195_groupi_n_2162, csa_tree_add_190_195_groupi_n_2163, csa_tree_add_190_195_groupi_n_2164, csa_tree_add_190_195_groupi_n_2165, csa_tree_add_190_195_groupi_n_2166;
  wire csa_tree_add_190_195_groupi_n_2167, csa_tree_add_190_195_groupi_n_2168, csa_tree_add_190_195_groupi_n_2169, csa_tree_add_190_195_groupi_n_2170, csa_tree_add_190_195_groupi_n_2171, csa_tree_add_190_195_groupi_n_2172, csa_tree_add_190_195_groupi_n_2173, csa_tree_add_190_195_groupi_n_2174;
  wire csa_tree_add_190_195_groupi_n_2175, csa_tree_add_190_195_groupi_n_2176, csa_tree_add_190_195_groupi_n_2177, csa_tree_add_190_195_groupi_n_2178, csa_tree_add_190_195_groupi_n_2179, csa_tree_add_190_195_groupi_n_2180, csa_tree_add_190_195_groupi_n_2181, csa_tree_add_190_195_groupi_n_2182;
  wire csa_tree_add_190_195_groupi_n_2183, csa_tree_add_190_195_groupi_n_2184, csa_tree_add_190_195_groupi_n_2185, csa_tree_add_190_195_groupi_n_2186, csa_tree_add_190_195_groupi_n_2187, csa_tree_add_190_195_groupi_n_2188, csa_tree_add_190_195_groupi_n_2189, csa_tree_add_190_195_groupi_n_2190;
  wire csa_tree_add_190_195_groupi_n_2191, csa_tree_add_190_195_groupi_n_2192, csa_tree_add_190_195_groupi_n_2193, csa_tree_add_190_195_groupi_n_2194, csa_tree_add_190_195_groupi_n_2195, csa_tree_add_190_195_groupi_n_2196, csa_tree_add_190_195_groupi_n_2197, csa_tree_add_190_195_groupi_n_2198;
  wire csa_tree_add_190_195_groupi_n_2199, csa_tree_add_190_195_groupi_n_2200, csa_tree_add_190_195_groupi_n_2201, csa_tree_add_190_195_groupi_n_2202, csa_tree_add_190_195_groupi_n_2203, csa_tree_add_190_195_groupi_n_2204, csa_tree_add_190_195_groupi_n_2205, csa_tree_add_190_195_groupi_n_2206;
  wire csa_tree_add_190_195_groupi_n_2207, csa_tree_add_190_195_groupi_n_2208, csa_tree_add_190_195_groupi_n_2209, csa_tree_add_190_195_groupi_n_2210, csa_tree_add_190_195_groupi_n_2211, csa_tree_add_190_195_groupi_n_2212, csa_tree_add_190_195_groupi_n_2213, csa_tree_add_190_195_groupi_n_2214;
  wire csa_tree_add_190_195_groupi_n_2215, csa_tree_add_190_195_groupi_n_2216, csa_tree_add_190_195_groupi_n_2217, csa_tree_add_190_195_groupi_n_2218, csa_tree_add_190_195_groupi_n_2219, csa_tree_add_190_195_groupi_n_2220, csa_tree_add_190_195_groupi_n_2221, csa_tree_add_190_195_groupi_n_2222;
  wire csa_tree_add_190_195_groupi_n_2223, csa_tree_add_190_195_groupi_n_2224, csa_tree_add_190_195_groupi_n_2225, csa_tree_add_190_195_groupi_n_2226, csa_tree_add_190_195_groupi_n_2227, csa_tree_add_190_195_groupi_n_2228, csa_tree_add_190_195_groupi_n_2229, csa_tree_add_190_195_groupi_n_2230;
  wire csa_tree_add_190_195_groupi_n_2231, csa_tree_add_190_195_groupi_n_2232, csa_tree_add_190_195_groupi_n_2233, csa_tree_add_190_195_groupi_n_2234, csa_tree_add_190_195_groupi_n_2235, csa_tree_add_190_195_groupi_n_2236, csa_tree_add_190_195_groupi_n_2237, csa_tree_add_190_195_groupi_n_2238;
  wire csa_tree_add_190_195_groupi_n_2239, csa_tree_add_190_195_groupi_n_2240, csa_tree_add_190_195_groupi_n_2241, csa_tree_add_190_195_groupi_n_2242, csa_tree_add_190_195_groupi_n_2243, csa_tree_add_190_195_groupi_n_2244, csa_tree_add_190_195_groupi_n_2245, csa_tree_add_190_195_groupi_n_2246;
  wire csa_tree_add_190_195_groupi_n_2247, csa_tree_add_190_195_groupi_n_2248, csa_tree_add_190_195_groupi_n_2249, csa_tree_add_190_195_groupi_n_2250, csa_tree_add_190_195_groupi_n_2251, csa_tree_add_190_195_groupi_n_2252, csa_tree_add_190_195_groupi_n_2253, csa_tree_add_190_195_groupi_n_2254;
  wire csa_tree_add_190_195_groupi_n_2255, csa_tree_add_190_195_groupi_n_2256, csa_tree_add_190_195_groupi_n_2257, csa_tree_add_190_195_groupi_n_2258, csa_tree_add_190_195_groupi_n_2259, csa_tree_add_190_195_groupi_n_2260, csa_tree_add_190_195_groupi_n_2261, csa_tree_add_190_195_groupi_n_2262;
  wire csa_tree_add_190_195_groupi_n_2263, csa_tree_add_190_195_groupi_n_2264, csa_tree_add_190_195_groupi_n_2265, csa_tree_add_190_195_groupi_n_2266, csa_tree_add_190_195_groupi_n_2267, csa_tree_add_190_195_groupi_n_2268, csa_tree_add_190_195_groupi_n_2269, csa_tree_add_190_195_groupi_n_2270;
  wire csa_tree_add_190_195_groupi_n_2271, csa_tree_add_190_195_groupi_n_2272, csa_tree_add_190_195_groupi_n_2273, csa_tree_add_190_195_groupi_n_2274, csa_tree_add_190_195_groupi_n_2275, csa_tree_add_190_195_groupi_n_2276, csa_tree_add_190_195_groupi_n_2277, csa_tree_add_190_195_groupi_n_2278;
  wire csa_tree_add_190_195_groupi_n_2279, csa_tree_add_190_195_groupi_n_2280, csa_tree_add_190_195_groupi_n_2281, csa_tree_add_190_195_groupi_n_2282, csa_tree_add_190_195_groupi_n_2283, csa_tree_add_190_195_groupi_n_2284, csa_tree_add_190_195_groupi_n_2285, csa_tree_add_190_195_groupi_n_2286;
  wire csa_tree_add_190_195_groupi_n_2287, csa_tree_add_190_195_groupi_n_2288, csa_tree_add_190_195_groupi_n_2289, csa_tree_add_190_195_groupi_n_2290, csa_tree_add_190_195_groupi_n_2291, csa_tree_add_190_195_groupi_n_2292, csa_tree_add_190_195_groupi_n_2293, csa_tree_add_190_195_groupi_n_2294;
  wire csa_tree_add_190_195_groupi_n_2295, csa_tree_add_190_195_groupi_n_2296, csa_tree_add_190_195_groupi_n_2297, csa_tree_add_190_195_groupi_n_2298, csa_tree_add_190_195_groupi_n_2299, csa_tree_add_190_195_groupi_n_2300, csa_tree_add_190_195_groupi_n_2301, csa_tree_add_190_195_groupi_n_2302;
  wire csa_tree_add_190_195_groupi_n_2303, csa_tree_add_190_195_groupi_n_2304, csa_tree_add_190_195_groupi_n_2305, csa_tree_add_190_195_groupi_n_2306, csa_tree_add_190_195_groupi_n_2307, csa_tree_add_190_195_groupi_n_2308, csa_tree_add_190_195_groupi_n_2309, csa_tree_add_190_195_groupi_n_2310;
  wire csa_tree_add_190_195_groupi_n_2311, csa_tree_add_190_195_groupi_n_2312, csa_tree_add_190_195_groupi_n_2313, csa_tree_add_190_195_groupi_n_2314, csa_tree_add_190_195_groupi_n_2315, csa_tree_add_190_195_groupi_n_2316, csa_tree_add_190_195_groupi_n_2317, csa_tree_add_190_195_groupi_n_2318;
  wire csa_tree_add_190_195_groupi_n_2319, csa_tree_add_190_195_groupi_n_2320, csa_tree_add_190_195_groupi_n_2321, csa_tree_add_190_195_groupi_n_2322, csa_tree_add_190_195_groupi_n_2323, csa_tree_add_190_195_groupi_n_2324, csa_tree_add_190_195_groupi_n_2325, csa_tree_add_190_195_groupi_n_2326;
  wire csa_tree_add_190_195_groupi_n_2327, csa_tree_add_190_195_groupi_n_2328, csa_tree_add_190_195_groupi_n_2329, csa_tree_add_190_195_groupi_n_2330, csa_tree_add_190_195_groupi_n_2331, csa_tree_add_190_195_groupi_n_2332, csa_tree_add_190_195_groupi_n_2333, csa_tree_add_190_195_groupi_n_2334;
  wire csa_tree_add_190_195_groupi_n_2335, csa_tree_add_190_195_groupi_n_2336, csa_tree_add_190_195_groupi_n_2337, csa_tree_add_190_195_groupi_n_2338, csa_tree_add_190_195_groupi_n_2339, csa_tree_add_190_195_groupi_n_2340, csa_tree_add_190_195_groupi_n_2341, csa_tree_add_190_195_groupi_n_2342;
  wire csa_tree_add_190_195_groupi_n_2343, csa_tree_add_190_195_groupi_n_2344, csa_tree_add_190_195_groupi_n_2345, csa_tree_add_190_195_groupi_n_2346, csa_tree_add_190_195_groupi_n_2347, csa_tree_add_190_195_groupi_n_2348, csa_tree_add_190_195_groupi_n_2349, csa_tree_add_190_195_groupi_n_2350;
  wire csa_tree_add_190_195_groupi_n_2351, csa_tree_add_190_195_groupi_n_2352, csa_tree_add_190_195_groupi_n_2353, csa_tree_add_190_195_groupi_n_2354, csa_tree_add_190_195_groupi_n_2355, csa_tree_add_190_195_groupi_n_2356, csa_tree_add_190_195_groupi_n_2357, csa_tree_add_190_195_groupi_n_2358;
  wire csa_tree_add_190_195_groupi_n_2359, csa_tree_add_190_195_groupi_n_2360, csa_tree_add_190_195_groupi_n_2361, csa_tree_add_190_195_groupi_n_2362, csa_tree_add_190_195_groupi_n_2363, csa_tree_add_190_195_groupi_n_2364, csa_tree_add_190_195_groupi_n_2365, csa_tree_add_190_195_groupi_n_2366;
  wire csa_tree_add_190_195_groupi_n_2367, csa_tree_add_190_195_groupi_n_2368, csa_tree_add_190_195_groupi_n_2369, csa_tree_add_190_195_groupi_n_2370, csa_tree_add_190_195_groupi_n_2371, csa_tree_add_190_195_groupi_n_2372, csa_tree_add_190_195_groupi_n_2373, csa_tree_add_190_195_groupi_n_2374;
  wire csa_tree_add_190_195_groupi_n_2375, csa_tree_add_190_195_groupi_n_2376, csa_tree_add_190_195_groupi_n_2377, csa_tree_add_190_195_groupi_n_2378, csa_tree_add_190_195_groupi_n_2379, csa_tree_add_190_195_groupi_n_2380, csa_tree_add_190_195_groupi_n_2381, csa_tree_add_190_195_groupi_n_2382;
  wire csa_tree_add_190_195_groupi_n_2383, csa_tree_add_190_195_groupi_n_2384, csa_tree_add_190_195_groupi_n_2385, csa_tree_add_190_195_groupi_n_2386, csa_tree_add_190_195_groupi_n_2387, csa_tree_add_190_195_groupi_n_2388, csa_tree_add_190_195_groupi_n_2389, csa_tree_add_190_195_groupi_n_2390;
  wire csa_tree_add_190_195_groupi_n_2391, csa_tree_add_190_195_groupi_n_2392, csa_tree_add_190_195_groupi_n_2393, csa_tree_add_190_195_groupi_n_2394, csa_tree_add_190_195_groupi_n_2395, csa_tree_add_190_195_groupi_n_2396, csa_tree_add_190_195_groupi_n_2397, csa_tree_add_190_195_groupi_n_2398;
  wire csa_tree_add_190_195_groupi_n_2399, csa_tree_add_190_195_groupi_n_2400, csa_tree_add_190_195_groupi_n_2401, csa_tree_add_190_195_groupi_n_2402, csa_tree_add_190_195_groupi_n_2403, csa_tree_add_190_195_groupi_n_2404, csa_tree_add_190_195_groupi_n_2405, csa_tree_add_190_195_groupi_n_2406;
  wire csa_tree_add_190_195_groupi_n_2407, csa_tree_add_190_195_groupi_n_2408, csa_tree_add_190_195_groupi_n_2409, csa_tree_add_190_195_groupi_n_2410, csa_tree_add_190_195_groupi_n_2411, csa_tree_add_190_195_groupi_n_2412, csa_tree_add_190_195_groupi_n_2413, csa_tree_add_190_195_groupi_n_2414;
  wire csa_tree_add_190_195_groupi_n_2415, csa_tree_add_190_195_groupi_n_2416, csa_tree_add_190_195_groupi_n_2417, csa_tree_add_190_195_groupi_n_2418, csa_tree_add_190_195_groupi_n_2419, csa_tree_add_190_195_groupi_n_2420, csa_tree_add_190_195_groupi_n_2421, csa_tree_add_190_195_groupi_n_2422;
  wire csa_tree_add_190_195_groupi_n_2423, csa_tree_add_190_195_groupi_n_2424, csa_tree_add_190_195_groupi_n_2425, csa_tree_add_190_195_groupi_n_2426, csa_tree_add_190_195_groupi_n_2427, csa_tree_add_190_195_groupi_n_2428, csa_tree_add_190_195_groupi_n_2429, csa_tree_add_190_195_groupi_n_2430;
  wire csa_tree_add_190_195_groupi_n_2431, csa_tree_add_190_195_groupi_n_2432, csa_tree_add_190_195_groupi_n_2433, csa_tree_add_190_195_groupi_n_2434, csa_tree_add_190_195_groupi_n_2435, csa_tree_add_190_195_groupi_n_2436, csa_tree_add_190_195_groupi_n_2437, csa_tree_add_190_195_groupi_n_2438;
  wire csa_tree_add_190_195_groupi_n_2439, csa_tree_add_190_195_groupi_n_2440, csa_tree_add_190_195_groupi_n_2441, csa_tree_add_190_195_groupi_n_2442, csa_tree_add_190_195_groupi_n_2443, csa_tree_add_190_195_groupi_n_2444, csa_tree_add_190_195_groupi_n_2445, csa_tree_add_190_195_groupi_n_2446;
  wire csa_tree_add_190_195_groupi_n_2447, csa_tree_add_190_195_groupi_n_2448, csa_tree_add_190_195_groupi_n_2449, csa_tree_add_190_195_groupi_n_2450, csa_tree_add_190_195_groupi_n_2451, csa_tree_add_190_195_groupi_n_2452, csa_tree_add_190_195_groupi_n_2453, csa_tree_add_190_195_groupi_n_2454;
  wire csa_tree_add_190_195_groupi_n_2455, csa_tree_add_190_195_groupi_n_2456, csa_tree_add_190_195_groupi_n_2457, csa_tree_add_190_195_groupi_n_2458, csa_tree_add_190_195_groupi_n_2459, csa_tree_add_190_195_groupi_n_2460, csa_tree_add_190_195_groupi_n_2461, csa_tree_add_190_195_groupi_n_2462;
  wire csa_tree_add_190_195_groupi_n_2463, csa_tree_add_190_195_groupi_n_2464, csa_tree_add_190_195_groupi_n_2465, csa_tree_add_190_195_groupi_n_2466, csa_tree_add_190_195_groupi_n_2467, csa_tree_add_190_195_groupi_n_2468, csa_tree_add_190_195_groupi_n_2469, csa_tree_add_190_195_groupi_n_2470;
  wire csa_tree_add_190_195_groupi_n_2471, csa_tree_add_190_195_groupi_n_2472, csa_tree_add_190_195_groupi_n_2473, csa_tree_add_190_195_groupi_n_2474, csa_tree_add_190_195_groupi_n_2475, csa_tree_add_190_195_groupi_n_2476, csa_tree_add_190_195_groupi_n_2477, csa_tree_add_190_195_groupi_n_2478;
  wire csa_tree_add_190_195_groupi_n_2479, csa_tree_add_190_195_groupi_n_2480, csa_tree_add_190_195_groupi_n_2481, csa_tree_add_190_195_groupi_n_2482, csa_tree_add_190_195_groupi_n_2483, csa_tree_add_190_195_groupi_n_2484, csa_tree_add_190_195_groupi_n_2485, csa_tree_add_190_195_groupi_n_2486;
  wire csa_tree_add_190_195_groupi_n_2487, csa_tree_add_190_195_groupi_n_2488, csa_tree_add_190_195_groupi_n_2489, csa_tree_add_190_195_groupi_n_2490, csa_tree_add_190_195_groupi_n_2491, csa_tree_add_190_195_groupi_n_2492, csa_tree_add_190_195_groupi_n_2493, csa_tree_add_190_195_groupi_n_2494;
  wire csa_tree_add_190_195_groupi_n_2495, csa_tree_add_190_195_groupi_n_2496, csa_tree_add_190_195_groupi_n_2497, csa_tree_add_190_195_groupi_n_2498, csa_tree_add_190_195_groupi_n_2499, csa_tree_add_190_195_groupi_n_2500, csa_tree_add_190_195_groupi_n_2501, csa_tree_add_190_195_groupi_n_2502;
  wire csa_tree_add_190_195_groupi_n_2503, csa_tree_add_190_195_groupi_n_2504, csa_tree_add_190_195_groupi_n_2505, csa_tree_add_190_195_groupi_n_2506, csa_tree_add_190_195_groupi_n_2507, csa_tree_add_190_195_groupi_n_2508, csa_tree_add_190_195_groupi_n_2509, csa_tree_add_190_195_groupi_n_2510;
  wire csa_tree_add_190_195_groupi_n_2511, csa_tree_add_190_195_groupi_n_2512, csa_tree_add_190_195_groupi_n_2513, csa_tree_add_190_195_groupi_n_2514, csa_tree_add_190_195_groupi_n_2515, csa_tree_add_190_195_groupi_n_2516, csa_tree_add_190_195_groupi_n_2517, csa_tree_add_190_195_groupi_n_2518;
  wire csa_tree_add_190_195_groupi_n_2519, csa_tree_add_190_195_groupi_n_2520, csa_tree_add_190_195_groupi_n_2521, csa_tree_add_190_195_groupi_n_2522, csa_tree_add_190_195_groupi_n_2523, csa_tree_add_190_195_groupi_n_2524, csa_tree_add_190_195_groupi_n_2525, csa_tree_add_190_195_groupi_n_2526;
  wire csa_tree_add_190_195_groupi_n_2527, csa_tree_add_190_195_groupi_n_2528, csa_tree_add_190_195_groupi_n_2529, csa_tree_add_190_195_groupi_n_2530, csa_tree_add_190_195_groupi_n_2531, csa_tree_add_190_195_groupi_n_2532, csa_tree_add_190_195_groupi_n_2533, csa_tree_add_190_195_groupi_n_2534;
  wire csa_tree_add_190_195_groupi_n_2535, csa_tree_add_190_195_groupi_n_2536, csa_tree_add_190_195_groupi_n_2537, csa_tree_add_190_195_groupi_n_2538, csa_tree_add_190_195_groupi_n_2539, csa_tree_add_190_195_groupi_n_2540, csa_tree_add_190_195_groupi_n_2541, csa_tree_add_190_195_groupi_n_2542;
  wire csa_tree_add_190_195_groupi_n_2543, csa_tree_add_190_195_groupi_n_2544, csa_tree_add_190_195_groupi_n_2545, csa_tree_add_190_195_groupi_n_2546, csa_tree_add_190_195_groupi_n_2547, csa_tree_add_190_195_groupi_n_2548, csa_tree_add_190_195_groupi_n_2549, csa_tree_add_190_195_groupi_n_2550;
  wire csa_tree_add_190_195_groupi_n_2551, csa_tree_add_190_195_groupi_n_2552, csa_tree_add_190_195_groupi_n_2553, csa_tree_add_190_195_groupi_n_2554, csa_tree_add_190_195_groupi_n_2555, csa_tree_add_190_195_groupi_n_2556, csa_tree_add_190_195_groupi_n_2557, csa_tree_add_190_195_groupi_n_2558;
  wire csa_tree_add_190_195_groupi_n_2559, csa_tree_add_190_195_groupi_n_2560, csa_tree_add_190_195_groupi_n_2561, csa_tree_add_190_195_groupi_n_2562, csa_tree_add_190_195_groupi_n_2563, csa_tree_add_190_195_groupi_n_2564, csa_tree_add_190_195_groupi_n_2565, csa_tree_add_190_195_groupi_n_2566;
  wire csa_tree_add_190_195_groupi_n_2567, csa_tree_add_190_195_groupi_n_2568, csa_tree_add_190_195_groupi_n_2569, csa_tree_add_190_195_groupi_n_2570, csa_tree_add_190_195_groupi_n_2571, csa_tree_add_190_195_groupi_n_2572, csa_tree_add_190_195_groupi_n_2573, csa_tree_add_190_195_groupi_n_2574;
  wire csa_tree_add_190_195_groupi_n_2575, csa_tree_add_190_195_groupi_n_2576, csa_tree_add_190_195_groupi_n_2577, csa_tree_add_190_195_groupi_n_2578, csa_tree_add_190_195_groupi_n_2579, csa_tree_add_190_195_groupi_n_2580, csa_tree_add_190_195_groupi_n_2581, csa_tree_add_190_195_groupi_n_2582;
  wire csa_tree_add_190_195_groupi_n_2583, csa_tree_add_190_195_groupi_n_2584, csa_tree_add_190_195_groupi_n_2585, csa_tree_add_190_195_groupi_n_2586, csa_tree_add_190_195_groupi_n_2587, csa_tree_add_190_195_groupi_n_2588, csa_tree_add_190_195_groupi_n_2589, csa_tree_add_190_195_groupi_n_2590;
  wire csa_tree_add_190_195_groupi_n_2591, csa_tree_add_190_195_groupi_n_2592, csa_tree_add_190_195_groupi_n_2593, csa_tree_add_190_195_groupi_n_2594, csa_tree_add_190_195_groupi_n_2595, csa_tree_add_190_195_groupi_n_2596, csa_tree_add_190_195_groupi_n_2597, csa_tree_add_190_195_groupi_n_2598;
  wire csa_tree_add_190_195_groupi_n_2599, csa_tree_add_190_195_groupi_n_2600, csa_tree_add_190_195_groupi_n_2601, csa_tree_add_190_195_groupi_n_2602, csa_tree_add_190_195_groupi_n_2603, csa_tree_add_190_195_groupi_n_2604, csa_tree_add_190_195_groupi_n_2605, csa_tree_add_190_195_groupi_n_2606;
  wire csa_tree_add_190_195_groupi_n_2607, csa_tree_add_190_195_groupi_n_2608, csa_tree_add_190_195_groupi_n_2609, csa_tree_add_190_195_groupi_n_2610, csa_tree_add_190_195_groupi_n_2611, csa_tree_add_190_195_groupi_n_2612, csa_tree_add_190_195_groupi_n_2613, csa_tree_add_190_195_groupi_n_2614;
  wire csa_tree_add_190_195_groupi_n_2615, csa_tree_add_190_195_groupi_n_2616, csa_tree_add_190_195_groupi_n_2617, csa_tree_add_190_195_groupi_n_2618, csa_tree_add_190_195_groupi_n_2619, csa_tree_add_190_195_groupi_n_2620, csa_tree_add_190_195_groupi_n_2621, csa_tree_add_190_195_groupi_n_2622;
  wire csa_tree_add_190_195_groupi_n_2623, csa_tree_add_190_195_groupi_n_2624, csa_tree_add_190_195_groupi_n_2625, csa_tree_add_190_195_groupi_n_2626, csa_tree_add_190_195_groupi_n_2627, csa_tree_add_190_195_groupi_n_2628, csa_tree_add_190_195_groupi_n_2629, csa_tree_add_190_195_groupi_n_2630;
  wire csa_tree_add_190_195_groupi_n_2631, csa_tree_add_190_195_groupi_n_2632, csa_tree_add_190_195_groupi_n_2633, csa_tree_add_190_195_groupi_n_2634, csa_tree_add_190_195_groupi_n_2635, csa_tree_add_190_195_groupi_n_2636, csa_tree_add_190_195_groupi_n_2637, csa_tree_add_190_195_groupi_n_2638;
  wire csa_tree_add_190_195_groupi_n_2639, csa_tree_add_190_195_groupi_n_2640, csa_tree_add_190_195_groupi_n_2641, csa_tree_add_190_195_groupi_n_2642, csa_tree_add_190_195_groupi_n_2643, csa_tree_add_190_195_groupi_n_2644, csa_tree_add_190_195_groupi_n_2645, csa_tree_add_190_195_groupi_n_2646;
  wire csa_tree_add_190_195_groupi_n_2647, csa_tree_add_190_195_groupi_n_2648, csa_tree_add_190_195_groupi_n_2649, csa_tree_add_190_195_groupi_n_2650, csa_tree_add_190_195_groupi_n_2651, csa_tree_add_190_195_groupi_n_2652, csa_tree_add_190_195_groupi_n_2653, csa_tree_add_190_195_groupi_n_2654;
  wire csa_tree_add_190_195_groupi_n_2655, csa_tree_add_190_195_groupi_n_2656, csa_tree_add_190_195_groupi_n_2657, csa_tree_add_190_195_groupi_n_2658, csa_tree_add_190_195_groupi_n_2659, csa_tree_add_190_195_groupi_n_2660, csa_tree_add_190_195_groupi_n_2661, csa_tree_add_190_195_groupi_n_2662;
  wire csa_tree_add_190_195_groupi_n_2663, csa_tree_add_190_195_groupi_n_2664, csa_tree_add_190_195_groupi_n_2665, csa_tree_add_190_195_groupi_n_2666, csa_tree_add_190_195_groupi_n_2667, csa_tree_add_190_195_groupi_n_2668, csa_tree_add_190_195_groupi_n_2669, csa_tree_add_190_195_groupi_n_2670;
  wire csa_tree_add_190_195_groupi_n_2671, csa_tree_add_190_195_groupi_n_2672, csa_tree_add_190_195_groupi_n_2673, csa_tree_add_190_195_groupi_n_2674, csa_tree_add_190_195_groupi_n_2675, csa_tree_add_190_195_groupi_n_2676, csa_tree_add_190_195_groupi_n_2677, csa_tree_add_190_195_groupi_n_2678;
  wire csa_tree_add_190_195_groupi_n_2679, csa_tree_add_190_195_groupi_n_2680, csa_tree_add_190_195_groupi_n_2681, csa_tree_add_190_195_groupi_n_2682, csa_tree_add_190_195_groupi_n_2683, csa_tree_add_190_195_groupi_n_2684, csa_tree_add_190_195_groupi_n_2685, csa_tree_add_190_195_groupi_n_2686;
  wire csa_tree_add_190_195_groupi_n_2687, csa_tree_add_190_195_groupi_n_2688, csa_tree_add_190_195_groupi_n_2689, csa_tree_add_190_195_groupi_n_2690, csa_tree_add_190_195_groupi_n_2691, csa_tree_add_190_195_groupi_n_2692, csa_tree_add_190_195_groupi_n_2693, csa_tree_add_190_195_groupi_n_2694;
  wire csa_tree_add_190_195_groupi_n_2695, csa_tree_add_190_195_groupi_n_2696, csa_tree_add_190_195_groupi_n_2697, csa_tree_add_190_195_groupi_n_2698, csa_tree_add_190_195_groupi_n_2699, csa_tree_add_190_195_groupi_n_2700, csa_tree_add_190_195_groupi_n_2701, csa_tree_add_190_195_groupi_n_2702;
  wire csa_tree_add_190_195_groupi_n_2703, csa_tree_add_190_195_groupi_n_2704, csa_tree_add_190_195_groupi_n_2705, csa_tree_add_190_195_groupi_n_2706, csa_tree_add_190_195_groupi_n_2707, csa_tree_add_190_195_groupi_n_2708, csa_tree_add_190_195_groupi_n_2709, csa_tree_add_190_195_groupi_n_2710;
  wire csa_tree_add_190_195_groupi_n_2711, csa_tree_add_190_195_groupi_n_2712, csa_tree_add_190_195_groupi_n_2713, csa_tree_add_190_195_groupi_n_2714, csa_tree_add_190_195_groupi_n_2715, csa_tree_add_190_195_groupi_n_2716, csa_tree_add_190_195_groupi_n_2717, csa_tree_add_190_195_groupi_n_2718;
  wire csa_tree_add_190_195_groupi_n_2719, csa_tree_add_190_195_groupi_n_2720, csa_tree_add_190_195_groupi_n_2721, csa_tree_add_190_195_groupi_n_2722, csa_tree_add_190_195_groupi_n_2723, csa_tree_add_190_195_groupi_n_2724, csa_tree_add_190_195_groupi_n_2725, csa_tree_add_190_195_groupi_n_2726;
  wire csa_tree_add_190_195_groupi_n_2727, csa_tree_add_190_195_groupi_n_2728, csa_tree_add_190_195_groupi_n_2729, csa_tree_add_190_195_groupi_n_2730, csa_tree_add_190_195_groupi_n_2731, csa_tree_add_190_195_groupi_n_2732, csa_tree_add_190_195_groupi_n_2733, csa_tree_add_190_195_groupi_n_2734;
  wire csa_tree_add_190_195_groupi_n_2735, csa_tree_add_190_195_groupi_n_2736, csa_tree_add_190_195_groupi_n_2737, csa_tree_add_190_195_groupi_n_2738, csa_tree_add_190_195_groupi_n_2739, csa_tree_add_190_195_groupi_n_2740, csa_tree_add_190_195_groupi_n_2741, csa_tree_add_190_195_groupi_n_2742;
  wire csa_tree_add_190_195_groupi_n_2743, csa_tree_add_190_195_groupi_n_2744, csa_tree_add_190_195_groupi_n_2745, csa_tree_add_190_195_groupi_n_2746, csa_tree_add_190_195_groupi_n_2747, csa_tree_add_190_195_groupi_n_2748, csa_tree_add_190_195_groupi_n_2749, csa_tree_add_190_195_groupi_n_2750;
  wire csa_tree_add_190_195_groupi_n_2751, csa_tree_add_190_195_groupi_n_2752, csa_tree_add_190_195_groupi_n_2753, csa_tree_add_190_195_groupi_n_2754, csa_tree_add_190_195_groupi_n_2755, csa_tree_add_190_195_groupi_n_2756, csa_tree_add_190_195_groupi_n_2757, csa_tree_add_190_195_groupi_n_2758;
  wire csa_tree_add_190_195_groupi_n_2759, csa_tree_add_190_195_groupi_n_2760, csa_tree_add_190_195_groupi_n_2761, csa_tree_add_190_195_groupi_n_2762, csa_tree_add_190_195_groupi_n_2763, csa_tree_add_190_195_groupi_n_2764, csa_tree_add_190_195_groupi_n_2765, csa_tree_add_190_195_groupi_n_2766;
  wire csa_tree_add_190_195_groupi_n_2767, csa_tree_add_190_195_groupi_n_2768, csa_tree_add_190_195_groupi_n_2769, csa_tree_add_190_195_groupi_n_2770, csa_tree_add_190_195_groupi_n_2771, csa_tree_add_190_195_groupi_n_2772, csa_tree_add_190_195_groupi_n_2773, csa_tree_add_190_195_groupi_n_2774;
  wire csa_tree_add_190_195_groupi_n_2775, csa_tree_add_190_195_groupi_n_2776, csa_tree_add_190_195_groupi_n_2777, csa_tree_add_190_195_groupi_n_2778, csa_tree_add_190_195_groupi_n_2779, csa_tree_add_190_195_groupi_n_2780, csa_tree_add_190_195_groupi_n_2781, csa_tree_add_190_195_groupi_n_2782;
  wire csa_tree_add_190_195_groupi_n_2783, csa_tree_add_190_195_groupi_n_2784, csa_tree_add_190_195_groupi_n_2785, csa_tree_add_190_195_groupi_n_2786, csa_tree_add_190_195_groupi_n_2787, csa_tree_add_190_195_groupi_n_2788, csa_tree_add_190_195_groupi_n_2789, csa_tree_add_190_195_groupi_n_2790;
  wire csa_tree_add_190_195_groupi_n_2791, csa_tree_add_190_195_groupi_n_2792, csa_tree_add_190_195_groupi_n_2793, csa_tree_add_190_195_groupi_n_2794, csa_tree_add_190_195_groupi_n_2795, csa_tree_add_190_195_groupi_n_2796, csa_tree_add_190_195_groupi_n_2797, csa_tree_add_190_195_groupi_n_2798;
  wire csa_tree_add_190_195_groupi_n_2799, csa_tree_add_190_195_groupi_n_2800, csa_tree_add_190_195_groupi_n_2801, csa_tree_add_190_195_groupi_n_2802, csa_tree_add_190_195_groupi_n_2803, csa_tree_add_190_195_groupi_n_2804, csa_tree_add_190_195_groupi_n_2805, csa_tree_add_190_195_groupi_n_2806;
  wire csa_tree_add_190_195_groupi_n_2807, csa_tree_add_190_195_groupi_n_2808, csa_tree_add_190_195_groupi_n_2809, csa_tree_add_190_195_groupi_n_2810, csa_tree_add_190_195_groupi_n_2811, csa_tree_add_190_195_groupi_n_2812, csa_tree_add_190_195_groupi_n_2813, csa_tree_add_190_195_groupi_n_2814;
  wire csa_tree_add_190_195_groupi_n_2815, csa_tree_add_190_195_groupi_n_2816, csa_tree_add_190_195_groupi_n_2817, csa_tree_add_190_195_groupi_n_2818, csa_tree_add_190_195_groupi_n_2819, csa_tree_add_190_195_groupi_n_2820, csa_tree_add_190_195_groupi_n_2821, csa_tree_add_190_195_groupi_n_2822;
  wire csa_tree_add_190_195_groupi_n_2823, csa_tree_add_190_195_groupi_n_2824, csa_tree_add_190_195_groupi_n_2825, csa_tree_add_190_195_groupi_n_2826, csa_tree_add_190_195_groupi_n_2827, csa_tree_add_190_195_groupi_n_2828, csa_tree_add_190_195_groupi_n_2829, csa_tree_add_190_195_groupi_n_2830;
  wire csa_tree_add_190_195_groupi_n_2831, csa_tree_add_190_195_groupi_n_2832, csa_tree_add_190_195_groupi_n_2833, csa_tree_add_190_195_groupi_n_2834, csa_tree_add_190_195_groupi_n_2835, csa_tree_add_190_195_groupi_n_2836, csa_tree_add_190_195_groupi_n_2837, csa_tree_add_190_195_groupi_n_2838;
  wire csa_tree_add_190_195_groupi_n_2839, csa_tree_add_190_195_groupi_n_2840, csa_tree_add_190_195_groupi_n_2841, csa_tree_add_190_195_groupi_n_2842, csa_tree_add_190_195_groupi_n_2843, csa_tree_add_190_195_groupi_n_2844, csa_tree_add_190_195_groupi_n_2845, csa_tree_add_190_195_groupi_n_2846;
  wire csa_tree_add_190_195_groupi_n_2847, csa_tree_add_190_195_groupi_n_2848, csa_tree_add_190_195_groupi_n_2849, csa_tree_add_190_195_groupi_n_2850, csa_tree_add_190_195_groupi_n_2851, csa_tree_add_190_195_groupi_n_2852, csa_tree_add_190_195_groupi_n_2853, csa_tree_add_190_195_groupi_n_2854;
  wire csa_tree_add_190_195_groupi_n_2855, csa_tree_add_190_195_groupi_n_2856, csa_tree_add_190_195_groupi_n_2857, csa_tree_add_190_195_groupi_n_2858, csa_tree_add_190_195_groupi_n_2859, csa_tree_add_190_195_groupi_n_2860, csa_tree_add_190_195_groupi_n_2861, csa_tree_add_190_195_groupi_n_2862;
  wire csa_tree_add_190_195_groupi_n_2863, csa_tree_add_190_195_groupi_n_2864, csa_tree_add_190_195_groupi_n_2865, csa_tree_add_190_195_groupi_n_2866, csa_tree_add_190_195_groupi_n_2867, csa_tree_add_190_195_groupi_n_2868, csa_tree_add_190_195_groupi_n_2869, csa_tree_add_190_195_groupi_n_2870;
  wire csa_tree_add_190_195_groupi_n_2871, csa_tree_add_190_195_groupi_n_2872, csa_tree_add_190_195_groupi_n_2873, csa_tree_add_190_195_groupi_n_2874, csa_tree_add_190_195_groupi_n_2875, csa_tree_add_190_195_groupi_n_2876, csa_tree_add_190_195_groupi_n_2877, csa_tree_add_190_195_groupi_n_2878;
  wire csa_tree_add_190_195_groupi_n_2879, csa_tree_add_190_195_groupi_n_2880, csa_tree_add_190_195_groupi_n_2881, csa_tree_add_190_195_groupi_n_2882, csa_tree_add_190_195_groupi_n_2883, csa_tree_add_190_195_groupi_n_2884, csa_tree_add_190_195_groupi_n_2885, csa_tree_add_190_195_groupi_n_2886;
  wire csa_tree_add_190_195_groupi_n_2887, csa_tree_add_190_195_groupi_n_2888, csa_tree_add_190_195_groupi_n_2889, csa_tree_add_190_195_groupi_n_2890, csa_tree_add_190_195_groupi_n_2891, csa_tree_add_190_195_groupi_n_2892, csa_tree_add_190_195_groupi_n_2893, csa_tree_add_190_195_groupi_n_2894;
  wire csa_tree_add_190_195_groupi_n_2895, csa_tree_add_190_195_groupi_n_2896, csa_tree_add_190_195_groupi_n_2897, csa_tree_add_190_195_groupi_n_2898, csa_tree_add_190_195_groupi_n_2899, csa_tree_add_190_195_groupi_n_2900, csa_tree_add_190_195_groupi_n_2901, csa_tree_add_190_195_groupi_n_2902;
  wire csa_tree_add_190_195_groupi_n_2903, csa_tree_add_190_195_groupi_n_2904, csa_tree_add_190_195_groupi_n_2905, csa_tree_add_190_195_groupi_n_2906, csa_tree_add_190_195_groupi_n_2907, csa_tree_add_190_195_groupi_n_2908, csa_tree_add_190_195_groupi_n_2909, csa_tree_add_190_195_groupi_n_2910;
  wire csa_tree_add_190_195_groupi_n_2911, csa_tree_add_190_195_groupi_n_2912, csa_tree_add_190_195_groupi_n_2913, csa_tree_add_190_195_groupi_n_2914, csa_tree_add_190_195_groupi_n_2915, csa_tree_add_190_195_groupi_n_2916, csa_tree_add_190_195_groupi_n_2917, csa_tree_add_190_195_groupi_n_2918;
  wire csa_tree_add_190_195_groupi_n_2919, csa_tree_add_190_195_groupi_n_2920, csa_tree_add_190_195_groupi_n_2921, csa_tree_add_190_195_groupi_n_2922, csa_tree_add_190_195_groupi_n_2923, csa_tree_add_190_195_groupi_n_2924, csa_tree_add_190_195_groupi_n_2925, csa_tree_add_190_195_groupi_n_2926;
  wire csa_tree_add_190_195_groupi_n_2927, csa_tree_add_190_195_groupi_n_2928, csa_tree_add_190_195_groupi_n_2929, csa_tree_add_190_195_groupi_n_2930, csa_tree_add_190_195_groupi_n_2931, csa_tree_add_190_195_groupi_n_2932, csa_tree_add_190_195_groupi_n_2933, csa_tree_add_190_195_groupi_n_2934;
  wire csa_tree_add_190_195_groupi_n_2935, csa_tree_add_190_195_groupi_n_2936, csa_tree_add_190_195_groupi_n_2937, csa_tree_add_190_195_groupi_n_2938, csa_tree_add_190_195_groupi_n_2939, csa_tree_add_190_195_groupi_n_2940, csa_tree_add_190_195_groupi_n_2941, csa_tree_add_190_195_groupi_n_2942;
  wire csa_tree_add_190_195_groupi_n_2943, csa_tree_add_190_195_groupi_n_2944, csa_tree_add_190_195_groupi_n_2945, csa_tree_add_190_195_groupi_n_2946, csa_tree_add_190_195_groupi_n_2947, csa_tree_add_190_195_groupi_n_2948, csa_tree_add_190_195_groupi_n_2949, csa_tree_add_190_195_groupi_n_2950;
  wire csa_tree_add_190_195_groupi_n_2951, csa_tree_add_190_195_groupi_n_2952, csa_tree_add_190_195_groupi_n_2953, csa_tree_add_190_195_groupi_n_2954, csa_tree_add_190_195_groupi_n_2955, csa_tree_add_190_195_groupi_n_2956, csa_tree_add_190_195_groupi_n_2957, csa_tree_add_190_195_groupi_n_2958;
  wire csa_tree_add_190_195_groupi_n_2959, csa_tree_add_190_195_groupi_n_2960, csa_tree_add_190_195_groupi_n_2961, csa_tree_add_190_195_groupi_n_2962, csa_tree_add_190_195_groupi_n_2963, csa_tree_add_190_195_groupi_n_2964, csa_tree_add_190_195_groupi_n_2965, csa_tree_add_190_195_groupi_n_2966;
  wire csa_tree_add_190_195_groupi_n_2967, csa_tree_add_190_195_groupi_n_2968, csa_tree_add_190_195_groupi_n_2969, csa_tree_add_190_195_groupi_n_2970, csa_tree_add_190_195_groupi_n_2971, csa_tree_add_190_195_groupi_n_2972, csa_tree_add_190_195_groupi_n_2973, csa_tree_add_190_195_groupi_n_2975;
  wire csa_tree_add_190_195_groupi_n_2976, csa_tree_add_190_195_groupi_n_2977, csa_tree_add_190_195_groupi_n_2978, csa_tree_add_190_195_groupi_n_2979, csa_tree_add_190_195_groupi_n_2980, csa_tree_add_190_195_groupi_n_2981, csa_tree_add_190_195_groupi_n_2982, csa_tree_add_190_195_groupi_n_2983;
  wire csa_tree_add_190_195_groupi_n_2984, csa_tree_add_190_195_groupi_n_2985, csa_tree_add_190_195_groupi_n_2986, csa_tree_add_190_195_groupi_n_2987, csa_tree_add_190_195_groupi_n_2988, csa_tree_add_190_195_groupi_n_2989, csa_tree_add_190_195_groupi_n_2990, csa_tree_add_190_195_groupi_n_2991;
  wire csa_tree_add_190_195_groupi_n_2992, csa_tree_add_190_195_groupi_n_2993, csa_tree_add_190_195_groupi_n_2994, csa_tree_add_190_195_groupi_n_2995, csa_tree_add_190_195_groupi_n_2996, csa_tree_add_190_195_groupi_n_2997, csa_tree_add_190_195_groupi_n_2998, csa_tree_add_190_195_groupi_n_2999;
  wire csa_tree_add_190_195_groupi_n_3000, csa_tree_add_190_195_groupi_n_3001, csa_tree_add_190_195_groupi_n_3002, csa_tree_add_190_195_groupi_n_3003, csa_tree_add_190_195_groupi_n_3004, csa_tree_add_190_195_groupi_n_3005, csa_tree_add_190_195_groupi_n_3006, csa_tree_add_190_195_groupi_n_3007;
  wire csa_tree_add_190_195_groupi_n_3008, csa_tree_add_190_195_groupi_n_3009, csa_tree_add_190_195_groupi_n_3010, csa_tree_add_190_195_groupi_n_3011, csa_tree_add_190_195_groupi_n_3012, csa_tree_add_190_195_groupi_n_3013, csa_tree_add_190_195_groupi_n_3014, csa_tree_add_190_195_groupi_n_3015;
  wire csa_tree_add_190_195_groupi_n_3016, csa_tree_add_190_195_groupi_n_3017, csa_tree_add_190_195_groupi_n_3018, csa_tree_add_190_195_groupi_n_3019, csa_tree_add_190_195_groupi_n_3020, csa_tree_add_190_195_groupi_n_3021, csa_tree_add_190_195_groupi_n_3022, csa_tree_add_190_195_groupi_n_3023;
  wire csa_tree_add_190_195_groupi_n_3024, csa_tree_add_190_195_groupi_n_3025, csa_tree_add_190_195_groupi_n_3026, csa_tree_add_190_195_groupi_n_3027, csa_tree_add_190_195_groupi_n_3028, csa_tree_add_190_195_groupi_n_3029, csa_tree_add_190_195_groupi_n_3030, csa_tree_add_190_195_groupi_n_3031;
  wire csa_tree_add_190_195_groupi_n_3032, csa_tree_add_190_195_groupi_n_3033, csa_tree_add_190_195_groupi_n_3034, csa_tree_add_190_195_groupi_n_3035, csa_tree_add_190_195_groupi_n_3036, csa_tree_add_190_195_groupi_n_3037, csa_tree_add_190_195_groupi_n_3038, csa_tree_add_190_195_groupi_n_3039;
  wire csa_tree_add_190_195_groupi_n_3040, csa_tree_add_190_195_groupi_n_3041, csa_tree_add_190_195_groupi_n_3042, csa_tree_add_190_195_groupi_n_3043, csa_tree_add_190_195_groupi_n_3044, csa_tree_add_190_195_groupi_n_3045, csa_tree_add_190_195_groupi_n_3046, csa_tree_add_190_195_groupi_n_3047;
  wire csa_tree_add_190_195_groupi_n_3048, csa_tree_add_190_195_groupi_n_3049, csa_tree_add_190_195_groupi_n_3050, csa_tree_add_190_195_groupi_n_3051, csa_tree_add_190_195_groupi_n_3052, csa_tree_add_190_195_groupi_n_3053, csa_tree_add_190_195_groupi_n_3054, csa_tree_add_190_195_groupi_n_3055;
  wire csa_tree_add_190_195_groupi_n_3056, csa_tree_add_190_195_groupi_n_3057, csa_tree_add_190_195_groupi_n_3058, csa_tree_add_190_195_groupi_n_3059, csa_tree_add_190_195_groupi_n_3060, csa_tree_add_190_195_groupi_n_3061, csa_tree_add_190_195_groupi_n_3062, csa_tree_add_190_195_groupi_n_3063;
  wire csa_tree_add_190_195_groupi_n_3064, csa_tree_add_190_195_groupi_n_3065, csa_tree_add_190_195_groupi_n_3066, csa_tree_add_190_195_groupi_n_3067, csa_tree_add_190_195_groupi_n_3068, csa_tree_add_190_195_groupi_n_3069, csa_tree_add_190_195_groupi_n_3070, csa_tree_add_190_195_groupi_n_3071;
  wire csa_tree_add_190_195_groupi_n_3072, csa_tree_add_190_195_groupi_n_3073, csa_tree_add_190_195_groupi_n_3074, csa_tree_add_190_195_groupi_n_3075, csa_tree_add_190_195_groupi_n_3076, csa_tree_add_190_195_groupi_n_3077, csa_tree_add_190_195_groupi_n_3078, csa_tree_add_190_195_groupi_n_3079;
  wire csa_tree_add_190_195_groupi_n_3080, csa_tree_add_190_195_groupi_n_3081, csa_tree_add_190_195_groupi_n_3082, csa_tree_add_190_195_groupi_n_3083, csa_tree_add_190_195_groupi_n_3084, csa_tree_add_190_195_groupi_n_3085, csa_tree_add_190_195_groupi_n_3086, csa_tree_add_190_195_groupi_n_3087;
  wire csa_tree_add_190_195_groupi_n_3088, csa_tree_add_190_195_groupi_n_3089, csa_tree_add_190_195_groupi_n_3090, csa_tree_add_190_195_groupi_n_3091, csa_tree_add_190_195_groupi_n_3092, csa_tree_add_190_195_groupi_n_3093, csa_tree_add_190_195_groupi_n_3094, csa_tree_add_190_195_groupi_n_3095;
  wire csa_tree_add_190_195_groupi_n_3096, csa_tree_add_190_195_groupi_n_3097, csa_tree_add_190_195_groupi_n_3098, csa_tree_add_190_195_groupi_n_3099, csa_tree_add_190_195_groupi_n_3100, csa_tree_add_190_195_groupi_n_3101, csa_tree_add_190_195_groupi_n_3102, csa_tree_add_190_195_groupi_n_3103;
  wire csa_tree_add_190_195_groupi_n_3104, csa_tree_add_190_195_groupi_n_3105, csa_tree_add_190_195_groupi_n_3106, csa_tree_add_190_195_groupi_n_3107, csa_tree_add_190_195_groupi_n_3108, csa_tree_add_190_195_groupi_n_3109, csa_tree_add_190_195_groupi_n_3110, csa_tree_add_190_195_groupi_n_3111;
  wire csa_tree_add_190_195_groupi_n_3112, csa_tree_add_190_195_groupi_n_3113, csa_tree_add_190_195_groupi_n_3114, csa_tree_add_190_195_groupi_n_3115, csa_tree_add_190_195_groupi_n_3116, csa_tree_add_190_195_groupi_n_3117, csa_tree_add_190_195_groupi_n_3118, csa_tree_add_190_195_groupi_n_3119;
  wire csa_tree_add_190_195_groupi_n_3120, csa_tree_add_190_195_groupi_n_3121, csa_tree_add_190_195_groupi_n_3122, csa_tree_add_190_195_groupi_n_3123, csa_tree_add_190_195_groupi_n_3124, csa_tree_add_190_195_groupi_n_3125, csa_tree_add_190_195_groupi_n_3126, csa_tree_add_190_195_groupi_n_3127;
  wire csa_tree_add_190_195_groupi_n_3128, csa_tree_add_190_195_groupi_n_3129, csa_tree_add_190_195_groupi_n_3130, csa_tree_add_190_195_groupi_n_3131, csa_tree_add_190_195_groupi_n_3132, csa_tree_add_190_195_groupi_n_3133, csa_tree_add_190_195_groupi_n_3134, csa_tree_add_190_195_groupi_n_3135;
  wire csa_tree_add_190_195_groupi_n_3136, csa_tree_add_190_195_groupi_n_3137, csa_tree_add_190_195_groupi_n_3138, csa_tree_add_190_195_groupi_n_3139, csa_tree_add_190_195_groupi_n_3140, csa_tree_add_190_195_groupi_n_3141, csa_tree_add_190_195_groupi_n_3142, csa_tree_add_190_195_groupi_n_3143;
  wire csa_tree_add_190_195_groupi_n_3144, csa_tree_add_190_195_groupi_n_3145, csa_tree_add_190_195_groupi_n_3146, csa_tree_add_190_195_groupi_n_3147, csa_tree_add_190_195_groupi_n_3148, csa_tree_add_190_195_groupi_n_3149, csa_tree_add_190_195_groupi_n_3150, csa_tree_add_190_195_groupi_n_3151;
  wire csa_tree_add_190_195_groupi_n_3152, csa_tree_add_190_195_groupi_n_3153, csa_tree_add_190_195_groupi_n_3154, csa_tree_add_190_195_groupi_n_3155, csa_tree_add_190_195_groupi_n_3156, csa_tree_add_190_195_groupi_n_3157, csa_tree_add_190_195_groupi_n_3158, csa_tree_add_190_195_groupi_n_3159;
  wire csa_tree_add_190_195_groupi_n_3160, csa_tree_add_190_195_groupi_n_3161, csa_tree_add_190_195_groupi_n_3162, csa_tree_add_190_195_groupi_n_3163, csa_tree_add_190_195_groupi_n_3164, csa_tree_add_190_195_groupi_n_3165, csa_tree_add_190_195_groupi_n_3166, csa_tree_add_190_195_groupi_n_3167;
  wire csa_tree_add_190_195_groupi_n_3168, csa_tree_add_190_195_groupi_n_3169, csa_tree_add_190_195_groupi_n_3170, csa_tree_add_190_195_groupi_n_3171, csa_tree_add_190_195_groupi_n_3172, csa_tree_add_190_195_groupi_n_3173, csa_tree_add_190_195_groupi_n_3174, csa_tree_add_190_195_groupi_n_3175;
  wire csa_tree_add_190_195_groupi_n_3176, csa_tree_add_190_195_groupi_n_3177, csa_tree_add_190_195_groupi_n_3178, csa_tree_add_190_195_groupi_n_3179, csa_tree_add_190_195_groupi_n_3180, csa_tree_add_190_195_groupi_n_3181, csa_tree_add_190_195_groupi_n_3182, csa_tree_add_190_195_groupi_n_3183;
  wire csa_tree_add_190_195_groupi_n_3184, csa_tree_add_190_195_groupi_n_3185, csa_tree_add_190_195_groupi_n_3186, csa_tree_add_190_195_groupi_n_3187, csa_tree_add_190_195_groupi_n_3188, csa_tree_add_190_195_groupi_n_3189, csa_tree_add_190_195_groupi_n_3190, csa_tree_add_190_195_groupi_n_3191;
  wire csa_tree_add_190_195_groupi_n_3192, csa_tree_add_190_195_groupi_n_3193, csa_tree_add_190_195_groupi_n_3194, csa_tree_add_190_195_groupi_n_3195, csa_tree_add_190_195_groupi_n_3196, csa_tree_add_190_195_groupi_n_3197, csa_tree_add_190_195_groupi_n_3198, csa_tree_add_190_195_groupi_n_3199;
  wire csa_tree_add_190_195_groupi_n_3200, csa_tree_add_190_195_groupi_n_3201, csa_tree_add_190_195_groupi_n_3202, csa_tree_add_190_195_groupi_n_3203, csa_tree_add_190_195_groupi_n_3204, csa_tree_add_190_195_groupi_n_3205, csa_tree_add_190_195_groupi_n_3206, csa_tree_add_190_195_groupi_n_3207;
  wire csa_tree_add_190_195_groupi_n_3208, csa_tree_add_190_195_groupi_n_3209, csa_tree_add_190_195_groupi_n_3210, csa_tree_add_190_195_groupi_n_3211, csa_tree_add_190_195_groupi_n_3212, csa_tree_add_190_195_groupi_n_3213, csa_tree_add_190_195_groupi_n_3214, csa_tree_add_190_195_groupi_n_3215;
  wire csa_tree_add_190_195_groupi_n_3216, csa_tree_add_190_195_groupi_n_3217, csa_tree_add_190_195_groupi_n_3218, csa_tree_add_190_195_groupi_n_3219, csa_tree_add_190_195_groupi_n_3220, csa_tree_add_190_195_groupi_n_3221, csa_tree_add_190_195_groupi_n_3222, csa_tree_add_190_195_groupi_n_3223;
  wire csa_tree_add_190_195_groupi_n_3224, csa_tree_add_190_195_groupi_n_3225, csa_tree_add_190_195_groupi_n_3226, csa_tree_add_190_195_groupi_n_3227, csa_tree_add_190_195_groupi_n_3228, csa_tree_add_190_195_groupi_n_3229, csa_tree_add_190_195_groupi_n_3230, csa_tree_add_190_195_groupi_n_3231;
  wire csa_tree_add_190_195_groupi_n_3232, csa_tree_add_190_195_groupi_n_3233, csa_tree_add_190_195_groupi_n_3234, csa_tree_add_190_195_groupi_n_3235, csa_tree_add_190_195_groupi_n_3236, csa_tree_add_190_195_groupi_n_3237, csa_tree_add_190_195_groupi_n_3238, csa_tree_add_190_195_groupi_n_3239;
  wire csa_tree_add_190_195_groupi_n_3240, csa_tree_add_190_195_groupi_n_3241, csa_tree_add_190_195_groupi_n_3242, csa_tree_add_190_195_groupi_n_3243, csa_tree_add_190_195_groupi_n_3244, csa_tree_add_190_195_groupi_n_3245, csa_tree_add_190_195_groupi_n_3246, csa_tree_add_190_195_groupi_n_3247;
  wire csa_tree_add_190_195_groupi_n_3248, csa_tree_add_190_195_groupi_n_3249, csa_tree_add_190_195_groupi_n_3250, csa_tree_add_190_195_groupi_n_3251, csa_tree_add_190_195_groupi_n_3252, csa_tree_add_190_195_groupi_n_3253, csa_tree_add_190_195_groupi_n_3254, csa_tree_add_190_195_groupi_n_3255;
  wire csa_tree_add_190_195_groupi_n_3256, csa_tree_add_190_195_groupi_n_3257, csa_tree_add_190_195_groupi_n_3258, csa_tree_add_190_195_groupi_n_3259, csa_tree_add_190_195_groupi_n_3260, csa_tree_add_190_195_groupi_n_3261, csa_tree_add_190_195_groupi_n_3262, csa_tree_add_190_195_groupi_n_3263;
  wire csa_tree_add_190_195_groupi_n_3264, csa_tree_add_190_195_groupi_n_3265, csa_tree_add_190_195_groupi_n_3266, csa_tree_add_190_195_groupi_n_3267, csa_tree_add_190_195_groupi_n_3268, csa_tree_add_190_195_groupi_n_3269, csa_tree_add_190_195_groupi_n_3270, csa_tree_add_190_195_groupi_n_3271;
  wire csa_tree_add_190_195_groupi_n_3272, csa_tree_add_190_195_groupi_n_3273, csa_tree_add_190_195_groupi_n_3274, csa_tree_add_190_195_groupi_n_3275, csa_tree_add_190_195_groupi_n_3276, csa_tree_add_190_195_groupi_n_3277, csa_tree_add_190_195_groupi_n_3278, csa_tree_add_190_195_groupi_n_3279;
  wire csa_tree_add_190_195_groupi_n_3280, csa_tree_add_190_195_groupi_n_3281, csa_tree_add_190_195_groupi_n_3282, csa_tree_add_190_195_groupi_n_3283, csa_tree_add_190_195_groupi_n_3284, csa_tree_add_190_195_groupi_n_3285, csa_tree_add_190_195_groupi_n_3286, csa_tree_add_190_195_groupi_n_3287;
  wire csa_tree_add_190_195_groupi_n_3288, csa_tree_add_190_195_groupi_n_3289, csa_tree_add_190_195_groupi_n_3290, csa_tree_add_190_195_groupi_n_3291, csa_tree_add_190_195_groupi_n_3292, csa_tree_add_190_195_groupi_n_3293, csa_tree_add_190_195_groupi_n_3294, csa_tree_add_190_195_groupi_n_3295;
  wire csa_tree_add_190_195_groupi_n_3296, csa_tree_add_190_195_groupi_n_3297, csa_tree_add_190_195_groupi_n_3298, csa_tree_add_190_195_groupi_n_3299, csa_tree_add_190_195_groupi_n_3300, csa_tree_add_190_195_groupi_n_3301, csa_tree_add_190_195_groupi_n_3302, csa_tree_add_190_195_groupi_n_3303;
  wire csa_tree_add_190_195_groupi_n_3304, csa_tree_add_190_195_groupi_n_3305, csa_tree_add_190_195_groupi_n_3306, csa_tree_add_190_195_groupi_n_3307, csa_tree_add_190_195_groupi_n_3308, csa_tree_add_190_195_groupi_n_3309, csa_tree_add_190_195_groupi_n_3310, csa_tree_add_190_195_groupi_n_3311;
  wire csa_tree_add_190_195_groupi_n_3312, csa_tree_add_190_195_groupi_n_3313, csa_tree_add_190_195_groupi_n_3314, csa_tree_add_190_195_groupi_n_3315, csa_tree_add_190_195_groupi_n_3316, csa_tree_add_190_195_groupi_n_3317, csa_tree_add_190_195_groupi_n_3318, csa_tree_add_190_195_groupi_n_3319;
  wire csa_tree_add_190_195_groupi_n_3320, csa_tree_add_190_195_groupi_n_3321, csa_tree_add_190_195_groupi_n_3322, csa_tree_add_190_195_groupi_n_3323, csa_tree_add_190_195_groupi_n_3324, csa_tree_add_190_195_groupi_n_3325, csa_tree_add_190_195_groupi_n_3326, csa_tree_add_190_195_groupi_n_3327;
  wire csa_tree_add_190_195_groupi_n_3328, csa_tree_add_190_195_groupi_n_3329, csa_tree_add_190_195_groupi_n_3330, csa_tree_add_190_195_groupi_n_3331, csa_tree_add_190_195_groupi_n_3332, csa_tree_add_190_195_groupi_n_3333, csa_tree_add_190_195_groupi_n_3334, csa_tree_add_190_195_groupi_n_3335;
  wire csa_tree_add_190_195_groupi_n_3336, csa_tree_add_190_195_groupi_n_3337, csa_tree_add_190_195_groupi_n_3338, csa_tree_add_190_195_groupi_n_3339, csa_tree_add_190_195_groupi_n_3340, csa_tree_add_190_195_groupi_n_3341, csa_tree_add_190_195_groupi_n_3342, csa_tree_add_190_195_groupi_n_3343;
  wire csa_tree_add_190_195_groupi_n_3344, csa_tree_add_190_195_groupi_n_3345, csa_tree_add_190_195_groupi_n_3346, csa_tree_add_190_195_groupi_n_3347, csa_tree_add_190_195_groupi_n_3348, csa_tree_add_190_195_groupi_n_3349, csa_tree_add_190_195_groupi_n_3350, csa_tree_add_190_195_groupi_n_3351;
  wire csa_tree_add_190_195_groupi_n_3352, csa_tree_add_190_195_groupi_n_3353, csa_tree_add_190_195_groupi_n_3354, csa_tree_add_190_195_groupi_n_3355, csa_tree_add_190_195_groupi_n_3356, csa_tree_add_190_195_groupi_n_3357, csa_tree_add_190_195_groupi_n_3358, csa_tree_add_190_195_groupi_n_3359;
  wire csa_tree_add_190_195_groupi_n_3360, csa_tree_add_190_195_groupi_n_3361, csa_tree_add_190_195_groupi_n_3362, csa_tree_add_190_195_groupi_n_3363, csa_tree_add_190_195_groupi_n_3364, csa_tree_add_190_195_groupi_n_3365, csa_tree_add_190_195_groupi_n_3366, csa_tree_add_190_195_groupi_n_3367;
  wire csa_tree_add_190_195_groupi_n_3368, csa_tree_add_190_195_groupi_n_3369, csa_tree_add_190_195_groupi_n_3370, csa_tree_add_190_195_groupi_n_3371, csa_tree_add_190_195_groupi_n_3372, csa_tree_add_190_195_groupi_n_3373, csa_tree_add_190_195_groupi_n_3374, csa_tree_add_190_195_groupi_n_3375;
  wire csa_tree_add_190_195_groupi_n_3376, csa_tree_add_190_195_groupi_n_3377, csa_tree_add_190_195_groupi_n_3378, csa_tree_add_190_195_groupi_n_3379, csa_tree_add_190_195_groupi_n_3380, csa_tree_add_190_195_groupi_n_3381, csa_tree_add_190_195_groupi_n_3382, csa_tree_add_190_195_groupi_n_3383;
  wire csa_tree_add_190_195_groupi_n_3384, csa_tree_add_190_195_groupi_n_3385, csa_tree_add_190_195_groupi_n_3386, csa_tree_add_190_195_groupi_n_3387, csa_tree_add_190_195_groupi_n_3388, csa_tree_add_190_195_groupi_n_3389, csa_tree_add_190_195_groupi_n_3390, csa_tree_add_190_195_groupi_n_3391;
  wire csa_tree_add_190_195_groupi_n_3392, csa_tree_add_190_195_groupi_n_3393, csa_tree_add_190_195_groupi_n_3394, csa_tree_add_190_195_groupi_n_3395, csa_tree_add_190_195_groupi_n_3396, csa_tree_add_190_195_groupi_n_3397, csa_tree_add_190_195_groupi_n_3398, csa_tree_add_190_195_groupi_n_3399;
  wire csa_tree_add_190_195_groupi_n_3400, csa_tree_add_190_195_groupi_n_3401, csa_tree_add_190_195_groupi_n_3402, csa_tree_add_190_195_groupi_n_3403, csa_tree_add_190_195_groupi_n_3404, csa_tree_add_190_195_groupi_n_3405, csa_tree_add_190_195_groupi_n_3406, csa_tree_add_190_195_groupi_n_3407;
  wire csa_tree_add_190_195_groupi_n_3408, csa_tree_add_190_195_groupi_n_3409, csa_tree_add_190_195_groupi_n_3410, csa_tree_add_190_195_groupi_n_3411, csa_tree_add_190_195_groupi_n_3412, csa_tree_add_190_195_groupi_n_3413, csa_tree_add_190_195_groupi_n_3414, csa_tree_add_190_195_groupi_n_3415;
  wire csa_tree_add_190_195_groupi_n_3416, csa_tree_add_190_195_groupi_n_3417, csa_tree_add_190_195_groupi_n_3418, csa_tree_add_190_195_groupi_n_3419, csa_tree_add_190_195_groupi_n_3420, csa_tree_add_190_195_groupi_n_3421, csa_tree_add_190_195_groupi_n_3422, csa_tree_add_190_195_groupi_n_3423;
  wire csa_tree_add_190_195_groupi_n_3424, csa_tree_add_190_195_groupi_n_3425, csa_tree_add_190_195_groupi_n_3426, csa_tree_add_190_195_groupi_n_3427, csa_tree_add_190_195_groupi_n_3428, csa_tree_add_190_195_groupi_n_3429, csa_tree_add_190_195_groupi_n_3430, csa_tree_add_190_195_groupi_n_3431;
  wire csa_tree_add_190_195_groupi_n_3432, csa_tree_add_190_195_groupi_n_3433, csa_tree_add_190_195_groupi_n_3434, csa_tree_add_190_195_groupi_n_3435, csa_tree_add_190_195_groupi_n_3436, csa_tree_add_190_195_groupi_n_3437, csa_tree_add_190_195_groupi_n_3438, csa_tree_add_190_195_groupi_n_3439;
  wire csa_tree_add_190_195_groupi_n_3440, csa_tree_add_190_195_groupi_n_3441, csa_tree_add_190_195_groupi_n_3442, csa_tree_add_190_195_groupi_n_3443, csa_tree_add_190_195_groupi_n_3444, csa_tree_add_190_195_groupi_n_3445, csa_tree_add_190_195_groupi_n_3446, csa_tree_add_190_195_groupi_n_3447;
  wire csa_tree_add_190_195_groupi_n_3448, csa_tree_add_190_195_groupi_n_3449, csa_tree_add_190_195_groupi_n_3450, csa_tree_add_190_195_groupi_n_3451, csa_tree_add_190_195_groupi_n_3452, csa_tree_add_190_195_groupi_n_3453, csa_tree_add_190_195_groupi_n_3454, csa_tree_add_190_195_groupi_n_3455;
  wire csa_tree_add_190_195_groupi_n_3456, csa_tree_add_190_195_groupi_n_3457, csa_tree_add_190_195_groupi_n_3458, csa_tree_add_190_195_groupi_n_3459, csa_tree_add_190_195_groupi_n_3460, csa_tree_add_190_195_groupi_n_3461, csa_tree_add_190_195_groupi_n_3462, csa_tree_add_190_195_groupi_n_3463;
  wire csa_tree_add_190_195_groupi_n_3464, csa_tree_add_190_195_groupi_n_3465, csa_tree_add_190_195_groupi_n_3466, csa_tree_add_190_195_groupi_n_3467, csa_tree_add_190_195_groupi_n_3468, csa_tree_add_190_195_groupi_n_3469, csa_tree_add_190_195_groupi_n_3470, csa_tree_add_190_195_groupi_n_3471;
  wire csa_tree_add_190_195_groupi_n_3472, csa_tree_add_190_195_groupi_n_3473, csa_tree_add_190_195_groupi_n_3474, csa_tree_add_190_195_groupi_n_3475, csa_tree_add_190_195_groupi_n_3476, csa_tree_add_190_195_groupi_n_3477, csa_tree_add_190_195_groupi_n_3478, csa_tree_add_190_195_groupi_n_3479;
  wire csa_tree_add_190_195_groupi_n_3480, csa_tree_add_190_195_groupi_n_3481, csa_tree_add_190_195_groupi_n_3482, csa_tree_add_190_195_groupi_n_3483, csa_tree_add_190_195_groupi_n_3484, csa_tree_add_190_195_groupi_n_3485, csa_tree_add_190_195_groupi_n_3486, csa_tree_add_190_195_groupi_n_3487;
  wire csa_tree_add_190_195_groupi_n_3488, csa_tree_add_190_195_groupi_n_3489, csa_tree_add_190_195_groupi_n_3490, csa_tree_add_190_195_groupi_n_3491, csa_tree_add_190_195_groupi_n_3492, csa_tree_add_190_195_groupi_n_3493, csa_tree_add_190_195_groupi_n_3494, csa_tree_add_190_195_groupi_n_3495;
  wire csa_tree_add_190_195_groupi_n_3496, csa_tree_add_190_195_groupi_n_3497, csa_tree_add_190_195_groupi_n_3498, csa_tree_add_190_195_groupi_n_3499, csa_tree_add_190_195_groupi_n_3500, csa_tree_add_190_195_groupi_n_3501, csa_tree_add_190_195_groupi_n_3502, csa_tree_add_190_195_groupi_n_3503;
  wire csa_tree_add_190_195_groupi_n_3504, csa_tree_add_190_195_groupi_n_3505, csa_tree_add_190_195_groupi_n_3506, csa_tree_add_190_195_groupi_n_3507, csa_tree_add_190_195_groupi_n_3508, csa_tree_add_190_195_groupi_n_3509, csa_tree_add_190_195_groupi_n_3510, csa_tree_add_190_195_groupi_n_3511;
  wire csa_tree_add_190_195_groupi_n_3512, csa_tree_add_190_195_groupi_n_3513, csa_tree_add_190_195_groupi_n_3514, csa_tree_add_190_195_groupi_n_3515, csa_tree_add_190_195_groupi_n_3516, csa_tree_add_190_195_groupi_n_3517, csa_tree_add_190_195_groupi_n_3518, csa_tree_add_190_195_groupi_n_3519;
  wire csa_tree_add_190_195_groupi_n_3520, csa_tree_add_190_195_groupi_n_3521, csa_tree_add_190_195_groupi_n_3522, csa_tree_add_190_195_groupi_n_3523, csa_tree_add_190_195_groupi_n_3524, csa_tree_add_190_195_groupi_n_3525, csa_tree_add_190_195_groupi_n_3526, csa_tree_add_190_195_groupi_n_3527;
  wire csa_tree_add_190_195_groupi_n_3528, csa_tree_add_190_195_groupi_n_3529, csa_tree_add_190_195_groupi_n_3530, csa_tree_add_190_195_groupi_n_3531, csa_tree_add_190_195_groupi_n_3532, csa_tree_add_190_195_groupi_n_3533, csa_tree_add_190_195_groupi_n_3534, csa_tree_add_190_195_groupi_n_3535;
  wire csa_tree_add_190_195_groupi_n_3536, csa_tree_add_190_195_groupi_n_3537, csa_tree_add_190_195_groupi_n_3538, csa_tree_add_190_195_groupi_n_3539, csa_tree_add_190_195_groupi_n_3540, csa_tree_add_190_195_groupi_n_3541, csa_tree_add_190_195_groupi_n_3542, csa_tree_add_190_195_groupi_n_3543;
  wire csa_tree_add_190_195_groupi_n_3544, csa_tree_add_190_195_groupi_n_3545, csa_tree_add_190_195_groupi_n_3546, csa_tree_add_190_195_groupi_n_3547, csa_tree_add_190_195_groupi_n_3548, csa_tree_add_190_195_groupi_n_3549, csa_tree_add_190_195_groupi_n_3550, csa_tree_add_190_195_groupi_n_3551;
  wire csa_tree_add_190_195_groupi_n_3552, csa_tree_add_190_195_groupi_n_3553, csa_tree_add_190_195_groupi_n_3554, csa_tree_add_190_195_groupi_n_3555, csa_tree_add_190_195_groupi_n_3556, csa_tree_add_190_195_groupi_n_3557, csa_tree_add_190_195_groupi_n_3558, csa_tree_add_190_195_groupi_n_3559;
  wire csa_tree_add_190_195_groupi_n_3560, csa_tree_add_190_195_groupi_n_3561, csa_tree_add_190_195_groupi_n_3562, csa_tree_add_190_195_groupi_n_3563, csa_tree_add_190_195_groupi_n_3564, csa_tree_add_190_195_groupi_n_3565, csa_tree_add_190_195_groupi_n_3566, csa_tree_add_190_195_groupi_n_3567;
  wire csa_tree_add_190_195_groupi_n_3568, csa_tree_add_190_195_groupi_n_3569, csa_tree_add_190_195_groupi_n_3570, csa_tree_add_190_195_groupi_n_3571, csa_tree_add_190_195_groupi_n_3572, csa_tree_add_190_195_groupi_n_3573, csa_tree_add_190_195_groupi_n_3574, csa_tree_add_190_195_groupi_n_3575;
  wire csa_tree_add_190_195_groupi_n_3576, csa_tree_add_190_195_groupi_n_3577, csa_tree_add_190_195_groupi_n_3578, csa_tree_add_190_195_groupi_n_3579, csa_tree_add_190_195_groupi_n_3580, csa_tree_add_190_195_groupi_n_3581, csa_tree_add_190_195_groupi_n_3582, csa_tree_add_190_195_groupi_n_3583;
  wire csa_tree_add_190_195_groupi_n_3584, csa_tree_add_190_195_groupi_n_3585, csa_tree_add_190_195_groupi_n_3586, csa_tree_add_190_195_groupi_n_3587, csa_tree_add_190_195_groupi_n_3588, csa_tree_add_190_195_groupi_n_3589, csa_tree_add_190_195_groupi_n_3590, csa_tree_add_190_195_groupi_n_3591;
  wire csa_tree_add_190_195_groupi_n_3592, csa_tree_add_190_195_groupi_n_3593, csa_tree_add_190_195_groupi_n_3594, csa_tree_add_190_195_groupi_n_3595, csa_tree_add_190_195_groupi_n_3596, csa_tree_add_190_195_groupi_n_3597, csa_tree_add_190_195_groupi_n_3598, csa_tree_add_190_195_groupi_n_3599;
  wire csa_tree_add_190_195_groupi_n_3600, csa_tree_add_190_195_groupi_n_3601, csa_tree_add_190_195_groupi_n_3602, csa_tree_add_190_195_groupi_n_3603, csa_tree_add_190_195_groupi_n_3604, csa_tree_add_190_195_groupi_n_3605, csa_tree_add_190_195_groupi_n_3606, csa_tree_add_190_195_groupi_n_3607;
  wire csa_tree_add_190_195_groupi_n_3608, csa_tree_add_190_195_groupi_n_3609, csa_tree_add_190_195_groupi_n_3610, csa_tree_add_190_195_groupi_n_3611, csa_tree_add_190_195_groupi_n_3612, csa_tree_add_190_195_groupi_n_3613, csa_tree_add_190_195_groupi_n_3614, csa_tree_add_190_195_groupi_n_3615;
  wire csa_tree_add_190_195_groupi_n_3616, csa_tree_add_190_195_groupi_n_3617, csa_tree_add_190_195_groupi_n_3618, csa_tree_add_190_195_groupi_n_3619, csa_tree_add_190_195_groupi_n_3620, csa_tree_add_190_195_groupi_n_3621, csa_tree_add_190_195_groupi_n_3622, csa_tree_add_190_195_groupi_n_3623;
  wire csa_tree_add_190_195_groupi_n_3624, csa_tree_add_190_195_groupi_n_3625, csa_tree_add_190_195_groupi_n_3626, csa_tree_add_190_195_groupi_n_3627, csa_tree_add_190_195_groupi_n_3628, csa_tree_add_190_195_groupi_n_3629, csa_tree_add_190_195_groupi_n_3630, csa_tree_add_190_195_groupi_n_3631;
  wire csa_tree_add_190_195_groupi_n_3632, csa_tree_add_190_195_groupi_n_3633, csa_tree_add_190_195_groupi_n_3634, csa_tree_add_190_195_groupi_n_3635, csa_tree_add_190_195_groupi_n_3636, csa_tree_add_190_195_groupi_n_3637, csa_tree_add_190_195_groupi_n_3638, csa_tree_add_190_195_groupi_n_3639;
  wire csa_tree_add_190_195_groupi_n_3640, csa_tree_add_190_195_groupi_n_3641, csa_tree_add_190_195_groupi_n_3642, csa_tree_add_190_195_groupi_n_3643, csa_tree_add_190_195_groupi_n_3644, csa_tree_add_190_195_groupi_n_3645, csa_tree_add_190_195_groupi_n_3646, csa_tree_add_190_195_groupi_n_3647;
  wire csa_tree_add_190_195_groupi_n_3648, csa_tree_add_190_195_groupi_n_3649, csa_tree_add_190_195_groupi_n_3650, csa_tree_add_190_195_groupi_n_3651, csa_tree_add_190_195_groupi_n_3652, csa_tree_add_190_195_groupi_n_3653, csa_tree_add_190_195_groupi_n_3654, csa_tree_add_190_195_groupi_n_3655;
  wire csa_tree_add_190_195_groupi_n_3656, csa_tree_add_190_195_groupi_n_3657, csa_tree_add_190_195_groupi_n_3658, csa_tree_add_190_195_groupi_n_3659, csa_tree_add_190_195_groupi_n_3660, csa_tree_add_190_195_groupi_n_3661, csa_tree_add_190_195_groupi_n_3662, csa_tree_add_190_195_groupi_n_3663;
  wire csa_tree_add_190_195_groupi_n_3664, csa_tree_add_190_195_groupi_n_3665, csa_tree_add_190_195_groupi_n_3666, csa_tree_add_190_195_groupi_n_3667, csa_tree_add_190_195_groupi_n_3668, csa_tree_add_190_195_groupi_n_3669, csa_tree_add_190_195_groupi_n_3670, csa_tree_add_190_195_groupi_n_3671;
  wire csa_tree_add_190_195_groupi_n_3672, csa_tree_add_190_195_groupi_n_3673, csa_tree_add_190_195_groupi_n_3674, csa_tree_add_190_195_groupi_n_3675, csa_tree_add_190_195_groupi_n_3676, csa_tree_add_190_195_groupi_n_3677, csa_tree_add_190_195_groupi_n_3678, csa_tree_add_190_195_groupi_n_3679;
  wire csa_tree_add_190_195_groupi_n_3680, csa_tree_add_190_195_groupi_n_3681, csa_tree_add_190_195_groupi_n_3682, csa_tree_add_190_195_groupi_n_3683, csa_tree_add_190_195_groupi_n_3684, csa_tree_add_190_195_groupi_n_3685, csa_tree_add_190_195_groupi_n_3686, csa_tree_add_190_195_groupi_n_3687;
  wire csa_tree_add_190_195_groupi_n_3688, csa_tree_add_190_195_groupi_n_3689, csa_tree_add_190_195_groupi_n_3690, csa_tree_add_190_195_groupi_n_3691, csa_tree_add_190_195_groupi_n_3692, csa_tree_add_190_195_groupi_n_3693, csa_tree_add_190_195_groupi_n_3694, csa_tree_add_190_195_groupi_n_3695;
  wire csa_tree_add_190_195_groupi_n_3696, csa_tree_add_190_195_groupi_n_3697, csa_tree_add_190_195_groupi_n_3698, csa_tree_add_190_195_groupi_n_3699, csa_tree_add_190_195_groupi_n_3700, csa_tree_add_190_195_groupi_n_3701, csa_tree_add_190_195_groupi_n_3702, csa_tree_add_190_195_groupi_n_3703;
  wire csa_tree_add_190_195_groupi_n_3704, csa_tree_add_190_195_groupi_n_3705, csa_tree_add_190_195_groupi_n_3706, csa_tree_add_190_195_groupi_n_3707, csa_tree_add_190_195_groupi_n_3708, csa_tree_add_190_195_groupi_n_3709, csa_tree_add_190_195_groupi_n_3710, csa_tree_add_190_195_groupi_n_3711;
  wire csa_tree_add_190_195_groupi_n_3712, csa_tree_add_190_195_groupi_n_3713, csa_tree_add_190_195_groupi_n_3714, csa_tree_add_190_195_groupi_n_3715, csa_tree_add_190_195_groupi_n_3716, csa_tree_add_190_195_groupi_n_3717, csa_tree_add_190_195_groupi_n_3718, csa_tree_add_190_195_groupi_n_3719;
  wire csa_tree_add_190_195_groupi_n_3720, csa_tree_add_190_195_groupi_n_3721, csa_tree_add_190_195_groupi_n_3722, csa_tree_add_190_195_groupi_n_3723, csa_tree_add_190_195_groupi_n_3724, csa_tree_add_190_195_groupi_n_3725, csa_tree_add_190_195_groupi_n_3726, csa_tree_add_190_195_groupi_n_3727;
  wire csa_tree_add_190_195_groupi_n_3728, csa_tree_add_190_195_groupi_n_3729, csa_tree_add_190_195_groupi_n_3730, csa_tree_add_190_195_groupi_n_3731, csa_tree_add_190_195_groupi_n_3732, csa_tree_add_190_195_groupi_n_3733, csa_tree_add_190_195_groupi_n_3734, csa_tree_add_190_195_groupi_n_3735;
  wire csa_tree_add_190_195_groupi_n_3736, csa_tree_add_190_195_groupi_n_3737, csa_tree_add_190_195_groupi_n_3738, csa_tree_add_190_195_groupi_n_3739, csa_tree_add_190_195_groupi_n_3740, csa_tree_add_190_195_groupi_n_3741, csa_tree_add_190_195_groupi_n_3742, csa_tree_add_190_195_groupi_n_3743;
  wire csa_tree_add_190_195_groupi_n_3744, csa_tree_add_190_195_groupi_n_3745, csa_tree_add_190_195_groupi_n_3746, csa_tree_add_190_195_groupi_n_3747, csa_tree_add_190_195_groupi_n_3748, csa_tree_add_190_195_groupi_n_3749, csa_tree_add_190_195_groupi_n_3750, csa_tree_add_190_195_groupi_n_3751;
  wire csa_tree_add_190_195_groupi_n_3752, csa_tree_add_190_195_groupi_n_3753, csa_tree_add_190_195_groupi_n_3754, csa_tree_add_190_195_groupi_n_3755, csa_tree_add_190_195_groupi_n_3756, csa_tree_add_190_195_groupi_n_3757, csa_tree_add_190_195_groupi_n_3758, csa_tree_add_190_195_groupi_n_3759;
  wire csa_tree_add_190_195_groupi_n_3760, csa_tree_add_190_195_groupi_n_3761, csa_tree_add_190_195_groupi_n_3762, csa_tree_add_190_195_groupi_n_3763, csa_tree_add_190_195_groupi_n_3764, csa_tree_add_190_195_groupi_n_3765, csa_tree_add_190_195_groupi_n_3766, csa_tree_add_190_195_groupi_n_3767;
  wire csa_tree_add_190_195_groupi_n_3768, csa_tree_add_190_195_groupi_n_3769, csa_tree_add_190_195_groupi_n_3770, csa_tree_add_190_195_groupi_n_3771, csa_tree_add_190_195_groupi_n_3772, csa_tree_add_190_195_groupi_n_3773, csa_tree_add_190_195_groupi_n_3774, csa_tree_add_190_195_groupi_n_3775;
  wire csa_tree_add_190_195_groupi_n_3776, csa_tree_add_190_195_groupi_n_3777, csa_tree_add_190_195_groupi_n_3778, csa_tree_add_190_195_groupi_n_3779, csa_tree_add_190_195_groupi_n_3780, csa_tree_add_190_195_groupi_n_3781, csa_tree_add_190_195_groupi_n_3782, csa_tree_add_190_195_groupi_n_3783;
  wire csa_tree_add_190_195_groupi_n_3784, csa_tree_add_190_195_groupi_n_3785, csa_tree_add_190_195_groupi_n_3786, csa_tree_add_190_195_groupi_n_3787, csa_tree_add_190_195_groupi_n_3788, csa_tree_add_190_195_groupi_n_3789, csa_tree_add_190_195_groupi_n_3790, csa_tree_add_190_195_groupi_n_3791;
  wire csa_tree_add_190_195_groupi_n_3792, csa_tree_add_190_195_groupi_n_3793, csa_tree_add_190_195_groupi_n_3794, csa_tree_add_190_195_groupi_n_3795, csa_tree_add_190_195_groupi_n_3796, csa_tree_add_190_195_groupi_n_3797, csa_tree_add_190_195_groupi_n_3798, csa_tree_add_190_195_groupi_n_3799;
  wire csa_tree_add_190_195_groupi_n_3800, csa_tree_add_190_195_groupi_n_3801, csa_tree_add_190_195_groupi_n_3802, csa_tree_add_190_195_groupi_n_3803, csa_tree_add_190_195_groupi_n_3804, csa_tree_add_190_195_groupi_n_3805, csa_tree_add_190_195_groupi_n_3806, csa_tree_add_190_195_groupi_n_3807;
  wire csa_tree_add_190_195_groupi_n_3808, csa_tree_add_190_195_groupi_n_3809, csa_tree_add_190_195_groupi_n_3810, csa_tree_add_190_195_groupi_n_3811, csa_tree_add_190_195_groupi_n_3812, csa_tree_add_190_195_groupi_n_3813, csa_tree_add_190_195_groupi_n_3814, csa_tree_add_190_195_groupi_n_3815;
  wire csa_tree_add_190_195_groupi_n_3816, csa_tree_add_190_195_groupi_n_3817, csa_tree_add_190_195_groupi_n_3818, csa_tree_add_190_195_groupi_n_3819, csa_tree_add_190_195_groupi_n_3820, csa_tree_add_190_195_groupi_n_3821, csa_tree_add_190_195_groupi_n_3822, csa_tree_add_190_195_groupi_n_3823;
  wire csa_tree_add_190_195_groupi_n_3824, csa_tree_add_190_195_groupi_n_3825, csa_tree_add_190_195_groupi_n_3826, csa_tree_add_190_195_groupi_n_3827, csa_tree_add_190_195_groupi_n_3828, csa_tree_add_190_195_groupi_n_3829, csa_tree_add_190_195_groupi_n_3830, csa_tree_add_190_195_groupi_n_3831;
  wire csa_tree_add_190_195_groupi_n_3832, csa_tree_add_190_195_groupi_n_3833, csa_tree_add_190_195_groupi_n_3834, csa_tree_add_190_195_groupi_n_3835, csa_tree_add_190_195_groupi_n_3836, csa_tree_add_190_195_groupi_n_3837, csa_tree_add_190_195_groupi_n_3838, csa_tree_add_190_195_groupi_n_3839;
  wire csa_tree_add_190_195_groupi_n_3840, csa_tree_add_190_195_groupi_n_3841, csa_tree_add_190_195_groupi_n_3842, csa_tree_add_190_195_groupi_n_3843, csa_tree_add_190_195_groupi_n_3844, csa_tree_add_190_195_groupi_n_3845, csa_tree_add_190_195_groupi_n_3846, csa_tree_add_190_195_groupi_n_3847;
  wire csa_tree_add_190_195_groupi_n_3848, csa_tree_add_190_195_groupi_n_3849, csa_tree_add_190_195_groupi_n_3850, csa_tree_add_190_195_groupi_n_3851, csa_tree_add_190_195_groupi_n_3852, csa_tree_add_190_195_groupi_n_3853, csa_tree_add_190_195_groupi_n_3854, csa_tree_add_190_195_groupi_n_3855;
  wire csa_tree_add_190_195_groupi_n_3856, csa_tree_add_190_195_groupi_n_3857, csa_tree_add_190_195_groupi_n_3858, csa_tree_add_190_195_groupi_n_3859, csa_tree_add_190_195_groupi_n_3860, csa_tree_add_190_195_groupi_n_3861, csa_tree_add_190_195_groupi_n_3862, csa_tree_add_190_195_groupi_n_3863;
  wire csa_tree_add_190_195_groupi_n_3864, csa_tree_add_190_195_groupi_n_3865, csa_tree_add_190_195_groupi_n_3866, csa_tree_add_190_195_groupi_n_3867, csa_tree_add_190_195_groupi_n_3868, csa_tree_add_190_195_groupi_n_3869, csa_tree_add_190_195_groupi_n_3870, csa_tree_add_190_195_groupi_n_3871;
  wire csa_tree_add_190_195_groupi_n_3872, csa_tree_add_190_195_groupi_n_3873, csa_tree_add_190_195_groupi_n_3874, csa_tree_add_190_195_groupi_n_3875, csa_tree_add_190_195_groupi_n_3876, csa_tree_add_190_195_groupi_n_3877, csa_tree_add_190_195_groupi_n_3878, csa_tree_add_190_195_groupi_n_3879;
  wire csa_tree_add_190_195_groupi_n_3880, csa_tree_add_190_195_groupi_n_3881, csa_tree_add_190_195_groupi_n_3882, csa_tree_add_190_195_groupi_n_3883, csa_tree_add_190_195_groupi_n_3884, csa_tree_add_190_195_groupi_n_3885, csa_tree_add_190_195_groupi_n_3886, csa_tree_add_190_195_groupi_n_3887;
  wire csa_tree_add_190_195_groupi_n_3888, csa_tree_add_190_195_groupi_n_3889, csa_tree_add_190_195_groupi_n_3890, csa_tree_add_190_195_groupi_n_3891, csa_tree_add_190_195_groupi_n_3892, csa_tree_add_190_195_groupi_n_3893, csa_tree_add_190_195_groupi_n_3894, csa_tree_add_190_195_groupi_n_3895;
  wire csa_tree_add_190_195_groupi_n_3896, csa_tree_add_190_195_groupi_n_3897, csa_tree_add_190_195_groupi_n_3898, csa_tree_add_190_195_groupi_n_3899, csa_tree_add_190_195_groupi_n_3900, csa_tree_add_190_195_groupi_n_3901, csa_tree_add_190_195_groupi_n_3902, csa_tree_add_190_195_groupi_n_3903;
  wire csa_tree_add_190_195_groupi_n_3904, csa_tree_add_190_195_groupi_n_3905, csa_tree_add_190_195_groupi_n_3906, csa_tree_add_190_195_groupi_n_3907, csa_tree_add_190_195_groupi_n_3908, csa_tree_add_190_195_groupi_n_3909, csa_tree_add_190_195_groupi_n_3910, csa_tree_add_190_195_groupi_n_3911;
  wire csa_tree_add_190_195_groupi_n_3912, csa_tree_add_190_195_groupi_n_3913, csa_tree_add_190_195_groupi_n_3914, csa_tree_add_190_195_groupi_n_3915, csa_tree_add_190_195_groupi_n_3916, csa_tree_add_190_195_groupi_n_3917, csa_tree_add_190_195_groupi_n_3918, csa_tree_add_190_195_groupi_n_3919;
  wire csa_tree_add_190_195_groupi_n_3920, csa_tree_add_190_195_groupi_n_3921, csa_tree_add_190_195_groupi_n_3922, csa_tree_add_190_195_groupi_n_3923, csa_tree_add_190_195_groupi_n_3924, csa_tree_add_190_195_groupi_n_3925, csa_tree_add_190_195_groupi_n_3926, csa_tree_add_190_195_groupi_n_3927;
  wire csa_tree_add_190_195_groupi_n_3928, csa_tree_add_190_195_groupi_n_3929, csa_tree_add_190_195_groupi_n_3930, csa_tree_add_190_195_groupi_n_3931, csa_tree_add_190_195_groupi_n_3932, csa_tree_add_190_195_groupi_n_3933, csa_tree_add_190_195_groupi_n_3934, csa_tree_add_190_195_groupi_n_3935;
  wire csa_tree_add_190_195_groupi_n_3936, csa_tree_add_190_195_groupi_n_3937, csa_tree_add_190_195_groupi_n_3938, csa_tree_add_190_195_groupi_n_3939, csa_tree_add_190_195_groupi_n_3940, csa_tree_add_190_195_groupi_n_3941, csa_tree_add_190_195_groupi_n_3942, csa_tree_add_190_195_groupi_n_3943;
  wire csa_tree_add_190_195_groupi_n_3944, csa_tree_add_190_195_groupi_n_3945, csa_tree_add_190_195_groupi_n_3946, csa_tree_add_190_195_groupi_n_3947, csa_tree_add_190_195_groupi_n_3948, csa_tree_add_190_195_groupi_n_3949, csa_tree_add_190_195_groupi_n_3950, csa_tree_add_190_195_groupi_n_3951;
  wire csa_tree_add_190_195_groupi_n_3952, csa_tree_add_190_195_groupi_n_3953, csa_tree_add_190_195_groupi_n_3954, csa_tree_add_190_195_groupi_n_3955, csa_tree_add_190_195_groupi_n_3956, csa_tree_add_190_195_groupi_n_3957, csa_tree_add_190_195_groupi_n_3958, csa_tree_add_190_195_groupi_n_3959;
  wire csa_tree_add_190_195_groupi_n_3960, csa_tree_add_190_195_groupi_n_3961, csa_tree_add_190_195_groupi_n_3962, csa_tree_add_190_195_groupi_n_3963, csa_tree_add_190_195_groupi_n_3964, csa_tree_add_190_195_groupi_n_3965, csa_tree_add_190_195_groupi_n_3966, csa_tree_add_190_195_groupi_n_3967;
  wire csa_tree_add_190_195_groupi_n_3968, csa_tree_add_190_195_groupi_n_3969, csa_tree_add_190_195_groupi_n_3970, csa_tree_add_190_195_groupi_n_3971, csa_tree_add_190_195_groupi_n_3972, csa_tree_add_190_195_groupi_n_3973, csa_tree_add_190_195_groupi_n_3974, csa_tree_add_190_195_groupi_n_3975;
  wire csa_tree_add_190_195_groupi_n_3976, csa_tree_add_190_195_groupi_n_3977, csa_tree_add_190_195_groupi_n_3978, csa_tree_add_190_195_groupi_n_3979, csa_tree_add_190_195_groupi_n_3980, csa_tree_add_190_195_groupi_n_3981, csa_tree_add_190_195_groupi_n_3982, csa_tree_add_190_195_groupi_n_3983;
  wire csa_tree_add_190_195_groupi_n_3984, csa_tree_add_190_195_groupi_n_3985, csa_tree_add_190_195_groupi_n_3986, csa_tree_add_190_195_groupi_n_3987, csa_tree_add_190_195_groupi_n_3988, csa_tree_add_190_195_groupi_n_3989, csa_tree_add_190_195_groupi_n_3990, csa_tree_add_190_195_groupi_n_3991;
  wire csa_tree_add_190_195_groupi_n_3992, csa_tree_add_190_195_groupi_n_3993, csa_tree_add_190_195_groupi_n_3994, csa_tree_add_190_195_groupi_n_3995, csa_tree_add_190_195_groupi_n_3996, csa_tree_add_190_195_groupi_n_3997, csa_tree_add_190_195_groupi_n_3998, csa_tree_add_190_195_groupi_n_3999;
  wire csa_tree_add_190_195_groupi_n_4000, csa_tree_add_190_195_groupi_n_4001, csa_tree_add_190_195_groupi_n_4002, csa_tree_add_190_195_groupi_n_4003, csa_tree_add_190_195_groupi_n_4004, csa_tree_add_190_195_groupi_n_4005, csa_tree_add_190_195_groupi_n_4006, csa_tree_add_190_195_groupi_n_4007;
  wire csa_tree_add_190_195_groupi_n_4008, csa_tree_add_190_195_groupi_n_4009, csa_tree_add_190_195_groupi_n_4010, csa_tree_add_190_195_groupi_n_4011, csa_tree_add_190_195_groupi_n_4012, csa_tree_add_190_195_groupi_n_4013, csa_tree_add_190_195_groupi_n_4014, csa_tree_add_190_195_groupi_n_4015;
  wire csa_tree_add_190_195_groupi_n_4016, csa_tree_add_190_195_groupi_n_4017, csa_tree_add_190_195_groupi_n_4018, csa_tree_add_190_195_groupi_n_4019, csa_tree_add_190_195_groupi_n_4020, csa_tree_add_190_195_groupi_n_4021, csa_tree_add_190_195_groupi_n_4022, csa_tree_add_190_195_groupi_n_4023;
  wire csa_tree_add_190_195_groupi_n_4024, csa_tree_add_190_195_groupi_n_4025, csa_tree_add_190_195_groupi_n_4026, csa_tree_add_190_195_groupi_n_4027, csa_tree_add_190_195_groupi_n_4028, csa_tree_add_190_195_groupi_n_4029, csa_tree_add_190_195_groupi_n_4030, csa_tree_add_190_195_groupi_n_4031;
  wire csa_tree_add_190_195_groupi_n_4032, csa_tree_add_190_195_groupi_n_4033, csa_tree_add_190_195_groupi_n_4034, csa_tree_add_190_195_groupi_n_4035, csa_tree_add_190_195_groupi_n_4036, csa_tree_add_190_195_groupi_n_4037, csa_tree_add_190_195_groupi_n_4038, csa_tree_add_190_195_groupi_n_4039;
  wire csa_tree_add_190_195_groupi_n_4040, csa_tree_add_190_195_groupi_n_4041, csa_tree_add_190_195_groupi_n_4042, csa_tree_add_190_195_groupi_n_4043, csa_tree_add_190_195_groupi_n_4044, csa_tree_add_190_195_groupi_n_4045, csa_tree_add_190_195_groupi_n_4046, csa_tree_add_190_195_groupi_n_4047;
  wire csa_tree_add_190_195_groupi_n_4048, csa_tree_add_190_195_groupi_n_4049, csa_tree_add_190_195_groupi_n_4050, csa_tree_add_190_195_groupi_n_4051, csa_tree_add_190_195_groupi_n_4052, csa_tree_add_190_195_groupi_n_4053, csa_tree_add_190_195_groupi_n_4054, csa_tree_add_190_195_groupi_n_4055;
  wire csa_tree_add_190_195_groupi_n_4056, csa_tree_add_190_195_groupi_n_4057, csa_tree_add_190_195_groupi_n_4058, csa_tree_add_190_195_groupi_n_4059, csa_tree_add_190_195_groupi_n_4060, csa_tree_add_190_195_groupi_n_4061, csa_tree_add_190_195_groupi_n_4062, csa_tree_add_190_195_groupi_n_4063;
  wire csa_tree_add_190_195_groupi_n_4064, csa_tree_add_190_195_groupi_n_4065, csa_tree_add_190_195_groupi_n_4066, csa_tree_add_190_195_groupi_n_4067, csa_tree_add_190_195_groupi_n_4068, csa_tree_add_190_195_groupi_n_4069, csa_tree_add_190_195_groupi_n_4070, csa_tree_add_190_195_groupi_n_4071;
  wire csa_tree_add_190_195_groupi_n_4072, csa_tree_add_190_195_groupi_n_4073, csa_tree_add_190_195_groupi_n_4074, csa_tree_add_190_195_groupi_n_4075, csa_tree_add_190_195_groupi_n_4076, csa_tree_add_190_195_groupi_n_4077, csa_tree_add_190_195_groupi_n_4078, csa_tree_add_190_195_groupi_n_4079;
  wire csa_tree_add_190_195_groupi_n_4080, csa_tree_add_190_195_groupi_n_4081, csa_tree_add_190_195_groupi_n_4082, csa_tree_add_190_195_groupi_n_4083, csa_tree_add_190_195_groupi_n_4084, csa_tree_add_190_195_groupi_n_4085, csa_tree_add_190_195_groupi_n_4086, csa_tree_add_190_195_groupi_n_4087;
  wire csa_tree_add_190_195_groupi_n_4088, csa_tree_add_190_195_groupi_n_4089, csa_tree_add_190_195_groupi_n_4090, csa_tree_add_190_195_groupi_n_4091, csa_tree_add_190_195_groupi_n_4092, csa_tree_add_190_195_groupi_n_4093, csa_tree_add_190_195_groupi_n_4094, csa_tree_add_190_195_groupi_n_4095;
  wire csa_tree_add_190_195_groupi_n_4096, csa_tree_add_190_195_groupi_n_4097, csa_tree_add_190_195_groupi_n_4098, csa_tree_add_190_195_groupi_n_4099, csa_tree_add_190_195_groupi_n_4100, csa_tree_add_190_195_groupi_n_4101, csa_tree_add_190_195_groupi_n_4102, csa_tree_add_190_195_groupi_n_4103;
  wire csa_tree_add_190_195_groupi_n_4104, csa_tree_add_190_195_groupi_n_4105, csa_tree_add_190_195_groupi_n_4106, csa_tree_add_190_195_groupi_n_4107, csa_tree_add_190_195_groupi_n_4108, csa_tree_add_190_195_groupi_n_4109, csa_tree_add_190_195_groupi_n_4110, csa_tree_add_190_195_groupi_n_4111;
  wire csa_tree_add_190_195_groupi_n_4112, csa_tree_add_190_195_groupi_n_4113, csa_tree_add_190_195_groupi_n_4114, csa_tree_add_190_195_groupi_n_4115, csa_tree_add_190_195_groupi_n_4116, csa_tree_add_190_195_groupi_n_4117, csa_tree_add_190_195_groupi_n_4118, csa_tree_add_190_195_groupi_n_4119;
  wire csa_tree_add_190_195_groupi_n_4120, csa_tree_add_190_195_groupi_n_4121, csa_tree_add_190_195_groupi_n_4122, csa_tree_add_190_195_groupi_n_4123, csa_tree_add_190_195_groupi_n_4124, csa_tree_add_190_195_groupi_n_4125, csa_tree_add_190_195_groupi_n_4126, csa_tree_add_190_195_groupi_n_4127;
  wire csa_tree_add_190_195_groupi_n_4128, csa_tree_add_190_195_groupi_n_4129, csa_tree_add_190_195_groupi_n_4130, csa_tree_add_190_195_groupi_n_4131, csa_tree_add_190_195_groupi_n_4132, csa_tree_add_190_195_groupi_n_4133, csa_tree_add_190_195_groupi_n_4134, csa_tree_add_190_195_groupi_n_4135;
  wire csa_tree_add_190_195_groupi_n_4136, csa_tree_add_190_195_groupi_n_4137, csa_tree_add_190_195_groupi_n_4138, csa_tree_add_190_195_groupi_n_4139, csa_tree_add_190_195_groupi_n_4140, csa_tree_add_190_195_groupi_n_4141, csa_tree_add_190_195_groupi_n_4142, csa_tree_add_190_195_groupi_n_4143;
  wire csa_tree_add_190_195_groupi_n_4144, csa_tree_add_190_195_groupi_n_4145, csa_tree_add_190_195_groupi_n_4146, csa_tree_add_190_195_groupi_n_4147, csa_tree_add_190_195_groupi_n_4148, csa_tree_add_190_195_groupi_n_4149, csa_tree_add_190_195_groupi_n_4150, csa_tree_add_190_195_groupi_n_4151;
  wire csa_tree_add_190_195_groupi_n_4152, csa_tree_add_190_195_groupi_n_4153, csa_tree_add_190_195_groupi_n_4154, csa_tree_add_190_195_groupi_n_4155, csa_tree_add_190_195_groupi_n_4156, csa_tree_add_190_195_groupi_n_4157, csa_tree_add_190_195_groupi_n_4158, csa_tree_add_190_195_groupi_n_4159;
  wire csa_tree_add_190_195_groupi_n_4160, csa_tree_add_190_195_groupi_n_4161, csa_tree_add_190_195_groupi_n_4162, csa_tree_add_190_195_groupi_n_4163, csa_tree_add_190_195_groupi_n_4164, csa_tree_add_190_195_groupi_n_4165, csa_tree_add_190_195_groupi_n_4166, csa_tree_add_190_195_groupi_n_4167;
  wire csa_tree_add_190_195_groupi_n_4168, csa_tree_add_190_195_groupi_n_4169, csa_tree_add_190_195_groupi_n_4170, csa_tree_add_190_195_groupi_n_4171, csa_tree_add_190_195_groupi_n_4172, csa_tree_add_190_195_groupi_n_4173, csa_tree_add_190_195_groupi_n_4174, csa_tree_add_190_195_groupi_n_4175;
  wire csa_tree_add_190_195_groupi_n_4176, csa_tree_add_190_195_groupi_n_4177, csa_tree_add_190_195_groupi_n_4178, csa_tree_add_190_195_groupi_n_4179, csa_tree_add_190_195_groupi_n_4180, csa_tree_add_190_195_groupi_n_4181, csa_tree_add_190_195_groupi_n_4182, csa_tree_add_190_195_groupi_n_4183;
  wire csa_tree_add_190_195_groupi_n_4184, csa_tree_add_190_195_groupi_n_4185, csa_tree_add_190_195_groupi_n_4186, csa_tree_add_190_195_groupi_n_4187, csa_tree_add_190_195_groupi_n_4188, csa_tree_add_190_195_groupi_n_4189, csa_tree_add_190_195_groupi_n_4190, csa_tree_add_190_195_groupi_n_4191;
  wire csa_tree_add_190_195_groupi_n_4192, csa_tree_add_190_195_groupi_n_4193, csa_tree_add_190_195_groupi_n_4194, csa_tree_add_190_195_groupi_n_4195, csa_tree_add_190_195_groupi_n_4196, csa_tree_add_190_195_groupi_n_4197, csa_tree_add_190_195_groupi_n_4198, csa_tree_add_190_195_groupi_n_4199;
  wire csa_tree_add_190_195_groupi_n_4200, csa_tree_add_190_195_groupi_n_4201, csa_tree_add_190_195_groupi_n_4202, csa_tree_add_190_195_groupi_n_4203, csa_tree_add_190_195_groupi_n_4204, csa_tree_add_190_195_groupi_n_4205, csa_tree_add_190_195_groupi_n_4206, csa_tree_add_190_195_groupi_n_4207;
  wire csa_tree_add_190_195_groupi_n_4208, csa_tree_add_190_195_groupi_n_4209, csa_tree_add_190_195_groupi_n_4210, csa_tree_add_190_195_groupi_n_4211, csa_tree_add_190_195_groupi_n_4212, csa_tree_add_190_195_groupi_n_4213, csa_tree_add_190_195_groupi_n_4214, csa_tree_add_190_195_groupi_n_4215;
  wire csa_tree_add_190_195_groupi_n_4216, csa_tree_add_190_195_groupi_n_4217, csa_tree_add_190_195_groupi_n_4218, csa_tree_add_190_195_groupi_n_4219, csa_tree_add_190_195_groupi_n_4220, csa_tree_add_190_195_groupi_n_4221, csa_tree_add_190_195_groupi_n_4222, csa_tree_add_190_195_groupi_n_4223;
  wire csa_tree_add_190_195_groupi_n_4224, csa_tree_add_190_195_groupi_n_4225, csa_tree_add_190_195_groupi_n_4226, csa_tree_add_190_195_groupi_n_4227, csa_tree_add_190_195_groupi_n_4228, csa_tree_add_190_195_groupi_n_4229, csa_tree_add_190_195_groupi_n_4230, csa_tree_add_190_195_groupi_n_4231;
  wire csa_tree_add_190_195_groupi_n_4232, csa_tree_add_190_195_groupi_n_4233, csa_tree_add_190_195_groupi_n_4234, csa_tree_add_190_195_groupi_n_4235, csa_tree_add_190_195_groupi_n_4236, csa_tree_add_190_195_groupi_n_4237, csa_tree_add_190_195_groupi_n_4238, csa_tree_add_190_195_groupi_n_4239;
  wire csa_tree_add_190_195_groupi_n_4240, csa_tree_add_190_195_groupi_n_4241, csa_tree_add_190_195_groupi_n_4242, csa_tree_add_190_195_groupi_n_4243, csa_tree_add_190_195_groupi_n_4244, csa_tree_add_190_195_groupi_n_4245, csa_tree_add_190_195_groupi_n_4246, csa_tree_add_190_195_groupi_n_4247;
  wire csa_tree_add_190_195_groupi_n_4248, csa_tree_add_190_195_groupi_n_4249, csa_tree_add_190_195_groupi_n_4250, csa_tree_add_190_195_groupi_n_4251, csa_tree_add_190_195_groupi_n_4252, csa_tree_add_190_195_groupi_n_4253, csa_tree_add_190_195_groupi_n_4254, csa_tree_add_190_195_groupi_n_4255;
  wire csa_tree_add_190_195_groupi_n_4256, csa_tree_add_190_195_groupi_n_4257, csa_tree_add_190_195_groupi_n_4258, csa_tree_add_190_195_groupi_n_4259, csa_tree_add_190_195_groupi_n_4260, csa_tree_add_190_195_groupi_n_4261, csa_tree_add_190_195_groupi_n_4262, csa_tree_add_190_195_groupi_n_4263;
  wire csa_tree_add_190_195_groupi_n_4264, csa_tree_add_190_195_groupi_n_4265, csa_tree_add_190_195_groupi_n_4266, csa_tree_add_190_195_groupi_n_4267, csa_tree_add_190_195_groupi_n_4268, csa_tree_add_190_195_groupi_n_4269, csa_tree_add_190_195_groupi_n_4270, csa_tree_add_190_195_groupi_n_4271;
  wire csa_tree_add_190_195_groupi_n_4272, csa_tree_add_190_195_groupi_n_4273, csa_tree_add_190_195_groupi_n_4274, csa_tree_add_190_195_groupi_n_4275, csa_tree_add_190_195_groupi_n_4276, csa_tree_add_190_195_groupi_n_4277, csa_tree_add_190_195_groupi_n_4278, csa_tree_add_190_195_groupi_n_4279;
  wire csa_tree_add_190_195_groupi_n_4280, csa_tree_add_190_195_groupi_n_4281, csa_tree_add_190_195_groupi_n_4282, csa_tree_add_190_195_groupi_n_4283, csa_tree_add_190_195_groupi_n_4284, csa_tree_add_190_195_groupi_n_4285, csa_tree_add_190_195_groupi_n_4286, csa_tree_add_190_195_groupi_n_4287;
  wire csa_tree_add_190_195_groupi_n_4288, csa_tree_add_190_195_groupi_n_4289, csa_tree_add_190_195_groupi_n_4290, csa_tree_add_190_195_groupi_n_4291, csa_tree_add_190_195_groupi_n_4292, csa_tree_add_190_195_groupi_n_4293, csa_tree_add_190_195_groupi_n_4294, csa_tree_add_190_195_groupi_n_4295;
  wire csa_tree_add_190_195_groupi_n_4296, csa_tree_add_190_195_groupi_n_4297, csa_tree_add_190_195_groupi_n_4298, csa_tree_add_190_195_groupi_n_4299, csa_tree_add_190_195_groupi_n_4300, csa_tree_add_190_195_groupi_n_4301, csa_tree_add_190_195_groupi_n_4302, csa_tree_add_190_195_groupi_n_4303;
  wire csa_tree_add_190_195_groupi_n_4304, csa_tree_add_190_195_groupi_n_4305, csa_tree_add_190_195_groupi_n_4306, csa_tree_add_190_195_groupi_n_4307, csa_tree_add_190_195_groupi_n_4308, csa_tree_add_190_195_groupi_n_4309, csa_tree_add_190_195_groupi_n_4310, csa_tree_add_190_195_groupi_n_4311;
  wire csa_tree_add_190_195_groupi_n_4312, csa_tree_add_190_195_groupi_n_4313, csa_tree_add_190_195_groupi_n_4314, csa_tree_add_190_195_groupi_n_4315, csa_tree_add_190_195_groupi_n_4316, csa_tree_add_190_195_groupi_n_4317, csa_tree_add_190_195_groupi_n_4318, csa_tree_add_190_195_groupi_n_4319;
  wire csa_tree_add_190_195_groupi_n_4320, csa_tree_add_190_195_groupi_n_4321, csa_tree_add_190_195_groupi_n_4322, csa_tree_add_190_195_groupi_n_4323, csa_tree_add_190_195_groupi_n_4324, csa_tree_add_190_195_groupi_n_4325, csa_tree_add_190_195_groupi_n_4326, csa_tree_add_190_195_groupi_n_4327;
  wire csa_tree_add_190_195_groupi_n_4328, csa_tree_add_190_195_groupi_n_4329, csa_tree_add_190_195_groupi_n_4330, csa_tree_add_190_195_groupi_n_4331, csa_tree_add_190_195_groupi_n_4332, csa_tree_add_190_195_groupi_n_4333, csa_tree_add_190_195_groupi_n_4334, csa_tree_add_190_195_groupi_n_4335;
  wire csa_tree_add_190_195_groupi_n_4336, csa_tree_add_190_195_groupi_n_4337, csa_tree_add_190_195_groupi_n_4338, csa_tree_add_190_195_groupi_n_4339, csa_tree_add_190_195_groupi_n_4340, csa_tree_add_190_195_groupi_n_4341, csa_tree_add_190_195_groupi_n_4342, csa_tree_add_190_195_groupi_n_4343;
  wire csa_tree_add_190_195_groupi_n_4344, csa_tree_add_190_195_groupi_n_4345, csa_tree_add_190_195_groupi_n_4346, csa_tree_add_190_195_groupi_n_4347, csa_tree_add_190_195_groupi_n_4348, csa_tree_add_190_195_groupi_n_4349, csa_tree_add_190_195_groupi_n_4350, csa_tree_add_190_195_groupi_n_4351;
  wire csa_tree_add_190_195_groupi_n_4352, csa_tree_add_190_195_groupi_n_4353, csa_tree_add_190_195_groupi_n_4354, csa_tree_add_190_195_groupi_n_4355, csa_tree_add_190_195_groupi_n_4356, csa_tree_add_190_195_groupi_n_4357, csa_tree_add_190_195_groupi_n_4358, csa_tree_add_190_195_groupi_n_4359;
  wire csa_tree_add_190_195_groupi_n_4360, csa_tree_add_190_195_groupi_n_4361, csa_tree_add_190_195_groupi_n_4362, csa_tree_add_190_195_groupi_n_4363, csa_tree_add_190_195_groupi_n_4364, csa_tree_add_190_195_groupi_n_4365, csa_tree_add_190_195_groupi_n_4366, csa_tree_add_190_195_groupi_n_4367;
  wire csa_tree_add_190_195_groupi_n_4368, csa_tree_add_190_195_groupi_n_4369, csa_tree_add_190_195_groupi_n_4370, csa_tree_add_190_195_groupi_n_4371, csa_tree_add_190_195_groupi_n_4372, csa_tree_add_190_195_groupi_n_4373, csa_tree_add_190_195_groupi_n_4374, csa_tree_add_190_195_groupi_n_4375;
  wire csa_tree_add_190_195_groupi_n_4376, csa_tree_add_190_195_groupi_n_4377, csa_tree_add_190_195_groupi_n_4378, csa_tree_add_190_195_groupi_n_4379, csa_tree_add_190_195_groupi_n_4380, csa_tree_add_190_195_groupi_n_4381, csa_tree_add_190_195_groupi_n_4382, csa_tree_add_190_195_groupi_n_4383;
  wire csa_tree_add_190_195_groupi_n_4384, csa_tree_add_190_195_groupi_n_4385, csa_tree_add_190_195_groupi_n_4386, csa_tree_add_190_195_groupi_n_4387, csa_tree_add_190_195_groupi_n_4388, csa_tree_add_190_195_groupi_n_4389, csa_tree_add_190_195_groupi_n_4390, csa_tree_add_190_195_groupi_n_4391;
  wire csa_tree_add_190_195_groupi_n_4392, csa_tree_add_190_195_groupi_n_4393, csa_tree_add_190_195_groupi_n_4394, csa_tree_add_190_195_groupi_n_4395, csa_tree_add_190_195_groupi_n_4396, csa_tree_add_190_195_groupi_n_4397, csa_tree_add_190_195_groupi_n_4398, csa_tree_add_190_195_groupi_n_4399;
  wire csa_tree_add_190_195_groupi_n_4400, csa_tree_add_190_195_groupi_n_4401, csa_tree_add_190_195_groupi_n_4402, csa_tree_add_190_195_groupi_n_4403, csa_tree_add_190_195_groupi_n_4404, csa_tree_add_190_195_groupi_n_4405, csa_tree_add_190_195_groupi_n_4406, csa_tree_add_190_195_groupi_n_4407;
  wire csa_tree_add_190_195_groupi_n_4408, csa_tree_add_190_195_groupi_n_4409, csa_tree_add_190_195_groupi_n_4410, csa_tree_add_190_195_groupi_n_4411, csa_tree_add_190_195_groupi_n_4412, csa_tree_add_190_195_groupi_n_4413, csa_tree_add_190_195_groupi_n_4414, csa_tree_add_190_195_groupi_n_4415;
  wire csa_tree_add_190_195_groupi_n_4416, csa_tree_add_190_195_groupi_n_4417, csa_tree_add_190_195_groupi_n_4418, csa_tree_add_190_195_groupi_n_4419, csa_tree_add_190_195_groupi_n_4420, csa_tree_add_190_195_groupi_n_4421, csa_tree_add_190_195_groupi_n_4422, csa_tree_add_190_195_groupi_n_4423;
  wire csa_tree_add_190_195_groupi_n_4424, csa_tree_add_190_195_groupi_n_4425, csa_tree_add_190_195_groupi_n_4426, csa_tree_add_190_195_groupi_n_4427, csa_tree_add_190_195_groupi_n_4428, csa_tree_add_190_195_groupi_n_4429, csa_tree_add_190_195_groupi_n_4430, csa_tree_add_190_195_groupi_n_4431;
  wire csa_tree_add_190_195_groupi_n_4432, csa_tree_add_190_195_groupi_n_4433, csa_tree_add_190_195_groupi_n_4434, csa_tree_add_190_195_groupi_n_4435, csa_tree_add_190_195_groupi_n_4436, csa_tree_add_190_195_groupi_n_4437, csa_tree_add_190_195_groupi_n_4438, csa_tree_add_190_195_groupi_n_4439;
  wire csa_tree_add_190_195_groupi_n_4440, csa_tree_add_190_195_groupi_n_4441, csa_tree_add_190_195_groupi_n_4442, csa_tree_add_190_195_groupi_n_4443, csa_tree_add_190_195_groupi_n_4444, csa_tree_add_190_195_groupi_n_4445, csa_tree_add_190_195_groupi_n_4446, csa_tree_add_190_195_groupi_n_4447;
  wire csa_tree_add_190_195_groupi_n_4448, csa_tree_add_190_195_groupi_n_4449, csa_tree_add_190_195_groupi_n_4450, csa_tree_add_190_195_groupi_n_4451, csa_tree_add_190_195_groupi_n_4452, csa_tree_add_190_195_groupi_n_4453, csa_tree_add_190_195_groupi_n_4454, csa_tree_add_190_195_groupi_n_4455;
  wire csa_tree_add_190_195_groupi_n_4456, csa_tree_add_190_195_groupi_n_4457, csa_tree_add_190_195_groupi_n_4458, csa_tree_add_190_195_groupi_n_4459, csa_tree_add_190_195_groupi_n_4460, csa_tree_add_190_195_groupi_n_4461, csa_tree_add_190_195_groupi_n_4462, csa_tree_add_190_195_groupi_n_4463;
  wire csa_tree_add_190_195_groupi_n_4464, csa_tree_add_190_195_groupi_n_4465, csa_tree_add_190_195_groupi_n_4466, csa_tree_add_190_195_groupi_n_4467, csa_tree_add_190_195_groupi_n_4468, csa_tree_add_190_195_groupi_n_4469, csa_tree_add_190_195_groupi_n_4470, csa_tree_add_190_195_groupi_n_4471;
  wire csa_tree_add_190_195_groupi_n_4472, csa_tree_add_190_195_groupi_n_4473, csa_tree_add_190_195_groupi_n_4474, csa_tree_add_190_195_groupi_n_4475, csa_tree_add_190_195_groupi_n_4476, csa_tree_add_190_195_groupi_n_4477, csa_tree_add_190_195_groupi_n_4478, csa_tree_add_190_195_groupi_n_4479;
  wire csa_tree_add_190_195_groupi_n_4480, csa_tree_add_190_195_groupi_n_4481, csa_tree_add_190_195_groupi_n_4482, csa_tree_add_190_195_groupi_n_4483, csa_tree_add_190_195_groupi_n_4484, csa_tree_add_190_195_groupi_n_4485, csa_tree_add_190_195_groupi_n_4486, csa_tree_add_190_195_groupi_n_4487;
  wire csa_tree_add_190_195_groupi_n_4488, csa_tree_add_190_195_groupi_n_4489, csa_tree_add_190_195_groupi_n_4490, csa_tree_add_190_195_groupi_n_4491, csa_tree_add_190_195_groupi_n_4492, csa_tree_add_190_195_groupi_n_4493, csa_tree_add_190_195_groupi_n_4494, csa_tree_add_190_195_groupi_n_4495;
  wire csa_tree_add_190_195_groupi_n_4496, csa_tree_add_190_195_groupi_n_4497, csa_tree_add_190_195_groupi_n_4498, csa_tree_add_190_195_groupi_n_4499, csa_tree_add_190_195_groupi_n_4500, csa_tree_add_190_195_groupi_n_4501, csa_tree_add_190_195_groupi_n_4502, csa_tree_add_190_195_groupi_n_4503;
  wire csa_tree_add_190_195_groupi_n_4504, csa_tree_add_190_195_groupi_n_4505, csa_tree_add_190_195_groupi_n_4506, csa_tree_add_190_195_groupi_n_4507, csa_tree_add_190_195_groupi_n_4508, csa_tree_add_190_195_groupi_n_4509, csa_tree_add_190_195_groupi_n_4510, csa_tree_add_190_195_groupi_n_4511;
  wire csa_tree_add_190_195_groupi_n_4512, csa_tree_add_190_195_groupi_n_4513, csa_tree_add_190_195_groupi_n_4514, csa_tree_add_190_195_groupi_n_4515, csa_tree_add_190_195_groupi_n_4516, csa_tree_add_190_195_groupi_n_4517, csa_tree_add_190_195_groupi_n_4518, csa_tree_add_190_195_groupi_n_4519;
  wire csa_tree_add_190_195_groupi_n_4520, csa_tree_add_190_195_groupi_n_4521, csa_tree_add_190_195_groupi_n_4522, csa_tree_add_190_195_groupi_n_4523, csa_tree_add_190_195_groupi_n_4524, csa_tree_add_190_195_groupi_n_4525, csa_tree_add_190_195_groupi_n_4526, csa_tree_add_190_195_groupi_n_4527;
  wire csa_tree_add_190_195_groupi_n_4528, csa_tree_add_190_195_groupi_n_4529, csa_tree_add_190_195_groupi_n_4530, csa_tree_add_190_195_groupi_n_4531, csa_tree_add_190_195_groupi_n_4532, csa_tree_add_190_195_groupi_n_4533, csa_tree_add_190_195_groupi_n_4534, csa_tree_add_190_195_groupi_n_4535;
  wire csa_tree_add_190_195_groupi_n_4536, csa_tree_add_190_195_groupi_n_4537, csa_tree_add_190_195_groupi_n_4538, csa_tree_add_190_195_groupi_n_4539, csa_tree_add_190_195_groupi_n_4540, csa_tree_add_190_195_groupi_n_4541, csa_tree_add_190_195_groupi_n_4542, csa_tree_add_190_195_groupi_n_4543;
  wire csa_tree_add_190_195_groupi_n_4544, csa_tree_add_190_195_groupi_n_4545, csa_tree_add_190_195_groupi_n_4546, csa_tree_add_190_195_groupi_n_4547, csa_tree_add_190_195_groupi_n_4548, csa_tree_add_190_195_groupi_n_4549, csa_tree_add_190_195_groupi_n_4550, csa_tree_add_190_195_groupi_n_4551;
  wire csa_tree_add_190_195_groupi_n_4552, csa_tree_add_190_195_groupi_n_4553, csa_tree_add_190_195_groupi_n_4554, csa_tree_add_190_195_groupi_n_4555, csa_tree_add_190_195_groupi_n_4556, csa_tree_add_190_195_groupi_n_4557, csa_tree_add_190_195_groupi_n_4558, csa_tree_add_190_195_groupi_n_4559;
  wire csa_tree_add_190_195_groupi_n_4560, csa_tree_add_190_195_groupi_n_4561, csa_tree_add_190_195_groupi_n_4562, csa_tree_add_190_195_groupi_n_4563, csa_tree_add_190_195_groupi_n_4564, csa_tree_add_190_195_groupi_n_4565, csa_tree_add_190_195_groupi_n_4566, csa_tree_add_190_195_groupi_n_4567;
  wire csa_tree_add_190_195_groupi_n_4568, csa_tree_add_190_195_groupi_n_4569, csa_tree_add_190_195_groupi_n_4570, csa_tree_add_190_195_groupi_n_4571, csa_tree_add_190_195_groupi_n_4572, csa_tree_add_190_195_groupi_n_4573, csa_tree_add_190_195_groupi_n_4574, csa_tree_add_190_195_groupi_n_4575;
  wire csa_tree_add_190_195_groupi_n_4576, csa_tree_add_190_195_groupi_n_4577, csa_tree_add_190_195_groupi_n_4578, csa_tree_add_190_195_groupi_n_4579, csa_tree_add_190_195_groupi_n_4580, csa_tree_add_190_195_groupi_n_4581, csa_tree_add_190_195_groupi_n_4582, csa_tree_add_190_195_groupi_n_4583;
  wire csa_tree_add_190_195_groupi_n_4584, csa_tree_add_190_195_groupi_n_4585, csa_tree_add_190_195_groupi_n_4586, csa_tree_add_190_195_groupi_n_4587, csa_tree_add_190_195_groupi_n_4588, csa_tree_add_190_195_groupi_n_4589, csa_tree_add_190_195_groupi_n_4590, csa_tree_add_190_195_groupi_n_4591;
  wire csa_tree_add_190_195_groupi_n_4592, csa_tree_add_190_195_groupi_n_4593, csa_tree_add_190_195_groupi_n_4594, csa_tree_add_190_195_groupi_n_4595, csa_tree_add_190_195_groupi_n_4596, csa_tree_add_190_195_groupi_n_4597, csa_tree_add_190_195_groupi_n_4598, csa_tree_add_190_195_groupi_n_4599;
  wire csa_tree_add_190_195_groupi_n_4600, csa_tree_add_190_195_groupi_n_4601, csa_tree_add_190_195_groupi_n_4602, csa_tree_add_190_195_groupi_n_4603, csa_tree_add_190_195_groupi_n_4604, csa_tree_add_190_195_groupi_n_4605, csa_tree_add_190_195_groupi_n_4606, csa_tree_add_190_195_groupi_n_4607;
  wire csa_tree_add_190_195_groupi_n_4608, csa_tree_add_190_195_groupi_n_4609, csa_tree_add_190_195_groupi_n_4610, csa_tree_add_190_195_groupi_n_4611, csa_tree_add_190_195_groupi_n_4612, csa_tree_add_190_195_groupi_n_4613, csa_tree_add_190_195_groupi_n_4614, csa_tree_add_190_195_groupi_n_4615;
  wire csa_tree_add_190_195_groupi_n_4616, csa_tree_add_190_195_groupi_n_4617, csa_tree_add_190_195_groupi_n_4618, csa_tree_add_190_195_groupi_n_4619, csa_tree_add_190_195_groupi_n_4620, csa_tree_add_190_195_groupi_n_4621, csa_tree_add_190_195_groupi_n_4622, csa_tree_add_190_195_groupi_n_4623;
  wire csa_tree_add_190_195_groupi_n_4624, csa_tree_add_190_195_groupi_n_4625, csa_tree_add_190_195_groupi_n_4626, csa_tree_add_190_195_groupi_n_4627, csa_tree_add_190_195_groupi_n_4628, csa_tree_add_190_195_groupi_n_4629, csa_tree_add_190_195_groupi_n_4630, csa_tree_add_190_195_groupi_n_4631;
  wire csa_tree_add_190_195_groupi_n_4632, csa_tree_add_190_195_groupi_n_4633, csa_tree_add_190_195_groupi_n_4634, csa_tree_add_190_195_groupi_n_4635, csa_tree_add_190_195_groupi_n_4636, csa_tree_add_190_195_groupi_n_4637, csa_tree_add_190_195_groupi_n_4638, csa_tree_add_190_195_groupi_n_4639;
  wire csa_tree_add_190_195_groupi_n_4640, csa_tree_add_190_195_groupi_n_4641, csa_tree_add_190_195_groupi_n_4642, csa_tree_add_190_195_groupi_n_4643, csa_tree_add_190_195_groupi_n_4644, csa_tree_add_190_195_groupi_n_4645, csa_tree_add_190_195_groupi_n_4646, csa_tree_add_190_195_groupi_n_4647;
  wire csa_tree_add_190_195_groupi_n_4648, csa_tree_add_190_195_groupi_n_4649, csa_tree_add_190_195_groupi_n_4650, csa_tree_add_190_195_groupi_n_4651, csa_tree_add_190_195_groupi_n_4652, csa_tree_add_190_195_groupi_n_4653, csa_tree_add_190_195_groupi_n_4654, csa_tree_add_190_195_groupi_n_4655;
  wire csa_tree_add_190_195_groupi_n_4656, csa_tree_add_190_195_groupi_n_4657, csa_tree_add_190_195_groupi_n_4658, csa_tree_add_190_195_groupi_n_4659, csa_tree_add_190_195_groupi_n_4660, csa_tree_add_190_195_groupi_n_4661, csa_tree_add_190_195_groupi_n_4662, csa_tree_add_190_195_groupi_n_4663;
  wire csa_tree_add_190_195_groupi_n_4664, csa_tree_add_190_195_groupi_n_4665, csa_tree_add_190_195_groupi_n_4666, csa_tree_add_190_195_groupi_n_4667, csa_tree_add_190_195_groupi_n_4668, csa_tree_add_190_195_groupi_n_4669, csa_tree_add_190_195_groupi_n_4670, csa_tree_add_190_195_groupi_n_4671;
  wire csa_tree_add_190_195_groupi_n_4672, csa_tree_add_190_195_groupi_n_4673, csa_tree_add_190_195_groupi_n_4674, csa_tree_add_190_195_groupi_n_4675, csa_tree_add_190_195_groupi_n_4676, csa_tree_add_190_195_groupi_n_4677, csa_tree_add_190_195_groupi_n_4678, csa_tree_add_190_195_groupi_n_4679;
  wire csa_tree_add_190_195_groupi_n_4680, csa_tree_add_190_195_groupi_n_4681, csa_tree_add_190_195_groupi_n_4682, csa_tree_add_190_195_groupi_n_4683, csa_tree_add_190_195_groupi_n_4684, csa_tree_add_190_195_groupi_n_4685, csa_tree_add_190_195_groupi_n_4686, csa_tree_add_190_195_groupi_n_4687;
  wire csa_tree_add_190_195_groupi_n_4688, csa_tree_add_190_195_groupi_n_4689, csa_tree_add_190_195_groupi_n_4690, csa_tree_add_190_195_groupi_n_4691, csa_tree_add_190_195_groupi_n_4692, csa_tree_add_190_195_groupi_n_4693, csa_tree_add_190_195_groupi_n_4694, csa_tree_add_190_195_groupi_n_4695;
  wire csa_tree_add_190_195_groupi_n_4696, csa_tree_add_190_195_groupi_n_4697, csa_tree_add_190_195_groupi_n_4698, csa_tree_add_190_195_groupi_n_4699, csa_tree_add_190_195_groupi_n_4700, csa_tree_add_190_195_groupi_n_4701, csa_tree_add_190_195_groupi_n_4702, csa_tree_add_190_195_groupi_n_4703;
  wire csa_tree_add_190_195_groupi_n_4704, csa_tree_add_190_195_groupi_n_4705, csa_tree_add_190_195_groupi_n_4706, csa_tree_add_190_195_groupi_n_4707, csa_tree_add_190_195_groupi_n_4708, csa_tree_add_190_195_groupi_n_4709, csa_tree_add_190_195_groupi_n_4710, csa_tree_add_190_195_groupi_n_4711;
  wire csa_tree_add_190_195_groupi_n_4712, csa_tree_add_190_195_groupi_n_4713, csa_tree_add_190_195_groupi_n_4714, csa_tree_add_190_195_groupi_n_4715, csa_tree_add_190_195_groupi_n_4716, csa_tree_add_190_195_groupi_n_4717, csa_tree_add_190_195_groupi_n_4718, csa_tree_add_190_195_groupi_n_4719;
  wire csa_tree_add_190_195_groupi_n_4720, csa_tree_add_190_195_groupi_n_4721, csa_tree_add_190_195_groupi_n_4722, csa_tree_add_190_195_groupi_n_4723, csa_tree_add_190_195_groupi_n_4724, csa_tree_add_190_195_groupi_n_4725, csa_tree_add_190_195_groupi_n_4726, csa_tree_add_190_195_groupi_n_4727;
  wire csa_tree_add_190_195_groupi_n_4728, csa_tree_add_190_195_groupi_n_4729, csa_tree_add_190_195_groupi_n_4730, csa_tree_add_190_195_groupi_n_4731, csa_tree_add_190_195_groupi_n_4732, csa_tree_add_190_195_groupi_n_4733, csa_tree_add_190_195_groupi_n_4734, csa_tree_add_190_195_groupi_n_4735;
  wire csa_tree_add_190_195_groupi_n_4736, csa_tree_add_190_195_groupi_n_4737, csa_tree_add_190_195_groupi_n_4738, csa_tree_add_190_195_groupi_n_4739, csa_tree_add_190_195_groupi_n_4740, csa_tree_add_190_195_groupi_n_4741, csa_tree_add_190_195_groupi_n_4742, csa_tree_add_190_195_groupi_n_4743;
  wire csa_tree_add_190_195_groupi_n_4744, csa_tree_add_190_195_groupi_n_4745, csa_tree_add_190_195_groupi_n_4746, csa_tree_add_190_195_groupi_n_4747, csa_tree_add_190_195_groupi_n_4748, csa_tree_add_190_195_groupi_n_4749, csa_tree_add_190_195_groupi_n_4750, csa_tree_add_190_195_groupi_n_4751;
  wire csa_tree_add_190_195_groupi_n_4752, csa_tree_add_190_195_groupi_n_4753, csa_tree_add_190_195_groupi_n_4754, csa_tree_add_190_195_groupi_n_4755, csa_tree_add_190_195_groupi_n_4756, csa_tree_add_190_195_groupi_n_4757, csa_tree_add_190_195_groupi_n_4758, csa_tree_add_190_195_groupi_n_4759;
  wire csa_tree_add_190_195_groupi_n_4760, csa_tree_add_190_195_groupi_n_4761, csa_tree_add_190_195_groupi_n_4762, csa_tree_add_190_195_groupi_n_4763, csa_tree_add_190_195_groupi_n_4764, csa_tree_add_190_195_groupi_n_4765, csa_tree_add_190_195_groupi_n_4766, csa_tree_add_190_195_groupi_n_4767;
  wire csa_tree_add_190_195_groupi_n_4768, csa_tree_add_190_195_groupi_n_4769, csa_tree_add_190_195_groupi_n_4770, csa_tree_add_190_195_groupi_n_4771, csa_tree_add_190_195_groupi_n_4772, csa_tree_add_190_195_groupi_n_4773, csa_tree_add_190_195_groupi_n_4774, csa_tree_add_190_195_groupi_n_4775;
  wire csa_tree_add_190_195_groupi_n_4776, csa_tree_add_190_195_groupi_n_4777, csa_tree_add_190_195_groupi_n_4778, csa_tree_add_190_195_groupi_n_4779, csa_tree_add_190_195_groupi_n_4780, csa_tree_add_190_195_groupi_n_4781, csa_tree_add_190_195_groupi_n_4782, csa_tree_add_190_195_groupi_n_4783;
  wire csa_tree_add_190_195_groupi_n_4784, csa_tree_add_190_195_groupi_n_4785, csa_tree_add_190_195_groupi_n_4786, csa_tree_add_190_195_groupi_n_4787, csa_tree_add_190_195_groupi_n_4788, csa_tree_add_190_195_groupi_n_4789, csa_tree_add_190_195_groupi_n_4790, csa_tree_add_190_195_groupi_n_4791;
  wire csa_tree_add_190_195_groupi_n_4792, csa_tree_add_190_195_groupi_n_4793, csa_tree_add_190_195_groupi_n_4794, csa_tree_add_190_195_groupi_n_4795, csa_tree_add_190_195_groupi_n_4796, csa_tree_add_190_195_groupi_n_4797, csa_tree_add_190_195_groupi_n_4798, csa_tree_add_190_195_groupi_n_4799;
  wire csa_tree_add_190_195_groupi_n_4800, csa_tree_add_190_195_groupi_n_4801, csa_tree_add_190_195_groupi_n_4802, csa_tree_add_190_195_groupi_n_4803, csa_tree_add_190_195_groupi_n_4804, csa_tree_add_190_195_groupi_n_4805, csa_tree_add_190_195_groupi_n_4806, csa_tree_add_190_195_groupi_n_4807;
  wire csa_tree_add_190_195_groupi_n_4808, csa_tree_add_190_195_groupi_n_4809, csa_tree_add_190_195_groupi_n_4810, csa_tree_add_190_195_groupi_n_4811, csa_tree_add_190_195_groupi_n_4812, csa_tree_add_190_195_groupi_n_4813, csa_tree_add_190_195_groupi_n_4814, csa_tree_add_190_195_groupi_n_4815;
  wire csa_tree_add_190_195_groupi_n_4816, csa_tree_add_190_195_groupi_n_4817, csa_tree_add_190_195_groupi_n_4818, csa_tree_add_190_195_groupi_n_4819, csa_tree_add_190_195_groupi_n_4820, csa_tree_add_190_195_groupi_n_4821, csa_tree_add_190_195_groupi_n_4822, csa_tree_add_190_195_groupi_n_4823;
  wire csa_tree_add_190_195_groupi_n_4824, csa_tree_add_190_195_groupi_n_4825, csa_tree_add_190_195_groupi_n_4826, csa_tree_add_190_195_groupi_n_4827, csa_tree_add_190_195_groupi_n_4828, csa_tree_add_190_195_groupi_n_4829, csa_tree_add_190_195_groupi_n_4830, csa_tree_add_190_195_groupi_n_4831;
  wire csa_tree_add_190_195_groupi_n_4832, csa_tree_add_190_195_groupi_n_4833, csa_tree_add_190_195_groupi_n_4834, csa_tree_add_190_195_groupi_n_4835, csa_tree_add_190_195_groupi_n_4836, csa_tree_add_190_195_groupi_n_4837, csa_tree_add_190_195_groupi_n_4838, csa_tree_add_190_195_groupi_n_4839;
  wire csa_tree_add_190_195_groupi_n_4840, csa_tree_add_190_195_groupi_n_4841, csa_tree_add_190_195_groupi_n_4842, csa_tree_add_190_195_groupi_n_4843, csa_tree_add_190_195_groupi_n_4844, csa_tree_add_190_195_groupi_n_4845, csa_tree_add_190_195_groupi_n_4846, csa_tree_add_190_195_groupi_n_4847;
  wire csa_tree_add_190_195_groupi_n_4848, csa_tree_add_190_195_groupi_n_4849, csa_tree_add_190_195_groupi_n_4850, csa_tree_add_190_195_groupi_n_4851, csa_tree_add_190_195_groupi_n_4852, csa_tree_add_190_195_groupi_n_4853, csa_tree_add_190_195_groupi_n_4854, csa_tree_add_190_195_groupi_n_4855;
  wire csa_tree_add_190_195_groupi_n_4856, csa_tree_add_190_195_groupi_n_4857, csa_tree_add_190_195_groupi_n_4858, csa_tree_add_190_195_groupi_n_4859, csa_tree_add_190_195_groupi_n_4860, csa_tree_add_190_195_groupi_n_4861, csa_tree_add_190_195_groupi_n_4862, csa_tree_add_190_195_groupi_n_4863;
  wire csa_tree_add_190_195_groupi_n_4864, csa_tree_add_190_195_groupi_n_4865, csa_tree_add_190_195_groupi_n_4866, csa_tree_add_190_195_groupi_n_4867, csa_tree_add_190_195_groupi_n_4868, csa_tree_add_190_195_groupi_n_4869, csa_tree_add_190_195_groupi_n_4870, csa_tree_add_190_195_groupi_n_4871;
  wire csa_tree_add_190_195_groupi_n_4872, csa_tree_add_190_195_groupi_n_4873, csa_tree_add_190_195_groupi_n_4874, csa_tree_add_190_195_groupi_n_4875, csa_tree_add_190_195_groupi_n_4876, csa_tree_add_190_195_groupi_n_4877, csa_tree_add_190_195_groupi_n_4878, csa_tree_add_190_195_groupi_n_4879;
  wire csa_tree_add_190_195_groupi_n_4880, csa_tree_add_190_195_groupi_n_4881, csa_tree_add_190_195_groupi_n_4882, csa_tree_add_190_195_groupi_n_4883, csa_tree_add_190_195_groupi_n_4884, csa_tree_add_190_195_groupi_n_4885, csa_tree_add_190_195_groupi_n_4886, csa_tree_add_190_195_groupi_n_4887;
  wire csa_tree_add_190_195_groupi_n_4888, csa_tree_add_190_195_groupi_n_4889, csa_tree_add_190_195_groupi_n_4890, csa_tree_add_190_195_groupi_n_4891, csa_tree_add_190_195_groupi_n_4892, csa_tree_add_190_195_groupi_n_4893, csa_tree_add_190_195_groupi_n_4894, csa_tree_add_190_195_groupi_n_4895;
  wire csa_tree_add_190_195_groupi_n_4896, csa_tree_add_190_195_groupi_n_4897, csa_tree_add_190_195_groupi_n_4898, csa_tree_add_190_195_groupi_n_4899, csa_tree_add_190_195_groupi_n_4900, csa_tree_add_190_195_groupi_n_4901, csa_tree_add_190_195_groupi_n_4902, csa_tree_add_190_195_groupi_n_4903;
  wire csa_tree_add_190_195_groupi_n_4904, csa_tree_add_190_195_groupi_n_4905, csa_tree_add_190_195_groupi_n_4906, csa_tree_add_190_195_groupi_n_4907, csa_tree_add_190_195_groupi_n_4908, csa_tree_add_190_195_groupi_n_4909, csa_tree_add_190_195_groupi_n_4910, csa_tree_add_190_195_groupi_n_4911;
  wire csa_tree_add_190_195_groupi_n_4912, csa_tree_add_190_195_groupi_n_4913, csa_tree_add_190_195_groupi_n_4914, csa_tree_add_190_195_groupi_n_4915, csa_tree_add_190_195_groupi_n_4916, csa_tree_add_190_195_groupi_n_4917, csa_tree_add_190_195_groupi_n_4918, csa_tree_add_190_195_groupi_n_4919;
  wire csa_tree_add_190_195_groupi_n_4920, csa_tree_add_190_195_groupi_n_4921, csa_tree_add_190_195_groupi_n_4922, csa_tree_add_190_195_groupi_n_4923, csa_tree_add_190_195_groupi_n_4924, csa_tree_add_190_195_groupi_n_4925, csa_tree_add_190_195_groupi_n_4926, csa_tree_add_190_195_groupi_n_4927;
  wire csa_tree_add_190_195_groupi_n_4928, csa_tree_add_190_195_groupi_n_4929, csa_tree_add_190_195_groupi_n_4930, csa_tree_add_190_195_groupi_n_4931, csa_tree_add_190_195_groupi_n_4932, csa_tree_add_190_195_groupi_n_4933, csa_tree_add_190_195_groupi_n_4934, csa_tree_add_190_195_groupi_n_4935;
  wire csa_tree_add_190_195_groupi_n_4936, csa_tree_add_190_195_groupi_n_4937, csa_tree_add_190_195_groupi_n_4938, csa_tree_add_190_195_groupi_n_4939, csa_tree_add_190_195_groupi_n_4940, csa_tree_add_190_195_groupi_n_4941, csa_tree_add_190_195_groupi_n_4942, csa_tree_add_190_195_groupi_n_4943;
  wire csa_tree_add_190_195_groupi_n_4944, csa_tree_add_190_195_groupi_n_4945, csa_tree_add_190_195_groupi_n_4946, csa_tree_add_190_195_groupi_n_4947, csa_tree_add_190_195_groupi_n_4948, csa_tree_add_190_195_groupi_n_4949, csa_tree_add_190_195_groupi_n_4950, csa_tree_add_190_195_groupi_n_4951;
  wire csa_tree_add_190_195_groupi_n_4952, csa_tree_add_190_195_groupi_n_4953, csa_tree_add_190_195_groupi_n_4954, csa_tree_add_190_195_groupi_n_4955, csa_tree_add_190_195_groupi_n_4956, csa_tree_add_190_195_groupi_n_4957, csa_tree_add_190_195_groupi_n_4958, csa_tree_add_190_195_groupi_n_4959;
  wire csa_tree_add_190_195_groupi_n_4960, csa_tree_add_190_195_groupi_n_4961, csa_tree_add_190_195_groupi_n_4962, csa_tree_add_190_195_groupi_n_4963, csa_tree_add_190_195_groupi_n_4964, csa_tree_add_190_195_groupi_n_4965, csa_tree_add_190_195_groupi_n_4966, csa_tree_add_190_195_groupi_n_4967;
  wire csa_tree_add_190_195_groupi_n_4968, csa_tree_add_190_195_groupi_n_4969, csa_tree_add_190_195_groupi_n_4970, csa_tree_add_190_195_groupi_n_4971, csa_tree_add_190_195_groupi_n_4972, csa_tree_add_190_195_groupi_n_4973, csa_tree_add_190_195_groupi_n_4974, csa_tree_add_190_195_groupi_n_4975;
  wire csa_tree_add_190_195_groupi_n_4976, csa_tree_add_190_195_groupi_n_4977, csa_tree_add_190_195_groupi_n_4978, csa_tree_add_190_195_groupi_n_4979, csa_tree_add_190_195_groupi_n_4980, csa_tree_add_190_195_groupi_n_4981, csa_tree_add_190_195_groupi_n_4982, csa_tree_add_190_195_groupi_n_4983;
  wire csa_tree_add_190_195_groupi_n_4984, csa_tree_add_190_195_groupi_n_4985, csa_tree_add_190_195_groupi_n_4986, csa_tree_add_190_195_groupi_n_4987, csa_tree_add_190_195_groupi_n_4988, csa_tree_add_190_195_groupi_n_4989, csa_tree_add_190_195_groupi_n_4990, csa_tree_add_190_195_groupi_n_4991;
  wire csa_tree_add_190_195_groupi_n_4992, csa_tree_add_190_195_groupi_n_4993, csa_tree_add_190_195_groupi_n_4994, csa_tree_add_190_195_groupi_n_4995, csa_tree_add_190_195_groupi_n_4996, csa_tree_add_190_195_groupi_n_4997, csa_tree_add_190_195_groupi_n_4998, csa_tree_add_190_195_groupi_n_4999;
  wire csa_tree_add_190_195_groupi_n_5000, csa_tree_add_190_195_groupi_n_5001, csa_tree_add_190_195_groupi_n_5002, csa_tree_add_190_195_groupi_n_5003, csa_tree_add_190_195_groupi_n_5004, csa_tree_add_190_195_groupi_n_5005, csa_tree_add_190_195_groupi_n_5006, csa_tree_add_190_195_groupi_n_5007;
  wire csa_tree_add_190_195_groupi_n_5008, csa_tree_add_190_195_groupi_n_5009, csa_tree_add_190_195_groupi_n_5010, csa_tree_add_190_195_groupi_n_5011, csa_tree_add_190_195_groupi_n_5012, csa_tree_add_190_195_groupi_n_5013, csa_tree_add_190_195_groupi_n_5014, csa_tree_add_190_195_groupi_n_5015;
  wire csa_tree_add_190_195_groupi_n_5016, csa_tree_add_190_195_groupi_n_5017, csa_tree_add_190_195_groupi_n_5018, csa_tree_add_190_195_groupi_n_5019, csa_tree_add_190_195_groupi_n_5020, csa_tree_add_190_195_groupi_n_5021, csa_tree_add_190_195_groupi_n_5022, csa_tree_add_190_195_groupi_n_5023;
  wire csa_tree_add_190_195_groupi_n_5024, csa_tree_add_190_195_groupi_n_5025, csa_tree_add_190_195_groupi_n_5026, csa_tree_add_190_195_groupi_n_5027, csa_tree_add_190_195_groupi_n_5028, csa_tree_add_190_195_groupi_n_5029, csa_tree_add_190_195_groupi_n_5030, csa_tree_add_190_195_groupi_n_5031;
  wire csa_tree_add_190_195_groupi_n_5032, csa_tree_add_190_195_groupi_n_5033, csa_tree_add_190_195_groupi_n_5034, csa_tree_add_190_195_groupi_n_5035, csa_tree_add_190_195_groupi_n_5036, csa_tree_add_190_195_groupi_n_5037, csa_tree_add_190_195_groupi_n_5038, csa_tree_add_190_195_groupi_n_5039;
  wire csa_tree_add_190_195_groupi_n_5040, csa_tree_add_190_195_groupi_n_5041, csa_tree_add_190_195_groupi_n_5042, csa_tree_add_190_195_groupi_n_5043, csa_tree_add_190_195_groupi_n_5044, csa_tree_add_190_195_groupi_n_5045, csa_tree_add_190_195_groupi_n_5046, csa_tree_add_190_195_groupi_n_5047;
  wire csa_tree_add_190_195_groupi_n_5048, csa_tree_add_190_195_groupi_n_5049, csa_tree_add_190_195_groupi_n_5050, csa_tree_add_190_195_groupi_n_5051, csa_tree_add_190_195_groupi_n_5052, csa_tree_add_190_195_groupi_n_5053, csa_tree_add_190_195_groupi_n_5054, csa_tree_add_190_195_groupi_n_5055;
  wire csa_tree_add_190_195_groupi_n_5056, csa_tree_add_190_195_groupi_n_5057, csa_tree_add_190_195_groupi_n_5058, csa_tree_add_190_195_groupi_n_5059, csa_tree_add_190_195_groupi_n_5060, csa_tree_add_190_195_groupi_n_5061, csa_tree_add_190_195_groupi_n_5062, csa_tree_add_190_195_groupi_n_5063;
  wire csa_tree_add_190_195_groupi_n_5064, csa_tree_add_190_195_groupi_n_5065, csa_tree_add_190_195_groupi_n_5066, csa_tree_add_190_195_groupi_n_5067, csa_tree_add_190_195_groupi_n_5068, csa_tree_add_190_195_groupi_n_5069, csa_tree_add_190_195_groupi_n_5070, csa_tree_add_190_195_groupi_n_5071;
  wire csa_tree_add_190_195_groupi_n_5072, csa_tree_add_190_195_groupi_n_5073, csa_tree_add_190_195_groupi_n_5074, csa_tree_add_190_195_groupi_n_5075, csa_tree_add_190_195_groupi_n_5076, csa_tree_add_190_195_groupi_n_5077, csa_tree_add_190_195_groupi_n_5078, csa_tree_add_190_195_groupi_n_5079;
  wire csa_tree_add_190_195_groupi_n_5080, csa_tree_add_190_195_groupi_n_5081, csa_tree_add_190_195_groupi_n_5082, csa_tree_add_190_195_groupi_n_5083, csa_tree_add_190_195_groupi_n_5084, csa_tree_add_190_195_groupi_n_5085, csa_tree_add_190_195_groupi_n_5086, csa_tree_add_190_195_groupi_n_5087;
  wire csa_tree_add_190_195_groupi_n_5088, csa_tree_add_190_195_groupi_n_5089, csa_tree_add_190_195_groupi_n_5090, csa_tree_add_190_195_groupi_n_5091, csa_tree_add_190_195_groupi_n_5092, csa_tree_add_190_195_groupi_n_5093, csa_tree_add_190_195_groupi_n_5094, csa_tree_add_190_195_groupi_n_5095;
  wire csa_tree_add_190_195_groupi_n_5096, csa_tree_add_190_195_groupi_n_5097, csa_tree_add_190_195_groupi_n_5098, csa_tree_add_190_195_groupi_n_5099, csa_tree_add_190_195_groupi_n_5100, csa_tree_add_190_195_groupi_n_5101, csa_tree_add_190_195_groupi_n_5102, csa_tree_add_190_195_groupi_n_5103;
  wire csa_tree_add_190_195_groupi_n_5104, csa_tree_add_190_195_groupi_n_5105, csa_tree_add_190_195_groupi_n_5106, csa_tree_add_190_195_groupi_n_5107, csa_tree_add_190_195_groupi_n_5108, csa_tree_add_190_195_groupi_n_5109, csa_tree_add_190_195_groupi_n_5110, csa_tree_add_190_195_groupi_n_5111;
  wire csa_tree_add_190_195_groupi_n_5112, csa_tree_add_190_195_groupi_n_5113, csa_tree_add_190_195_groupi_n_5114, csa_tree_add_190_195_groupi_n_5115, csa_tree_add_190_195_groupi_n_5116, csa_tree_add_190_195_groupi_n_5117, csa_tree_add_190_195_groupi_n_5118, csa_tree_add_190_195_groupi_n_5119;
  wire csa_tree_add_190_195_groupi_n_5120, csa_tree_add_190_195_groupi_n_5121, csa_tree_add_190_195_groupi_n_5122, csa_tree_add_190_195_groupi_n_5123, csa_tree_add_190_195_groupi_n_5124, csa_tree_add_190_195_groupi_n_5125, csa_tree_add_190_195_groupi_n_5126, csa_tree_add_190_195_groupi_n_5127;
  wire csa_tree_add_190_195_groupi_n_5128, csa_tree_add_190_195_groupi_n_5129, csa_tree_add_190_195_groupi_n_5130, csa_tree_add_190_195_groupi_n_5131, csa_tree_add_190_195_groupi_n_5132, csa_tree_add_190_195_groupi_n_5133, csa_tree_add_190_195_groupi_n_5134, csa_tree_add_190_195_groupi_n_5135;
  wire csa_tree_add_190_195_groupi_n_5136, csa_tree_add_190_195_groupi_n_5137, csa_tree_add_190_195_groupi_n_5138, csa_tree_add_190_195_groupi_n_5139, csa_tree_add_190_195_groupi_n_5140, csa_tree_add_190_195_groupi_n_5141, csa_tree_add_190_195_groupi_n_5142, csa_tree_add_190_195_groupi_n_5143;
  wire csa_tree_add_190_195_groupi_n_5144, csa_tree_add_190_195_groupi_n_5145, csa_tree_add_190_195_groupi_n_5146, csa_tree_add_190_195_groupi_n_5147, csa_tree_add_190_195_groupi_n_5148, csa_tree_add_190_195_groupi_n_5149, csa_tree_add_190_195_groupi_n_5150, csa_tree_add_190_195_groupi_n_5151;
  wire csa_tree_add_190_195_groupi_n_5152, csa_tree_add_190_195_groupi_n_5153, csa_tree_add_190_195_groupi_n_5154, csa_tree_add_190_195_groupi_n_5155, csa_tree_add_190_195_groupi_n_5156, csa_tree_add_190_195_groupi_n_5157, csa_tree_add_190_195_groupi_n_5158, csa_tree_add_190_195_groupi_n_5159;
  wire csa_tree_add_190_195_groupi_n_5160, csa_tree_add_190_195_groupi_n_5161, csa_tree_add_190_195_groupi_n_5162, csa_tree_add_190_195_groupi_n_5163, csa_tree_add_190_195_groupi_n_5164, csa_tree_add_190_195_groupi_n_5165, csa_tree_add_190_195_groupi_n_5166, csa_tree_add_190_195_groupi_n_5167;
  wire csa_tree_add_190_195_groupi_n_5168, csa_tree_add_190_195_groupi_n_5169, csa_tree_add_190_195_groupi_n_5170, csa_tree_add_190_195_groupi_n_5171, csa_tree_add_190_195_groupi_n_5172, csa_tree_add_190_195_groupi_n_5173, csa_tree_add_190_195_groupi_n_5174, csa_tree_add_190_195_groupi_n_5175;
  wire csa_tree_add_190_195_groupi_n_5176, csa_tree_add_190_195_groupi_n_5177, csa_tree_add_190_195_groupi_n_5178, csa_tree_add_190_195_groupi_n_5179, csa_tree_add_190_195_groupi_n_5180, csa_tree_add_190_195_groupi_n_5181, csa_tree_add_190_195_groupi_n_5182, csa_tree_add_190_195_groupi_n_5183;
  wire csa_tree_add_190_195_groupi_n_5184, csa_tree_add_190_195_groupi_n_5185, csa_tree_add_190_195_groupi_n_5186, csa_tree_add_190_195_groupi_n_5187, csa_tree_add_190_195_groupi_n_5188, csa_tree_add_190_195_groupi_n_5189, csa_tree_add_190_195_groupi_n_5190, csa_tree_add_190_195_groupi_n_5191;
  wire csa_tree_add_190_195_groupi_n_5192, csa_tree_add_190_195_groupi_n_5193, csa_tree_add_190_195_groupi_n_5194, csa_tree_add_190_195_groupi_n_5195, csa_tree_add_190_195_groupi_n_5196, csa_tree_add_190_195_groupi_n_5197, csa_tree_add_190_195_groupi_n_5198, csa_tree_add_190_195_groupi_n_5199;
  wire csa_tree_add_190_195_groupi_n_5200, csa_tree_add_190_195_groupi_n_5201, csa_tree_add_190_195_groupi_n_5202, csa_tree_add_190_195_groupi_n_5203, csa_tree_add_190_195_groupi_n_5204, csa_tree_add_190_195_groupi_n_5205, csa_tree_add_190_195_groupi_n_5206, csa_tree_add_190_195_groupi_n_5207;
  wire csa_tree_add_190_195_groupi_n_5208, csa_tree_add_190_195_groupi_n_5209, csa_tree_add_190_195_groupi_n_5210, csa_tree_add_190_195_groupi_n_5211, csa_tree_add_190_195_groupi_n_5212, csa_tree_add_190_195_groupi_n_5213, csa_tree_add_190_195_groupi_n_5214, csa_tree_add_190_195_groupi_n_5215;
  wire csa_tree_add_190_195_groupi_n_5216, csa_tree_add_190_195_groupi_n_5217, csa_tree_add_190_195_groupi_n_5218, csa_tree_add_190_195_groupi_n_5219, csa_tree_add_190_195_groupi_n_5220, csa_tree_add_190_195_groupi_n_5221, csa_tree_add_190_195_groupi_n_5222, csa_tree_add_190_195_groupi_n_5223;
  wire csa_tree_add_190_195_groupi_n_5224, csa_tree_add_190_195_groupi_n_5225, csa_tree_add_190_195_groupi_n_5226, csa_tree_add_190_195_groupi_n_5227, csa_tree_add_190_195_groupi_n_5228, csa_tree_add_190_195_groupi_n_5229, csa_tree_add_190_195_groupi_n_5230, csa_tree_add_190_195_groupi_n_5231;
  wire csa_tree_add_190_195_groupi_n_5232, csa_tree_add_190_195_groupi_n_5233, csa_tree_add_190_195_groupi_n_5234, csa_tree_add_190_195_groupi_n_5235, csa_tree_add_190_195_groupi_n_5236, csa_tree_add_190_195_groupi_n_5237, csa_tree_add_190_195_groupi_n_5238, csa_tree_add_190_195_groupi_n_5239;
  wire csa_tree_add_190_195_groupi_n_5240, csa_tree_add_190_195_groupi_n_5241, csa_tree_add_190_195_groupi_n_5242, csa_tree_add_190_195_groupi_n_5243, csa_tree_add_190_195_groupi_n_5244, csa_tree_add_190_195_groupi_n_5245, csa_tree_add_190_195_groupi_n_5246, csa_tree_add_190_195_groupi_n_5247;
  wire csa_tree_add_190_195_groupi_n_5248, csa_tree_add_190_195_groupi_n_5249, csa_tree_add_190_195_groupi_n_5250, csa_tree_add_190_195_groupi_n_5251, csa_tree_add_190_195_groupi_n_5252, csa_tree_add_190_195_groupi_n_5253, csa_tree_add_190_195_groupi_n_5254, csa_tree_add_190_195_groupi_n_5255;
  wire csa_tree_add_190_195_groupi_n_5256, csa_tree_add_190_195_groupi_n_5257, csa_tree_add_190_195_groupi_n_5258, csa_tree_add_190_195_groupi_n_5259, csa_tree_add_190_195_groupi_n_5260, csa_tree_add_190_195_groupi_n_5261, csa_tree_add_190_195_groupi_n_5262, csa_tree_add_190_195_groupi_n_5263;
  wire csa_tree_add_190_195_groupi_n_5264, csa_tree_add_190_195_groupi_n_5265, csa_tree_add_190_195_groupi_n_5266, csa_tree_add_190_195_groupi_n_5267, csa_tree_add_190_195_groupi_n_5268, csa_tree_add_190_195_groupi_n_5269, csa_tree_add_190_195_groupi_n_5270, csa_tree_add_190_195_groupi_n_5271;
  wire csa_tree_add_190_195_groupi_n_5272, csa_tree_add_190_195_groupi_n_5273, csa_tree_add_190_195_groupi_n_5274, csa_tree_add_190_195_groupi_n_5275, csa_tree_add_190_195_groupi_n_5276, csa_tree_add_190_195_groupi_n_5277, csa_tree_add_190_195_groupi_n_5278, csa_tree_add_190_195_groupi_n_5279;
  wire csa_tree_add_190_195_groupi_n_5280, csa_tree_add_190_195_groupi_n_5281, csa_tree_add_190_195_groupi_n_5282, csa_tree_add_190_195_groupi_n_5283, csa_tree_add_190_195_groupi_n_5284, csa_tree_add_190_195_groupi_n_5285, csa_tree_add_190_195_groupi_n_5286, csa_tree_add_190_195_groupi_n_5287;
  wire csa_tree_add_190_195_groupi_n_5288, csa_tree_add_190_195_groupi_n_5289, csa_tree_add_190_195_groupi_n_5290, csa_tree_add_190_195_groupi_n_5291, csa_tree_add_190_195_groupi_n_5292, csa_tree_add_190_195_groupi_n_5293, csa_tree_add_190_195_groupi_n_5294, csa_tree_add_190_195_groupi_n_5295;
  wire csa_tree_add_190_195_groupi_n_5296, csa_tree_add_190_195_groupi_n_5297, csa_tree_add_190_195_groupi_n_5298, csa_tree_add_190_195_groupi_n_5299, csa_tree_add_190_195_groupi_n_5300, csa_tree_add_190_195_groupi_n_5301, csa_tree_add_190_195_groupi_n_5302, csa_tree_add_190_195_groupi_n_5303;
  wire csa_tree_add_190_195_groupi_n_5304, csa_tree_add_190_195_groupi_n_5305, csa_tree_add_190_195_groupi_n_5306, csa_tree_add_190_195_groupi_n_5307, csa_tree_add_190_195_groupi_n_5308, csa_tree_add_190_195_groupi_n_5309, csa_tree_add_190_195_groupi_n_5310, csa_tree_add_190_195_groupi_n_5311;
  wire csa_tree_add_190_195_groupi_n_5312, csa_tree_add_190_195_groupi_n_5313, csa_tree_add_190_195_groupi_n_5314, csa_tree_add_190_195_groupi_n_5315, csa_tree_add_190_195_groupi_n_5316, csa_tree_add_190_195_groupi_n_5317, csa_tree_add_190_195_groupi_n_5318, csa_tree_add_190_195_groupi_n_5319;
  wire csa_tree_add_190_195_groupi_n_5320, csa_tree_add_190_195_groupi_n_5321, csa_tree_add_190_195_groupi_n_5322, csa_tree_add_190_195_groupi_n_5323, csa_tree_add_190_195_groupi_n_5324, csa_tree_add_190_195_groupi_n_5325, csa_tree_add_190_195_groupi_n_5326, csa_tree_add_190_195_groupi_n_5327;
  wire csa_tree_add_190_195_groupi_n_5328, csa_tree_add_190_195_groupi_n_5329, csa_tree_add_190_195_groupi_n_5330, csa_tree_add_190_195_groupi_n_5331, csa_tree_add_190_195_groupi_n_5332, csa_tree_add_190_195_groupi_n_5333, csa_tree_add_190_195_groupi_n_5334, csa_tree_add_190_195_groupi_n_5335;
  wire csa_tree_add_190_195_groupi_n_5336, csa_tree_add_190_195_groupi_n_5337, csa_tree_add_190_195_groupi_n_5338, csa_tree_add_190_195_groupi_n_5339, csa_tree_add_190_195_groupi_n_5340, csa_tree_add_190_195_groupi_n_5341, csa_tree_add_190_195_groupi_n_5342, csa_tree_add_190_195_groupi_n_5343;
  wire csa_tree_add_190_195_groupi_n_5344, csa_tree_add_190_195_groupi_n_5345, csa_tree_add_190_195_groupi_n_5346, csa_tree_add_190_195_groupi_n_5347, csa_tree_add_190_195_groupi_n_5348, csa_tree_add_190_195_groupi_n_5349, csa_tree_add_190_195_groupi_n_5350, csa_tree_add_190_195_groupi_n_5351;
  wire csa_tree_add_190_195_groupi_n_5352, csa_tree_add_190_195_groupi_n_5353, csa_tree_add_190_195_groupi_n_5354, csa_tree_add_190_195_groupi_n_5355, csa_tree_add_190_195_groupi_n_5356, csa_tree_add_190_195_groupi_n_5357, csa_tree_add_190_195_groupi_n_5358, csa_tree_add_190_195_groupi_n_5359;
  wire csa_tree_add_190_195_groupi_n_5360, csa_tree_add_190_195_groupi_n_5361, csa_tree_add_190_195_groupi_n_5362, csa_tree_add_190_195_groupi_n_5363, csa_tree_add_190_195_groupi_n_5364, csa_tree_add_190_195_groupi_n_5365, csa_tree_add_190_195_groupi_n_5366, csa_tree_add_190_195_groupi_n_5367;
  wire csa_tree_add_190_195_groupi_n_5368, csa_tree_add_190_195_groupi_n_5369, csa_tree_add_190_195_groupi_n_5370, csa_tree_add_190_195_groupi_n_5371, csa_tree_add_190_195_groupi_n_5372, csa_tree_add_190_195_groupi_n_5373, csa_tree_add_190_195_groupi_n_5374, csa_tree_add_190_195_groupi_n_5375;
  wire csa_tree_add_190_195_groupi_n_5376, csa_tree_add_190_195_groupi_n_5377, csa_tree_add_190_195_groupi_n_5378, csa_tree_add_190_195_groupi_n_5379, csa_tree_add_190_195_groupi_n_5380, csa_tree_add_190_195_groupi_n_5381, csa_tree_add_190_195_groupi_n_5382, csa_tree_add_190_195_groupi_n_5383;
  wire csa_tree_add_190_195_groupi_n_5384, csa_tree_add_190_195_groupi_n_5385, csa_tree_add_190_195_groupi_n_5386, csa_tree_add_190_195_groupi_n_5387, csa_tree_add_190_195_groupi_n_5388, csa_tree_add_190_195_groupi_n_5389, csa_tree_add_190_195_groupi_n_5390, csa_tree_add_190_195_groupi_n_5391;
  wire csa_tree_add_190_195_groupi_n_5392, csa_tree_add_190_195_groupi_n_5393, csa_tree_add_190_195_groupi_n_5394, csa_tree_add_190_195_groupi_n_5395, csa_tree_add_190_195_groupi_n_5396, csa_tree_add_190_195_groupi_n_5397, csa_tree_add_190_195_groupi_n_5398, csa_tree_add_190_195_groupi_n_5399;
  wire csa_tree_add_190_195_groupi_n_5400, csa_tree_add_190_195_groupi_n_5401, csa_tree_add_190_195_groupi_n_5402, csa_tree_add_190_195_groupi_n_5403, csa_tree_add_190_195_groupi_n_5404, csa_tree_add_190_195_groupi_n_5405, csa_tree_add_190_195_groupi_n_5406, csa_tree_add_190_195_groupi_n_5407;
  wire csa_tree_add_190_195_groupi_n_5408, csa_tree_add_190_195_groupi_n_5409, csa_tree_add_190_195_groupi_n_5410, csa_tree_add_190_195_groupi_n_5411, csa_tree_add_190_195_groupi_n_5412, csa_tree_add_190_195_groupi_n_5413, csa_tree_add_190_195_groupi_n_5414, csa_tree_add_190_195_groupi_n_5415;
  wire csa_tree_add_190_195_groupi_n_5416, csa_tree_add_190_195_groupi_n_5417, csa_tree_add_190_195_groupi_n_5418, csa_tree_add_190_195_groupi_n_5419, csa_tree_add_190_195_groupi_n_5420, csa_tree_add_190_195_groupi_n_5421, csa_tree_add_190_195_groupi_n_5422, csa_tree_add_190_195_groupi_n_5423;
  wire csa_tree_add_190_195_groupi_n_5424, csa_tree_add_190_195_groupi_n_5425, csa_tree_add_190_195_groupi_n_5426, csa_tree_add_190_195_groupi_n_5427, csa_tree_add_190_195_groupi_n_5428, csa_tree_add_190_195_groupi_n_5429, csa_tree_add_190_195_groupi_n_5430, csa_tree_add_190_195_groupi_n_5431;
  wire csa_tree_add_190_195_groupi_n_5432, csa_tree_add_190_195_groupi_n_5433, csa_tree_add_190_195_groupi_n_5434, csa_tree_add_190_195_groupi_n_5435, csa_tree_add_190_195_groupi_n_5436, csa_tree_add_190_195_groupi_n_5437, csa_tree_add_190_195_groupi_n_5438, csa_tree_add_190_195_groupi_n_5439;
  wire csa_tree_add_190_195_groupi_n_5440, csa_tree_add_190_195_groupi_n_5441, csa_tree_add_190_195_groupi_n_5442, csa_tree_add_190_195_groupi_n_5443, csa_tree_add_190_195_groupi_n_5444, csa_tree_add_190_195_groupi_n_5445, csa_tree_add_190_195_groupi_n_5446, csa_tree_add_190_195_groupi_n_5447;
  wire csa_tree_add_190_195_groupi_n_5448, csa_tree_add_190_195_groupi_n_5449, csa_tree_add_190_195_groupi_n_5450, csa_tree_add_190_195_groupi_n_5451, csa_tree_add_190_195_groupi_n_5452, csa_tree_add_190_195_groupi_n_5453, csa_tree_add_190_195_groupi_n_5454, csa_tree_add_190_195_groupi_n_5455;
  wire csa_tree_add_190_195_groupi_n_5456, csa_tree_add_190_195_groupi_n_5457, csa_tree_add_190_195_groupi_n_5458, csa_tree_add_190_195_groupi_n_5459, csa_tree_add_190_195_groupi_n_5460, csa_tree_add_190_195_groupi_n_5461, csa_tree_add_190_195_groupi_n_5462, csa_tree_add_190_195_groupi_n_5463;
  wire csa_tree_add_190_195_groupi_n_5464, csa_tree_add_190_195_groupi_n_5465, csa_tree_add_190_195_groupi_n_5466, csa_tree_add_190_195_groupi_n_5467, csa_tree_add_190_195_groupi_n_5468, csa_tree_add_190_195_groupi_n_5469, csa_tree_add_190_195_groupi_n_5470, csa_tree_add_190_195_groupi_n_5471;
  wire csa_tree_add_190_195_groupi_n_5472, csa_tree_add_190_195_groupi_n_5473, csa_tree_add_190_195_groupi_n_5474, csa_tree_add_190_195_groupi_n_5475, csa_tree_add_190_195_groupi_n_5476, csa_tree_add_190_195_groupi_n_5477, csa_tree_add_190_195_groupi_n_5478, csa_tree_add_190_195_groupi_n_5479;
  wire csa_tree_add_190_195_groupi_n_5480, csa_tree_add_190_195_groupi_n_5481, csa_tree_add_190_195_groupi_n_5482, csa_tree_add_190_195_groupi_n_5483, csa_tree_add_190_195_groupi_n_5484, csa_tree_add_190_195_groupi_n_5485, csa_tree_add_190_195_groupi_n_5486, csa_tree_add_190_195_groupi_n_5487;
  wire csa_tree_add_190_195_groupi_n_5488, csa_tree_add_190_195_groupi_n_5489, csa_tree_add_190_195_groupi_n_5490, csa_tree_add_190_195_groupi_n_5491, csa_tree_add_190_195_groupi_n_5492, csa_tree_add_190_195_groupi_n_5493, csa_tree_add_190_195_groupi_n_5494, csa_tree_add_190_195_groupi_n_5495;
  wire csa_tree_add_190_195_groupi_n_5496, csa_tree_add_190_195_groupi_n_5497, csa_tree_add_190_195_groupi_n_5498, csa_tree_add_190_195_groupi_n_5499, csa_tree_add_190_195_groupi_n_5500, csa_tree_add_190_195_groupi_n_5501, csa_tree_add_190_195_groupi_n_5502, csa_tree_add_190_195_groupi_n_5503;
  wire csa_tree_add_190_195_groupi_n_5504, csa_tree_add_190_195_groupi_n_5505, csa_tree_add_190_195_groupi_n_5506, csa_tree_add_190_195_groupi_n_5507, csa_tree_add_190_195_groupi_n_5508, csa_tree_add_190_195_groupi_n_5509, csa_tree_add_190_195_groupi_n_5510, csa_tree_add_190_195_groupi_n_5511;
  wire csa_tree_add_190_195_groupi_n_5512, csa_tree_add_190_195_groupi_n_5513, csa_tree_add_190_195_groupi_n_5514, csa_tree_add_190_195_groupi_n_5515, csa_tree_add_190_195_groupi_n_5516, csa_tree_add_190_195_groupi_n_5517, csa_tree_add_190_195_groupi_n_5518, csa_tree_add_190_195_groupi_n_5519;
  wire csa_tree_add_190_195_groupi_n_5520, csa_tree_add_190_195_groupi_n_5521, csa_tree_add_190_195_groupi_n_5522, csa_tree_add_190_195_groupi_n_5523, csa_tree_add_190_195_groupi_n_5524, csa_tree_add_190_195_groupi_n_5525, csa_tree_add_190_195_groupi_n_5526, csa_tree_add_190_195_groupi_n_5527;
  wire csa_tree_add_190_195_groupi_n_5528, csa_tree_add_190_195_groupi_n_5529, csa_tree_add_190_195_groupi_n_5530, csa_tree_add_190_195_groupi_n_5531, csa_tree_add_190_195_groupi_n_5532, csa_tree_add_190_195_groupi_n_5533, csa_tree_add_190_195_groupi_n_5534, csa_tree_add_190_195_groupi_n_5535;
  wire csa_tree_add_190_195_groupi_n_5536, csa_tree_add_190_195_groupi_n_5537, csa_tree_add_190_195_groupi_n_5538, csa_tree_add_190_195_groupi_n_5539, csa_tree_add_190_195_groupi_n_5540, csa_tree_add_190_195_groupi_n_5541, csa_tree_add_190_195_groupi_n_5542, csa_tree_add_190_195_groupi_n_5543;
  wire csa_tree_add_190_195_groupi_n_5544, csa_tree_add_190_195_groupi_n_5545, csa_tree_add_190_195_groupi_n_5546, csa_tree_add_190_195_groupi_n_5547, csa_tree_add_190_195_groupi_n_5548, csa_tree_add_190_195_groupi_n_5549, csa_tree_add_190_195_groupi_n_5550, csa_tree_add_190_195_groupi_n_5551;
  wire csa_tree_add_190_195_groupi_n_5552, csa_tree_add_190_195_groupi_n_5553, csa_tree_add_190_195_groupi_n_5554, csa_tree_add_190_195_groupi_n_5555, csa_tree_add_190_195_groupi_n_5556, csa_tree_add_190_195_groupi_n_5557, csa_tree_add_190_195_groupi_n_5558, csa_tree_add_190_195_groupi_n_5559;
  wire csa_tree_add_190_195_groupi_n_5560, csa_tree_add_190_195_groupi_n_5561, csa_tree_add_190_195_groupi_n_5562, csa_tree_add_190_195_groupi_n_5563, csa_tree_add_190_195_groupi_n_5564, csa_tree_add_190_195_groupi_n_5565, csa_tree_add_190_195_groupi_n_5566, csa_tree_add_190_195_groupi_n_5567;
  wire csa_tree_add_190_195_groupi_n_5568, csa_tree_add_190_195_groupi_n_5569, csa_tree_add_190_195_groupi_n_5570, csa_tree_add_190_195_groupi_n_5571, csa_tree_add_190_195_groupi_n_5572, csa_tree_add_190_195_groupi_n_5573, csa_tree_add_190_195_groupi_n_5574, csa_tree_add_190_195_groupi_n_5575;
  wire csa_tree_add_190_195_groupi_n_5576, csa_tree_add_190_195_groupi_n_5577, csa_tree_add_190_195_groupi_n_5578, csa_tree_add_190_195_groupi_n_5579, csa_tree_add_190_195_groupi_n_5580, csa_tree_add_190_195_groupi_n_5581, csa_tree_add_190_195_groupi_n_5582, csa_tree_add_190_195_groupi_n_5583;
  wire csa_tree_add_190_195_groupi_n_5584, csa_tree_add_190_195_groupi_n_5585, csa_tree_add_190_195_groupi_n_5586, csa_tree_add_190_195_groupi_n_5587, csa_tree_add_190_195_groupi_n_5588, csa_tree_add_190_195_groupi_n_5589, csa_tree_add_190_195_groupi_n_5590, csa_tree_add_190_195_groupi_n_5591;
  wire csa_tree_add_190_195_groupi_n_5592, csa_tree_add_190_195_groupi_n_5593, csa_tree_add_190_195_groupi_n_5594, csa_tree_add_190_195_groupi_n_5595, csa_tree_add_190_195_groupi_n_5596, csa_tree_add_190_195_groupi_n_5597, csa_tree_add_190_195_groupi_n_5598, csa_tree_add_190_195_groupi_n_5599;
  wire csa_tree_add_190_195_groupi_n_5600, csa_tree_add_190_195_groupi_n_5601, csa_tree_add_190_195_groupi_n_5602, csa_tree_add_190_195_groupi_n_5603, csa_tree_add_190_195_groupi_n_5604, csa_tree_add_190_195_groupi_n_5605, csa_tree_add_190_195_groupi_n_5606, csa_tree_add_190_195_groupi_n_5607;
  wire csa_tree_add_190_195_groupi_n_5608, csa_tree_add_190_195_groupi_n_5609, csa_tree_add_190_195_groupi_n_5610, csa_tree_add_190_195_groupi_n_5611, csa_tree_add_190_195_groupi_n_5612, csa_tree_add_190_195_groupi_n_5613, csa_tree_add_190_195_groupi_n_5614, csa_tree_add_190_195_groupi_n_5615;
  wire csa_tree_add_190_195_groupi_n_5616, csa_tree_add_190_195_groupi_n_5617, csa_tree_add_190_195_groupi_n_5618, csa_tree_add_190_195_groupi_n_5619, csa_tree_add_190_195_groupi_n_5620, csa_tree_add_190_195_groupi_n_5621, csa_tree_add_190_195_groupi_n_5622, csa_tree_add_190_195_groupi_n_5623;
  wire csa_tree_add_190_195_groupi_n_5624, csa_tree_add_190_195_groupi_n_5625, csa_tree_add_190_195_groupi_n_5626, csa_tree_add_190_195_groupi_n_5627, csa_tree_add_190_195_groupi_n_5628, csa_tree_add_190_195_groupi_n_5629, csa_tree_add_190_195_groupi_n_5630, csa_tree_add_190_195_groupi_n_5631;
  wire csa_tree_add_190_195_groupi_n_5632, csa_tree_add_190_195_groupi_n_5633, csa_tree_add_190_195_groupi_n_5634, csa_tree_add_190_195_groupi_n_5635, csa_tree_add_190_195_groupi_n_5636, csa_tree_add_190_195_groupi_n_5637, csa_tree_add_190_195_groupi_n_5638, csa_tree_add_190_195_groupi_n_5639;
  wire csa_tree_add_190_195_groupi_n_5640, csa_tree_add_190_195_groupi_n_5641, csa_tree_add_190_195_groupi_n_5642, csa_tree_add_190_195_groupi_n_5643, csa_tree_add_190_195_groupi_n_5644, csa_tree_add_190_195_groupi_n_5645, csa_tree_add_190_195_groupi_n_5646, csa_tree_add_190_195_groupi_n_5647;
  wire csa_tree_add_190_195_groupi_n_5648, csa_tree_add_190_195_groupi_n_5649, csa_tree_add_190_195_groupi_n_5650, csa_tree_add_190_195_groupi_n_5651, csa_tree_add_190_195_groupi_n_5652, csa_tree_add_190_195_groupi_n_5653, csa_tree_add_190_195_groupi_n_5654, csa_tree_add_190_195_groupi_n_5655;
  wire csa_tree_add_190_195_groupi_n_5656, csa_tree_add_190_195_groupi_n_5657, csa_tree_add_190_195_groupi_n_5658, csa_tree_add_190_195_groupi_n_5659, csa_tree_add_190_195_groupi_n_5660, csa_tree_add_190_195_groupi_n_5661, csa_tree_add_190_195_groupi_n_5662, csa_tree_add_190_195_groupi_n_5663;
  wire csa_tree_add_190_195_groupi_n_5664, csa_tree_add_190_195_groupi_n_5665, csa_tree_add_190_195_groupi_n_5666, csa_tree_add_190_195_groupi_n_5667, csa_tree_add_190_195_groupi_n_5668, csa_tree_add_190_195_groupi_n_5669, csa_tree_add_190_195_groupi_n_5670, csa_tree_add_190_195_groupi_n_5671;
  wire csa_tree_add_190_195_groupi_n_5672, csa_tree_add_190_195_groupi_n_5673, csa_tree_add_190_195_groupi_n_5674, csa_tree_add_190_195_groupi_n_5675, csa_tree_add_190_195_groupi_n_5676, csa_tree_add_190_195_groupi_n_5677, csa_tree_add_190_195_groupi_n_5678, csa_tree_add_190_195_groupi_n_5679;
  wire csa_tree_add_190_195_groupi_n_5680, csa_tree_add_190_195_groupi_n_5681, csa_tree_add_190_195_groupi_n_5682, csa_tree_add_190_195_groupi_n_5683, csa_tree_add_190_195_groupi_n_5684, csa_tree_add_190_195_groupi_n_5685, csa_tree_add_190_195_groupi_n_5686, csa_tree_add_190_195_groupi_n_5687;
  wire csa_tree_add_190_195_groupi_n_5688, csa_tree_add_190_195_groupi_n_5689, csa_tree_add_190_195_groupi_n_5690, csa_tree_add_190_195_groupi_n_5691, csa_tree_add_190_195_groupi_n_5692, csa_tree_add_190_195_groupi_n_5693, csa_tree_add_190_195_groupi_n_5694, csa_tree_add_190_195_groupi_n_5695;
  wire csa_tree_add_190_195_groupi_n_5696, csa_tree_add_190_195_groupi_n_5697, csa_tree_add_190_195_groupi_n_5698, csa_tree_add_190_195_groupi_n_5699, csa_tree_add_190_195_groupi_n_5700, csa_tree_add_190_195_groupi_n_5701, csa_tree_add_190_195_groupi_n_5702, csa_tree_add_190_195_groupi_n_5703;
  wire csa_tree_add_190_195_groupi_n_5704, csa_tree_add_190_195_groupi_n_5705, csa_tree_add_190_195_groupi_n_5706, csa_tree_add_190_195_groupi_n_5707, csa_tree_add_190_195_groupi_n_5708, csa_tree_add_190_195_groupi_n_5709, csa_tree_add_190_195_groupi_n_5710, csa_tree_add_190_195_groupi_n_5711;
  wire csa_tree_add_190_195_groupi_n_5712, csa_tree_add_190_195_groupi_n_5713, csa_tree_add_190_195_groupi_n_5714, csa_tree_add_190_195_groupi_n_5715, csa_tree_add_190_195_groupi_n_5716, csa_tree_add_190_195_groupi_n_5717, csa_tree_add_190_195_groupi_n_5718, csa_tree_add_190_195_groupi_n_5719;
  wire csa_tree_add_190_195_groupi_n_5720, csa_tree_add_190_195_groupi_n_5721, csa_tree_add_190_195_groupi_n_5722, csa_tree_add_190_195_groupi_n_5723, csa_tree_add_190_195_groupi_n_5724, csa_tree_add_190_195_groupi_n_5725, csa_tree_add_190_195_groupi_n_5726, csa_tree_add_190_195_groupi_n_5727;
  wire csa_tree_add_190_195_groupi_n_5728, csa_tree_add_190_195_groupi_n_5729, csa_tree_add_190_195_groupi_n_5730, csa_tree_add_190_195_groupi_n_5731, csa_tree_add_190_195_groupi_n_5732, csa_tree_add_190_195_groupi_n_5733, csa_tree_add_190_195_groupi_n_5734, csa_tree_add_190_195_groupi_n_5735;
  wire csa_tree_add_190_195_groupi_n_5736, csa_tree_add_190_195_groupi_n_5737, csa_tree_add_190_195_groupi_n_5738, csa_tree_add_190_195_groupi_n_5739, csa_tree_add_190_195_groupi_n_5740, csa_tree_add_190_195_groupi_n_5741, csa_tree_add_190_195_groupi_n_5742, csa_tree_add_190_195_groupi_n_5743;
  wire csa_tree_add_190_195_groupi_n_5744, csa_tree_add_190_195_groupi_n_5745, csa_tree_add_190_195_groupi_n_5746, csa_tree_add_190_195_groupi_n_5747, csa_tree_add_190_195_groupi_n_5748, csa_tree_add_190_195_groupi_n_5749, csa_tree_add_190_195_groupi_n_5750, csa_tree_add_190_195_groupi_n_5751;
  wire csa_tree_add_190_195_groupi_n_5752, csa_tree_add_190_195_groupi_n_5753, csa_tree_add_190_195_groupi_n_5754, csa_tree_add_190_195_groupi_n_5755, csa_tree_add_190_195_groupi_n_5756, csa_tree_add_190_195_groupi_n_5757, csa_tree_add_190_195_groupi_n_5758, csa_tree_add_190_195_groupi_n_5759;
  wire csa_tree_add_190_195_groupi_n_5760, csa_tree_add_190_195_groupi_n_5761, csa_tree_add_190_195_groupi_n_5762, csa_tree_add_190_195_groupi_n_5763, csa_tree_add_190_195_groupi_n_5764, csa_tree_add_190_195_groupi_n_5765, csa_tree_add_190_195_groupi_n_5766, csa_tree_add_190_195_groupi_n_5767;
  wire csa_tree_add_190_195_groupi_n_5768, csa_tree_add_190_195_groupi_n_5769, csa_tree_add_190_195_groupi_n_5770, csa_tree_add_190_195_groupi_n_5771, csa_tree_add_190_195_groupi_n_5772, csa_tree_add_190_195_groupi_n_5773, csa_tree_add_190_195_groupi_n_5774, csa_tree_add_190_195_groupi_n_5775;
  wire csa_tree_add_190_195_groupi_n_5776, csa_tree_add_190_195_groupi_n_5777, csa_tree_add_190_195_groupi_n_5778, csa_tree_add_190_195_groupi_n_5779, csa_tree_add_190_195_groupi_n_5780, csa_tree_add_190_195_groupi_n_5781, csa_tree_add_190_195_groupi_n_5782, csa_tree_add_190_195_groupi_n_5783;
  wire csa_tree_add_190_195_groupi_n_5784, csa_tree_add_190_195_groupi_n_5785, csa_tree_add_190_195_groupi_n_5786, csa_tree_add_190_195_groupi_n_5787, csa_tree_add_190_195_groupi_n_5788, csa_tree_add_190_195_groupi_n_5789, csa_tree_add_190_195_groupi_n_5790, csa_tree_add_190_195_groupi_n_5791;
  wire csa_tree_add_190_195_groupi_n_5792, csa_tree_add_190_195_groupi_n_5793, csa_tree_add_190_195_groupi_n_5794, csa_tree_add_190_195_groupi_n_5795, csa_tree_add_190_195_groupi_n_5796, csa_tree_add_190_195_groupi_n_5797, csa_tree_add_190_195_groupi_n_5798, csa_tree_add_190_195_groupi_n_5799;
  wire csa_tree_add_190_195_groupi_n_5800, csa_tree_add_190_195_groupi_n_5801, csa_tree_add_190_195_groupi_n_5802, csa_tree_add_190_195_groupi_n_5803, csa_tree_add_190_195_groupi_n_5804, csa_tree_add_190_195_groupi_n_5805, csa_tree_add_190_195_groupi_n_5806, csa_tree_add_190_195_groupi_n_5807;
  wire csa_tree_add_190_195_groupi_n_5808, csa_tree_add_190_195_groupi_n_5809, csa_tree_add_190_195_groupi_n_5810, csa_tree_add_190_195_groupi_n_5811, csa_tree_add_190_195_groupi_n_5812, csa_tree_add_190_195_groupi_n_5813, csa_tree_add_190_195_groupi_n_5814, csa_tree_add_190_195_groupi_n_5815;
  wire csa_tree_add_190_195_groupi_n_5816, csa_tree_add_190_195_groupi_n_5817, csa_tree_add_190_195_groupi_n_5818, csa_tree_add_190_195_groupi_n_5819, csa_tree_add_190_195_groupi_n_5820, csa_tree_add_190_195_groupi_n_5821, csa_tree_add_190_195_groupi_n_5822, csa_tree_add_190_195_groupi_n_5823;
  wire csa_tree_add_190_195_groupi_n_5824, csa_tree_add_190_195_groupi_n_5825, csa_tree_add_190_195_groupi_n_5826, csa_tree_add_190_195_groupi_n_5827, csa_tree_add_190_195_groupi_n_5828, csa_tree_add_190_195_groupi_n_5829, csa_tree_add_190_195_groupi_n_5830, csa_tree_add_190_195_groupi_n_5831;
  wire csa_tree_add_190_195_groupi_n_5832, csa_tree_add_190_195_groupi_n_5833, csa_tree_add_190_195_groupi_n_5834, csa_tree_add_190_195_groupi_n_5835, csa_tree_add_190_195_groupi_n_5836, csa_tree_add_190_195_groupi_n_5837, csa_tree_add_190_195_groupi_n_5838, csa_tree_add_190_195_groupi_n_5839;
  wire csa_tree_add_190_195_groupi_n_5840, csa_tree_add_190_195_groupi_n_5841, csa_tree_add_190_195_groupi_n_5842, csa_tree_add_190_195_groupi_n_5843, csa_tree_add_190_195_groupi_n_5844, csa_tree_add_190_195_groupi_n_5845, csa_tree_add_190_195_groupi_n_5846, csa_tree_add_190_195_groupi_n_5847;
  wire csa_tree_add_190_195_groupi_n_5848, csa_tree_add_190_195_groupi_n_5849, csa_tree_add_190_195_groupi_n_5850, csa_tree_add_190_195_groupi_n_5851, csa_tree_add_190_195_groupi_n_5852, csa_tree_add_190_195_groupi_n_5853, csa_tree_add_190_195_groupi_n_5854, csa_tree_add_190_195_groupi_n_5855;
  wire csa_tree_add_190_195_groupi_n_5856, csa_tree_add_190_195_groupi_n_5857, csa_tree_add_190_195_groupi_n_5858, csa_tree_add_190_195_groupi_n_5859, csa_tree_add_190_195_groupi_n_5860, csa_tree_add_190_195_groupi_n_5861, csa_tree_add_190_195_groupi_n_5862, csa_tree_add_190_195_groupi_n_5863;
  wire csa_tree_add_190_195_groupi_n_5864, csa_tree_add_190_195_groupi_n_5865, csa_tree_add_190_195_groupi_n_5866, csa_tree_add_190_195_groupi_n_5867, csa_tree_add_190_195_groupi_n_5868, csa_tree_add_190_195_groupi_n_5869, csa_tree_add_190_195_groupi_n_5870, csa_tree_add_190_195_groupi_n_5871;
  wire csa_tree_add_190_195_groupi_n_5872, csa_tree_add_190_195_groupi_n_5873, csa_tree_add_190_195_groupi_n_5874, csa_tree_add_190_195_groupi_n_5875, csa_tree_add_190_195_groupi_n_5876, csa_tree_add_190_195_groupi_n_5877, csa_tree_add_190_195_groupi_n_5878, csa_tree_add_190_195_groupi_n_5879;
  wire csa_tree_add_190_195_groupi_n_5880, csa_tree_add_190_195_groupi_n_5881, csa_tree_add_190_195_groupi_n_5882, csa_tree_add_190_195_groupi_n_5883, csa_tree_add_190_195_groupi_n_5884, csa_tree_add_190_195_groupi_n_5885, csa_tree_add_190_195_groupi_n_5886, csa_tree_add_190_195_groupi_n_5887;
  wire csa_tree_add_190_195_groupi_n_5888, csa_tree_add_190_195_groupi_n_5889, csa_tree_add_190_195_groupi_n_5890, csa_tree_add_190_195_groupi_n_5891, csa_tree_add_190_195_groupi_n_5892, csa_tree_add_190_195_groupi_n_5893, csa_tree_add_190_195_groupi_n_5894, csa_tree_add_190_195_groupi_n_5895;
  wire csa_tree_add_190_195_groupi_n_5896, csa_tree_add_190_195_groupi_n_5897, csa_tree_add_190_195_groupi_n_5898, csa_tree_add_190_195_groupi_n_5899, csa_tree_add_190_195_groupi_n_5900, csa_tree_add_190_195_groupi_n_5901, csa_tree_add_190_195_groupi_n_5902, csa_tree_add_190_195_groupi_n_5903;
  wire csa_tree_add_190_195_groupi_n_5904, csa_tree_add_190_195_groupi_n_5905, csa_tree_add_190_195_groupi_n_5906, csa_tree_add_190_195_groupi_n_5907, csa_tree_add_190_195_groupi_n_5908, csa_tree_add_190_195_groupi_n_5909, csa_tree_add_190_195_groupi_n_5910, csa_tree_add_190_195_groupi_n_5911;
  wire csa_tree_add_190_195_groupi_n_5912, csa_tree_add_190_195_groupi_n_5913, csa_tree_add_190_195_groupi_n_5914, csa_tree_add_190_195_groupi_n_5915, csa_tree_add_190_195_groupi_n_5916, csa_tree_add_190_195_groupi_n_5917, csa_tree_add_190_195_groupi_n_5918, csa_tree_add_190_195_groupi_n_5919;
  wire csa_tree_add_190_195_groupi_n_5920, csa_tree_add_190_195_groupi_n_5921, csa_tree_add_190_195_groupi_n_5922, csa_tree_add_190_195_groupi_n_5923, csa_tree_add_190_195_groupi_n_5924, csa_tree_add_190_195_groupi_n_5925, csa_tree_add_190_195_groupi_n_5926, csa_tree_add_190_195_groupi_n_5927;
  wire csa_tree_add_190_195_groupi_n_5928, csa_tree_add_190_195_groupi_n_5929, csa_tree_add_190_195_groupi_n_5930, csa_tree_add_190_195_groupi_n_5931, csa_tree_add_190_195_groupi_n_5932, csa_tree_add_190_195_groupi_n_5933, csa_tree_add_190_195_groupi_n_5934, csa_tree_add_190_195_groupi_n_5935;
  wire csa_tree_add_190_195_groupi_n_5936, csa_tree_add_190_195_groupi_n_5937, csa_tree_add_190_195_groupi_n_5938, csa_tree_add_190_195_groupi_n_5939, csa_tree_add_190_195_groupi_n_5940, csa_tree_add_190_195_groupi_n_5941, csa_tree_add_190_195_groupi_n_5942, csa_tree_add_190_195_groupi_n_5943;
  wire csa_tree_add_190_195_groupi_n_5944, csa_tree_add_190_195_groupi_n_5945, csa_tree_add_190_195_groupi_n_5946, csa_tree_add_190_195_groupi_n_5947, csa_tree_add_190_195_groupi_n_5948, csa_tree_add_190_195_groupi_n_5949, csa_tree_add_190_195_groupi_n_5950, csa_tree_add_190_195_groupi_n_5951;
  wire csa_tree_add_190_195_groupi_n_5952, csa_tree_add_190_195_groupi_n_5953, csa_tree_add_190_195_groupi_n_5954, csa_tree_add_190_195_groupi_n_5955, csa_tree_add_190_195_groupi_n_5956, csa_tree_add_190_195_groupi_n_5957, csa_tree_add_190_195_groupi_n_5958, csa_tree_add_190_195_groupi_n_5959;
  wire csa_tree_add_190_195_groupi_n_5960, csa_tree_add_190_195_groupi_n_5961, csa_tree_add_190_195_groupi_n_5962, csa_tree_add_190_195_groupi_n_5963, csa_tree_add_190_195_groupi_n_5964, csa_tree_add_190_195_groupi_n_5965, csa_tree_add_190_195_groupi_n_5966, csa_tree_add_190_195_groupi_n_5967;
  wire csa_tree_add_190_195_groupi_n_5968, csa_tree_add_190_195_groupi_n_5969, csa_tree_add_190_195_groupi_n_5970, csa_tree_add_190_195_groupi_n_5971, csa_tree_add_190_195_groupi_n_5972, csa_tree_add_190_195_groupi_n_5973, csa_tree_add_190_195_groupi_n_5974, csa_tree_add_190_195_groupi_n_5975;
  wire csa_tree_add_190_195_groupi_n_5976, csa_tree_add_190_195_groupi_n_5977, csa_tree_add_190_195_groupi_n_5978, csa_tree_add_190_195_groupi_n_5979, csa_tree_add_190_195_groupi_n_5980, csa_tree_add_190_195_groupi_n_5981, csa_tree_add_190_195_groupi_n_5982, csa_tree_add_190_195_groupi_n_5983;
  wire csa_tree_add_190_195_groupi_n_5984, csa_tree_add_190_195_groupi_n_5985, csa_tree_add_190_195_groupi_n_5986, csa_tree_add_190_195_groupi_n_5987, csa_tree_add_190_195_groupi_n_5988, csa_tree_add_190_195_groupi_n_5989, csa_tree_add_190_195_groupi_n_5990, csa_tree_add_190_195_groupi_n_5991;
  wire csa_tree_add_190_195_groupi_n_5992, csa_tree_add_190_195_groupi_n_5993, csa_tree_add_190_195_groupi_n_5994, csa_tree_add_190_195_groupi_n_5995, csa_tree_add_190_195_groupi_n_5996, csa_tree_add_190_195_groupi_n_5997, csa_tree_add_190_195_groupi_n_5998, csa_tree_add_190_195_groupi_n_5999;
  wire csa_tree_add_190_195_groupi_n_6000, csa_tree_add_190_195_groupi_n_6001, csa_tree_add_190_195_groupi_n_6002, csa_tree_add_190_195_groupi_n_6003, csa_tree_add_190_195_groupi_n_6004, csa_tree_add_190_195_groupi_n_6005, csa_tree_add_190_195_groupi_n_6006, csa_tree_add_190_195_groupi_n_6007;
  wire csa_tree_add_190_195_groupi_n_6008, csa_tree_add_190_195_groupi_n_6009, csa_tree_add_190_195_groupi_n_6010, csa_tree_add_190_195_groupi_n_6011, csa_tree_add_190_195_groupi_n_6012, csa_tree_add_190_195_groupi_n_6013, csa_tree_add_190_195_groupi_n_6014, csa_tree_add_190_195_groupi_n_6015;
  wire csa_tree_add_190_195_groupi_n_6016, csa_tree_add_190_195_groupi_n_6017, csa_tree_add_190_195_groupi_n_6018, csa_tree_add_190_195_groupi_n_6019, csa_tree_add_190_195_groupi_n_6020, csa_tree_add_190_195_groupi_n_6021, csa_tree_add_190_195_groupi_n_6022, csa_tree_add_190_195_groupi_n_6023;
  wire csa_tree_add_190_195_groupi_n_6024, csa_tree_add_190_195_groupi_n_6025, csa_tree_add_190_195_groupi_n_6026, csa_tree_add_190_195_groupi_n_6027, csa_tree_add_190_195_groupi_n_6028, csa_tree_add_190_195_groupi_n_6029, csa_tree_add_190_195_groupi_n_6030, csa_tree_add_190_195_groupi_n_6031;
  wire csa_tree_add_190_195_groupi_n_6032, csa_tree_add_190_195_groupi_n_6033, csa_tree_add_190_195_groupi_n_6034, csa_tree_add_190_195_groupi_n_6035, csa_tree_add_190_195_groupi_n_6036, csa_tree_add_190_195_groupi_n_6037, csa_tree_add_190_195_groupi_n_6038, csa_tree_add_190_195_groupi_n_6039;
  wire csa_tree_add_190_195_groupi_n_6040, csa_tree_add_190_195_groupi_n_6041, csa_tree_add_190_195_groupi_n_6042, csa_tree_add_190_195_groupi_n_6043, csa_tree_add_190_195_groupi_n_6044, csa_tree_add_190_195_groupi_n_6045, csa_tree_add_190_195_groupi_n_6046, csa_tree_add_190_195_groupi_n_6047;
  wire csa_tree_add_190_195_groupi_n_6048, csa_tree_add_190_195_groupi_n_6049, csa_tree_add_190_195_groupi_n_6050, csa_tree_add_190_195_groupi_n_6051, csa_tree_add_190_195_groupi_n_6052, csa_tree_add_190_195_groupi_n_6053, csa_tree_add_190_195_groupi_n_6054, csa_tree_add_190_195_groupi_n_6055;
  wire csa_tree_add_190_195_groupi_n_6056, csa_tree_add_190_195_groupi_n_6057, csa_tree_add_190_195_groupi_n_6058, csa_tree_add_190_195_groupi_n_6059, csa_tree_add_190_195_groupi_n_6060, csa_tree_add_190_195_groupi_n_6061, csa_tree_add_190_195_groupi_n_6062, csa_tree_add_190_195_groupi_n_6063;
  wire csa_tree_add_190_195_groupi_n_6064, csa_tree_add_190_195_groupi_n_6065, csa_tree_add_190_195_groupi_n_6066, csa_tree_add_190_195_groupi_n_6067, csa_tree_add_190_195_groupi_n_6068, csa_tree_add_190_195_groupi_n_6069, csa_tree_add_190_195_groupi_n_6070, csa_tree_add_190_195_groupi_n_6071;
  wire csa_tree_add_190_195_groupi_n_6072, csa_tree_add_190_195_groupi_n_6073, csa_tree_add_190_195_groupi_n_6074, csa_tree_add_190_195_groupi_n_6075, csa_tree_add_190_195_groupi_n_6076, csa_tree_add_190_195_groupi_n_6077, csa_tree_add_190_195_groupi_n_6078, csa_tree_add_190_195_groupi_n_6079;
  wire csa_tree_add_190_195_groupi_n_6080, csa_tree_add_190_195_groupi_n_6081, csa_tree_add_190_195_groupi_n_6082, csa_tree_add_190_195_groupi_n_6083, csa_tree_add_190_195_groupi_n_6084, csa_tree_add_190_195_groupi_n_6085, csa_tree_add_190_195_groupi_n_6086, csa_tree_add_190_195_groupi_n_6087;
  wire csa_tree_add_190_195_groupi_n_6088, csa_tree_add_190_195_groupi_n_6089, csa_tree_add_190_195_groupi_n_6090, csa_tree_add_190_195_groupi_n_6091, csa_tree_add_190_195_groupi_n_6092, csa_tree_add_190_195_groupi_n_6093, csa_tree_add_190_195_groupi_n_6094, csa_tree_add_190_195_groupi_n_6095;
  wire csa_tree_add_190_195_groupi_n_6096, csa_tree_add_190_195_groupi_n_6097, csa_tree_add_190_195_groupi_n_6098, csa_tree_add_190_195_groupi_n_6099, csa_tree_add_190_195_groupi_n_6100, csa_tree_add_190_195_groupi_n_6101, csa_tree_add_190_195_groupi_n_6102, csa_tree_add_190_195_groupi_n_6103;
  wire csa_tree_add_190_195_groupi_n_6104, csa_tree_add_190_195_groupi_n_6105, csa_tree_add_190_195_groupi_n_6106, csa_tree_add_190_195_groupi_n_6107, csa_tree_add_190_195_groupi_n_6108, csa_tree_add_190_195_groupi_n_6109, csa_tree_add_190_195_groupi_n_6110, csa_tree_add_190_195_groupi_n_6111;
  wire csa_tree_add_190_195_groupi_n_6112, csa_tree_add_190_195_groupi_n_6113, csa_tree_add_190_195_groupi_n_6114, csa_tree_add_190_195_groupi_n_6115, csa_tree_add_190_195_groupi_n_6116, csa_tree_add_190_195_groupi_n_6117, csa_tree_add_190_195_groupi_n_6118, csa_tree_add_190_195_groupi_n_6119;
  wire csa_tree_add_190_195_groupi_n_6120, csa_tree_add_190_195_groupi_n_6121, csa_tree_add_190_195_groupi_n_6122, csa_tree_add_190_195_groupi_n_6123, csa_tree_add_190_195_groupi_n_6124, csa_tree_add_190_195_groupi_n_6125, csa_tree_add_190_195_groupi_n_6126, csa_tree_add_190_195_groupi_n_6127;
  wire csa_tree_add_190_195_groupi_n_6128, csa_tree_add_190_195_groupi_n_6129, csa_tree_add_190_195_groupi_n_6130, csa_tree_add_190_195_groupi_n_6131, csa_tree_add_190_195_groupi_n_6132, csa_tree_add_190_195_groupi_n_6133, csa_tree_add_190_195_groupi_n_6134, csa_tree_add_190_195_groupi_n_6135;
  wire csa_tree_add_190_195_groupi_n_6136, csa_tree_add_190_195_groupi_n_6137, csa_tree_add_190_195_groupi_n_6138, csa_tree_add_190_195_groupi_n_6139, csa_tree_add_190_195_groupi_n_6140, csa_tree_add_190_195_groupi_n_6141, csa_tree_add_190_195_groupi_n_6142, csa_tree_add_190_195_groupi_n_6143;
  wire csa_tree_add_190_195_groupi_n_6144, csa_tree_add_190_195_groupi_n_6145, csa_tree_add_190_195_groupi_n_6146, csa_tree_add_190_195_groupi_n_6147, csa_tree_add_190_195_groupi_n_6148, csa_tree_add_190_195_groupi_n_6149, csa_tree_add_190_195_groupi_n_6150, csa_tree_add_190_195_groupi_n_6151;
  wire csa_tree_add_190_195_groupi_n_6152, csa_tree_add_190_195_groupi_n_6153, csa_tree_add_190_195_groupi_n_6154, csa_tree_add_190_195_groupi_n_6155, csa_tree_add_190_195_groupi_n_6156, csa_tree_add_190_195_groupi_n_6157, csa_tree_add_190_195_groupi_n_6158, csa_tree_add_190_195_groupi_n_6159;
  wire csa_tree_add_190_195_groupi_n_6160, csa_tree_add_190_195_groupi_n_6161, csa_tree_add_190_195_groupi_n_6162, csa_tree_add_190_195_groupi_n_6163, csa_tree_add_190_195_groupi_n_6164, csa_tree_add_190_195_groupi_n_6165, csa_tree_add_190_195_groupi_n_6166, csa_tree_add_190_195_groupi_n_6167;
  wire csa_tree_add_190_195_groupi_n_6168, csa_tree_add_190_195_groupi_n_6169, csa_tree_add_190_195_groupi_n_6170, csa_tree_add_190_195_groupi_n_6171, csa_tree_add_190_195_groupi_n_6172, csa_tree_add_190_195_groupi_n_6173, csa_tree_add_190_195_groupi_n_6174, csa_tree_add_190_195_groupi_n_6175;
  wire csa_tree_add_190_195_groupi_n_6176, csa_tree_add_190_195_groupi_n_6177, csa_tree_add_190_195_groupi_n_6178, csa_tree_add_190_195_groupi_n_6179, csa_tree_add_190_195_groupi_n_6180, csa_tree_add_190_195_groupi_n_6181, csa_tree_add_190_195_groupi_n_6182, csa_tree_add_190_195_groupi_n_6183;
  wire csa_tree_add_190_195_groupi_n_6184, csa_tree_add_190_195_groupi_n_6185, csa_tree_add_190_195_groupi_n_6186, csa_tree_add_190_195_groupi_n_6187, csa_tree_add_190_195_groupi_n_6188, csa_tree_add_190_195_groupi_n_6189, csa_tree_add_190_195_groupi_n_6190, csa_tree_add_190_195_groupi_n_6191;
  wire csa_tree_add_190_195_groupi_n_6192, csa_tree_add_190_195_groupi_n_6193, csa_tree_add_190_195_groupi_n_6194, csa_tree_add_190_195_groupi_n_6195, csa_tree_add_190_195_groupi_n_6196, csa_tree_add_190_195_groupi_n_6197, csa_tree_add_190_195_groupi_n_6198, csa_tree_add_190_195_groupi_n_6199;
  wire csa_tree_add_190_195_groupi_n_6200, csa_tree_add_190_195_groupi_n_6201, csa_tree_add_190_195_groupi_n_6202, csa_tree_add_190_195_groupi_n_6203, csa_tree_add_190_195_groupi_n_6204, csa_tree_add_190_195_groupi_n_6205, csa_tree_add_190_195_groupi_n_6206, csa_tree_add_190_195_groupi_n_6207;
  wire csa_tree_add_190_195_groupi_n_6208, csa_tree_add_190_195_groupi_n_6209, csa_tree_add_190_195_groupi_n_6210, csa_tree_add_190_195_groupi_n_6211, csa_tree_add_190_195_groupi_n_6212, csa_tree_add_190_195_groupi_n_6213, csa_tree_add_190_195_groupi_n_6214, csa_tree_add_190_195_groupi_n_6215;
  wire csa_tree_add_190_195_groupi_n_6216, csa_tree_add_190_195_groupi_n_6217, csa_tree_add_190_195_groupi_n_6218, csa_tree_add_190_195_groupi_n_6219, csa_tree_add_190_195_groupi_n_6220, csa_tree_add_190_195_groupi_n_6221, csa_tree_add_190_195_groupi_n_6222, csa_tree_add_190_195_groupi_n_6223;
  wire csa_tree_add_190_195_groupi_n_6224, csa_tree_add_190_195_groupi_n_6225, csa_tree_add_190_195_groupi_n_6226, csa_tree_add_190_195_groupi_n_6227, csa_tree_add_190_195_groupi_n_6228, csa_tree_add_190_195_groupi_n_6229, csa_tree_add_190_195_groupi_n_6230, csa_tree_add_190_195_groupi_n_6231;
  wire csa_tree_add_190_195_groupi_n_6232, csa_tree_add_190_195_groupi_n_6233, csa_tree_add_190_195_groupi_n_6234, csa_tree_add_190_195_groupi_n_6235, csa_tree_add_190_195_groupi_n_6236, csa_tree_add_190_195_groupi_n_6237, csa_tree_add_190_195_groupi_n_6238, csa_tree_add_190_195_groupi_n_6239;
  wire csa_tree_add_190_195_groupi_n_6240, csa_tree_add_190_195_groupi_n_6241, csa_tree_add_190_195_groupi_n_6242, csa_tree_add_190_195_groupi_n_6243, csa_tree_add_190_195_groupi_n_6244, csa_tree_add_190_195_groupi_n_6245, csa_tree_add_190_195_groupi_n_6246, csa_tree_add_190_195_groupi_n_6247;
  wire csa_tree_add_190_195_groupi_n_6248, csa_tree_add_190_195_groupi_n_6249, csa_tree_add_190_195_groupi_n_6250, csa_tree_add_190_195_groupi_n_6251, csa_tree_add_190_195_groupi_n_6252, csa_tree_add_190_195_groupi_n_6253, csa_tree_add_190_195_groupi_n_6254, csa_tree_add_190_195_groupi_n_6255;
  wire csa_tree_add_190_195_groupi_n_6256, csa_tree_add_190_195_groupi_n_6257, csa_tree_add_190_195_groupi_n_6258, csa_tree_add_190_195_groupi_n_6259, csa_tree_add_190_195_groupi_n_6260, csa_tree_add_190_195_groupi_n_6261, csa_tree_add_190_195_groupi_n_6262, csa_tree_add_190_195_groupi_n_6263;
  wire csa_tree_add_190_195_groupi_n_6264, csa_tree_add_190_195_groupi_n_6265, csa_tree_add_190_195_groupi_n_6266, csa_tree_add_190_195_groupi_n_6267, csa_tree_add_190_195_groupi_n_6268, csa_tree_add_190_195_groupi_n_6269, csa_tree_add_190_195_groupi_n_6270, csa_tree_add_190_195_groupi_n_6271;
  wire csa_tree_add_190_195_groupi_n_6272, csa_tree_add_190_195_groupi_n_6273, csa_tree_add_190_195_groupi_n_6274, csa_tree_add_190_195_groupi_n_6275, csa_tree_add_190_195_groupi_n_6276, csa_tree_add_190_195_groupi_n_6277, csa_tree_add_190_195_groupi_n_6278, csa_tree_add_190_195_groupi_n_6279;
  wire csa_tree_add_190_195_groupi_n_6280, csa_tree_add_190_195_groupi_n_6281, csa_tree_add_190_195_groupi_n_6282, csa_tree_add_190_195_groupi_n_6283, csa_tree_add_190_195_groupi_n_6284, csa_tree_add_190_195_groupi_n_6285, csa_tree_add_190_195_groupi_n_6286, csa_tree_add_190_195_groupi_n_6287;
  wire csa_tree_add_190_195_groupi_n_6288, csa_tree_add_190_195_groupi_n_6289, csa_tree_add_190_195_groupi_n_6290, csa_tree_add_190_195_groupi_n_6291, csa_tree_add_190_195_groupi_n_6292, csa_tree_add_190_195_groupi_n_6293, csa_tree_add_190_195_groupi_n_6294, csa_tree_add_190_195_groupi_n_6295;
  wire csa_tree_add_190_195_groupi_n_6296, csa_tree_add_190_195_groupi_n_6297, csa_tree_add_190_195_groupi_n_6298, csa_tree_add_190_195_groupi_n_6299, csa_tree_add_190_195_groupi_n_6300, csa_tree_add_190_195_groupi_n_6301, csa_tree_add_190_195_groupi_n_6302, csa_tree_add_190_195_groupi_n_6303;
  wire csa_tree_add_190_195_groupi_n_6304, csa_tree_add_190_195_groupi_n_6305, csa_tree_add_190_195_groupi_n_6306, csa_tree_add_190_195_groupi_n_6307, csa_tree_add_190_195_groupi_n_6308, csa_tree_add_190_195_groupi_n_6309, csa_tree_add_190_195_groupi_n_6310, csa_tree_add_190_195_groupi_n_6311;
  wire csa_tree_add_190_195_groupi_n_6312, csa_tree_add_190_195_groupi_n_6313, csa_tree_add_190_195_groupi_n_6314, csa_tree_add_190_195_groupi_n_6315, csa_tree_add_190_195_groupi_n_6316, csa_tree_add_190_195_groupi_n_6317, csa_tree_add_190_195_groupi_n_6318, csa_tree_add_190_195_groupi_n_6319;
  wire csa_tree_add_190_195_groupi_n_6320, csa_tree_add_190_195_groupi_n_6321, csa_tree_add_190_195_groupi_n_6322, csa_tree_add_190_195_groupi_n_6323, csa_tree_add_190_195_groupi_n_6324, csa_tree_add_190_195_groupi_n_6325, csa_tree_add_190_195_groupi_n_6326, csa_tree_add_190_195_groupi_n_6327;
  wire csa_tree_add_190_195_groupi_n_6328, csa_tree_add_190_195_groupi_n_6329, csa_tree_add_190_195_groupi_n_6330, csa_tree_add_190_195_groupi_n_6331, csa_tree_add_190_195_groupi_n_6332, csa_tree_add_190_195_groupi_n_6333, csa_tree_add_190_195_groupi_n_6334, csa_tree_add_190_195_groupi_n_6335;
  wire csa_tree_add_190_195_groupi_n_6336, csa_tree_add_190_195_groupi_n_6337, csa_tree_add_190_195_groupi_n_6338, csa_tree_add_190_195_groupi_n_6339, csa_tree_add_190_195_groupi_n_6340, csa_tree_add_190_195_groupi_n_6341, csa_tree_add_190_195_groupi_n_6342, csa_tree_add_190_195_groupi_n_6343;
  wire csa_tree_add_190_195_groupi_n_6344, csa_tree_add_190_195_groupi_n_6345, csa_tree_add_190_195_groupi_n_6346, csa_tree_add_190_195_groupi_n_6347, csa_tree_add_190_195_groupi_n_6348, csa_tree_add_190_195_groupi_n_6349, csa_tree_add_190_195_groupi_n_6350, csa_tree_add_190_195_groupi_n_6351;
  wire csa_tree_add_190_195_groupi_n_6352, csa_tree_add_190_195_groupi_n_6353, csa_tree_add_190_195_groupi_n_6354, csa_tree_add_190_195_groupi_n_6355, csa_tree_add_190_195_groupi_n_6356, csa_tree_add_190_195_groupi_n_6357, csa_tree_add_190_195_groupi_n_6358, csa_tree_add_190_195_groupi_n_6359;
  wire csa_tree_add_190_195_groupi_n_6360, csa_tree_add_190_195_groupi_n_6361, csa_tree_add_190_195_groupi_n_6362, csa_tree_add_190_195_groupi_n_6363, csa_tree_add_190_195_groupi_n_6364, csa_tree_add_190_195_groupi_n_6365, csa_tree_add_190_195_groupi_n_6366, csa_tree_add_190_195_groupi_n_6367;
  wire csa_tree_add_190_195_groupi_n_6368, csa_tree_add_190_195_groupi_n_6369, csa_tree_add_190_195_groupi_n_6370, csa_tree_add_190_195_groupi_n_6371, csa_tree_add_190_195_groupi_n_6372, csa_tree_add_190_195_groupi_n_6373, csa_tree_add_190_195_groupi_n_6374, csa_tree_add_190_195_groupi_n_6375;
  wire csa_tree_add_190_195_groupi_n_6376, csa_tree_add_190_195_groupi_n_6377, csa_tree_add_190_195_groupi_n_6378, csa_tree_add_190_195_groupi_n_6379, csa_tree_add_190_195_groupi_n_6380, csa_tree_add_190_195_groupi_n_6381, csa_tree_add_190_195_groupi_n_6382, csa_tree_add_190_195_groupi_n_6383;
  wire csa_tree_add_190_195_groupi_n_6384, csa_tree_add_190_195_groupi_n_6385, csa_tree_add_190_195_groupi_n_6386, csa_tree_add_190_195_groupi_n_6387, csa_tree_add_190_195_groupi_n_6388, csa_tree_add_190_195_groupi_n_6389, csa_tree_add_190_195_groupi_n_6390, csa_tree_add_190_195_groupi_n_6391;
  wire csa_tree_add_190_195_groupi_n_6392, csa_tree_add_190_195_groupi_n_6393, csa_tree_add_190_195_groupi_n_6394, csa_tree_add_190_195_groupi_n_6395, csa_tree_add_190_195_groupi_n_6396, csa_tree_add_190_195_groupi_n_6397, csa_tree_add_190_195_groupi_n_6398, csa_tree_add_190_195_groupi_n_6399;
  wire csa_tree_add_190_195_groupi_n_6400, csa_tree_add_190_195_groupi_n_6401, csa_tree_add_190_195_groupi_n_6402, csa_tree_add_190_195_groupi_n_6403, csa_tree_add_190_195_groupi_n_6404, csa_tree_add_190_195_groupi_n_6405, csa_tree_add_190_195_groupi_n_6406, csa_tree_add_190_195_groupi_n_6407;
  wire csa_tree_add_190_195_groupi_n_6408, csa_tree_add_190_195_groupi_n_6409, csa_tree_add_190_195_groupi_n_6410, csa_tree_add_190_195_groupi_n_6411, csa_tree_add_190_195_groupi_n_6412, csa_tree_add_190_195_groupi_n_6413, csa_tree_add_190_195_groupi_n_6414, csa_tree_add_190_195_groupi_n_6415;
  wire csa_tree_add_190_195_groupi_n_6416, csa_tree_add_190_195_groupi_n_6417, csa_tree_add_190_195_groupi_n_6418, csa_tree_add_190_195_groupi_n_6419, csa_tree_add_190_195_groupi_n_6420, csa_tree_add_190_195_groupi_n_6421, csa_tree_add_190_195_groupi_n_6422, csa_tree_add_190_195_groupi_n_6423;
  wire csa_tree_add_190_195_groupi_n_6424, csa_tree_add_190_195_groupi_n_6425, csa_tree_add_190_195_groupi_n_6426, csa_tree_add_190_195_groupi_n_6427, csa_tree_add_190_195_groupi_n_6428, csa_tree_add_190_195_groupi_n_6429, csa_tree_add_190_195_groupi_n_6430, csa_tree_add_190_195_groupi_n_6431;
  wire csa_tree_add_190_195_groupi_n_6432, csa_tree_add_190_195_groupi_n_6433, csa_tree_add_190_195_groupi_n_6434, csa_tree_add_190_195_groupi_n_6435, csa_tree_add_190_195_groupi_n_6436, csa_tree_add_190_195_groupi_n_6437, csa_tree_add_190_195_groupi_n_6438, csa_tree_add_190_195_groupi_n_6439;
  wire csa_tree_add_190_195_groupi_n_6440, csa_tree_add_190_195_groupi_n_6441, csa_tree_add_190_195_groupi_n_6442, csa_tree_add_190_195_groupi_n_6443, csa_tree_add_190_195_groupi_n_6444, csa_tree_add_190_195_groupi_n_6445, csa_tree_add_190_195_groupi_n_6446, csa_tree_add_190_195_groupi_n_6447;
  wire csa_tree_add_190_195_groupi_n_6448, csa_tree_add_190_195_groupi_n_6449, csa_tree_add_190_195_groupi_n_6450, csa_tree_add_190_195_groupi_n_6451, csa_tree_add_190_195_groupi_n_6452, csa_tree_add_190_195_groupi_n_6453, csa_tree_add_190_195_groupi_n_6454, csa_tree_add_190_195_groupi_n_6455;
  wire csa_tree_add_190_195_groupi_n_6456, csa_tree_add_190_195_groupi_n_6457, csa_tree_add_190_195_groupi_n_6458, csa_tree_add_190_195_groupi_n_6459, csa_tree_add_190_195_groupi_n_6460, csa_tree_add_190_195_groupi_n_6461, csa_tree_add_190_195_groupi_n_6462, csa_tree_add_190_195_groupi_n_6463;
  wire csa_tree_add_190_195_groupi_n_6464, csa_tree_add_190_195_groupi_n_6465, csa_tree_add_190_195_groupi_n_6466, csa_tree_add_190_195_groupi_n_6467, csa_tree_add_190_195_groupi_n_6468, csa_tree_add_190_195_groupi_n_6469, csa_tree_add_190_195_groupi_n_6470, csa_tree_add_190_195_groupi_n_6471;
  wire csa_tree_add_190_195_groupi_n_6472, csa_tree_add_190_195_groupi_n_6473, csa_tree_add_190_195_groupi_n_6474, csa_tree_add_190_195_groupi_n_6475, csa_tree_add_190_195_groupi_n_6476, csa_tree_add_190_195_groupi_n_6477, csa_tree_add_190_195_groupi_n_6478, csa_tree_add_190_195_groupi_n_6479;
  wire csa_tree_add_190_195_groupi_n_6480, csa_tree_add_190_195_groupi_n_6481, csa_tree_add_190_195_groupi_n_6482, csa_tree_add_190_195_groupi_n_6483, csa_tree_add_190_195_groupi_n_6484, csa_tree_add_190_195_groupi_n_6485, csa_tree_add_190_195_groupi_n_6486, csa_tree_add_190_195_groupi_n_6487;
  wire csa_tree_add_190_195_groupi_n_6488, csa_tree_add_190_195_groupi_n_6489, csa_tree_add_190_195_groupi_n_6490, csa_tree_add_190_195_groupi_n_6491, csa_tree_add_190_195_groupi_n_6492, csa_tree_add_190_195_groupi_n_6493, csa_tree_add_190_195_groupi_n_6494, csa_tree_add_190_195_groupi_n_6495;
  wire csa_tree_add_190_195_groupi_n_6496, csa_tree_add_190_195_groupi_n_6497, csa_tree_add_190_195_groupi_n_6498, csa_tree_add_190_195_groupi_n_6499, csa_tree_add_190_195_groupi_n_6500, csa_tree_add_190_195_groupi_n_6501, csa_tree_add_190_195_groupi_n_6502, csa_tree_add_190_195_groupi_n_6503;
  wire csa_tree_add_190_195_groupi_n_6504, csa_tree_add_190_195_groupi_n_6505, csa_tree_add_190_195_groupi_n_6506, csa_tree_add_190_195_groupi_n_6507, csa_tree_add_190_195_groupi_n_6508, csa_tree_add_190_195_groupi_n_6509, csa_tree_add_190_195_groupi_n_6510, csa_tree_add_190_195_groupi_n_6511;
  wire csa_tree_add_190_195_groupi_n_6512, csa_tree_add_190_195_groupi_n_6513, csa_tree_add_190_195_groupi_n_6514, csa_tree_add_190_195_groupi_n_6515, csa_tree_add_190_195_groupi_n_6516, csa_tree_add_190_195_groupi_n_6517, csa_tree_add_190_195_groupi_n_6518, csa_tree_add_190_195_groupi_n_6519;
  wire csa_tree_add_190_195_groupi_n_6520, csa_tree_add_190_195_groupi_n_6521, csa_tree_add_190_195_groupi_n_6522, csa_tree_add_190_195_groupi_n_6523, csa_tree_add_190_195_groupi_n_6524, csa_tree_add_190_195_groupi_n_6525, csa_tree_add_190_195_groupi_n_6526, csa_tree_add_190_195_groupi_n_6527;
  wire csa_tree_add_190_195_groupi_n_6528, csa_tree_add_190_195_groupi_n_6529, csa_tree_add_190_195_groupi_n_6530, csa_tree_add_190_195_groupi_n_6531, csa_tree_add_190_195_groupi_n_6532, csa_tree_add_190_195_groupi_n_6533, csa_tree_add_190_195_groupi_n_6534, csa_tree_add_190_195_groupi_n_6535;
  wire csa_tree_add_190_195_groupi_n_6536, csa_tree_add_190_195_groupi_n_6537, csa_tree_add_190_195_groupi_n_6538, csa_tree_add_190_195_groupi_n_6539, csa_tree_add_190_195_groupi_n_6540, csa_tree_add_190_195_groupi_n_6541, csa_tree_add_190_195_groupi_n_6542, csa_tree_add_190_195_groupi_n_6543;
  wire csa_tree_add_190_195_groupi_n_6544, csa_tree_add_190_195_groupi_n_6545, csa_tree_add_190_195_groupi_n_6546, csa_tree_add_190_195_groupi_n_6547, csa_tree_add_190_195_groupi_n_6548, csa_tree_add_190_195_groupi_n_6549, csa_tree_add_190_195_groupi_n_6550, csa_tree_add_190_195_groupi_n_6551;
  wire csa_tree_add_190_195_groupi_n_6552, csa_tree_add_190_195_groupi_n_6553, csa_tree_add_190_195_groupi_n_6554, csa_tree_add_190_195_groupi_n_6555, csa_tree_add_190_195_groupi_n_6556, csa_tree_add_190_195_groupi_n_6557, csa_tree_add_190_195_groupi_n_6558, csa_tree_add_190_195_groupi_n_6559;
  wire csa_tree_add_190_195_groupi_n_6560, csa_tree_add_190_195_groupi_n_6561, csa_tree_add_190_195_groupi_n_6562, csa_tree_add_190_195_groupi_n_6563, csa_tree_add_190_195_groupi_n_6564, csa_tree_add_190_195_groupi_n_6565, csa_tree_add_190_195_groupi_n_6566, csa_tree_add_190_195_groupi_n_6567;
  wire csa_tree_add_190_195_groupi_n_6568, csa_tree_add_190_195_groupi_n_6569, csa_tree_add_190_195_groupi_n_6570, csa_tree_add_190_195_groupi_n_6571, csa_tree_add_190_195_groupi_n_6572, csa_tree_add_190_195_groupi_n_6573, csa_tree_add_190_195_groupi_n_6574, csa_tree_add_190_195_groupi_n_6575;
  wire csa_tree_add_190_195_groupi_n_6576, csa_tree_add_190_195_groupi_n_6577, csa_tree_add_190_195_groupi_n_6578, csa_tree_add_190_195_groupi_n_6579, csa_tree_add_190_195_groupi_n_6580, csa_tree_add_190_195_groupi_n_6581, csa_tree_add_190_195_groupi_n_6582, csa_tree_add_190_195_groupi_n_6583;
  wire csa_tree_add_190_195_groupi_n_6584, csa_tree_add_190_195_groupi_n_6585, csa_tree_add_190_195_groupi_n_6586, csa_tree_add_190_195_groupi_n_6587, csa_tree_add_190_195_groupi_n_6588, csa_tree_add_190_195_groupi_n_6589, csa_tree_add_190_195_groupi_n_6590, csa_tree_add_190_195_groupi_n_6591;
  wire csa_tree_add_190_195_groupi_n_6592, csa_tree_add_190_195_groupi_n_6593, csa_tree_add_190_195_groupi_n_6594, csa_tree_add_190_195_groupi_n_6595, csa_tree_add_190_195_groupi_n_6596, csa_tree_add_190_195_groupi_n_6597, csa_tree_add_190_195_groupi_n_6598, csa_tree_add_190_195_groupi_n_6599;
  wire csa_tree_add_190_195_groupi_n_6600, csa_tree_add_190_195_groupi_n_6601, csa_tree_add_190_195_groupi_n_6602, csa_tree_add_190_195_groupi_n_6603, csa_tree_add_190_195_groupi_n_6604, csa_tree_add_190_195_groupi_n_6605, csa_tree_add_190_195_groupi_n_6606, csa_tree_add_190_195_groupi_n_6607;
  wire csa_tree_add_190_195_groupi_n_6608, csa_tree_add_190_195_groupi_n_6609, csa_tree_add_190_195_groupi_n_6610, csa_tree_add_190_195_groupi_n_6611, csa_tree_add_190_195_groupi_n_6612, csa_tree_add_190_195_groupi_n_6613, csa_tree_add_190_195_groupi_n_6614, csa_tree_add_190_195_groupi_n_6615;
  wire csa_tree_add_190_195_groupi_n_6616, csa_tree_add_190_195_groupi_n_6617, csa_tree_add_190_195_groupi_n_6618, csa_tree_add_190_195_groupi_n_6619, csa_tree_add_190_195_groupi_n_6620, csa_tree_add_190_195_groupi_n_6621, csa_tree_add_190_195_groupi_n_6622, csa_tree_add_190_195_groupi_n_6623;
  wire csa_tree_add_190_195_groupi_n_6624, csa_tree_add_190_195_groupi_n_6625, csa_tree_add_190_195_groupi_n_6626, csa_tree_add_190_195_groupi_n_6627, csa_tree_add_190_195_groupi_n_6628, csa_tree_add_190_195_groupi_n_6629, csa_tree_add_190_195_groupi_n_6630, csa_tree_add_190_195_groupi_n_6631;
  wire csa_tree_add_190_195_groupi_n_6632, csa_tree_add_190_195_groupi_n_6633, csa_tree_add_190_195_groupi_n_6634, csa_tree_add_190_195_groupi_n_6635, csa_tree_add_190_195_groupi_n_6636, csa_tree_add_190_195_groupi_n_6637, csa_tree_add_190_195_groupi_n_6638, csa_tree_add_190_195_groupi_n_6639;
  wire csa_tree_add_190_195_groupi_n_6640, csa_tree_add_190_195_groupi_n_6641, csa_tree_add_190_195_groupi_n_6642, csa_tree_add_190_195_groupi_n_6643, csa_tree_add_190_195_groupi_n_6644, csa_tree_add_190_195_groupi_n_6645, csa_tree_add_190_195_groupi_n_6646, csa_tree_add_190_195_groupi_n_6647;
  wire csa_tree_add_190_195_groupi_n_6648, csa_tree_add_190_195_groupi_n_6649, csa_tree_add_190_195_groupi_n_6650, csa_tree_add_190_195_groupi_n_6651, csa_tree_add_190_195_groupi_n_6652, csa_tree_add_190_195_groupi_n_6653, csa_tree_add_190_195_groupi_n_6654, csa_tree_add_190_195_groupi_n_6655;
  wire csa_tree_add_190_195_groupi_n_6656, csa_tree_add_190_195_groupi_n_6657, csa_tree_add_190_195_groupi_n_6658, csa_tree_add_190_195_groupi_n_6659, csa_tree_add_190_195_groupi_n_6660, csa_tree_add_190_195_groupi_n_6661, csa_tree_add_190_195_groupi_n_6662, csa_tree_add_190_195_groupi_n_6663;
  wire csa_tree_add_190_195_groupi_n_6664, csa_tree_add_190_195_groupi_n_6665, csa_tree_add_190_195_groupi_n_6666, csa_tree_add_190_195_groupi_n_6667, csa_tree_add_190_195_groupi_n_6668, csa_tree_add_190_195_groupi_n_6669, csa_tree_add_190_195_groupi_n_6670, csa_tree_add_190_195_groupi_n_6671;
  wire csa_tree_add_190_195_groupi_n_6672, csa_tree_add_190_195_groupi_n_6673, csa_tree_add_190_195_groupi_n_6674, csa_tree_add_190_195_groupi_n_6675, csa_tree_add_190_195_groupi_n_6676, csa_tree_add_190_195_groupi_n_6677, csa_tree_add_190_195_groupi_n_6678, csa_tree_add_190_195_groupi_n_6679;
  wire csa_tree_add_190_195_groupi_n_6680, csa_tree_add_190_195_groupi_n_6681, csa_tree_add_190_195_groupi_n_6682, csa_tree_add_190_195_groupi_n_6683, csa_tree_add_190_195_groupi_n_6684, csa_tree_add_190_195_groupi_n_6685, csa_tree_add_190_195_groupi_n_6686, csa_tree_add_190_195_groupi_n_6687;
  wire csa_tree_add_190_195_groupi_n_6688, csa_tree_add_190_195_groupi_n_6689, csa_tree_add_190_195_groupi_n_6690, csa_tree_add_190_195_groupi_n_6691, csa_tree_add_190_195_groupi_n_6692, csa_tree_add_190_195_groupi_n_6693, csa_tree_add_190_195_groupi_n_6694, csa_tree_add_190_195_groupi_n_6695;
  wire csa_tree_add_190_195_groupi_n_6696, csa_tree_add_190_195_groupi_n_6697, csa_tree_add_190_195_groupi_n_6698, csa_tree_add_190_195_groupi_n_6699, csa_tree_add_190_195_groupi_n_6700, csa_tree_add_190_195_groupi_n_6701, csa_tree_add_190_195_groupi_n_6702, csa_tree_add_190_195_groupi_n_6703;
  wire csa_tree_add_190_195_groupi_n_6704, csa_tree_add_190_195_groupi_n_6705, csa_tree_add_190_195_groupi_n_6706, csa_tree_add_190_195_groupi_n_6707, csa_tree_add_190_195_groupi_n_6708, csa_tree_add_190_195_groupi_n_6709, csa_tree_add_190_195_groupi_n_6710, csa_tree_add_190_195_groupi_n_6711;
  wire csa_tree_add_190_195_groupi_n_6712, csa_tree_add_190_195_groupi_n_6713, csa_tree_add_190_195_groupi_n_6714, csa_tree_add_190_195_groupi_n_6715, csa_tree_add_190_195_groupi_n_6716, csa_tree_add_190_195_groupi_n_6717, csa_tree_add_190_195_groupi_n_6718, csa_tree_add_190_195_groupi_n_6719;
  wire csa_tree_add_190_195_groupi_n_6720, csa_tree_add_190_195_groupi_n_6721, csa_tree_add_190_195_groupi_n_6722, csa_tree_add_190_195_groupi_n_6723, csa_tree_add_190_195_groupi_n_6724, csa_tree_add_190_195_groupi_n_6725, csa_tree_add_190_195_groupi_n_6726, csa_tree_add_190_195_groupi_n_6727;
  wire csa_tree_add_190_195_groupi_n_6728, csa_tree_add_190_195_groupi_n_6729, csa_tree_add_190_195_groupi_n_6730, csa_tree_add_190_195_groupi_n_6731, csa_tree_add_190_195_groupi_n_6732, csa_tree_add_190_195_groupi_n_6733, csa_tree_add_190_195_groupi_n_6734, csa_tree_add_190_195_groupi_n_6735;
  wire csa_tree_add_190_195_groupi_n_6736, csa_tree_add_190_195_groupi_n_6737, csa_tree_add_190_195_groupi_n_6738, csa_tree_add_190_195_groupi_n_6739, csa_tree_add_190_195_groupi_n_6740, csa_tree_add_190_195_groupi_n_6741, csa_tree_add_190_195_groupi_n_6742, csa_tree_add_190_195_groupi_n_6743;
  wire csa_tree_add_190_195_groupi_n_6744, csa_tree_add_190_195_groupi_n_6745, csa_tree_add_190_195_groupi_n_6746, csa_tree_add_190_195_groupi_n_6747, csa_tree_add_190_195_groupi_n_6748, csa_tree_add_190_195_groupi_n_6749, csa_tree_add_190_195_groupi_n_6750, csa_tree_add_190_195_groupi_n_6751;
  wire csa_tree_add_190_195_groupi_n_6752, csa_tree_add_190_195_groupi_n_6753, csa_tree_add_190_195_groupi_n_6754, csa_tree_add_190_195_groupi_n_6755, csa_tree_add_190_195_groupi_n_6756, csa_tree_add_190_195_groupi_n_6757, csa_tree_add_190_195_groupi_n_6758, csa_tree_add_190_195_groupi_n_6759;
  wire csa_tree_add_190_195_groupi_n_6760, csa_tree_add_190_195_groupi_n_6761, csa_tree_add_190_195_groupi_n_6762, csa_tree_add_190_195_groupi_n_6763, csa_tree_add_190_195_groupi_n_6764, csa_tree_add_190_195_groupi_n_6765, csa_tree_add_190_195_groupi_n_6766, csa_tree_add_190_195_groupi_n_6767;
  wire csa_tree_add_190_195_groupi_n_6768, csa_tree_add_190_195_groupi_n_6769, csa_tree_add_190_195_groupi_n_6770, csa_tree_add_190_195_groupi_n_6771, csa_tree_add_190_195_groupi_n_6772, csa_tree_add_190_195_groupi_n_6773, csa_tree_add_190_195_groupi_n_6774, csa_tree_add_190_195_groupi_n_6775;
  wire csa_tree_add_190_195_groupi_n_6776, csa_tree_add_190_195_groupi_n_6777, csa_tree_add_190_195_groupi_n_6778, csa_tree_add_190_195_groupi_n_6779, csa_tree_add_190_195_groupi_n_6780, csa_tree_add_190_195_groupi_n_6781, csa_tree_add_190_195_groupi_n_6782, csa_tree_add_190_195_groupi_n_6783;
  wire csa_tree_add_190_195_groupi_n_6784, csa_tree_add_190_195_groupi_n_6785, csa_tree_add_190_195_groupi_n_6786, csa_tree_add_190_195_groupi_n_6787, csa_tree_add_190_195_groupi_n_6788, csa_tree_add_190_195_groupi_n_6789, csa_tree_add_190_195_groupi_n_6790, csa_tree_add_190_195_groupi_n_6791;
  wire csa_tree_add_190_195_groupi_n_6792, csa_tree_add_190_195_groupi_n_6793, csa_tree_add_190_195_groupi_n_6794, csa_tree_add_190_195_groupi_n_6795, csa_tree_add_190_195_groupi_n_6796, csa_tree_add_190_195_groupi_n_6797, csa_tree_add_190_195_groupi_n_6798, csa_tree_add_190_195_groupi_n_6799;
  wire csa_tree_add_190_195_groupi_n_6800, csa_tree_add_190_195_groupi_n_6801, csa_tree_add_190_195_groupi_n_6802, csa_tree_add_190_195_groupi_n_6803, csa_tree_add_190_195_groupi_n_6804, csa_tree_add_190_195_groupi_n_6805, csa_tree_add_190_195_groupi_n_6806, csa_tree_add_190_195_groupi_n_6807;
  wire csa_tree_add_190_195_groupi_n_6808, csa_tree_add_190_195_groupi_n_6809, csa_tree_add_190_195_groupi_n_6810, csa_tree_add_190_195_groupi_n_6811, csa_tree_add_190_195_groupi_n_6812, csa_tree_add_190_195_groupi_n_6813, csa_tree_add_190_195_groupi_n_6814, csa_tree_add_190_195_groupi_n_6815;
  wire csa_tree_add_190_195_groupi_n_6816, csa_tree_add_190_195_groupi_n_6817, csa_tree_add_190_195_groupi_n_6818, csa_tree_add_190_195_groupi_n_6819, csa_tree_add_190_195_groupi_n_6820, csa_tree_add_190_195_groupi_n_6821, csa_tree_add_190_195_groupi_n_6822, csa_tree_add_190_195_groupi_n_6823;
  wire csa_tree_add_190_195_groupi_n_6824, csa_tree_add_190_195_groupi_n_6825, csa_tree_add_190_195_groupi_n_6826, csa_tree_add_190_195_groupi_n_6827, csa_tree_add_190_195_groupi_n_6828, csa_tree_add_190_195_groupi_n_6829, csa_tree_add_190_195_groupi_n_6830, csa_tree_add_190_195_groupi_n_6831;
  wire csa_tree_add_190_195_groupi_n_6832, csa_tree_add_190_195_groupi_n_6833, csa_tree_add_190_195_groupi_n_6834, csa_tree_add_190_195_groupi_n_6835, csa_tree_add_190_195_groupi_n_6836, csa_tree_add_190_195_groupi_n_6837, csa_tree_add_190_195_groupi_n_6838, csa_tree_add_190_195_groupi_n_6839;
  wire csa_tree_add_190_195_groupi_n_6840, csa_tree_add_190_195_groupi_n_6841, csa_tree_add_190_195_groupi_n_6842, csa_tree_add_190_195_groupi_n_6843, csa_tree_add_190_195_groupi_n_6844, csa_tree_add_190_195_groupi_n_6845, csa_tree_add_190_195_groupi_n_6846, csa_tree_add_190_195_groupi_n_6847;
  wire csa_tree_add_190_195_groupi_n_6848, csa_tree_add_190_195_groupi_n_6849, csa_tree_add_190_195_groupi_n_6850, csa_tree_add_190_195_groupi_n_6851, csa_tree_add_190_195_groupi_n_6852, csa_tree_add_190_195_groupi_n_6853, csa_tree_add_190_195_groupi_n_6854, csa_tree_add_190_195_groupi_n_6855;
  wire csa_tree_add_190_195_groupi_n_6856, csa_tree_add_190_195_groupi_n_6857, csa_tree_add_190_195_groupi_n_6858, csa_tree_add_190_195_groupi_n_6859, csa_tree_add_190_195_groupi_n_6860, csa_tree_add_190_195_groupi_n_6861, csa_tree_add_190_195_groupi_n_6862, csa_tree_add_190_195_groupi_n_6863;
  wire csa_tree_add_190_195_groupi_n_6864, csa_tree_add_190_195_groupi_n_6865, csa_tree_add_190_195_groupi_n_6866, csa_tree_add_190_195_groupi_n_6867, csa_tree_add_190_195_groupi_n_6868, csa_tree_add_190_195_groupi_n_6869, csa_tree_add_190_195_groupi_n_6870, csa_tree_add_190_195_groupi_n_6871;
  wire csa_tree_add_190_195_groupi_n_6872, csa_tree_add_190_195_groupi_n_6873, csa_tree_add_190_195_groupi_n_6874, csa_tree_add_190_195_groupi_n_6875, csa_tree_add_190_195_groupi_n_6876, csa_tree_add_190_195_groupi_n_6877, csa_tree_add_190_195_groupi_n_6878, csa_tree_add_190_195_groupi_n_6879;
  wire csa_tree_add_190_195_groupi_n_6880, csa_tree_add_190_195_groupi_n_6881, csa_tree_add_190_195_groupi_n_6882, csa_tree_add_190_195_groupi_n_6883, csa_tree_add_190_195_groupi_n_6884, csa_tree_add_190_195_groupi_n_6885, csa_tree_add_190_195_groupi_n_6886, csa_tree_add_190_195_groupi_n_6887;
  wire csa_tree_add_190_195_groupi_n_6888, csa_tree_add_190_195_groupi_n_6889, csa_tree_add_190_195_groupi_n_6890, csa_tree_add_190_195_groupi_n_6891, csa_tree_add_190_195_groupi_n_6892, csa_tree_add_190_195_groupi_n_6893, csa_tree_add_190_195_groupi_n_6894, csa_tree_add_190_195_groupi_n_6895;
  wire csa_tree_add_190_195_groupi_n_6896, csa_tree_add_190_195_groupi_n_6897, csa_tree_add_190_195_groupi_n_6898, csa_tree_add_190_195_groupi_n_6899, csa_tree_add_190_195_groupi_n_6900, csa_tree_add_190_195_groupi_n_6901, csa_tree_add_190_195_groupi_n_6902, csa_tree_add_190_195_groupi_n_6903;
  wire csa_tree_add_190_195_groupi_n_6904, csa_tree_add_190_195_groupi_n_6905, csa_tree_add_190_195_groupi_n_6906, csa_tree_add_190_195_groupi_n_6907, csa_tree_add_190_195_groupi_n_6908, csa_tree_add_190_195_groupi_n_6909, csa_tree_add_190_195_groupi_n_6910, csa_tree_add_190_195_groupi_n_6911;
  wire csa_tree_add_190_195_groupi_n_6912, csa_tree_add_190_195_groupi_n_6913, csa_tree_add_190_195_groupi_n_6914, csa_tree_add_190_195_groupi_n_6915, csa_tree_add_190_195_groupi_n_6916, csa_tree_add_190_195_groupi_n_6917, csa_tree_add_190_195_groupi_n_6918, csa_tree_add_190_195_groupi_n_6919;
  wire csa_tree_add_190_195_groupi_n_6920, csa_tree_add_190_195_groupi_n_6921, csa_tree_add_190_195_groupi_n_6922, csa_tree_add_190_195_groupi_n_6923, csa_tree_add_190_195_groupi_n_6924, csa_tree_add_190_195_groupi_n_6925, csa_tree_add_190_195_groupi_n_6926, csa_tree_add_190_195_groupi_n_6927;
  wire csa_tree_add_190_195_groupi_n_6928, csa_tree_add_190_195_groupi_n_6929, csa_tree_add_190_195_groupi_n_6930, csa_tree_add_190_195_groupi_n_6931, csa_tree_add_190_195_groupi_n_6932, csa_tree_add_190_195_groupi_n_6933, csa_tree_add_190_195_groupi_n_6934, csa_tree_add_190_195_groupi_n_6935;
  wire csa_tree_add_190_195_groupi_n_6936, csa_tree_add_190_195_groupi_n_6937, csa_tree_add_190_195_groupi_n_6938, csa_tree_add_190_195_groupi_n_6939, csa_tree_add_190_195_groupi_n_6940, csa_tree_add_190_195_groupi_n_6941, csa_tree_add_190_195_groupi_n_6942, csa_tree_add_190_195_groupi_n_6943;
  wire csa_tree_add_190_195_groupi_n_6944, csa_tree_add_190_195_groupi_n_6945, csa_tree_add_190_195_groupi_n_6946, csa_tree_add_190_195_groupi_n_6947, csa_tree_add_190_195_groupi_n_6948, csa_tree_add_190_195_groupi_n_6949, csa_tree_add_190_195_groupi_n_6950, csa_tree_add_190_195_groupi_n_6951;
  wire csa_tree_add_190_195_groupi_n_6952, csa_tree_add_190_195_groupi_n_6953, csa_tree_add_190_195_groupi_n_6954, csa_tree_add_190_195_groupi_n_6955, csa_tree_add_190_195_groupi_n_6956, csa_tree_add_190_195_groupi_n_6957, csa_tree_add_190_195_groupi_n_6958, csa_tree_add_190_195_groupi_n_6959;
  wire csa_tree_add_190_195_groupi_n_6960, csa_tree_add_190_195_groupi_n_6961, csa_tree_add_190_195_groupi_n_6962, csa_tree_add_190_195_groupi_n_6963, csa_tree_add_190_195_groupi_n_6964, csa_tree_add_190_195_groupi_n_6965, csa_tree_add_190_195_groupi_n_6966, csa_tree_add_190_195_groupi_n_6967;
  wire csa_tree_add_190_195_groupi_n_6968, csa_tree_add_190_195_groupi_n_6969, csa_tree_add_190_195_groupi_n_6970, csa_tree_add_190_195_groupi_n_6971, csa_tree_add_190_195_groupi_n_6972, csa_tree_add_190_195_groupi_n_6973, csa_tree_add_190_195_groupi_n_6974, csa_tree_add_190_195_groupi_n_6975;
  wire csa_tree_add_190_195_groupi_n_6976, csa_tree_add_190_195_groupi_n_6977, csa_tree_add_190_195_groupi_n_6978, csa_tree_add_190_195_groupi_n_6979, csa_tree_add_190_195_groupi_n_6980, csa_tree_add_190_195_groupi_n_6981, csa_tree_add_190_195_groupi_n_6982, csa_tree_add_190_195_groupi_n_6983;
  wire csa_tree_add_190_195_groupi_n_6984, csa_tree_add_190_195_groupi_n_6985, csa_tree_add_190_195_groupi_n_6986, csa_tree_add_190_195_groupi_n_6987, csa_tree_add_190_195_groupi_n_6988, csa_tree_add_190_195_groupi_n_6989, csa_tree_add_190_195_groupi_n_6990, csa_tree_add_190_195_groupi_n_6991;
  wire csa_tree_add_190_195_groupi_n_6992, csa_tree_add_190_195_groupi_n_6993, csa_tree_add_190_195_groupi_n_6994, csa_tree_add_190_195_groupi_n_6995, csa_tree_add_190_195_groupi_n_6996, csa_tree_add_190_195_groupi_n_6997, csa_tree_add_190_195_groupi_n_6998, csa_tree_add_190_195_groupi_n_6999;
  wire csa_tree_add_190_195_groupi_n_7000, csa_tree_add_190_195_groupi_n_7001, csa_tree_add_190_195_groupi_n_7002, csa_tree_add_190_195_groupi_n_7003, csa_tree_add_190_195_groupi_n_7004, csa_tree_add_190_195_groupi_n_7005, csa_tree_add_190_195_groupi_n_7006, csa_tree_add_190_195_groupi_n_7007;
  wire csa_tree_add_190_195_groupi_n_7008, csa_tree_add_190_195_groupi_n_7009, csa_tree_add_190_195_groupi_n_7010, csa_tree_add_190_195_groupi_n_7011, csa_tree_add_190_195_groupi_n_7012, csa_tree_add_190_195_groupi_n_7013, csa_tree_add_190_195_groupi_n_7014, csa_tree_add_190_195_groupi_n_7015;
  wire csa_tree_add_190_195_groupi_n_7016, csa_tree_add_190_195_groupi_n_7017, csa_tree_add_190_195_groupi_n_7018, csa_tree_add_190_195_groupi_n_7019, csa_tree_add_190_195_groupi_n_7020, csa_tree_add_190_195_groupi_n_7021, csa_tree_add_190_195_groupi_n_7022, csa_tree_add_190_195_groupi_n_7023;
  wire csa_tree_add_190_195_groupi_n_7024, csa_tree_add_190_195_groupi_n_7025, csa_tree_add_190_195_groupi_n_7026, csa_tree_add_190_195_groupi_n_7027, csa_tree_add_190_195_groupi_n_7028, csa_tree_add_190_195_groupi_n_7029, csa_tree_add_190_195_groupi_n_7030, csa_tree_add_190_195_groupi_n_7031;
  wire csa_tree_add_190_195_groupi_n_7032, csa_tree_add_190_195_groupi_n_7033, csa_tree_add_190_195_groupi_n_7034, csa_tree_add_190_195_groupi_n_7035, csa_tree_add_190_195_groupi_n_7036, csa_tree_add_190_195_groupi_n_7037, csa_tree_add_190_195_groupi_n_7038, csa_tree_add_190_195_groupi_n_7039;
  wire csa_tree_add_190_195_groupi_n_7040, csa_tree_add_190_195_groupi_n_7041, csa_tree_add_190_195_groupi_n_7042, csa_tree_add_190_195_groupi_n_7043, csa_tree_add_190_195_groupi_n_7044, csa_tree_add_190_195_groupi_n_7045, csa_tree_add_190_195_groupi_n_7046, csa_tree_add_190_195_groupi_n_7047;
  wire csa_tree_add_190_195_groupi_n_7048, csa_tree_add_190_195_groupi_n_7049, csa_tree_add_190_195_groupi_n_7050, csa_tree_add_190_195_groupi_n_7051, csa_tree_add_190_195_groupi_n_7052, csa_tree_add_190_195_groupi_n_7053, csa_tree_add_190_195_groupi_n_7054, csa_tree_add_190_195_groupi_n_7055;
  wire csa_tree_add_190_195_groupi_n_7056, csa_tree_add_190_195_groupi_n_7057, csa_tree_add_190_195_groupi_n_7058, csa_tree_add_190_195_groupi_n_7059, csa_tree_add_190_195_groupi_n_7060, csa_tree_add_190_195_groupi_n_7061, csa_tree_add_190_195_groupi_n_7062, csa_tree_add_190_195_groupi_n_7063;
  wire csa_tree_add_190_195_groupi_n_7064, csa_tree_add_190_195_groupi_n_7065, csa_tree_add_190_195_groupi_n_7066, csa_tree_add_190_195_groupi_n_7067, csa_tree_add_190_195_groupi_n_7068, csa_tree_add_190_195_groupi_n_7069, csa_tree_add_190_195_groupi_n_7070, csa_tree_add_190_195_groupi_n_7071;
  wire csa_tree_add_190_195_groupi_n_7072, csa_tree_add_190_195_groupi_n_7073, csa_tree_add_190_195_groupi_n_7074, csa_tree_add_190_195_groupi_n_7075, csa_tree_add_190_195_groupi_n_7076, csa_tree_add_190_195_groupi_n_7077, csa_tree_add_190_195_groupi_n_7078, csa_tree_add_190_195_groupi_n_7079;
  wire csa_tree_add_190_195_groupi_n_7080, csa_tree_add_190_195_groupi_n_7081, csa_tree_add_190_195_groupi_n_7082, csa_tree_add_190_195_groupi_n_7083, csa_tree_add_190_195_groupi_n_7084, csa_tree_add_190_195_groupi_n_7085, csa_tree_add_190_195_groupi_n_7086, csa_tree_add_190_195_groupi_n_7087;
  wire csa_tree_add_190_195_groupi_n_7088, csa_tree_add_190_195_groupi_n_7089, csa_tree_add_190_195_groupi_n_7090, csa_tree_add_190_195_groupi_n_7091, csa_tree_add_190_195_groupi_n_7092, csa_tree_add_190_195_groupi_n_7093, csa_tree_add_190_195_groupi_n_7094, csa_tree_add_190_195_groupi_n_7095;
  wire csa_tree_add_190_195_groupi_n_7096, csa_tree_add_190_195_groupi_n_7097, csa_tree_add_190_195_groupi_n_7098, csa_tree_add_190_195_groupi_n_7099, csa_tree_add_190_195_groupi_n_7100, csa_tree_add_190_195_groupi_n_7101, csa_tree_add_190_195_groupi_n_7102, csa_tree_add_190_195_groupi_n_7103;
  wire csa_tree_add_190_195_groupi_n_7104, csa_tree_add_190_195_groupi_n_7105, csa_tree_add_190_195_groupi_n_7106, csa_tree_add_190_195_groupi_n_7107, csa_tree_add_190_195_groupi_n_7108, csa_tree_add_190_195_groupi_n_7109, csa_tree_add_190_195_groupi_n_7110, csa_tree_add_190_195_groupi_n_7111;
  wire csa_tree_add_190_195_groupi_n_7112, csa_tree_add_190_195_groupi_n_7113, csa_tree_add_190_195_groupi_n_7114, csa_tree_add_190_195_groupi_n_7115, csa_tree_add_190_195_groupi_n_7116, csa_tree_add_190_195_groupi_n_7117, csa_tree_add_190_195_groupi_n_7118, csa_tree_add_190_195_groupi_n_7119;
  wire csa_tree_add_190_195_groupi_n_7120, csa_tree_add_190_195_groupi_n_7121, csa_tree_add_190_195_groupi_n_7122, csa_tree_add_190_195_groupi_n_7123, csa_tree_add_190_195_groupi_n_7124, csa_tree_add_190_195_groupi_n_7125, csa_tree_add_190_195_groupi_n_7126, csa_tree_add_190_195_groupi_n_7127;
  wire csa_tree_add_190_195_groupi_n_7128, csa_tree_add_190_195_groupi_n_7129, csa_tree_add_190_195_groupi_n_7130, csa_tree_add_190_195_groupi_n_7131, csa_tree_add_190_195_groupi_n_7132, csa_tree_add_190_195_groupi_n_7133, csa_tree_add_190_195_groupi_n_7134, csa_tree_add_190_195_groupi_n_7135;
  wire csa_tree_add_190_195_groupi_n_7136, csa_tree_add_190_195_groupi_n_7137, csa_tree_add_190_195_groupi_n_7138, csa_tree_add_190_195_groupi_n_7139, csa_tree_add_190_195_groupi_n_7140, csa_tree_add_190_195_groupi_n_7141, csa_tree_add_190_195_groupi_n_7142, csa_tree_add_190_195_groupi_n_7143;
  wire csa_tree_add_190_195_groupi_n_7144, csa_tree_add_190_195_groupi_n_7145, csa_tree_add_190_195_groupi_n_7146, csa_tree_add_190_195_groupi_n_7147, csa_tree_add_190_195_groupi_n_7148, csa_tree_add_190_195_groupi_n_7149, csa_tree_add_190_195_groupi_n_7150, csa_tree_add_190_195_groupi_n_7151;
  wire csa_tree_add_190_195_groupi_n_7152, csa_tree_add_190_195_groupi_n_7153, csa_tree_add_190_195_groupi_n_7154, csa_tree_add_190_195_groupi_n_7155, csa_tree_add_190_195_groupi_n_7156, csa_tree_add_190_195_groupi_n_7157, csa_tree_add_190_195_groupi_n_7158, csa_tree_add_190_195_groupi_n_7159;
  wire csa_tree_add_190_195_groupi_n_7160, csa_tree_add_190_195_groupi_n_7161, csa_tree_add_190_195_groupi_n_7162, csa_tree_add_190_195_groupi_n_7163, csa_tree_add_190_195_groupi_n_7164, csa_tree_add_190_195_groupi_n_7165, csa_tree_add_190_195_groupi_n_7166, csa_tree_add_190_195_groupi_n_7167;
  wire csa_tree_add_190_195_groupi_n_7168, csa_tree_add_190_195_groupi_n_7169, csa_tree_add_190_195_groupi_n_7170, csa_tree_add_190_195_groupi_n_7171, csa_tree_add_190_195_groupi_n_7172, csa_tree_add_190_195_groupi_n_7173, csa_tree_add_190_195_groupi_n_7174, csa_tree_add_190_195_groupi_n_7175;
  wire csa_tree_add_190_195_groupi_n_7176, csa_tree_add_190_195_groupi_n_7177, csa_tree_add_190_195_groupi_n_7178, csa_tree_add_190_195_groupi_n_7179, csa_tree_add_190_195_groupi_n_7180, csa_tree_add_190_195_groupi_n_7181, csa_tree_add_190_195_groupi_n_7182, csa_tree_add_190_195_groupi_n_7183;
  wire csa_tree_add_190_195_groupi_n_7184, csa_tree_add_190_195_groupi_n_7185, csa_tree_add_190_195_groupi_n_7186, csa_tree_add_190_195_groupi_n_7187, csa_tree_add_190_195_groupi_n_7188, csa_tree_add_190_195_groupi_n_7189, csa_tree_add_190_195_groupi_n_7190, csa_tree_add_190_195_groupi_n_7191;
  wire csa_tree_add_190_195_groupi_n_7192, csa_tree_add_190_195_groupi_n_7193, csa_tree_add_190_195_groupi_n_7194, csa_tree_add_190_195_groupi_n_7195, csa_tree_add_190_195_groupi_n_7196, csa_tree_add_190_195_groupi_n_7197, csa_tree_add_190_195_groupi_n_7198, csa_tree_add_190_195_groupi_n_7199;
  wire csa_tree_add_190_195_groupi_n_7200, csa_tree_add_190_195_groupi_n_7201, csa_tree_add_190_195_groupi_n_7202, csa_tree_add_190_195_groupi_n_7203, csa_tree_add_190_195_groupi_n_7204, csa_tree_add_190_195_groupi_n_7205, csa_tree_add_190_195_groupi_n_7206, csa_tree_add_190_195_groupi_n_7207;
  wire csa_tree_add_190_195_groupi_n_7208, csa_tree_add_190_195_groupi_n_7209, csa_tree_add_190_195_groupi_n_7210, csa_tree_add_190_195_groupi_n_7211, csa_tree_add_190_195_groupi_n_7212, csa_tree_add_190_195_groupi_n_7213, csa_tree_add_190_195_groupi_n_7214, csa_tree_add_190_195_groupi_n_7215;
  wire csa_tree_add_190_195_groupi_n_7216, csa_tree_add_190_195_groupi_n_7217, csa_tree_add_190_195_groupi_n_7218, csa_tree_add_190_195_groupi_n_7219, csa_tree_add_190_195_groupi_n_7220, csa_tree_add_190_195_groupi_n_7221, csa_tree_add_190_195_groupi_n_7222, csa_tree_add_190_195_groupi_n_7223;
  wire csa_tree_add_190_195_groupi_n_7224, csa_tree_add_190_195_groupi_n_7225, csa_tree_add_190_195_groupi_n_7226, csa_tree_add_190_195_groupi_n_7227, csa_tree_add_190_195_groupi_n_7228, csa_tree_add_190_195_groupi_n_7229, csa_tree_add_190_195_groupi_n_7230, csa_tree_add_190_195_groupi_n_7231;
  wire csa_tree_add_190_195_groupi_n_7232, csa_tree_add_190_195_groupi_n_7233, csa_tree_add_190_195_groupi_n_7234, csa_tree_add_190_195_groupi_n_7235, csa_tree_add_190_195_groupi_n_7236, csa_tree_add_190_195_groupi_n_7237, csa_tree_add_190_195_groupi_n_7238, csa_tree_add_190_195_groupi_n_7239;
  wire csa_tree_add_190_195_groupi_n_7240, csa_tree_add_190_195_groupi_n_7241, csa_tree_add_190_195_groupi_n_7242, csa_tree_add_190_195_groupi_n_7243, csa_tree_add_190_195_groupi_n_7244, csa_tree_add_190_195_groupi_n_7245, csa_tree_add_190_195_groupi_n_7246, csa_tree_add_190_195_groupi_n_7247;
  wire csa_tree_add_190_195_groupi_n_7248, csa_tree_add_190_195_groupi_n_7249, csa_tree_add_190_195_groupi_n_7250, csa_tree_add_190_195_groupi_n_7251, csa_tree_add_190_195_groupi_n_7252, csa_tree_add_190_195_groupi_n_7253, csa_tree_add_190_195_groupi_n_7254, csa_tree_add_190_195_groupi_n_7255;
  wire csa_tree_add_190_195_groupi_n_7256, csa_tree_add_190_195_groupi_n_7257, csa_tree_add_190_195_groupi_n_7258, csa_tree_add_190_195_groupi_n_7259, csa_tree_add_190_195_groupi_n_7260, csa_tree_add_190_195_groupi_n_7261, csa_tree_add_190_195_groupi_n_7262, csa_tree_add_190_195_groupi_n_7263;
  wire csa_tree_add_190_195_groupi_n_7264, csa_tree_add_190_195_groupi_n_7265, csa_tree_add_190_195_groupi_n_7266, csa_tree_add_190_195_groupi_n_7267, csa_tree_add_190_195_groupi_n_7268, csa_tree_add_190_195_groupi_n_7269, csa_tree_add_190_195_groupi_n_7270, csa_tree_add_190_195_groupi_n_7271;
  wire csa_tree_add_190_195_groupi_n_7272, csa_tree_add_190_195_groupi_n_7273, csa_tree_add_190_195_groupi_n_7274, csa_tree_add_190_195_groupi_n_7275, csa_tree_add_190_195_groupi_n_7276, csa_tree_add_190_195_groupi_n_7277, csa_tree_add_190_195_groupi_n_7278, csa_tree_add_190_195_groupi_n_7279;
  wire csa_tree_add_190_195_groupi_n_7280, csa_tree_add_190_195_groupi_n_7281, csa_tree_add_190_195_groupi_n_7282, csa_tree_add_190_195_groupi_n_7283, csa_tree_add_190_195_groupi_n_7284, csa_tree_add_190_195_groupi_n_7285, csa_tree_add_190_195_groupi_n_7286, csa_tree_add_190_195_groupi_n_7287;
  wire csa_tree_add_190_195_groupi_n_7288, csa_tree_add_190_195_groupi_n_7289, csa_tree_add_190_195_groupi_n_7290, csa_tree_add_190_195_groupi_n_7291, csa_tree_add_190_195_groupi_n_7292, csa_tree_add_190_195_groupi_n_7293, csa_tree_add_190_195_groupi_n_7294, csa_tree_add_190_195_groupi_n_7295;
  wire csa_tree_add_190_195_groupi_n_7296, csa_tree_add_190_195_groupi_n_7297, csa_tree_add_190_195_groupi_n_7298, csa_tree_add_190_195_groupi_n_7299, csa_tree_add_190_195_groupi_n_7300, csa_tree_add_190_195_groupi_n_7301, csa_tree_add_190_195_groupi_n_7302, csa_tree_add_190_195_groupi_n_7303;
  wire csa_tree_add_190_195_groupi_n_7304, csa_tree_add_190_195_groupi_n_7305, csa_tree_add_190_195_groupi_n_7306, csa_tree_add_190_195_groupi_n_7307, csa_tree_add_190_195_groupi_n_7308, csa_tree_add_190_195_groupi_n_7309, csa_tree_add_190_195_groupi_n_7310, csa_tree_add_190_195_groupi_n_7311;
  wire csa_tree_add_190_195_groupi_n_7312, csa_tree_add_190_195_groupi_n_7313, csa_tree_add_190_195_groupi_n_7314, csa_tree_add_190_195_groupi_n_7315, csa_tree_add_190_195_groupi_n_7316, csa_tree_add_190_195_groupi_n_7317, csa_tree_add_190_195_groupi_n_7318, csa_tree_add_190_195_groupi_n_7319;
  wire csa_tree_add_190_195_groupi_n_7320, csa_tree_add_190_195_groupi_n_7321, csa_tree_add_190_195_groupi_n_7322, csa_tree_add_190_195_groupi_n_7323, csa_tree_add_190_195_groupi_n_7324, csa_tree_add_190_195_groupi_n_7325, csa_tree_add_190_195_groupi_n_7326, csa_tree_add_190_195_groupi_n_7327;
  wire csa_tree_add_190_195_groupi_n_7328, csa_tree_add_190_195_groupi_n_7329, csa_tree_add_190_195_groupi_n_7330, csa_tree_add_190_195_groupi_n_7331, csa_tree_add_190_195_groupi_n_7332, csa_tree_add_190_195_groupi_n_7333, csa_tree_add_190_195_groupi_n_7334, csa_tree_add_190_195_groupi_n_7335;
  wire csa_tree_add_190_195_groupi_n_7336, csa_tree_add_190_195_groupi_n_7337, csa_tree_add_190_195_groupi_n_7338, csa_tree_add_190_195_groupi_n_7339, csa_tree_add_190_195_groupi_n_7340, csa_tree_add_190_195_groupi_n_7341, csa_tree_add_190_195_groupi_n_7342, csa_tree_add_190_195_groupi_n_7343;
  wire csa_tree_add_190_195_groupi_n_7344, csa_tree_add_190_195_groupi_n_7345, csa_tree_add_190_195_groupi_n_7346, csa_tree_add_190_195_groupi_n_7347, csa_tree_add_190_195_groupi_n_7348, csa_tree_add_190_195_groupi_n_7349, csa_tree_add_190_195_groupi_n_7350, csa_tree_add_190_195_groupi_n_7351;
  wire csa_tree_add_190_195_groupi_n_7352, csa_tree_add_190_195_groupi_n_7353, csa_tree_add_190_195_groupi_n_7354, csa_tree_add_190_195_groupi_n_7355, csa_tree_add_190_195_groupi_n_7356, csa_tree_add_190_195_groupi_n_7357, csa_tree_add_190_195_groupi_n_7358, csa_tree_add_190_195_groupi_n_7359;
  wire csa_tree_add_190_195_groupi_n_7360, csa_tree_add_190_195_groupi_n_7361, csa_tree_add_190_195_groupi_n_7362, csa_tree_add_190_195_groupi_n_7363, csa_tree_add_190_195_groupi_n_7364, csa_tree_add_190_195_groupi_n_7365, csa_tree_add_190_195_groupi_n_7366, csa_tree_add_190_195_groupi_n_7367;
  wire csa_tree_add_190_195_groupi_n_7368, csa_tree_add_190_195_groupi_n_7369, csa_tree_add_190_195_groupi_n_7370, csa_tree_add_190_195_groupi_n_7371, csa_tree_add_190_195_groupi_n_7372, csa_tree_add_190_195_groupi_n_7373, csa_tree_add_190_195_groupi_n_7374, csa_tree_add_190_195_groupi_n_7375;
  wire csa_tree_add_190_195_groupi_n_7376, csa_tree_add_190_195_groupi_n_7377, csa_tree_add_190_195_groupi_n_7378, csa_tree_add_190_195_groupi_n_7379, csa_tree_add_190_195_groupi_n_7380, csa_tree_add_190_195_groupi_n_7381, csa_tree_add_190_195_groupi_n_7382, csa_tree_add_190_195_groupi_n_7383;
  wire csa_tree_add_190_195_groupi_n_7384, csa_tree_add_190_195_groupi_n_7385, csa_tree_add_190_195_groupi_n_7386, csa_tree_add_190_195_groupi_n_7387, csa_tree_add_190_195_groupi_n_7388, csa_tree_add_190_195_groupi_n_7389, csa_tree_add_190_195_groupi_n_7390, csa_tree_add_190_195_groupi_n_7391;
  wire csa_tree_add_190_195_groupi_n_7392, csa_tree_add_190_195_groupi_n_7393, csa_tree_add_190_195_groupi_n_7394, csa_tree_add_190_195_groupi_n_7395, csa_tree_add_190_195_groupi_n_7396, csa_tree_add_190_195_groupi_n_7397, csa_tree_add_190_195_groupi_n_7398, csa_tree_add_190_195_groupi_n_7399;
  wire csa_tree_add_190_195_groupi_n_7400, csa_tree_add_190_195_groupi_n_7401, csa_tree_add_190_195_groupi_n_7402, csa_tree_add_190_195_groupi_n_7403, csa_tree_add_190_195_groupi_n_7404, csa_tree_add_190_195_groupi_n_7405, csa_tree_add_190_195_groupi_n_7406, csa_tree_add_190_195_groupi_n_7407;
  wire csa_tree_add_190_195_groupi_n_7408, csa_tree_add_190_195_groupi_n_7409, csa_tree_add_190_195_groupi_n_7410, csa_tree_add_190_195_groupi_n_7411, csa_tree_add_190_195_groupi_n_7412, csa_tree_add_190_195_groupi_n_7413, csa_tree_add_190_195_groupi_n_7414, csa_tree_add_190_195_groupi_n_7415;
  wire csa_tree_add_190_195_groupi_n_7416, csa_tree_add_190_195_groupi_n_7417, csa_tree_add_190_195_groupi_n_7418, csa_tree_add_190_195_groupi_n_7419, csa_tree_add_190_195_groupi_n_7420, csa_tree_add_190_195_groupi_n_7421, csa_tree_add_190_195_groupi_n_7422, csa_tree_add_190_195_groupi_n_7423;
  wire csa_tree_add_190_195_groupi_n_7424, csa_tree_add_190_195_groupi_n_7425, csa_tree_add_190_195_groupi_n_7426, csa_tree_add_190_195_groupi_n_7427, csa_tree_add_190_195_groupi_n_7428, csa_tree_add_190_195_groupi_n_7429, csa_tree_add_190_195_groupi_n_7430, csa_tree_add_190_195_groupi_n_7431;
  wire csa_tree_add_190_195_groupi_n_7432, csa_tree_add_190_195_groupi_n_7433, csa_tree_add_190_195_groupi_n_7434, csa_tree_add_190_195_groupi_n_7435, csa_tree_add_190_195_groupi_n_7436, csa_tree_add_190_195_groupi_n_7437, csa_tree_add_190_195_groupi_n_7438, csa_tree_add_190_195_groupi_n_7439;
  wire csa_tree_add_190_195_groupi_n_7440, csa_tree_add_190_195_groupi_n_7441, csa_tree_add_190_195_groupi_n_7442, csa_tree_add_190_195_groupi_n_7443, csa_tree_add_190_195_groupi_n_7444, csa_tree_add_190_195_groupi_n_7445, csa_tree_add_190_195_groupi_n_7446, csa_tree_add_190_195_groupi_n_7447;
  wire csa_tree_add_190_195_groupi_n_7448, csa_tree_add_190_195_groupi_n_7449, csa_tree_add_190_195_groupi_n_7450, csa_tree_add_190_195_groupi_n_7451, csa_tree_add_190_195_groupi_n_7452, csa_tree_add_190_195_groupi_n_7453, csa_tree_add_190_195_groupi_n_7454, csa_tree_add_190_195_groupi_n_7455;
  wire csa_tree_add_190_195_groupi_n_7456, csa_tree_add_190_195_groupi_n_7457, csa_tree_add_190_195_groupi_n_7458, csa_tree_add_190_195_groupi_n_7459, csa_tree_add_190_195_groupi_n_7460, csa_tree_add_190_195_groupi_n_7461, csa_tree_add_190_195_groupi_n_7462, csa_tree_add_190_195_groupi_n_7463;
  wire csa_tree_add_190_195_groupi_n_7464, csa_tree_add_190_195_groupi_n_7465, csa_tree_add_190_195_groupi_n_7466, csa_tree_add_190_195_groupi_n_7467, csa_tree_add_190_195_groupi_n_7468, csa_tree_add_190_195_groupi_n_7469, csa_tree_add_190_195_groupi_n_7470, csa_tree_add_190_195_groupi_n_7471;
  wire csa_tree_add_190_195_groupi_n_7472, csa_tree_add_190_195_groupi_n_7473, csa_tree_add_190_195_groupi_n_7474, csa_tree_add_190_195_groupi_n_7475, csa_tree_add_190_195_groupi_n_7476, csa_tree_add_190_195_groupi_n_7477, csa_tree_add_190_195_groupi_n_7478, csa_tree_add_190_195_groupi_n_7479;
  wire csa_tree_add_190_195_groupi_n_7480, csa_tree_add_190_195_groupi_n_7481, csa_tree_add_190_195_groupi_n_7482, csa_tree_add_190_195_groupi_n_7483, csa_tree_add_190_195_groupi_n_7484, csa_tree_add_190_195_groupi_n_7485, csa_tree_add_190_195_groupi_n_7486, csa_tree_add_190_195_groupi_n_7487;
  wire csa_tree_add_190_195_groupi_n_7488, csa_tree_add_190_195_groupi_n_7489, csa_tree_add_190_195_groupi_n_7490, csa_tree_add_190_195_groupi_n_7491, csa_tree_add_190_195_groupi_n_7492, csa_tree_add_190_195_groupi_n_7493, csa_tree_add_190_195_groupi_n_7494, csa_tree_add_190_195_groupi_n_7495;
  wire csa_tree_add_190_195_groupi_n_7496, csa_tree_add_190_195_groupi_n_7497, csa_tree_add_190_195_groupi_n_7498, csa_tree_add_190_195_groupi_n_7499, csa_tree_add_190_195_groupi_n_7500, csa_tree_add_190_195_groupi_n_7501, csa_tree_add_190_195_groupi_n_7502, csa_tree_add_190_195_groupi_n_7503;
  wire csa_tree_add_190_195_groupi_n_7504, csa_tree_add_190_195_groupi_n_7505, csa_tree_add_190_195_groupi_n_7506, csa_tree_add_190_195_groupi_n_7507, csa_tree_add_190_195_groupi_n_7508, csa_tree_add_190_195_groupi_n_7509, csa_tree_add_190_195_groupi_n_7510, csa_tree_add_190_195_groupi_n_7511;
  wire csa_tree_add_190_195_groupi_n_7512, csa_tree_add_190_195_groupi_n_7513, csa_tree_add_190_195_groupi_n_7514, csa_tree_add_190_195_groupi_n_7515, csa_tree_add_190_195_groupi_n_7516, csa_tree_add_190_195_groupi_n_7517, csa_tree_add_190_195_groupi_n_7518, csa_tree_add_190_195_groupi_n_7519;
  wire csa_tree_add_190_195_groupi_n_7520, csa_tree_add_190_195_groupi_n_7521, csa_tree_add_190_195_groupi_n_7522, csa_tree_add_190_195_groupi_n_7523, csa_tree_add_190_195_groupi_n_7524, csa_tree_add_190_195_groupi_n_7525, csa_tree_add_190_195_groupi_n_7526, csa_tree_add_190_195_groupi_n_7527;
  wire csa_tree_add_190_195_groupi_n_7528, csa_tree_add_190_195_groupi_n_7529, csa_tree_add_190_195_groupi_n_7530, csa_tree_add_190_195_groupi_n_7531, csa_tree_add_190_195_groupi_n_7532, csa_tree_add_190_195_groupi_n_7533, csa_tree_add_190_195_groupi_n_7534, csa_tree_add_190_195_groupi_n_7535;
  wire csa_tree_add_190_195_groupi_n_7536, csa_tree_add_190_195_groupi_n_7537, csa_tree_add_190_195_groupi_n_7538, csa_tree_add_190_195_groupi_n_7539, csa_tree_add_190_195_groupi_n_7540, csa_tree_add_190_195_groupi_n_7541, csa_tree_add_190_195_groupi_n_7542, csa_tree_add_190_195_groupi_n_7543;
  wire csa_tree_add_190_195_groupi_n_7544, csa_tree_add_190_195_groupi_n_7545, csa_tree_add_190_195_groupi_n_7546, csa_tree_add_190_195_groupi_n_7547, csa_tree_add_190_195_groupi_n_7548, csa_tree_add_190_195_groupi_n_7549, csa_tree_add_190_195_groupi_n_7550, csa_tree_add_190_195_groupi_n_7551;
  wire csa_tree_add_190_195_groupi_n_7552, csa_tree_add_190_195_groupi_n_7553, csa_tree_add_190_195_groupi_n_7554, csa_tree_add_190_195_groupi_n_7555, csa_tree_add_190_195_groupi_n_7556, csa_tree_add_190_195_groupi_n_7557, csa_tree_add_190_195_groupi_n_7558, csa_tree_add_190_195_groupi_n_7559;
  wire csa_tree_add_190_195_groupi_n_7560, csa_tree_add_190_195_groupi_n_7561, csa_tree_add_190_195_groupi_n_7562, csa_tree_add_190_195_groupi_n_7563, csa_tree_add_190_195_groupi_n_7564, csa_tree_add_190_195_groupi_n_7565, csa_tree_add_190_195_groupi_n_7566, csa_tree_add_190_195_groupi_n_7567;
  wire csa_tree_add_190_195_groupi_n_7568, csa_tree_add_190_195_groupi_n_7569, csa_tree_add_190_195_groupi_n_7570, csa_tree_add_190_195_groupi_n_7571, csa_tree_add_190_195_groupi_n_7572, csa_tree_add_190_195_groupi_n_7573, csa_tree_add_190_195_groupi_n_7574, csa_tree_add_190_195_groupi_n_7575;
  wire csa_tree_add_190_195_groupi_n_7576, csa_tree_add_190_195_groupi_n_7577, csa_tree_add_190_195_groupi_n_7578, csa_tree_add_190_195_groupi_n_7579, csa_tree_add_190_195_groupi_n_7580, csa_tree_add_190_195_groupi_n_7581, csa_tree_add_190_195_groupi_n_7582, csa_tree_add_190_195_groupi_n_7583;
  wire csa_tree_add_190_195_groupi_n_7584, csa_tree_add_190_195_groupi_n_7585, csa_tree_add_190_195_groupi_n_7586, csa_tree_add_190_195_groupi_n_7587, csa_tree_add_190_195_groupi_n_7588, csa_tree_add_190_195_groupi_n_7589, csa_tree_add_190_195_groupi_n_7590, csa_tree_add_190_195_groupi_n_7591;
  wire csa_tree_add_190_195_groupi_n_7592, csa_tree_add_190_195_groupi_n_7593, csa_tree_add_190_195_groupi_n_7594, csa_tree_add_190_195_groupi_n_7595, csa_tree_add_190_195_groupi_n_7596, csa_tree_add_190_195_groupi_n_7597, csa_tree_add_190_195_groupi_n_7598, csa_tree_add_190_195_groupi_n_7599;
  wire csa_tree_add_190_195_groupi_n_7600, csa_tree_add_190_195_groupi_n_7601, csa_tree_add_190_195_groupi_n_7602, csa_tree_add_190_195_groupi_n_7603, csa_tree_add_190_195_groupi_n_7604, csa_tree_add_190_195_groupi_n_7605, csa_tree_add_190_195_groupi_n_7606, csa_tree_add_190_195_groupi_n_7607;
  wire csa_tree_add_190_195_groupi_n_7608, csa_tree_add_190_195_groupi_n_7609, csa_tree_add_190_195_groupi_n_7610, csa_tree_add_190_195_groupi_n_7611, csa_tree_add_190_195_groupi_n_7612, csa_tree_add_190_195_groupi_n_7613, csa_tree_add_190_195_groupi_n_7614, csa_tree_add_190_195_groupi_n_7615;
  wire csa_tree_add_190_195_groupi_n_7616, csa_tree_add_190_195_groupi_n_7617, csa_tree_add_190_195_groupi_n_7618, csa_tree_add_190_195_groupi_n_7619, csa_tree_add_190_195_groupi_n_7620, csa_tree_add_190_195_groupi_n_7621, csa_tree_add_190_195_groupi_n_7622, csa_tree_add_190_195_groupi_n_7623;
  wire csa_tree_add_190_195_groupi_n_7624, csa_tree_add_190_195_groupi_n_7625, csa_tree_add_190_195_groupi_n_7626, csa_tree_add_190_195_groupi_n_7627, csa_tree_add_190_195_groupi_n_7628, csa_tree_add_190_195_groupi_n_7629, csa_tree_add_190_195_groupi_n_7630, csa_tree_add_190_195_groupi_n_7631;
  wire csa_tree_add_190_195_groupi_n_7632, csa_tree_add_190_195_groupi_n_7633, csa_tree_add_190_195_groupi_n_7634, csa_tree_add_190_195_groupi_n_7635, csa_tree_add_190_195_groupi_n_7636, csa_tree_add_190_195_groupi_n_7637, csa_tree_add_190_195_groupi_n_7638, csa_tree_add_190_195_groupi_n_7639;
  wire csa_tree_add_190_195_groupi_n_7640, csa_tree_add_190_195_groupi_n_7641, csa_tree_add_190_195_groupi_n_7642, csa_tree_add_190_195_groupi_n_7643, csa_tree_add_190_195_groupi_n_7644, csa_tree_add_190_195_groupi_n_7645, csa_tree_add_190_195_groupi_n_7646, csa_tree_add_190_195_groupi_n_7647;
  wire csa_tree_add_190_195_groupi_n_7648, csa_tree_add_190_195_groupi_n_7649, csa_tree_add_190_195_groupi_n_7650, csa_tree_add_190_195_groupi_n_7651, csa_tree_add_190_195_groupi_n_7652, csa_tree_add_190_195_groupi_n_7653, csa_tree_add_190_195_groupi_n_7654, csa_tree_add_190_195_groupi_n_7655;
  wire csa_tree_add_190_195_groupi_n_7656, csa_tree_add_190_195_groupi_n_7657, csa_tree_add_190_195_groupi_n_7658, csa_tree_add_190_195_groupi_n_7659, csa_tree_add_190_195_groupi_n_7660, csa_tree_add_190_195_groupi_n_7661, csa_tree_add_190_195_groupi_n_7662, csa_tree_add_190_195_groupi_n_7663;
  wire csa_tree_add_190_195_groupi_n_7664, csa_tree_add_190_195_groupi_n_7665, csa_tree_add_190_195_groupi_n_7666, csa_tree_add_190_195_groupi_n_7667, csa_tree_add_190_195_groupi_n_7668, csa_tree_add_190_195_groupi_n_7669, csa_tree_add_190_195_groupi_n_7670, csa_tree_add_190_195_groupi_n_7671;
  wire csa_tree_add_190_195_groupi_n_7672, csa_tree_add_190_195_groupi_n_7673, csa_tree_add_190_195_groupi_n_7674, csa_tree_add_190_195_groupi_n_7675, csa_tree_add_190_195_groupi_n_7676, csa_tree_add_190_195_groupi_n_7677, csa_tree_add_190_195_groupi_n_7678, csa_tree_add_190_195_groupi_n_7679;
  wire csa_tree_add_190_195_groupi_n_7680, csa_tree_add_190_195_groupi_n_7681, csa_tree_add_190_195_groupi_n_7682, csa_tree_add_190_195_groupi_n_7683, csa_tree_add_190_195_groupi_n_7684, csa_tree_add_190_195_groupi_n_7685, csa_tree_add_190_195_groupi_n_7686, csa_tree_add_190_195_groupi_n_7687;
  wire csa_tree_add_190_195_groupi_n_7688, csa_tree_add_190_195_groupi_n_7689, csa_tree_add_190_195_groupi_n_7690, csa_tree_add_190_195_groupi_n_7691, csa_tree_add_190_195_groupi_n_7692, csa_tree_add_190_195_groupi_n_7693, csa_tree_add_190_195_groupi_n_7694, csa_tree_add_190_195_groupi_n_7695;
  wire csa_tree_add_190_195_groupi_n_7696, csa_tree_add_190_195_groupi_n_7697, csa_tree_add_190_195_groupi_n_7698, csa_tree_add_190_195_groupi_n_7699, csa_tree_add_190_195_groupi_n_7700, csa_tree_add_190_195_groupi_n_7701, csa_tree_add_190_195_groupi_n_7702, csa_tree_add_190_195_groupi_n_7703;
  wire csa_tree_add_190_195_groupi_n_7704, csa_tree_add_190_195_groupi_n_7705, csa_tree_add_190_195_groupi_n_7706, csa_tree_add_190_195_groupi_n_7707, csa_tree_add_190_195_groupi_n_7708, csa_tree_add_190_195_groupi_n_7709, csa_tree_add_190_195_groupi_n_7710, csa_tree_add_190_195_groupi_n_7711;
  wire csa_tree_add_190_195_groupi_n_7712, csa_tree_add_190_195_groupi_n_7713, csa_tree_add_190_195_groupi_n_7714, csa_tree_add_190_195_groupi_n_7715, csa_tree_add_190_195_groupi_n_7716, csa_tree_add_190_195_groupi_n_7717, csa_tree_add_190_195_groupi_n_7718, csa_tree_add_190_195_groupi_n_7719;
  wire csa_tree_add_190_195_groupi_n_7720, csa_tree_add_190_195_groupi_n_7721, csa_tree_add_190_195_groupi_n_7722, csa_tree_add_190_195_groupi_n_7723, csa_tree_add_190_195_groupi_n_7724, csa_tree_add_190_195_groupi_n_7725, csa_tree_add_190_195_groupi_n_7726, csa_tree_add_190_195_groupi_n_7727;
  wire csa_tree_add_190_195_groupi_n_7728, csa_tree_add_190_195_groupi_n_7729, csa_tree_add_190_195_groupi_n_7730, csa_tree_add_190_195_groupi_n_7731, csa_tree_add_190_195_groupi_n_7732, csa_tree_add_190_195_groupi_n_7733, csa_tree_add_190_195_groupi_n_7734, csa_tree_add_190_195_groupi_n_7735;
  wire csa_tree_add_190_195_groupi_n_7736, csa_tree_add_190_195_groupi_n_7737, csa_tree_add_190_195_groupi_n_7738, csa_tree_add_190_195_groupi_n_7739, csa_tree_add_190_195_groupi_n_7740, csa_tree_add_190_195_groupi_n_7741, csa_tree_add_190_195_groupi_n_7742, csa_tree_add_190_195_groupi_n_7743;
  wire csa_tree_add_190_195_groupi_n_7744, csa_tree_add_190_195_groupi_n_7745, csa_tree_add_190_195_groupi_n_7746, csa_tree_add_190_195_groupi_n_7747, csa_tree_add_190_195_groupi_n_7748, csa_tree_add_190_195_groupi_n_7749, csa_tree_add_190_195_groupi_n_7750, csa_tree_add_190_195_groupi_n_7751;
  wire csa_tree_add_190_195_groupi_n_7752, csa_tree_add_190_195_groupi_n_7753, csa_tree_add_190_195_groupi_n_7754, csa_tree_add_190_195_groupi_n_7755, csa_tree_add_190_195_groupi_n_7756, csa_tree_add_190_195_groupi_n_7757, csa_tree_add_190_195_groupi_n_7758, csa_tree_add_190_195_groupi_n_7759;
  wire csa_tree_add_190_195_groupi_n_7760, csa_tree_add_190_195_groupi_n_7761, csa_tree_add_190_195_groupi_n_7762, csa_tree_add_190_195_groupi_n_7763, csa_tree_add_190_195_groupi_n_7764, csa_tree_add_190_195_groupi_n_7765, csa_tree_add_190_195_groupi_n_7766, csa_tree_add_190_195_groupi_n_7767;
  wire csa_tree_add_190_195_groupi_n_7768, csa_tree_add_190_195_groupi_n_7769, csa_tree_add_190_195_groupi_n_7770, csa_tree_add_190_195_groupi_n_7771, csa_tree_add_190_195_groupi_n_7772, csa_tree_add_190_195_groupi_n_7773, csa_tree_add_190_195_groupi_n_7774, csa_tree_add_190_195_groupi_n_7775;
  wire csa_tree_add_190_195_groupi_n_7776, csa_tree_add_190_195_groupi_n_7777, csa_tree_add_190_195_groupi_n_7778, csa_tree_add_190_195_groupi_n_7779, csa_tree_add_190_195_groupi_n_7780, csa_tree_add_190_195_groupi_n_7781, csa_tree_add_190_195_groupi_n_7782, csa_tree_add_190_195_groupi_n_7783;
  wire csa_tree_add_190_195_groupi_n_7784, csa_tree_add_190_195_groupi_n_7785, csa_tree_add_190_195_groupi_n_7786, csa_tree_add_190_195_groupi_n_7787, csa_tree_add_190_195_groupi_n_7788, csa_tree_add_190_195_groupi_n_7789, csa_tree_add_190_195_groupi_n_7790, csa_tree_add_190_195_groupi_n_7791;
  wire csa_tree_add_190_195_groupi_n_7792, csa_tree_add_190_195_groupi_n_7793, csa_tree_add_190_195_groupi_n_7794, csa_tree_add_190_195_groupi_n_7795, csa_tree_add_190_195_groupi_n_7796, csa_tree_add_190_195_groupi_n_7797, csa_tree_add_190_195_groupi_n_7798, csa_tree_add_190_195_groupi_n_7799;
  wire csa_tree_add_190_195_groupi_n_7800, csa_tree_add_190_195_groupi_n_7801, csa_tree_add_190_195_groupi_n_7802, csa_tree_add_190_195_groupi_n_7803, csa_tree_add_190_195_groupi_n_7804, csa_tree_add_190_195_groupi_n_7805, csa_tree_add_190_195_groupi_n_7806, csa_tree_add_190_195_groupi_n_7807;
  wire csa_tree_add_190_195_groupi_n_7808, csa_tree_add_190_195_groupi_n_7809, csa_tree_add_190_195_groupi_n_7810, csa_tree_add_190_195_groupi_n_7811, csa_tree_add_190_195_groupi_n_7812, csa_tree_add_190_195_groupi_n_7813, csa_tree_add_190_195_groupi_n_7814, csa_tree_add_190_195_groupi_n_7815;
  wire csa_tree_add_190_195_groupi_n_7816, csa_tree_add_190_195_groupi_n_7817, csa_tree_add_190_195_groupi_n_7818, csa_tree_add_190_195_groupi_n_7819, csa_tree_add_190_195_groupi_n_7820, csa_tree_add_190_195_groupi_n_7821, csa_tree_add_190_195_groupi_n_7822, csa_tree_add_190_195_groupi_n_7823;
  wire csa_tree_add_190_195_groupi_n_7824, csa_tree_add_190_195_groupi_n_7825, csa_tree_add_190_195_groupi_n_7826, csa_tree_add_190_195_groupi_n_7827, csa_tree_add_190_195_groupi_n_7828, csa_tree_add_190_195_groupi_n_7829, csa_tree_add_190_195_groupi_n_7830, csa_tree_add_190_195_groupi_n_7831;
  wire csa_tree_add_190_195_groupi_n_7832, csa_tree_add_190_195_groupi_n_7833, csa_tree_add_190_195_groupi_n_7834, csa_tree_add_190_195_groupi_n_7835, csa_tree_add_190_195_groupi_n_7836, csa_tree_add_190_195_groupi_n_7837, csa_tree_add_190_195_groupi_n_7838, csa_tree_add_190_195_groupi_n_7839;
  wire csa_tree_add_190_195_groupi_n_7840, csa_tree_add_190_195_groupi_n_7841, csa_tree_add_190_195_groupi_n_7842, csa_tree_add_190_195_groupi_n_7843, csa_tree_add_190_195_groupi_n_7844, csa_tree_add_190_195_groupi_n_7845, csa_tree_add_190_195_groupi_n_7846, csa_tree_add_190_195_groupi_n_7847;
  wire csa_tree_add_190_195_groupi_n_7848, csa_tree_add_190_195_groupi_n_7849, csa_tree_add_190_195_groupi_n_7850, csa_tree_add_190_195_groupi_n_7851, csa_tree_add_190_195_groupi_n_7852, csa_tree_add_190_195_groupi_n_7853, csa_tree_add_190_195_groupi_n_7854, csa_tree_add_190_195_groupi_n_7855;
  wire csa_tree_add_190_195_groupi_n_7856, csa_tree_add_190_195_groupi_n_7857, csa_tree_add_190_195_groupi_n_7858, csa_tree_add_190_195_groupi_n_7859, csa_tree_add_190_195_groupi_n_7860, csa_tree_add_190_195_groupi_n_7861, csa_tree_add_190_195_groupi_n_7862, csa_tree_add_190_195_groupi_n_7863;
  wire csa_tree_add_190_195_groupi_n_7864, csa_tree_add_190_195_groupi_n_7865, csa_tree_add_190_195_groupi_n_7866, csa_tree_add_190_195_groupi_n_7867, csa_tree_add_190_195_groupi_n_7868, csa_tree_add_190_195_groupi_n_7869, csa_tree_add_190_195_groupi_n_7870, csa_tree_add_190_195_groupi_n_7871;
  wire csa_tree_add_190_195_groupi_n_7872, csa_tree_add_190_195_groupi_n_7873, csa_tree_add_190_195_groupi_n_7874, csa_tree_add_190_195_groupi_n_7875, csa_tree_add_190_195_groupi_n_7876, csa_tree_add_190_195_groupi_n_7877, csa_tree_add_190_195_groupi_n_7878, csa_tree_add_190_195_groupi_n_7879;
  wire csa_tree_add_190_195_groupi_n_7880, csa_tree_add_190_195_groupi_n_7881, csa_tree_add_190_195_groupi_n_7882, csa_tree_add_190_195_groupi_n_7883, csa_tree_add_190_195_groupi_n_7884, csa_tree_add_190_195_groupi_n_7885, csa_tree_add_190_195_groupi_n_7886, csa_tree_add_190_195_groupi_n_7887;
  wire csa_tree_add_190_195_groupi_n_7888, csa_tree_add_190_195_groupi_n_7889, csa_tree_add_190_195_groupi_n_7890, csa_tree_add_190_195_groupi_n_7891, csa_tree_add_190_195_groupi_n_7892, csa_tree_add_190_195_groupi_n_7893, csa_tree_add_190_195_groupi_n_7894, csa_tree_add_190_195_groupi_n_7895;
  wire csa_tree_add_190_195_groupi_n_7896, csa_tree_add_190_195_groupi_n_7897, csa_tree_add_190_195_groupi_n_7898, csa_tree_add_190_195_groupi_n_7899, csa_tree_add_190_195_groupi_n_7900, csa_tree_add_190_195_groupi_n_7901, csa_tree_add_190_195_groupi_n_7902, csa_tree_add_190_195_groupi_n_7903;
  wire csa_tree_add_190_195_groupi_n_7904, csa_tree_add_190_195_groupi_n_7905, csa_tree_add_190_195_groupi_n_7906, csa_tree_add_190_195_groupi_n_7907, csa_tree_add_190_195_groupi_n_7908, csa_tree_add_190_195_groupi_n_7909, csa_tree_add_190_195_groupi_n_7910, csa_tree_add_190_195_groupi_n_7911;
  wire csa_tree_add_190_195_groupi_n_7912, csa_tree_add_190_195_groupi_n_7913, csa_tree_add_190_195_groupi_n_7914, csa_tree_add_190_195_groupi_n_7915, csa_tree_add_190_195_groupi_n_7916, csa_tree_add_190_195_groupi_n_7917, csa_tree_add_190_195_groupi_n_7918, csa_tree_add_190_195_groupi_n_7919;
  wire csa_tree_add_190_195_groupi_n_7920, csa_tree_add_190_195_groupi_n_7921, csa_tree_add_190_195_groupi_n_7922, csa_tree_add_190_195_groupi_n_7923, csa_tree_add_190_195_groupi_n_7924, csa_tree_add_190_195_groupi_n_7925, csa_tree_add_190_195_groupi_n_7926, csa_tree_add_190_195_groupi_n_7927;
  wire csa_tree_add_190_195_groupi_n_7928, csa_tree_add_190_195_groupi_n_7929, csa_tree_add_190_195_groupi_n_7930, csa_tree_add_190_195_groupi_n_7931, csa_tree_add_190_195_groupi_n_7932, csa_tree_add_190_195_groupi_n_7933, csa_tree_add_190_195_groupi_n_7934, csa_tree_add_190_195_groupi_n_7935;
  wire csa_tree_add_190_195_groupi_n_7936, csa_tree_add_190_195_groupi_n_7937, csa_tree_add_190_195_groupi_n_7938, csa_tree_add_190_195_groupi_n_7939, csa_tree_add_190_195_groupi_n_7940, csa_tree_add_190_195_groupi_n_7941, csa_tree_add_190_195_groupi_n_7942, csa_tree_add_190_195_groupi_n_7943;
  wire csa_tree_add_190_195_groupi_n_7944, csa_tree_add_190_195_groupi_n_7945, csa_tree_add_190_195_groupi_n_7946, csa_tree_add_190_195_groupi_n_7947, csa_tree_add_190_195_groupi_n_7948, csa_tree_add_190_195_groupi_n_7949, csa_tree_add_190_195_groupi_n_7950, csa_tree_add_190_195_groupi_n_7951;
  wire csa_tree_add_190_195_groupi_n_7952, csa_tree_add_190_195_groupi_n_7953, csa_tree_add_190_195_groupi_n_7954, csa_tree_add_190_195_groupi_n_7955, csa_tree_add_190_195_groupi_n_7956, csa_tree_add_190_195_groupi_n_7957, csa_tree_add_190_195_groupi_n_7958, csa_tree_add_190_195_groupi_n_7959;
  wire csa_tree_add_190_195_groupi_n_7960, csa_tree_add_190_195_groupi_n_7961, csa_tree_add_190_195_groupi_n_7962, csa_tree_add_190_195_groupi_n_7963, csa_tree_add_190_195_groupi_n_7964, csa_tree_add_190_195_groupi_n_7965, csa_tree_add_190_195_groupi_n_7966, csa_tree_add_190_195_groupi_n_7967;
  wire csa_tree_add_190_195_groupi_n_7968, csa_tree_add_190_195_groupi_n_7969, csa_tree_add_190_195_groupi_n_7970, csa_tree_add_190_195_groupi_n_7971, csa_tree_add_190_195_groupi_n_7972, csa_tree_add_190_195_groupi_n_7973, csa_tree_add_190_195_groupi_n_7974, csa_tree_add_190_195_groupi_n_7975;
  wire csa_tree_add_190_195_groupi_n_7976, csa_tree_add_190_195_groupi_n_7977, csa_tree_add_190_195_groupi_n_7978, csa_tree_add_190_195_groupi_n_7979, csa_tree_add_190_195_groupi_n_7980, csa_tree_add_190_195_groupi_n_7981, csa_tree_add_190_195_groupi_n_7982, csa_tree_add_190_195_groupi_n_7983;
  wire csa_tree_add_190_195_groupi_n_7984, csa_tree_add_190_195_groupi_n_7985, csa_tree_add_190_195_groupi_n_7986, csa_tree_add_190_195_groupi_n_7987, csa_tree_add_190_195_groupi_n_7988, csa_tree_add_190_195_groupi_n_7989, csa_tree_add_190_195_groupi_n_7990, csa_tree_add_190_195_groupi_n_7991;
  wire csa_tree_add_190_195_groupi_n_7992, csa_tree_add_190_195_groupi_n_7993, csa_tree_add_190_195_groupi_n_7994, csa_tree_add_190_195_groupi_n_7995, csa_tree_add_190_195_groupi_n_7996, csa_tree_add_190_195_groupi_n_7997, csa_tree_add_190_195_groupi_n_7998, csa_tree_add_190_195_groupi_n_7999;
  wire csa_tree_add_190_195_groupi_n_8000, csa_tree_add_190_195_groupi_n_8001, csa_tree_add_190_195_groupi_n_8002, csa_tree_add_190_195_groupi_n_8003, csa_tree_add_190_195_groupi_n_8004, csa_tree_add_190_195_groupi_n_8005, csa_tree_add_190_195_groupi_n_8006, csa_tree_add_190_195_groupi_n_8007;
  wire csa_tree_add_190_195_groupi_n_8008, csa_tree_add_190_195_groupi_n_8009, csa_tree_add_190_195_groupi_n_8010, csa_tree_add_190_195_groupi_n_8011, csa_tree_add_190_195_groupi_n_8012, csa_tree_add_190_195_groupi_n_8013, csa_tree_add_190_195_groupi_n_8014, csa_tree_add_190_195_groupi_n_8015;
  wire csa_tree_add_190_195_groupi_n_8016, csa_tree_add_190_195_groupi_n_8017, csa_tree_add_190_195_groupi_n_8018, csa_tree_add_190_195_groupi_n_8019, csa_tree_add_190_195_groupi_n_8020, csa_tree_add_190_195_groupi_n_8021, csa_tree_add_190_195_groupi_n_8022, csa_tree_add_190_195_groupi_n_8023;
  wire csa_tree_add_190_195_groupi_n_8024, csa_tree_add_190_195_groupi_n_8025, csa_tree_add_190_195_groupi_n_8026, csa_tree_add_190_195_groupi_n_8027, csa_tree_add_190_195_groupi_n_8028, csa_tree_add_190_195_groupi_n_8029, csa_tree_add_190_195_groupi_n_8030, csa_tree_add_190_195_groupi_n_8031;
  wire csa_tree_add_190_195_groupi_n_8032, csa_tree_add_190_195_groupi_n_8033, csa_tree_add_190_195_groupi_n_8034, csa_tree_add_190_195_groupi_n_8035, csa_tree_add_190_195_groupi_n_8036, csa_tree_add_190_195_groupi_n_8037, csa_tree_add_190_195_groupi_n_8038, csa_tree_add_190_195_groupi_n_8039;
  wire csa_tree_add_190_195_groupi_n_8040, csa_tree_add_190_195_groupi_n_8041, csa_tree_add_190_195_groupi_n_8042, csa_tree_add_190_195_groupi_n_8043, csa_tree_add_190_195_groupi_n_8044, csa_tree_add_190_195_groupi_n_8045, csa_tree_add_190_195_groupi_n_8046, csa_tree_add_190_195_groupi_n_8047;
  wire csa_tree_add_190_195_groupi_n_8048, csa_tree_add_190_195_groupi_n_8049, csa_tree_add_190_195_groupi_n_8050, csa_tree_add_190_195_groupi_n_8051, csa_tree_add_190_195_groupi_n_8052, csa_tree_add_190_195_groupi_n_8053, csa_tree_add_190_195_groupi_n_8054, csa_tree_add_190_195_groupi_n_8055;
  wire csa_tree_add_190_195_groupi_n_8056, csa_tree_add_190_195_groupi_n_8057, csa_tree_add_190_195_groupi_n_8058, csa_tree_add_190_195_groupi_n_8059, csa_tree_add_190_195_groupi_n_8060, csa_tree_add_190_195_groupi_n_8061, csa_tree_add_190_195_groupi_n_8062, csa_tree_add_190_195_groupi_n_8063;
  wire csa_tree_add_190_195_groupi_n_8064, csa_tree_add_190_195_groupi_n_8065, csa_tree_add_190_195_groupi_n_8066, csa_tree_add_190_195_groupi_n_8067, csa_tree_add_190_195_groupi_n_8068, csa_tree_add_190_195_groupi_n_8069, csa_tree_add_190_195_groupi_n_8070, csa_tree_add_190_195_groupi_n_8071;
  wire csa_tree_add_190_195_groupi_n_8072, csa_tree_add_190_195_groupi_n_8073, csa_tree_add_190_195_groupi_n_8074, csa_tree_add_190_195_groupi_n_8075, csa_tree_add_190_195_groupi_n_8076, csa_tree_add_190_195_groupi_n_8077, csa_tree_add_190_195_groupi_n_8078, csa_tree_add_190_195_groupi_n_8079;
  wire csa_tree_add_190_195_groupi_n_8080, csa_tree_add_190_195_groupi_n_8081, csa_tree_add_190_195_groupi_n_8082, csa_tree_add_190_195_groupi_n_8083, csa_tree_add_190_195_groupi_n_8084, csa_tree_add_190_195_groupi_n_8085, csa_tree_add_190_195_groupi_n_8086, csa_tree_add_190_195_groupi_n_8087;
  wire csa_tree_add_190_195_groupi_n_8088, csa_tree_add_190_195_groupi_n_8089, csa_tree_add_190_195_groupi_n_8090, csa_tree_add_190_195_groupi_n_8091, csa_tree_add_190_195_groupi_n_8092, csa_tree_add_190_195_groupi_n_8093, csa_tree_add_190_195_groupi_n_8094, csa_tree_add_190_195_groupi_n_8095;
  wire csa_tree_add_190_195_groupi_n_8096, csa_tree_add_190_195_groupi_n_8097, csa_tree_add_190_195_groupi_n_8098, csa_tree_add_190_195_groupi_n_8099, csa_tree_add_190_195_groupi_n_8100, csa_tree_add_190_195_groupi_n_8101, csa_tree_add_190_195_groupi_n_8102, csa_tree_add_190_195_groupi_n_8103;
  wire csa_tree_add_190_195_groupi_n_8104, csa_tree_add_190_195_groupi_n_8105, csa_tree_add_190_195_groupi_n_8106, csa_tree_add_190_195_groupi_n_8107, csa_tree_add_190_195_groupi_n_8108, csa_tree_add_190_195_groupi_n_8109, csa_tree_add_190_195_groupi_n_8110, csa_tree_add_190_195_groupi_n_8111;
  wire csa_tree_add_190_195_groupi_n_8112, csa_tree_add_190_195_groupi_n_8113, csa_tree_add_190_195_groupi_n_8114, csa_tree_add_190_195_groupi_n_8115, csa_tree_add_190_195_groupi_n_8116, csa_tree_add_190_195_groupi_n_8117, csa_tree_add_190_195_groupi_n_8118, csa_tree_add_190_195_groupi_n_8119;
  wire csa_tree_add_190_195_groupi_n_8120, csa_tree_add_190_195_groupi_n_8121, csa_tree_add_190_195_groupi_n_8122, csa_tree_add_190_195_groupi_n_8123, csa_tree_add_190_195_groupi_n_8124, csa_tree_add_190_195_groupi_n_8125, csa_tree_add_190_195_groupi_n_8126, csa_tree_add_190_195_groupi_n_8127;
  wire csa_tree_add_190_195_groupi_n_8128, csa_tree_add_190_195_groupi_n_8129, csa_tree_add_190_195_groupi_n_8130, csa_tree_add_190_195_groupi_n_8131, csa_tree_add_190_195_groupi_n_8132, csa_tree_add_190_195_groupi_n_8133, csa_tree_add_190_195_groupi_n_8134, csa_tree_add_190_195_groupi_n_8135;
  wire csa_tree_add_190_195_groupi_n_8136, csa_tree_add_190_195_groupi_n_8137, csa_tree_add_190_195_groupi_n_8138, csa_tree_add_190_195_groupi_n_8139, csa_tree_add_190_195_groupi_n_8140, csa_tree_add_190_195_groupi_n_8141, csa_tree_add_190_195_groupi_n_8142, csa_tree_add_190_195_groupi_n_8143;
  wire csa_tree_add_190_195_groupi_n_8144, csa_tree_add_190_195_groupi_n_8145, csa_tree_add_190_195_groupi_n_8146, csa_tree_add_190_195_groupi_n_8147, csa_tree_add_190_195_groupi_n_8148, csa_tree_add_190_195_groupi_n_8149, csa_tree_add_190_195_groupi_n_8150, csa_tree_add_190_195_groupi_n_8151;
  wire csa_tree_add_190_195_groupi_n_8152, csa_tree_add_190_195_groupi_n_8153, csa_tree_add_190_195_groupi_n_8154, csa_tree_add_190_195_groupi_n_8155, csa_tree_add_190_195_groupi_n_8156, csa_tree_add_190_195_groupi_n_8157, csa_tree_add_190_195_groupi_n_8158, csa_tree_add_190_195_groupi_n_8159;
  wire csa_tree_add_190_195_groupi_n_8160, csa_tree_add_190_195_groupi_n_8161, csa_tree_add_190_195_groupi_n_8162, csa_tree_add_190_195_groupi_n_8163, csa_tree_add_190_195_groupi_n_8164, csa_tree_add_190_195_groupi_n_8165, csa_tree_add_190_195_groupi_n_8166, csa_tree_add_190_195_groupi_n_8167;
  wire csa_tree_add_190_195_groupi_n_8168, csa_tree_add_190_195_groupi_n_8169, csa_tree_add_190_195_groupi_n_8170, csa_tree_add_190_195_groupi_n_8171, csa_tree_add_190_195_groupi_n_8172, csa_tree_add_190_195_groupi_n_8173, csa_tree_add_190_195_groupi_n_8174, csa_tree_add_190_195_groupi_n_8175;
  wire csa_tree_add_190_195_groupi_n_8176, csa_tree_add_190_195_groupi_n_8177, csa_tree_add_190_195_groupi_n_8178, csa_tree_add_190_195_groupi_n_8179, csa_tree_add_190_195_groupi_n_8180, csa_tree_add_190_195_groupi_n_8181, csa_tree_add_190_195_groupi_n_8182, csa_tree_add_190_195_groupi_n_8183;
  wire csa_tree_add_190_195_groupi_n_8184, csa_tree_add_190_195_groupi_n_8185, csa_tree_add_190_195_groupi_n_8186, csa_tree_add_190_195_groupi_n_8187, csa_tree_add_190_195_groupi_n_8188, csa_tree_add_190_195_groupi_n_8189, csa_tree_add_190_195_groupi_n_8190, csa_tree_add_190_195_groupi_n_8191;
  wire csa_tree_add_190_195_groupi_n_8192, csa_tree_add_190_195_groupi_n_8193, csa_tree_add_190_195_groupi_n_8194, csa_tree_add_190_195_groupi_n_8195, csa_tree_add_190_195_groupi_n_8196, csa_tree_add_190_195_groupi_n_8197, csa_tree_add_190_195_groupi_n_8198, csa_tree_add_190_195_groupi_n_8199;
  wire csa_tree_add_190_195_groupi_n_8200, csa_tree_add_190_195_groupi_n_8201, csa_tree_add_190_195_groupi_n_8202, csa_tree_add_190_195_groupi_n_8203, csa_tree_add_190_195_groupi_n_8204, csa_tree_add_190_195_groupi_n_8205, csa_tree_add_190_195_groupi_n_8206, csa_tree_add_190_195_groupi_n_8207;
  wire csa_tree_add_190_195_groupi_n_8208, csa_tree_add_190_195_groupi_n_8209, csa_tree_add_190_195_groupi_n_8210, csa_tree_add_190_195_groupi_n_8211, csa_tree_add_190_195_groupi_n_8212, csa_tree_add_190_195_groupi_n_8213, csa_tree_add_190_195_groupi_n_8214, csa_tree_add_190_195_groupi_n_8215;
  wire csa_tree_add_190_195_groupi_n_8216, csa_tree_add_190_195_groupi_n_8217, csa_tree_add_190_195_groupi_n_8218, csa_tree_add_190_195_groupi_n_8219, csa_tree_add_190_195_groupi_n_8220, csa_tree_add_190_195_groupi_n_8221, csa_tree_add_190_195_groupi_n_8222, csa_tree_add_190_195_groupi_n_8223;
  wire csa_tree_add_190_195_groupi_n_8224, csa_tree_add_190_195_groupi_n_8225, csa_tree_add_190_195_groupi_n_8226, csa_tree_add_190_195_groupi_n_8227, csa_tree_add_190_195_groupi_n_8228, csa_tree_add_190_195_groupi_n_8229, csa_tree_add_190_195_groupi_n_8230, csa_tree_add_190_195_groupi_n_8231;
  wire csa_tree_add_190_195_groupi_n_8232, csa_tree_add_190_195_groupi_n_8233, csa_tree_add_190_195_groupi_n_8234, csa_tree_add_190_195_groupi_n_8235, csa_tree_add_190_195_groupi_n_8236, csa_tree_add_190_195_groupi_n_8237, csa_tree_add_190_195_groupi_n_8238, csa_tree_add_190_195_groupi_n_8239;
  wire csa_tree_add_190_195_groupi_n_8240, csa_tree_add_190_195_groupi_n_8241, csa_tree_add_190_195_groupi_n_8242, csa_tree_add_190_195_groupi_n_8243, csa_tree_add_190_195_groupi_n_8244, csa_tree_add_190_195_groupi_n_8245, csa_tree_add_190_195_groupi_n_8246, csa_tree_add_190_195_groupi_n_8247;
  wire csa_tree_add_190_195_groupi_n_8248, csa_tree_add_190_195_groupi_n_8249, csa_tree_add_190_195_groupi_n_8250, csa_tree_add_190_195_groupi_n_8251, csa_tree_add_190_195_groupi_n_8252, csa_tree_add_190_195_groupi_n_8253, csa_tree_add_190_195_groupi_n_8254, csa_tree_add_190_195_groupi_n_8255;
  wire csa_tree_add_190_195_groupi_n_8256, csa_tree_add_190_195_groupi_n_8257, csa_tree_add_190_195_groupi_n_8258, csa_tree_add_190_195_groupi_n_8259, csa_tree_add_190_195_groupi_n_8260, csa_tree_add_190_195_groupi_n_8261, csa_tree_add_190_195_groupi_n_8262, csa_tree_add_190_195_groupi_n_8263;
  wire csa_tree_add_190_195_groupi_n_8264, csa_tree_add_190_195_groupi_n_8265, csa_tree_add_190_195_groupi_n_8266, csa_tree_add_190_195_groupi_n_8267, csa_tree_add_190_195_groupi_n_8268, csa_tree_add_190_195_groupi_n_8269, csa_tree_add_190_195_groupi_n_8270, csa_tree_add_190_195_groupi_n_8271;
  wire csa_tree_add_190_195_groupi_n_8272, csa_tree_add_190_195_groupi_n_8273, csa_tree_add_190_195_groupi_n_8274, csa_tree_add_190_195_groupi_n_8275, csa_tree_add_190_195_groupi_n_8276, csa_tree_add_190_195_groupi_n_8277, csa_tree_add_190_195_groupi_n_8278, csa_tree_add_190_195_groupi_n_8279;
  wire csa_tree_add_190_195_groupi_n_8280, csa_tree_add_190_195_groupi_n_8281, csa_tree_add_190_195_groupi_n_8282, csa_tree_add_190_195_groupi_n_8283, csa_tree_add_190_195_groupi_n_8284, csa_tree_add_190_195_groupi_n_8285, csa_tree_add_190_195_groupi_n_8286, csa_tree_add_190_195_groupi_n_8287;
  wire csa_tree_add_190_195_groupi_n_8288, csa_tree_add_190_195_groupi_n_8289, csa_tree_add_190_195_groupi_n_8290, csa_tree_add_190_195_groupi_n_8291, csa_tree_add_190_195_groupi_n_8292, csa_tree_add_190_195_groupi_n_8293, csa_tree_add_190_195_groupi_n_8294, csa_tree_add_190_195_groupi_n_8295;
  wire csa_tree_add_190_195_groupi_n_8296, csa_tree_add_190_195_groupi_n_8297, csa_tree_add_190_195_groupi_n_8298, csa_tree_add_190_195_groupi_n_8299, csa_tree_add_190_195_groupi_n_8300, csa_tree_add_190_195_groupi_n_8301, csa_tree_add_190_195_groupi_n_8302, csa_tree_add_190_195_groupi_n_8303;
  wire csa_tree_add_190_195_groupi_n_8304, csa_tree_add_190_195_groupi_n_8305, csa_tree_add_190_195_groupi_n_8306, csa_tree_add_190_195_groupi_n_8307, csa_tree_add_190_195_groupi_n_8308, csa_tree_add_190_195_groupi_n_8309, csa_tree_add_190_195_groupi_n_8310, csa_tree_add_190_195_groupi_n_8311;
  wire csa_tree_add_190_195_groupi_n_8312, csa_tree_add_190_195_groupi_n_8313, csa_tree_add_190_195_groupi_n_8314, csa_tree_add_190_195_groupi_n_8315, csa_tree_add_190_195_groupi_n_8316, csa_tree_add_190_195_groupi_n_8317, csa_tree_add_190_195_groupi_n_8318, csa_tree_add_190_195_groupi_n_8319;
  wire csa_tree_add_190_195_groupi_n_8320, csa_tree_add_190_195_groupi_n_8321, csa_tree_add_190_195_groupi_n_8322, csa_tree_add_190_195_groupi_n_8323, csa_tree_add_190_195_groupi_n_8324, csa_tree_add_190_195_groupi_n_8325, csa_tree_add_190_195_groupi_n_8326, csa_tree_add_190_195_groupi_n_8327;
  wire csa_tree_add_190_195_groupi_n_8328, csa_tree_add_190_195_groupi_n_8329, csa_tree_add_190_195_groupi_n_8330, csa_tree_add_190_195_groupi_n_8331, csa_tree_add_190_195_groupi_n_8332, csa_tree_add_190_195_groupi_n_8333, csa_tree_add_190_195_groupi_n_8334, csa_tree_add_190_195_groupi_n_8335;
  wire csa_tree_add_190_195_groupi_n_8336, csa_tree_add_190_195_groupi_n_8337, csa_tree_add_190_195_groupi_n_8338, csa_tree_add_190_195_groupi_n_8339, csa_tree_add_190_195_groupi_n_8340, csa_tree_add_190_195_groupi_n_8341, csa_tree_add_190_195_groupi_n_8342, csa_tree_add_190_195_groupi_n_8343;
  wire csa_tree_add_190_195_groupi_n_8344, csa_tree_add_190_195_groupi_n_8345, csa_tree_add_190_195_groupi_n_8346, csa_tree_add_190_195_groupi_n_8347, csa_tree_add_190_195_groupi_n_8348, csa_tree_add_190_195_groupi_n_8349, csa_tree_add_190_195_groupi_n_8350, csa_tree_add_190_195_groupi_n_8351;
  wire csa_tree_add_190_195_groupi_n_8352, csa_tree_add_190_195_groupi_n_8353, csa_tree_add_190_195_groupi_n_8354, csa_tree_add_190_195_groupi_n_8355, csa_tree_add_190_195_groupi_n_8356, csa_tree_add_190_195_groupi_n_8357, csa_tree_add_190_195_groupi_n_8358, csa_tree_add_190_195_groupi_n_8359;
  wire csa_tree_add_190_195_groupi_n_8360, csa_tree_add_190_195_groupi_n_8361, csa_tree_add_190_195_groupi_n_8362, csa_tree_add_190_195_groupi_n_8363, csa_tree_add_190_195_groupi_n_8364, csa_tree_add_190_195_groupi_n_8365, csa_tree_add_190_195_groupi_n_8366, csa_tree_add_190_195_groupi_n_8367;
  wire csa_tree_add_190_195_groupi_n_8368, csa_tree_add_190_195_groupi_n_8369, csa_tree_add_190_195_groupi_n_8370, csa_tree_add_190_195_groupi_n_8371, csa_tree_add_190_195_groupi_n_8372, csa_tree_add_190_195_groupi_n_8373, csa_tree_add_190_195_groupi_n_8374, csa_tree_add_190_195_groupi_n_8375;
  wire csa_tree_add_190_195_groupi_n_8376, csa_tree_add_190_195_groupi_n_8377, csa_tree_add_190_195_groupi_n_8378, csa_tree_add_190_195_groupi_n_8379, csa_tree_add_190_195_groupi_n_8380, csa_tree_add_190_195_groupi_n_8381, csa_tree_add_190_195_groupi_n_8382, csa_tree_add_190_195_groupi_n_8383;
  wire csa_tree_add_190_195_groupi_n_8384, csa_tree_add_190_195_groupi_n_8385, csa_tree_add_190_195_groupi_n_8386, csa_tree_add_190_195_groupi_n_8387, csa_tree_add_190_195_groupi_n_8388, csa_tree_add_190_195_groupi_n_8389, csa_tree_add_190_195_groupi_n_8390, csa_tree_add_190_195_groupi_n_8391;
  wire csa_tree_add_190_195_groupi_n_8392, csa_tree_add_190_195_groupi_n_8393, csa_tree_add_190_195_groupi_n_8394, csa_tree_add_190_195_groupi_n_8395, csa_tree_add_190_195_groupi_n_8396, csa_tree_add_190_195_groupi_n_8397, csa_tree_add_190_195_groupi_n_8398, csa_tree_add_190_195_groupi_n_8399;
  wire csa_tree_add_190_195_groupi_n_8400, csa_tree_add_190_195_groupi_n_8401, csa_tree_add_190_195_groupi_n_8402, csa_tree_add_190_195_groupi_n_8403, csa_tree_add_190_195_groupi_n_8404, csa_tree_add_190_195_groupi_n_8405, csa_tree_add_190_195_groupi_n_8406, csa_tree_add_190_195_groupi_n_8407;
  wire csa_tree_add_190_195_groupi_n_8408, csa_tree_add_190_195_groupi_n_8409, csa_tree_add_190_195_groupi_n_8410, csa_tree_add_190_195_groupi_n_8411, csa_tree_add_190_195_groupi_n_8412, csa_tree_add_190_195_groupi_n_8413, csa_tree_add_190_195_groupi_n_8414, csa_tree_add_190_195_groupi_n_8415;
  wire csa_tree_add_190_195_groupi_n_8416, csa_tree_add_190_195_groupi_n_8417, csa_tree_add_190_195_groupi_n_8418, csa_tree_add_190_195_groupi_n_8419, csa_tree_add_190_195_groupi_n_8420, csa_tree_add_190_195_groupi_n_8421, csa_tree_add_190_195_groupi_n_8422, csa_tree_add_190_195_groupi_n_8423;
  wire csa_tree_add_190_195_groupi_n_8424, csa_tree_add_190_195_groupi_n_8425, csa_tree_add_190_195_groupi_n_8426, csa_tree_add_190_195_groupi_n_8427, csa_tree_add_190_195_groupi_n_8428, csa_tree_add_190_195_groupi_n_8429, csa_tree_add_190_195_groupi_n_8430, csa_tree_add_190_195_groupi_n_8431;
  wire csa_tree_add_190_195_groupi_n_8432, csa_tree_add_190_195_groupi_n_8433, csa_tree_add_190_195_groupi_n_8434, csa_tree_add_190_195_groupi_n_8435, csa_tree_add_190_195_groupi_n_8436, csa_tree_add_190_195_groupi_n_8437, csa_tree_add_190_195_groupi_n_8438, csa_tree_add_190_195_groupi_n_8439;
  wire csa_tree_add_190_195_groupi_n_8440, csa_tree_add_190_195_groupi_n_8441, csa_tree_add_190_195_groupi_n_8442, csa_tree_add_190_195_groupi_n_8443, csa_tree_add_190_195_groupi_n_8444, csa_tree_add_190_195_groupi_n_8445, csa_tree_add_190_195_groupi_n_8446, csa_tree_add_190_195_groupi_n_8447;
  wire csa_tree_add_190_195_groupi_n_8448, csa_tree_add_190_195_groupi_n_8449, csa_tree_add_190_195_groupi_n_8450, csa_tree_add_190_195_groupi_n_8451, csa_tree_add_190_195_groupi_n_8452, csa_tree_add_190_195_groupi_n_8453, csa_tree_add_190_195_groupi_n_8454, csa_tree_add_190_195_groupi_n_8455;
  wire csa_tree_add_190_195_groupi_n_8456, csa_tree_add_190_195_groupi_n_8457, csa_tree_add_190_195_groupi_n_8458, csa_tree_add_190_195_groupi_n_8459, csa_tree_add_190_195_groupi_n_8460, csa_tree_add_190_195_groupi_n_8461, csa_tree_add_190_195_groupi_n_8462, csa_tree_add_190_195_groupi_n_8463;
  wire csa_tree_add_190_195_groupi_n_8464, csa_tree_add_190_195_groupi_n_8465, csa_tree_add_190_195_groupi_n_8466, csa_tree_add_190_195_groupi_n_8467, csa_tree_add_190_195_groupi_n_8468, csa_tree_add_190_195_groupi_n_8469, csa_tree_add_190_195_groupi_n_8470, csa_tree_add_190_195_groupi_n_8471;
  wire csa_tree_add_190_195_groupi_n_8472, csa_tree_add_190_195_groupi_n_8473, csa_tree_add_190_195_groupi_n_8474, csa_tree_add_190_195_groupi_n_8475, csa_tree_add_190_195_groupi_n_8476, csa_tree_add_190_195_groupi_n_8477, csa_tree_add_190_195_groupi_n_8478, csa_tree_add_190_195_groupi_n_8479;
  wire csa_tree_add_190_195_groupi_n_8480, csa_tree_add_190_195_groupi_n_8481, csa_tree_add_190_195_groupi_n_8482, csa_tree_add_190_195_groupi_n_8483, csa_tree_add_190_195_groupi_n_8484, csa_tree_add_190_195_groupi_n_8485, csa_tree_add_190_195_groupi_n_8486, csa_tree_add_190_195_groupi_n_8487;
  wire csa_tree_add_190_195_groupi_n_8488, csa_tree_add_190_195_groupi_n_8489, csa_tree_add_190_195_groupi_n_8490, csa_tree_add_190_195_groupi_n_8491, csa_tree_add_190_195_groupi_n_8492, csa_tree_add_190_195_groupi_n_8493, csa_tree_add_190_195_groupi_n_8494, csa_tree_add_190_195_groupi_n_8495;
  wire csa_tree_add_190_195_groupi_n_8496, csa_tree_add_190_195_groupi_n_8497, csa_tree_add_190_195_groupi_n_8498, csa_tree_add_190_195_groupi_n_8499, csa_tree_add_190_195_groupi_n_8500, csa_tree_add_190_195_groupi_n_8501, csa_tree_add_190_195_groupi_n_8502, csa_tree_add_190_195_groupi_n_8503;
  wire csa_tree_add_190_195_groupi_n_8504, csa_tree_add_190_195_groupi_n_8505, csa_tree_add_190_195_groupi_n_8506, csa_tree_add_190_195_groupi_n_8507, csa_tree_add_190_195_groupi_n_8508, csa_tree_add_190_195_groupi_n_8509, csa_tree_add_190_195_groupi_n_8510, csa_tree_add_190_195_groupi_n_8511;
  wire csa_tree_add_190_195_groupi_n_8512, csa_tree_add_190_195_groupi_n_8513, csa_tree_add_190_195_groupi_n_8514, csa_tree_add_190_195_groupi_n_8515, csa_tree_add_190_195_groupi_n_8516, csa_tree_add_190_195_groupi_n_8517, csa_tree_add_190_195_groupi_n_8518, csa_tree_add_190_195_groupi_n_8519;
  wire csa_tree_add_190_195_groupi_n_8520, csa_tree_add_190_195_groupi_n_8521, csa_tree_add_190_195_groupi_n_8522, csa_tree_add_190_195_groupi_n_8523, csa_tree_add_190_195_groupi_n_8524, csa_tree_add_190_195_groupi_n_8525, csa_tree_add_190_195_groupi_n_8526, csa_tree_add_190_195_groupi_n_8527;
  wire csa_tree_add_190_195_groupi_n_8528, csa_tree_add_190_195_groupi_n_8529, csa_tree_add_190_195_groupi_n_8530, csa_tree_add_190_195_groupi_n_8531, csa_tree_add_190_195_groupi_n_8532, csa_tree_add_190_195_groupi_n_8533, csa_tree_add_190_195_groupi_n_8534, csa_tree_add_190_195_groupi_n_8535;
  wire csa_tree_add_190_195_groupi_n_8536, csa_tree_add_190_195_groupi_n_8537, csa_tree_add_190_195_groupi_n_8538, csa_tree_add_190_195_groupi_n_8539, csa_tree_add_190_195_groupi_n_8540, csa_tree_add_190_195_groupi_n_8541, csa_tree_add_190_195_groupi_n_8542, csa_tree_add_190_195_groupi_n_8543;
  wire csa_tree_add_190_195_groupi_n_8544, csa_tree_add_190_195_groupi_n_8545, csa_tree_add_190_195_groupi_n_8546, csa_tree_add_190_195_groupi_n_8547, csa_tree_add_190_195_groupi_n_8548, csa_tree_add_190_195_groupi_n_8549, csa_tree_add_190_195_groupi_n_8550, csa_tree_add_190_195_groupi_n_8551;
  wire csa_tree_add_190_195_groupi_n_8552, csa_tree_add_190_195_groupi_n_8553, csa_tree_add_190_195_groupi_n_8554, csa_tree_add_190_195_groupi_n_8555, csa_tree_add_190_195_groupi_n_8556, csa_tree_add_190_195_groupi_n_8557, csa_tree_add_190_195_groupi_n_8558, csa_tree_add_190_195_groupi_n_8559;
  wire csa_tree_add_190_195_groupi_n_8560, csa_tree_add_190_195_groupi_n_8561, csa_tree_add_190_195_groupi_n_8562, csa_tree_add_190_195_groupi_n_8563, csa_tree_add_190_195_groupi_n_8564, csa_tree_add_190_195_groupi_n_8565, csa_tree_add_190_195_groupi_n_8566, csa_tree_add_190_195_groupi_n_8567;
  wire csa_tree_add_190_195_groupi_n_8568, csa_tree_add_190_195_groupi_n_8569, csa_tree_add_190_195_groupi_n_8570, csa_tree_add_190_195_groupi_n_8571, csa_tree_add_190_195_groupi_n_8572, csa_tree_add_190_195_groupi_n_8573, csa_tree_add_190_195_groupi_n_8574, csa_tree_add_190_195_groupi_n_8575;
  wire csa_tree_add_190_195_groupi_n_8576, csa_tree_add_190_195_groupi_n_8577, csa_tree_add_190_195_groupi_n_8578, csa_tree_add_190_195_groupi_n_8579, csa_tree_add_190_195_groupi_n_8580, csa_tree_add_190_195_groupi_n_8581, csa_tree_add_190_195_groupi_n_8582, csa_tree_add_190_195_groupi_n_8583;
  wire csa_tree_add_190_195_groupi_n_8584, csa_tree_add_190_195_groupi_n_8585, csa_tree_add_190_195_groupi_n_8586, csa_tree_add_190_195_groupi_n_8587, csa_tree_add_190_195_groupi_n_8588, csa_tree_add_190_195_groupi_n_8589, csa_tree_add_190_195_groupi_n_8590, csa_tree_add_190_195_groupi_n_8591;
  wire csa_tree_add_190_195_groupi_n_8592, csa_tree_add_190_195_groupi_n_8593, csa_tree_add_190_195_groupi_n_8594, csa_tree_add_190_195_groupi_n_8595, csa_tree_add_190_195_groupi_n_8596, csa_tree_add_190_195_groupi_n_8597, csa_tree_add_190_195_groupi_n_8598, csa_tree_add_190_195_groupi_n_8599;
  wire csa_tree_add_190_195_groupi_n_8600, csa_tree_add_190_195_groupi_n_8601, csa_tree_add_190_195_groupi_n_8602, csa_tree_add_190_195_groupi_n_8603, csa_tree_add_190_195_groupi_n_8604, csa_tree_add_190_195_groupi_n_8605, csa_tree_add_190_195_groupi_n_8606, csa_tree_add_190_195_groupi_n_8607;
  wire csa_tree_add_190_195_groupi_n_8608, csa_tree_add_190_195_groupi_n_8609, csa_tree_add_190_195_groupi_n_8610, csa_tree_add_190_195_groupi_n_8611, csa_tree_add_190_195_groupi_n_8612, csa_tree_add_190_195_groupi_n_8613, csa_tree_add_190_195_groupi_n_8614, csa_tree_add_190_195_groupi_n_8615;
  wire csa_tree_add_190_195_groupi_n_8616, csa_tree_add_190_195_groupi_n_8617, csa_tree_add_190_195_groupi_n_8618, csa_tree_add_190_195_groupi_n_8619, csa_tree_add_190_195_groupi_n_8620, csa_tree_add_190_195_groupi_n_8621, csa_tree_add_190_195_groupi_n_8622, csa_tree_add_190_195_groupi_n_8623;
  wire csa_tree_add_190_195_groupi_n_8624, csa_tree_add_190_195_groupi_n_8625, csa_tree_add_190_195_groupi_n_8626, csa_tree_add_190_195_groupi_n_8627, csa_tree_add_190_195_groupi_n_8628, csa_tree_add_190_195_groupi_n_8629, csa_tree_add_190_195_groupi_n_8630, csa_tree_add_190_195_groupi_n_8631;
  wire csa_tree_add_190_195_groupi_n_8632, csa_tree_add_190_195_groupi_n_8633, csa_tree_add_190_195_groupi_n_8634, csa_tree_add_190_195_groupi_n_8635, csa_tree_add_190_195_groupi_n_8636, csa_tree_add_190_195_groupi_n_8637, csa_tree_add_190_195_groupi_n_8638, csa_tree_add_190_195_groupi_n_8639;
  wire csa_tree_add_190_195_groupi_n_8640, csa_tree_add_190_195_groupi_n_8641, csa_tree_add_190_195_groupi_n_8642, csa_tree_add_190_195_groupi_n_8643, csa_tree_add_190_195_groupi_n_8644, csa_tree_add_190_195_groupi_n_8645, csa_tree_add_190_195_groupi_n_8646, csa_tree_add_190_195_groupi_n_8647;
  wire csa_tree_add_190_195_groupi_n_8648, csa_tree_add_190_195_groupi_n_8649, csa_tree_add_190_195_groupi_n_8650, csa_tree_add_190_195_groupi_n_8651, csa_tree_add_190_195_groupi_n_8652, csa_tree_add_190_195_groupi_n_8653, csa_tree_add_190_195_groupi_n_8654, csa_tree_add_190_195_groupi_n_8655;
  wire csa_tree_add_190_195_groupi_n_8656, csa_tree_add_190_195_groupi_n_8657, csa_tree_add_190_195_groupi_n_8658, csa_tree_add_190_195_groupi_n_8659, csa_tree_add_190_195_groupi_n_8660, csa_tree_add_190_195_groupi_n_8661, csa_tree_add_190_195_groupi_n_8662, csa_tree_add_190_195_groupi_n_8663;
  wire csa_tree_add_190_195_groupi_n_8664, csa_tree_add_190_195_groupi_n_8665, csa_tree_add_190_195_groupi_n_8666, csa_tree_add_190_195_groupi_n_8667, csa_tree_add_190_195_groupi_n_8668, csa_tree_add_190_195_groupi_n_8669, csa_tree_add_190_195_groupi_n_8670, csa_tree_add_190_195_groupi_n_8671;
  wire csa_tree_add_190_195_groupi_n_8672, csa_tree_add_190_195_groupi_n_8673, csa_tree_add_190_195_groupi_n_8674, csa_tree_add_190_195_groupi_n_8675, csa_tree_add_190_195_groupi_n_8676, csa_tree_add_190_195_groupi_n_8677, csa_tree_add_190_195_groupi_n_8678, csa_tree_add_190_195_groupi_n_8679;
  wire csa_tree_add_190_195_groupi_n_8680, csa_tree_add_190_195_groupi_n_8681, csa_tree_add_190_195_groupi_n_8682, csa_tree_add_190_195_groupi_n_8683, csa_tree_add_190_195_groupi_n_8684, csa_tree_add_190_195_groupi_n_8685, csa_tree_add_190_195_groupi_n_8686, csa_tree_add_190_195_groupi_n_8687;
  wire csa_tree_add_190_195_groupi_n_8688, csa_tree_add_190_195_groupi_n_8689, csa_tree_add_190_195_groupi_n_8690, csa_tree_add_190_195_groupi_n_8691, csa_tree_add_190_195_groupi_n_8692, csa_tree_add_190_195_groupi_n_8693, csa_tree_add_190_195_groupi_n_8694, csa_tree_add_190_195_groupi_n_8695;
  wire csa_tree_add_190_195_groupi_n_8696, csa_tree_add_190_195_groupi_n_8697, csa_tree_add_190_195_groupi_n_8698, csa_tree_add_190_195_groupi_n_8699, csa_tree_add_190_195_groupi_n_8700, csa_tree_add_190_195_groupi_n_8701, csa_tree_add_190_195_groupi_n_8702, csa_tree_add_190_195_groupi_n_8703;
  wire csa_tree_add_190_195_groupi_n_8704, csa_tree_add_190_195_groupi_n_8705, csa_tree_add_190_195_groupi_n_8706, csa_tree_add_190_195_groupi_n_8707, csa_tree_add_190_195_groupi_n_8708, csa_tree_add_190_195_groupi_n_8709, csa_tree_add_190_195_groupi_n_8710, csa_tree_add_190_195_groupi_n_8711;
  wire csa_tree_add_190_195_groupi_n_8712, csa_tree_add_190_195_groupi_n_8713, csa_tree_add_190_195_groupi_n_8714, csa_tree_add_190_195_groupi_n_8715, csa_tree_add_190_195_groupi_n_8716, csa_tree_add_190_195_groupi_n_8717, csa_tree_add_190_195_groupi_n_8718, csa_tree_add_190_195_groupi_n_8719;
  wire csa_tree_add_190_195_groupi_n_8720, csa_tree_add_190_195_groupi_n_8721, csa_tree_add_190_195_groupi_n_8722, csa_tree_add_190_195_groupi_n_8723, csa_tree_add_190_195_groupi_n_8724, csa_tree_add_190_195_groupi_n_8725, csa_tree_add_190_195_groupi_n_8726, csa_tree_add_190_195_groupi_n_8727;
  wire csa_tree_add_190_195_groupi_n_8728, csa_tree_add_190_195_groupi_n_8729, csa_tree_add_190_195_groupi_n_8730, csa_tree_add_190_195_groupi_n_8731, csa_tree_add_190_195_groupi_n_8732, csa_tree_add_190_195_groupi_n_8733, csa_tree_add_190_195_groupi_n_8734, csa_tree_add_190_195_groupi_n_8735;
  wire csa_tree_add_190_195_groupi_n_8736, csa_tree_add_190_195_groupi_n_8737, csa_tree_add_190_195_groupi_n_8738, csa_tree_add_190_195_groupi_n_8739, csa_tree_add_190_195_groupi_n_8740, csa_tree_add_190_195_groupi_n_8741, csa_tree_add_190_195_groupi_n_8742, csa_tree_add_190_195_groupi_n_8743;
  wire csa_tree_add_190_195_groupi_n_8744, csa_tree_add_190_195_groupi_n_8745, csa_tree_add_190_195_groupi_n_8746, csa_tree_add_190_195_groupi_n_8747, csa_tree_add_190_195_groupi_n_8748, csa_tree_add_190_195_groupi_n_8749, csa_tree_add_190_195_groupi_n_8750, csa_tree_add_190_195_groupi_n_8751;
  wire csa_tree_add_190_195_groupi_n_8752, csa_tree_add_190_195_groupi_n_8753, csa_tree_add_190_195_groupi_n_8754, csa_tree_add_190_195_groupi_n_8755, csa_tree_add_190_195_groupi_n_8756, csa_tree_add_190_195_groupi_n_8757, csa_tree_add_190_195_groupi_n_8758, csa_tree_add_190_195_groupi_n_8759;
  wire csa_tree_add_190_195_groupi_n_8760, csa_tree_add_190_195_groupi_n_8761, csa_tree_add_190_195_groupi_n_8762, csa_tree_add_190_195_groupi_n_8763, csa_tree_add_190_195_groupi_n_8764, csa_tree_add_190_195_groupi_n_8765, csa_tree_add_190_195_groupi_n_8766, csa_tree_add_190_195_groupi_n_8767;
  wire csa_tree_add_190_195_groupi_n_8768, csa_tree_add_190_195_groupi_n_8769, csa_tree_add_190_195_groupi_n_8770, csa_tree_add_190_195_groupi_n_8771, csa_tree_add_190_195_groupi_n_8772, csa_tree_add_190_195_groupi_n_8773, csa_tree_add_190_195_groupi_n_8774, csa_tree_add_190_195_groupi_n_8775;
  wire csa_tree_add_190_195_groupi_n_8776, csa_tree_add_190_195_groupi_n_8777, csa_tree_add_190_195_groupi_n_8778, csa_tree_add_190_195_groupi_n_8779, csa_tree_add_190_195_groupi_n_8780, csa_tree_add_190_195_groupi_n_8781, csa_tree_add_190_195_groupi_n_8782, csa_tree_add_190_195_groupi_n_8783;
  wire csa_tree_add_190_195_groupi_n_8784, csa_tree_add_190_195_groupi_n_8785, csa_tree_add_190_195_groupi_n_8786, csa_tree_add_190_195_groupi_n_8787, csa_tree_add_190_195_groupi_n_8788, csa_tree_add_190_195_groupi_n_8789, csa_tree_add_190_195_groupi_n_8790, csa_tree_add_190_195_groupi_n_8791;
  wire csa_tree_add_190_195_groupi_n_8792, csa_tree_add_190_195_groupi_n_8793, csa_tree_add_190_195_groupi_n_8794, csa_tree_add_190_195_groupi_n_8795, csa_tree_add_190_195_groupi_n_8796, csa_tree_add_190_195_groupi_n_8797, csa_tree_add_190_195_groupi_n_8798, csa_tree_add_190_195_groupi_n_8799;
  wire csa_tree_add_190_195_groupi_n_8800, csa_tree_add_190_195_groupi_n_8801, csa_tree_add_190_195_groupi_n_8802, csa_tree_add_190_195_groupi_n_8803, csa_tree_add_190_195_groupi_n_8804, csa_tree_add_190_195_groupi_n_8805, csa_tree_add_190_195_groupi_n_8806, csa_tree_add_190_195_groupi_n_8807;
  wire csa_tree_add_190_195_groupi_n_8808, csa_tree_add_190_195_groupi_n_8809, csa_tree_add_190_195_groupi_n_8810, csa_tree_add_190_195_groupi_n_8811, csa_tree_add_190_195_groupi_n_8812, csa_tree_add_190_195_groupi_n_8813, csa_tree_add_190_195_groupi_n_8814, csa_tree_add_190_195_groupi_n_8815;
  wire csa_tree_add_190_195_groupi_n_8816, csa_tree_add_190_195_groupi_n_8817, csa_tree_add_190_195_groupi_n_8818, csa_tree_add_190_195_groupi_n_8819, csa_tree_add_190_195_groupi_n_8820, csa_tree_add_190_195_groupi_n_8821, csa_tree_add_190_195_groupi_n_8822, csa_tree_add_190_195_groupi_n_8823;
  wire csa_tree_add_190_195_groupi_n_8824, csa_tree_add_190_195_groupi_n_8825, csa_tree_add_190_195_groupi_n_8826, csa_tree_add_190_195_groupi_n_8827, csa_tree_add_190_195_groupi_n_8828, csa_tree_add_190_195_groupi_n_8829, csa_tree_add_190_195_groupi_n_8830, csa_tree_add_190_195_groupi_n_8831;
  wire csa_tree_add_190_195_groupi_n_8832, csa_tree_add_190_195_groupi_n_8833, csa_tree_add_190_195_groupi_n_8834, csa_tree_add_190_195_groupi_n_8835, csa_tree_add_190_195_groupi_n_8836, csa_tree_add_190_195_groupi_n_8837, csa_tree_add_190_195_groupi_n_8838, csa_tree_add_190_195_groupi_n_8839;
  wire csa_tree_add_190_195_groupi_n_8840, csa_tree_add_190_195_groupi_n_8841, csa_tree_add_190_195_groupi_n_8842, csa_tree_add_190_195_groupi_n_8843, csa_tree_add_190_195_groupi_n_8844, csa_tree_add_190_195_groupi_n_8845, csa_tree_add_190_195_groupi_n_8846, csa_tree_add_190_195_groupi_n_8847;
  wire csa_tree_add_190_195_groupi_n_8848, csa_tree_add_190_195_groupi_n_8849, csa_tree_add_190_195_groupi_n_8850, csa_tree_add_190_195_groupi_n_8851, csa_tree_add_190_195_groupi_n_8852, csa_tree_add_190_195_groupi_n_8853, csa_tree_add_190_195_groupi_n_8854, csa_tree_add_190_195_groupi_n_8855;
  wire csa_tree_add_190_195_groupi_n_8856, csa_tree_add_190_195_groupi_n_8857, csa_tree_add_190_195_groupi_n_8858, csa_tree_add_190_195_groupi_n_8859, csa_tree_add_190_195_groupi_n_8860, csa_tree_add_190_195_groupi_n_8861, csa_tree_add_190_195_groupi_n_8862, csa_tree_add_190_195_groupi_n_8863;
  wire csa_tree_add_190_195_groupi_n_8864, csa_tree_add_190_195_groupi_n_8865, csa_tree_add_190_195_groupi_n_8866, csa_tree_add_190_195_groupi_n_8867, csa_tree_add_190_195_groupi_n_8868, csa_tree_add_190_195_groupi_n_8869, csa_tree_add_190_195_groupi_n_8870, csa_tree_add_190_195_groupi_n_8871;
  wire csa_tree_add_190_195_groupi_n_8872, csa_tree_add_190_195_groupi_n_8873, csa_tree_add_190_195_groupi_n_8874, csa_tree_add_190_195_groupi_n_8875, csa_tree_add_190_195_groupi_n_8876, csa_tree_add_190_195_groupi_n_8877, csa_tree_add_190_195_groupi_n_8878, csa_tree_add_190_195_groupi_n_8879;
  wire csa_tree_add_190_195_groupi_n_8880, csa_tree_add_190_195_groupi_n_8881, csa_tree_add_190_195_groupi_n_8882, csa_tree_add_190_195_groupi_n_8883, csa_tree_add_190_195_groupi_n_8884, csa_tree_add_190_195_groupi_n_8885, csa_tree_add_190_195_groupi_n_8886, csa_tree_add_190_195_groupi_n_8887;
  wire csa_tree_add_190_195_groupi_n_8888, csa_tree_add_190_195_groupi_n_8889, csa_tree_add_190_195_groupi_n_8890, csa_tree_add_190_195_groupi_n_8891, csa_tree_add_190_195_groupi_n_8892, csa_tree_add_190_195_groupi_n_8893, csa_tree_add_190_195_groupi_n_8894, csa_tree_add_190_195_groupi_n_8895;
  wire csa_tree_add_190_195_groupi_n_8896, csa_tree_add_190_195_groupi_n_8897, csa_tree_add_190_195_groupi_n_8898, csa_tree_add_190_195_groupi_n_8899, csa_tree_add_190_195_groupi_n_8900, csa_tree_add_190_195_groupi_n_8901, csa_tree_add_190_195_groupi_n_8902, csa_tree_add_190_195_groupi_n_8903;
  wire csa_tree_add_190_195_groupi_n_8904, csa_tree_add_190_195_groupi_n_8905, csa_tree_add_190_195_groupi_n_8906, csa_tree_add_190_195_groupi_n_8907, csa_tree_add_190_195_groupi_n_8908, csa_tree_add_190_195_groupi_n_8909, csa_tree_add_190_195_groupi_n_8910, csa_tree_add_190_195_groupi_n_8911;
  wire csa_tree_add_190_195_groupi_n_8912, csa_tree_add_190_195_groupi_n_8913, csa_tree_add_190_195_groupi_n_8914, csa_tree_add_190_195_groupi_n_8915, csa_tree_add_190_195_groupi_n_8916, csa_tree_add_190_195_groupi_n_8917, csa_tree_add_190_195_groupi_n_8918, csa_tree_add_190_195_groupi_n_8919;
  wire csa_tree_add_190_195_groupi_n_8920, csa_tree_add_190_195_groupi_n_8921, csa_tree_add_190_195_groupi_n_8922, csa_tree_add_190_195_groupi_n_8923, csa_tree_add_190_195_groupi_n_8924, csa_tree_add_190_195_groupi_n_8925, csa_tree_add_190_195_groupi_n_8926, csa_tree_add_190_195_groupi_n_8927;
  wire csa_tree_add_190_195_groupi_n_8928, csa_tree_add_190_195_groupi_n_8929, csa_tree_add_190_195_groupi_n_8930, csa_tree_add_190_195_groupi_n_8931, csa_tree_add_190_195_groupi_n_8932, csa_tree_add_190_195_groupi_n_8933, csa_tree_add_190_195_groupi_n_8934, csa_tree_add_190_195_groupi_n_8935;
  wire csa_tree_add_190_195_groupi_n_8936, csa_tree_add_190_195_groupi_n_8937, csa_tree_add_190_195_groupi_n_8938, csa_tree_add_190_195_groupi_n_8940, csa_tree_add_190_195_groupi_n_8941, csa_tree_add_190_195_groupi_n_8942, csa_tree_add_190_195_groupi_n_8943, csa_tree_add_190_195_groupi_n_8944;
  wire csa_tree_add_190_195_groupi_n_8945, csa_tree_add_190_195_groupi_n_8946, csa_tree_add_190_195_groupi_n_8947, csa_tree_add_190_195_groupi_n_8948, csa_tree_add_190_195_groupi_n_8949, csa_tree_add_190_195_groupi_n_8950, csa_tree_add_190_195_groupi_n_8951, csa_tree_add_190_195_groupi_n_8952;
  wire csa_tree_add_190_195_groupi_n_8953, csa_tree_add_190_195_groupi_n_8954, csa_tree_add_190_195_groupi_n_8955, csa_tree_add_190_195_groupi_n_8956, csa_tree_add_190_195_groupi_n_8957, csa_tree_add_190_195_groupi_n_8958, csa_tree_add_190_195_groupi_n_8959, csa_tree_add_190_195_groupi_n_8960;
  wire csa_tree_add_190_195_groupi_n_8961, csa_tree_add_190_195_groupi_n_8962, csa_tree_add_190_195_groupi_n_8963, csa_tree_add_190_195_groupi_n_8964, csa_tree_add_190_195_groupi_n_8965, csa_tree_add_190_195_groupi_n_8966, csa_tree_add_190_195_groupi_n_8967, csa_tree_add_190_195_groupi_n_8968;
  wire csa_tree_add_190_195_groupi_n_8969, csa_tree_add_190_195_groupi_n_8970, csa_tree_add_190_195_groupi_n_8971, csa_tree_add_190_195_groupi_n_8972, csa_tree_add_190_195_groupi_n_8973, csa_tree_add_190_195_groupi_n_8974, csa_tree_add_190_195_groupi_n_8975, csa_tree_add_190_195_groupi_n_8976;
  wire csa_tree_add_190_195_groupi_n_8977, csa_tree_add_190_195_groupi_n_8978, csa_tree_add_190_195_groupi_n_8979, csa_tree_add_190_195_groupi_n_8980, csa_tree_add_190_195_groupi_n_8981, csa_tree_add_190_195_groupi_n_8982, csa_tree_add_190_195_groupi_n_8983, csa_tree_add_190_195_groupi_n_8984;
  wire csa_tree_add_190_195_groupi_n_8985, csa_tree_add_190_195_groupi_n_8986, csa_tree_add_190_195_groupi_n_8987, csa_tree_add_190_195_groupi_n_8988, csa_tree_add_190_195_groupi_n_8989, csa_tree_add_190_195_groupi_n_8990, csa_tree_add_190_195_groupi_n_8991, csa_tree_add_190_195_groupi_n_8992;
  wire csa_tree_add_190_195_groupi_n_8993, csa_tree_add_190_195_groupi_n_8994, csa_tree_add_190_195_groupi_n_8995, csa_tree_add_190_195_groupi_n_8996, csa_tree_add_190_195_groupi_n_8997, csa_tree_add_190_195_groupi_n_8998, csa_tree_add_190_195_groupi_n_8999, csa_tree_add_190_195_groupi_n_9000;
  wire csa_tree_add_190_195_groupi_n_9001, csa_tree_add_190_195_groupi_n_9002, csa_tree_add_190_195_groupi_n_9003, csa_tree_add_190_195_groupi_n_9004, csa_tree_add_190_195_groupi_n_9005, csa_tree_add_190_195_groupi_n_9006, csa_tree_add_190_195_groupi_n_9007, csa_tree_add_190_195_groupi_n_9008;
  wire csa_tree_add_190_195_groupi_n_9009, csa_tree_add_190_195_groupi_n_9010, csa_tree_add_190_195_groupi_n_9011, csa_tree_add_190_195_groupi_n_9012, csa_tree_add_190_195_groupi_n_9013, csa_tree_add_190_195_groupi_n_9014, csa_tree_add_190_195_groupi_n_9015, csa_tree_add_190_195_groupi_n_9016;
  wire csa_tree_add_190_195_groupi_n_9017, csa_tree_add_190_195_groupi_n_9018, csa_tree_add_190_195_groupi_n_9019, csa_tree_add_190_195_groupi_n_9020, csa_tree_add_190_195_groupi_n_9021, csa_tree_add_190_195_groupi_n_9022, csa_tree_add_190_195_groupi_n_9023, csa_tree_add_190_195_groupi_n_9024;
  wire csa_tree_add_190_195_groupi_n_9025, csa_tree_add_190_195_groupi_n_9026, csa_tree_add_190_195_groupi_n_9027, csa_tree_add_190_195_groupi_n_9028, csa_tree_add_190_195_groupi_n_9029, csa_tree_add_190_195_groupi_n_9030, csa_tree_add_190_195_groupi_n_9031, csa_tree_add_190_195_groupi_n_9032;
  wire csa_tree_add_190_195_groupi_n_9033, csa_tree_add_190_195_groupi_n_9034, csa_tree_add_190_195_groupi_n_9035, csa_tree_add_190_195_groupi_n_9036, csa_tree_add_190_195_groupi_n_9037, csa_tree_add_190_195_groupi_n_9038, csa_tree_add_190_195_groupi_n_9039, csa_tree_add_190_195_groupi_n_9040;
  wire csa_tree_add_190_195_groupi_n_9041, csa_tree_add_190_195_groupi_n_9042, csa_tree_add_190_195_groupi_n_9043, csa_tree_add_190_195_groupi_n_9044, csa_tree_add_190_195_groupi_n_9045, csa_tree_add_190_195_groupi_n_9046, csa_tree_add_190_195_groupi_n_9047, csa_tree_add_190_195_groupi_n_9048;
  wire csa_tree_add_190_195_groupi_n_9049, csa_tree_add_190_195_groupi_n_9050, csa_tree_add_190_195_groupi_n_9051, csa_tree_add_190_195_groupi_n_9052, csa_tree_add_190_195_groupi_n_9053, csa_tree_add_190_195_groupi_n_9054, csa_tree_add_190_195_groupi_n_9055, csa_tree_add_190_195_groupi_n_9056;
  wire csa_tree_add_190_195_groupi_n_9057, csa_tree_add_190_195_groupi_n_9058, csa_tree_add_190_195_groupi_n_9059, csa_tree_add_190_195_groupi_n_9060, csa_tree_add_190_195_groupi_n_9061, csa_tree_add_190_195_groupi_n_9062, csa_tree_add_190_195_groupi_n_9063, csa_tree_add_190_195_groupi_n_9064;
  wire csa_tree_add_190_195_groupi_n_9065, csa_tree_add_190_195_groupi_n_9066, csa_tree_add_190_195_groupi_n_9067, csa_tree_add_190_195_groupi_n_9068, csa_tree_add_190_195_groupi_n_9069, csa_tree_add_190_195_groupi_n_9070, csa_tree_add_190_195_groupi_n_9071, csa_tree_add_190_195_groupi_n_9072;
  wire csa_tree_add_190_195_groupi_n_9073, csa_tree_add_190_195_groupi_n_9074, csa_tree_add_190_195_groupi_n_9075, csa_tree_add_190_195_groupi_n_9076, csa_tree_add_190_195_groupi_n_9077, csa_tree_add_190_195_groupi_n_9078, csa_tree_add_190_195_groupi_n_9079, csa_tree_add_190_195_groupi_n_9080;
  wire csa_tree_add_190_195_groupi_n_9081, csa_tree_add_190_195_groupi_n_9082, csa_tree_add_190_195_groupi_n_9083, csa_tree_add_190_195_groupi_n_9084, csa_tree_add_190_195_groupi_n_9085, csa_tree_add_190_195_groupi_n_9086, csa_tree_add_190_195_groupi_n_9087, csa_tree_add_190_195_groupi_n_9088;
  wire csa_tree_add_190_195_groupi_n_9089, csa_tree_add_190_195_groupi_n_9090, csa_tree_add_190_195_groupi_n_9091, csa_tree_add_190_195_groupi_n_9092, csa_tree_add_190_195_groupi_n_9093, csa_tree_add_190_195_groupi_n_9094, csa_tree_add_190_195_groupi_n_9095, csa_tree_add_190_195_groupi_n_9096;
  wire csa_tree_add_190_195_groupi_n_9097, csa_tree_add_190_195_groupi_n_9098, csa_tree_add_190_195_groupi_n_9099, csa_tree_add_190_195_groupi_n_9100, csa_tree_add_190_195_groupi_n_9101, csa_tree_add_190_195_groupi_n_9102, csa_tree_add_190_195_groupi_n_9103, csa_tree_add_190_195_groupi_n_9104;
  wire csa_tree_add_190_195_groupi_n_9105, csa_tree_add_190_195_groupi_n_9106, csa_tree_add_190_195_groupi_n_9107, csa_tree_add_190_195_groupi_n_9108, csa_tree_add_190_195_groupi_n_9109, csa_tree_add_190_195_groupi_n_9110, csa_tree_add_190_195_groupi_n_9111, csa_tree_add_190_195_groupi_n_9112;
  wire csa_tree_add_190_195_groupi_n_9113, csa_tree_add_190_195_groupi_n_9114, csa_tree_add_190_195_groupi_n_9115, csa_tree_add_190_195_groupi_n_9116, csa_tree_add_190_195_groupi_n_9117, csa_tree_add_190_195_groupi_n_9118, csa_tree_add_190_195_groupi_n_9119, csa_tree_add_190_195_groupi_n_9120;
  wire csa_tree_add_190_195_groupi_n_9121, csa_tree_add_190_195_groupi_n_9122, csa_tree_add_190_195_groupi_n_9123, csa_tree_add_190_195_groupi_n_9124, csa_tree_add_190_195_groupi_n_9125, csa_tree_add_190_195_groupi_n_9126, csa_tree_add_190_195_groupi_n_9127, csa_tree_add_190_195_groupi_n_9128;
  wire csa_tree_add_190_195_groupi_n_9129, csa_tree_add_190_195_groupi_n_9130, csa_tree_add_190_195_groupi_n_9131, csa_tree_add_190_195_groupi_n_9132, csa_tree_add_190_195_groupi_n_9133, csa_tree_add_190_195_groupi_n_9134, csa_tree_add_190_195_groupi_n_9135, csa_tree_add_190_195_groupi_n_9136;
  wire csa_tree_add_190_195_groupi_n_9137, csa_tree_add_190_195_groupi_n_9138, csa_tree_add_190_195_groupi_n_9139, csa_tree_add_190_195_groupi_n_9140, csa_tree_add_190_195_groupi_n_9141, csa_tree_add_190_195_groupi_n_9142, csa_tree_add_190_195_groupi_n_9143, csa_tree_add_190_195_groupi_n_9144;
  wire csa_tree_add_190_195_groupi_n_9145, csa_tree_add_190_195_groupi_n_9146, csa_tree_add_190_195_groupi_n_9147, csa_tree_add_190_195_groupi_n_9148, csa_tree_add_190_195_groupi_n_9149, csa_tree_add_190_195_groupi_n_9150, csa_tree_add_190_195_groupi_n_9151, csa_tree_add_190_195_groupi_n_9152;
  wire csa_tree_add_190_195_groupi_n_9153, csa_tree_add_190_195_groupi_n_9154, csa_tree_add_190_195_groupi_n_9155, csa_tree_add_190_195_groupi_n_9156, csa_tree_add_190_195_groupi_n_9157, csa_tree_add_190_195_groupi_n_9158, csa_tree_add_190_195_groupi_n_9159, csa_tree_add_190_195_groupi_n_9160;
  wire csa_tree_add_190_195_groupi_n_9161, csa_tree_add_190_195_groupi_n_9162, csa_tree_add_190_195_groupi_n_9163, csa_tree_add_190_195_groupi_n_9164, csa_tree_add_190_195_groupi_n_9165, csa_tree_add_190_195_groupi_n_9166, csa_tree_add_190_195_groupi_n_9167, csa_tree_add_190_195_groupi_n_9168;
  wire csa_tree_add_190_195_groupi_n_9169, csa_tree_add_190_195_groupi_n_9170, csa_tree_add_190_195_groupi_n_9171, csa_tree_add_190_195_groupi_n_9172, csa_tree_add_190_195_groupi_n_9173, csa_tree_add_190_195_groupi_n_9174, csa_tree_add_190_195_groupi_n_9175, csa_tree_add_190_195_groupi_n_9176;
  wire csa_tree_add_190_195_groupi_n_9177, csa_tree_add_190_195_groupi_n_9178, csa_tree_add_190_195_groupi_n_9179, csa_tree_add_190_195_groupi_n_9180, csa_tree_add_190_195_groupi_n_9181, csa_tree_add_190_195_groupi_n_9182, csa_tree_add_190_195_groupi_n_9183, csa_tree_add_190_195_groupi_n_9184;
  wire csa_tree_add_190_195_groupi_n_9185, csa_tree_add_190_195_groupi_n_9186, csa_tree_add_190_195_groupi_n_9187, csa_tree_add_190_195_groupi_n_9188, csa_tree_add_190_195_groupi_n_9189, csa_tree_add_190_195_groupi_n_9190, csa_tree_add_190_195_groupi_n_9191, csa_tree_add_190_195_groupi_n_9192;
  wire csa_tree_add_190_195_groupi_n_9193, csa_tree_add_190_195_groupi_n_9194, csa_tree_add_190_195_groupi_n_9195, csa_tree_add_190_195_groupi_n_9196, csa_tree_add_190_195_groupi_n_9197, csa_tree_add_190_195_groupi_n_9198, csa_tree_add_190_195_groupi_n_9199, csa_tree_add_190_195_groupi_n_9200;
  wire csa_tree_add_190_195_groupi_n_9201, csa_tree_add_190_195_groupi_n_9202, csa_tree_add_190_195_groupi_n_9203, csa_tree_add_190_195_groupi_n_9204, csa_tree_add_190_195_groupi_n_9205, csa_tree_add_190_195_groupi_n_9206, csa_tree_add_190_195_groupi_n_9207, csa_tree_add_190_195_groupi_n_9208;
  wire csa_tree_add_190_195_groupi_n_9209, csa_tree_add_190_195_groupi_n_9210, csa_tree_add_190_195_groupi_n_9211, csa_tree_add_190_195_groupi_n_9212, csa_tree_add_190_195_groupi_n_9213, csa_tree_add_190_195_groupi_n_9214, csa_tree_add_190_195_groupi_n_9215, csa_tree_add_190_195_groupi_n_9216;
  wire csa_tree_add_190_195_groupi_n_9217, csa_tree_add_190_195_groupi_n_9218, csa_tree_add_190_195_groupi_n_9219, csa_tree_add_190_195_groupi_n_9220, csa_tree_add_190_195_groupi_n_9221, csa_tree_add_190_195_groupi_n_9222, csa_tree_add_190_195_groupi_n_9223, csa_tree_add_190_195_groupi_n_9224;
  wire csa_tree_add_190_195_groupi_n_9225, csa_tree_add_190_195_groupi_n_9226, csa_tree_add_190_195_groupi_n_9227, csa_tree_add_190_195_groupi_n_9228, csa_tree_add_190_195_groupi_n_9229, csa_tree_add_190_195_groupi_n_9230, csa_tree_add_190_195_groupi_n_9231, csa_tree_add_190_195_groupi_n_9232;
  wire csa_tree_add_190_195_groupi_n_9233, csa_tree_add_190_195_groupi_n_9234, csa_tree_add_190_195_groupi_n_9235, csa_tree_add_190_195_groupi_n_9236, csa_tree_add_190_195_groupi_n_9237, csa_tree_add_190_195_groupi_n_9238, csa_tree_add_190_195_groupi_n_9239, csa_tree_add_190_195_groupi_n_9240;
  wire csa_tree_add_190_195_groupi_n_9241, csa_tree_add_190_195_groupi_n_9242, csa_tree_add_190_195_groupi_n_9243, csa_tree_add_190_195_groupi_n_9244, csa_tree_add_190_195_groupi_n_9245, csa_tree_add_190_195_groupi_n_9246, csa_tree_add_190_195_groupi_n_9247, csa_tree_add_190_195_groupi_n_9248;
  wire csa_tree_add_190_195_groupi_n_9249, csa_tree_add_190_195_groupi_n_9250, csa_tree_add_190_195_groupi_n_9251, csa_tree_add_190_195_groupi_n_9252, csa_tree_add_190_195_groupi_n_9253, csa_tree_add_190_195_groupi_n_9254, csa_tree_add_190_195_groupi_n_9255, csa_tree_add_190_195_groupi_n_9256;
  wire csa_tree_add_190_195_groupi_n_9257, csa_tree_add_190_195_groupi_n_9258, csa_tree_add_190_195_groupi_n_9259, csa_tree_add_190_195_groupi_n_9260, csa_tree_add_190_195_groupi_n_9261, csa_tree_add_190_195_groupi_n_9262, csa_tree_add_190_195_groupi_n_9263, csa_tree_add_190_195_groupi_n_9264;
  wire csa_tree_add_190_195_groupi_n_9265, csa_tree_add_190_195_groupi_n_9266, csa_tree_add_190_195_groupi_n_9267, csa_tree_add_190_195_groupi_n_9268, csa_tree_add_190_195_groupi_n_9269, csa_tree_add_190_195_groupi_n_9270, csa_tree_add_190_195_groupi_n_9271, csa_tree_add_190_195_groupi_n_9272;
  wire csa_tree_add_190_195_groupi_n_9273, csa_tree_add_190_195_groupi_n_9274, csa_tree_add_190_195_groupi_n_9275, csa_tree_add_190_195_groupi_n_9276, csa_tree_add_190_195_groupi_n_9277, csa_tree_add_190_195_groupi_n_9278, csa_tree_add_190_195_groupi_n_9279, csa_tree_add_190_195_groupi_n_9280;
  wire csa_tree_add_190_195_groupi_n_9281, csa_tree_add_190_195_groupi_n_9282, csa_tree_add_190_195_groupi_n_9283, csa_tree_add_190_195_groupi_n_9284, csa_tree_add_190_195_groupi_n_9285, csa_tree_add_190_195_groupi_n_9286, csa_tree_add_190_195_groupi_n_9287, csa_tree_add_190_195_groupi_n_9288;
  wire csa_tree_add_190_195_groupi_n_9289, csa_tree_add_190_195_groupi_n_9290, csa_tree_add_190_195_groupi_n_9291, csa_tree_add_190_195_groupi_n_9292, csa_tree_add_190_195_groupi_n_9293, csa_tree_add_190_195_groupi_n_9294, csa_tree_add_190_195_groupi_n_9295, csa_tree_add_190_195_groupi_n_9296;
  wire csa_tree_add_190_195_groupi_n_9297, csa_tree_add_190_195_groupi_n_9298, csa_tree_add_190_195_groupi_n_9299, csa_tree_add_190_195_groupi_n_9300, csa_tree_add_190_195_groupi_n_9301, csa_tree_add_190_195_groupi_n_9302, csa_tree_add_190_195_groupi_n_9303, csa_tree_add_190_195_groupi_n_9304;
  wire csa_tree_add_190_195_groupi_n_9305, csa_tree_add_190_195_groupi_n_9306, csa_tree_add_190_195_groupi_n_9307, csa_tree_add_190_195_groupi_n_9308, csa_tree_add_190_195_groupi_n_9309, csa_tree_add_190_195_groupi_n_9310, csa_tree_add_190_195_groupi_n_9311, csa_tree_add_190_195_groupi_n_9312;
  wire csa_tree_add_190_195_groupi_n_9313, csa_tree_add_190_195_groupi_n_9314, csa_tree_add_190_195_groupi_n_9315, csa_tree_add_190_195_groupi_n_9316, csa_tree_add_190_195_groupi_n_9317, csa_tree_add_190_195_groupi_n_9318, csa_tree_add_190_195_groupi_n_9319, csa_tree_add_190_195_groupi_n_9320;
  wire csa_tree_add_190_195_groupi_n_9321, csa_tree_add_190_195_groupi_n_9322, csa_tree_add_190_195_groupi_n_9323, csa_tree_add_190_195_groupi_n_9324, csa_tree_add_190_195_groupi_n_9325, csa_tree_add_190_195_groupi_n_9326, csa_tree_add_190_195_groupi_n_9327, csa_tree_add_190_195_groupi_n_9328;
  wire csa_tree_add_190_195_groupi_n_9329, csa_tree_add_190_195_groupi_n_9330, csa_tree_add_190_195_groupi_n_9331, csa_tree_add_190_195_groupi_n_9332, csa_tree_add_190_195_groupi_n_9333, csa_tree_add_190_195_groupi_n_9334, csa_tree_add_190_195_groupi_n_9335, csa_tree_add_190_195_groupi_n_9336;
  wire csa_tree_add_190_195_groupi_n_9337, csa_tree_add_190_195_groupi_n_9338, csa_tree_add_190_195_groupi_n_9339, csa_tree_add_190_195_groupi_n_9340, csa_tree_add_190_195_groupi_n_9341, csa_tree_add_190_195_groupi_n_9342, csa_tree_add_190_195_groupi_n_9343, csa_tree_add_190_195_groupi_n_9344;
  wire csa_tree_add_190_195_groupi_n_9345, csa_tree_add_190_195_groupi_n_9346, csa_tree_add_190_195_groupi_n_9347, csa_tree_add_190_195_groupi_n_9348, csa_tree_add_190_195_groupi_n_9349, csa_tree_add_190_195_groupi_n_9350, csa_tree_add_190_195_groupi_n_9351, csa_tree_add_190_195_groupi_n_9352;
  wire csa_tree_add_190_195_groupi_n_9353, csa_tree_add_190_195_groupi_n_9354, csa_tree_add_190_195_groupi_n_9355, csa_tree_add_190_195_groupi_n_9356, csa_tree_add_190_195_groupi_n_9357, csa_tree_add_190_195_groupi_n_9358, csa_tree_add_190_195_groupi_n_9359, csa_tree_add_190_195_groupi_n_9360;
  wire csa_tree_add_190_195_groupi_n_9361, csa_tree_add_190_195_groupi_n_9362, csa_tree_add_190_195_groupi_n_9363, csa_tree_add_190_195_groupi_n_9364, csa_tree_add_190_195_groupi_n_9365, csa_tree_add_190_195_groupi_n_9366, csa_tree_add_190_195_groupi_n_9367, csa_tree_add_190_195_groupi_n_9368;
  wire csa_tree_add_190_195_groupi_n_9369, csa_tree_add_190_195_groupi_n_9370, csa_tree_add_190_195_groupi_n_9371, csa_tree_add_190_195_groupi_n_9372, csa_tree_add_190_195_groupi_n_9373, csa_tree_add_190_195_groupi_n_9374, csa_tree_add_190_195_groupi_n_9375, csa_tree_add_190_195_groupi_n_9376;
  wire csa_tree_add_190_195_groupi_n_9377, csa_tree_add_190_195_groupi_n_9378, csa_tree_add_190_195_groupi_n_9379, csa_tree_add_190_195_groupi_n_9380, csa_tree_add_190_195_groupi_n_9381, csa_tree_add_190_195_groupi_n_9382, csa_tree_add_190_195_groupi_n_9383, csa_tree_add_190_195_groupi_n_9384;
  wire csa_tree_add_190_195_groupi_n_9385, csa_tree_add_190_195_groupi_n_9386, csa_tree_add_190_195_groupi_n_9387, csa_tree_add_190_195_groupi_n_9388, csa_tree_add_190_195_groupi_n_9389, csa_tree_add_190_195_groupi_n_9390, csa_tree_add_190_195_groupi_n_9391, csa_tree_add_190_195_groupi_n_9392;
  wire csa_tree_add_190_195_groupi_n_9393, csa_tree_add_190_195_groupi_n_9394, csa_tree_add_190_195_groupi_n_9395, csa_tree_add_190_195_groupi_n_9396, csa_tree_add_190_195_groupi_n_9397, csa_tree_add_190_195_groupi_n_9398, csa_tree_add_190_195_groupi_n_9399, csa_tree_add_190_195_groupi_n_9400;
  wire csa_tree_add_190_195_groupi_n_9401, csa_tree_add_190_195_groupi_n_9402, csa_tree_add_190_195_groupi_n_9403, csa_tree_add_190_195_groupi_n_9404, csa_tree_add_190_195_groupi_n_9405, csa_tree_add_190_195_groupi_n_9406, csa_tree_add_190_195_groupi_n_9407, csa_tree_add_190_195_groupi_n_9408;
  wire csa_tree_add_190_195_groupi_n_9409, csa_tree_add_190_195_groupi_n_9410, csa_tree_add_190_195_groupi_n_9411, csa_tree_add_190_195_groupi_n_9412, csa_tree_add_190_195_groupi_n_9413, csa_tree_add_190_195_groupi_n_9414, csa_tree_add_190_195_groupi_n_9415, csa_tree_add_190_195_groupi_n_9416;
  wire csa_tree_add_190_195_groupi_n_9417, csa_tree_add_190_195_groupi_n_9418, csa_tree_add_190_195_groupi_n_9419, csa_tree_add_190_195_groupi_n_9420, csa_tree_add_190_195_groupi_n_9421, csa_tree_add_190_195_groupi_n_9422, csa_tree_add_190_195_groupi_n_9423, csa_tree_add_190_195_groupi_n_9424;
  wire csa_tree_add_190_195_groupi_n_9425, csa_tree_add_190_195_groupi_n_9426, csa_tree_add_190_195_groupi_n_9427, csa_tree_add_190_195_groupi_n_9428, csa_tree_add_190_195_groupi_n_9429, csa_tree_add_190_195_groupi_n_9430, csa_tree_add_190_195_groupi_n_9431, csa_tree_add_190_195_groupi_n_9432;
  wire csa_tree_add_190_195_groupi_n_9433, csa_tree_add_190_195_groupi_n_9434, csa_tree_add_190_195_groupi_n_9435, csa_tree_add_190_195_groupi_n_9436, csa_tree_add_190_195_groupi_n_9437, csa_tree_add_190_195_groupi_n_9438, csa_tree_add_190_195_groupi_n_9439, csa_tree_add_190_195_groupi_n_9440;
  wire csa_tree_add_190_195_groupi_n_9441, csa_tree_add_190_195_groupi_n_9442, csa_tree_add_190_195_groupi_n_9443, csa_tree_add_190_195_groupi_n_9444, csa_tree_add_190_195_groupi_n_9445, csa_tree_add_190_195_groupi_n_9446, csa_tree_add_190_195_groupi_n_9447, csa_tree_add_190_195_groupi_n_9448;
  wire csa_tree_add_190_195_groupi_n_9449, csa_tree_add_190_195_groupi_n_9450, csa_tree_add_190_195_groupi_n_9451, csa_tree_add_190_195_groupi_n_9452, csa_tree_add_190_195_groupi_n_9453, csa_tree_add_190_195_groupi_n_9454, csa_tree_add_190_195_groupi_n_9455, csa_tree_add_190_195_groupi_n_9456;
  wire csa_tree_add_190_195_groupi_n_9457, csa_tree_add_190_195_groupi_n_9458, csa_tree_add_190_195_groupi_n_9459, csa_tree_add_190_195_groupi_n_9460, csa_tree_add_190_195_groupi_n_9461, csa_tree_add_190_195_groupi_n_9462, csa_tree_add_190_195_groupi_n_9463, csa_tree_add_190_195_groupi_n_9464;
  wire csa_tree_add_190_195_groupi_n_9465, csa_tree_add_190_195_groupi_n_9466, csa_tree_add_190_195_groupi_n_9467, csa_tree_add_190_195_groupi_n_9468, csa_tree_add_190_195_groupi_n_9469, csa_tree_add_190_195_groupi_n_9470, csa_tree_add_190_195_groupi_n_9471, csa_tree_add_190_195_groupi_n_9472;
  wire csa_tree_add_190_195_groupi_n_9473, csa_tree_add_190_195_groupi_n_9474, csa_tree_add_190_195_groupi_n_9475, csa_tree_add_190_195_groupi_n_9476, csa_tree_add_190_195_groupi_n_9477, csa_tree_add_190_195_groupi_n_9478, csa_tree_add_190_195_groupi_n_9479, csa_tree_add_190_195_groupi_n_9480;
  wire csa_tree_add_190_195_groupi_n_9481, csa_tree_add_190_195_groupi_n_9482, csa_tree_add_190_195_groupi_n_9483, csa_tree_add_190_195_groupi_n_9484, csa_tree_add_190_195_groupi_n_9485, csa_tree_add_190_195_groupi_n_9486, csa_tree_add_190_195_groupi_n_9487, csa_tree_add_190_195_groupi_n_9488;
  wire csa_tree_add_190_195_groupi_n_9489, csa_tree_add_190_195_groupi_n_9490, csa_tree_add_190_195_groupi_n_9491, csa_tree_add_190_195_groupi_n_9492, csa_tree_add_190_195_groupi_n_9493, csa_tree_add_190_195_groupi_n_9494, csa_tree_add_190_195_groupi_n_9495, csa_tree_add_190_195_groupi_n_9496;
  wire csa_tree_add_190_195_groupi_n_9497, csa_tree_add_190_195_groupi_n_9498, csa_tree_add_190_195_groupi_n_9499, csa_tree_add_190_195_groupi_n_9500, csa_tree_add_190_195_groupi_n_9501, csa_tree_add_190_195_groupi_n_9502, csa_tree_add_190_195_groupi_n_9503, csa_tree_add_190_195_groupi_n_9504;
  wire csa_tree_add_190_195_groupi_n_9505, csa_tree_add_190_195_groupi_n_9506, csa_tree_add_190_195_groupi_n_9507, csa_tree_add_190_195_groupi_n_9508, csa_tree_add_190_195_groupi_n_9509, csa_tree_add_190_195_groupi_n_9510, csa_tree_add_190_195_groupi_n_9511, csa_tree_add_190_195_groupi_n_9512;
  wire csa_tree_add_190_195_groupi_n_9513, csa_tree_add_190_195_groupi_n_9514, csa_tree_add_190_195_groupi_n_9515, csa_tree_add_190_195_groupi_n_9516, csa_tree_add_190_195_groupi_n_9517, csa_tree_add_190_195_groupi_n_9518, csa_tree_add_190_195_groupi_n_9519, csa_tree_add_190_195_groupi_n_9520;
  wire csa_tree_add_190_195_groupi_n_9521, csa_tree_add_190_195_groupi_n_9522, csa_tree_add_190_195_groupi_n_9523, csa_tree_add_190_195_groupi_n_9524, csa_tree_add_190_195_groupi_n_9525, csa_tree_add_190_195_groupi_n_9526, csa_tree_add_190_195_groupi_n_9527, csa_tree_add_190_195_groupi_n_9528;
  wire csa_tree_add_190_195_groupi_n_9529, csa_tree_add_190_195_groupi_n_9530, csa_tree_add_190_195_groupi_n_9531, csa_tree_add_190_195_groupi_n_9532, csa_tree_add_190_195_groupi_n_9533, csa_tree_add_190_195_groupi_n_9534, csa_tree_add_190_195_groupi_n_9535, csa_tree_add_190_195_groupi_n_9536;
  wire csa_tree_add_190_195_groupi_n_9537, csa_tree_add_190_195_groupi_n_9538, csa_tree_add_190_195_groupi_n_9539, csa_tree_add_190_195_groupi_n_9540, csa_tree_add_190_195_groupi_n_9541, csa_tree_add_190_195_groupi_n_9542, csa_tree_add_190_195_groupi_n_9543, csa_tree_add_190_195_groupi_n_9544;
  wire csa_tree_add_190_195_groupi_n_9545, csa_tree_add_190_195_groupi_n_9546, csa_tree_add_190_195_groupi_n_9547, csa_tree_add_190_195_groupi_n_9548, csa_tree_add_190_195_groupi_n_9549, csa_tree_add_190_195_groupi_n_9550, csa_tree_add_190_195_groupi_n_9551, csa_tree_add_190_195_groupi_n_9552;
  wire csa_tree_add_190_195_groupi_n_9553, csa_tree_add_190_195_groupi_n_9554, csa_tree_add_190_195_groupi_n_9555, csa_tree_add_190_195_groupi_n_9556, csa_tree_add_190_195_groupi_n_9557, csa_tree_add_190_195_groupi_n_9558, csa_tree_add_190_195_groupi_n_9559, csa_tree_add_190_195_groupi_n_9560;
  wire csa_tree_add_190_195_groupi_n_9561, csa_tree_add_190_195_groupi_n_9562, csa_tree_add_190_195_groupi_n_9563, csa_tree_add_190_195_groupi_n_9564, csa_tree_add_190_195_groupi_n_9565, csa_tree_add_190_195_groupi_n_9566, csa_tree_add_190_195_groupi_n_9567, csa_tree_add_190_195_groupi_n_9568;
  wire csa_tree_add_190_195_groupi_n_9569, csa_tree_add_190_195_groupi_n_9570, csa_tree_add_190_195_groupi_n_9571, csa_tree_add_190_195_groupi_n_9572, csa_tree_add_190_195_groupi_n_9573, csa_tree_add_190_195_groupi_n_9574, csa_tree_add_190_195_groupi_n_9575, csa_tree_add_190_195_groupi_n_9576;
  wire csa_tree_add_190_195_groupi_n_9577, csa_tree_add_190_195_groupi_n_9578, csa_tree_add_190_195_groupi_n_9579, csa_tree_add_190_195_groupi_n_9580, csa_tree_add_190_195_groupi_n_9581, csa_tree_add_190_195_groupi_n_9582, csa_tree_add_190_195_groupi_n_9583, csa_tree_add_190_195_groupi_n_9584;
  wire csa_tree_add_190_195_groupi_n_9585, csa_tree_add_190_195_groupi_n_9586, csa_tree_add_190_195_groupi_n_9587, csa_tree_add_190_195_groupi_n_9588, csa_tree_add_190_195_groupi_n_9589, csa_tree_add_190_195_groupi_n_9590, csa_tree_add_190_195_groupi_n_9591, csa_tree_add_190_195_groupi_n_9592;
  wire csa_tree_add_190_195_groupi_n_9593, csa_tree_add_190_195_groupi_n_9594, csa_tree_add_190_195_groupi_n_9595, csa_tree_add_190_195_groupi_n_9596, csa_tree_add_190_195_groupi_n_9597, csa_tree_add_190_195_groupi_n_9598, csa_tree_add_190_195_groupi_n_9599, csa_tree_add_190_195_groupi_n_9600;
  wire csa_tree_add_190_195_groupi_n_9601, csa_tree_add_190_195_groupi_n_9602, csa_tree_add_190_195_groupi_n_9603, csa_tree_add_190_195_groupi_n_9604, csa_tree_add_190_195_groupi_n_9605, csa_tree_add_190_195_groupi_n_9606, csa_tree_add_190_195_groupi_n_9607, csa_tree_add_190_195_groupi_n_9608;
  wire csa_tree_add_190_195_groupi_n_9609, csa_tree_add_190_195_groupi_n_9610, csa_tree_add_190_195_groupi_n_9611, csa_tree_add_190_195_groupi_n_9612, csa_tree_add_190_195_groupi_n_9613, csa_tree_add_190_195_groupi_n_9614, csa_tree_add_190_195_groupi_n_9615, csa_tree_add_190_195_groupi_n_9616;
  wire csa_tree_add_190_195_groupi_n_9617, csa_tree_add_190_195_groupi_n_9618, csa_tree_add_190_195_groupi_n_9619, csa_tree_add_190_195_groupi_n_9620, csa_tree_add_190_195_groupi_n_9621, csa_tree_add_190_195_groupi_n_9622, csa_tree_add_190_195_groupi_n_9623, csa_tree_add_190_195_groupi_n_9624;
  wire csa_tree_add_190_195_groupi_n_9625, csa_tree_add_190_195_groupi_n_9626, csa_tree_add_190_195_groupi_n_9627, csa_tree_add_190_195_groupi_n_9628, csa_tree_add_190_195_groupi_n_9629, csa_tree_add_190_195_groupi_n_9630, csa_tree_add_190_195_groupi_n_9631, csa_tree_add_190_195_groupi_n_9632;
  wire csa_tree_add_190_195_groupi_n_9633, csa_tree_add_190_195_groupi_n_9634, csa_tree_add_190_195_groupi_n_9635, csa_tree_add_190_195_groupi_n_9636, csa_tree_add_190_195_groupi_n_9637, csa_tree_add_190_195_groupi_n_9638, csa_tree_add_190_195_groupi_n_9639, csa_tree_add_190_195_groupi_n_9640;
  wire csa_tree_add_190_195_groupi_n_9641, csa_tree_add_190_195_groupi_n_9642, csa_tree_add_190_195_groupi_n_9643, csa_tree_add_190_195_groupi_n_9644, csa_tree_add_190_195_groupi_n_9645, csa_tree_add_190_195_groupi_n_9646, csa_tree_add_190_195_groupi_n_9647, csa_tree_add_190_195_groupi_n_9648;
  wire csa_tree_add_190_195_groupi_n_9649, csa_tree_add_190_195_groupi_n_9650, csa_tree_add_190_195_groupi_n_9651, csa_tree_add_190_195_groupi_n_9652, csa_tree_add_190_195_groupi_n_9653, csa_tree_add_190_195_groupi_n_9654, csa_tree_add_190_195_groupi_n_9655, csa_tree_add_190_195_groupi_n_9656;
  wire csa_tree_add_190_195_groupi_n_9657, csa_tree_add_190_195_groupi_n_9658, csa_tree_add_190_195_groupi_n_9659, csa_tree_add_190_195_groupi_n_9660, csa_tree_add_190_195_groupi_n_9661, csa_tree_add_190_195_groupi_n_9662, csa_tree_add_190_195_groupi_n_9663, csa_tree_add_190_195_groupi_n_9664;
  wire csa_tree_add_190_195_groupi_n_9665, csa_tree_add_190_195_groupi_n_9666, csa_tree_add_190_195_groupi_n_9667, csa_tree_add_190_195_groupi_n_9668, csa_tree_add_190_195_groupi_n_9669, csa_tree_add_190_195_groupi_n_9670, csa_tree_add_190_195_groupi_n_9671, csa_tree_add_190_195_groupi_n_9672;
  wire csa_tree_add_190_195_groupi_n_9673, csa_tree_add_190_195_groupi_n_9674, csa_tree_add_190_195_groupi_n_9675, csa_tree_add_190_195_groupi_n_9676, csa_tree_add_190_195_groupi_n_9677, csa_tree_add_190_195_groupi_n_9678, csa_tree_add_190_195_groupi_n_9679, csa_tree_add_190_195_groupi_n_9680;
  wire csa_tree_add_190_195_groupi_n_9681, csa_tree_add_190_195_groupi_n_9682, csa_tree_add_190_195_groupi_n_9683, csa_tree_add_190_195_groupi_n_9684, csa_tree_add_190_195_groupi_n_9685, csa_tree_add_190_195_groupi_n_9686, csa_tree_add_190_195_groupi_n_9687, csa_tree_add_190_195_groupi_n_9688;
  wire csa_tree_add_190_195_groupi_n_9689, csa_tree_add_190_195_groupi_n_9690, csa_tree_add_190_195_groupi_n_9691, csa_tree_add_190_195_groupi_n_9692, csa_tree_add_190_195_groupi_n_9693, csa_tree_add_190_195_groupi_n_9694, csa_tree_add_190_195_groupi_n_9695, csa_tree_add_190_195_groupi_n_9696;
  wire csa_tree_add_190_195_groupi_n_9697, csa_tree_add_190_195_groupi_n_9698, csa_tree_add_190_195_groupi_n_9699, csa_tree_add_190_195_groupi_n_9700, csa_tree_add_190_195_groupi_n_9701, csa_tree_add_190_195_groupi_n_9702, csa_tree_add_190_195_groupi_n_9703, csa_tree_add_190_195_groupi_n_9704;
  wire csa_tree_add_190_195_groupi_n_9705, csa_tree_add_190_195_groupi_n_9706, csa_tree_add_190_195_groupi_n_9707, csa_tree_add_190_195_groupi_n_9708, csa_tree_add_190_195_groupi_n_9709, csa_tree_add_190_195_groupi_n_9710, csa_tree_add_190_195_groupi_n_9711, csa_tree_add_190_195_groupi_n_9712;
  wire csa_tree_add_190_195_groupi_n_9713, csa_tree_add_190_195_groupi_n_9714, csa_tree_add_190_195_groupi_n_9715, csa_tree_add_190_195_groupi_n_9716, csa_tree_add_190_195_groupi_n_9717, csa_tree_add_190_195_groupi_n_9718, csa_tree_add_190_195_groupi_n_9719, csa_tree_add_190_195_groupi_n_9720;
  wire csa_tree_add_190_195_groupi_n_9721, csa_tree_add_190_195_groupi_n_9722, csa_tree_add_190_195_groupi_n_9723, csa_tree_add_190_195_groupi_n_9724, csa_tree_add_190_195_groupi_n_9725, csa_tree_add_190_195_groupi_n_9726, csa_tree_add_190_195_groupi_n_9727, csa_tree_add_190_195_groupi_n_9728;
  wire csa_tree_add_190_195_groupi_n_9729, csa_tree_add_190_195_groupi_n_9730, csa_tree_add_190_195_groupi_n_9731, csa_tree_add_190_195_groupi_n_9732, csa_tree_add_190_195_groupi_n_9733, csa_tree_add_190_195_groupi_n_9734, csa_tree_add_190_195_groupi_n_9735, csa_tree_add_190_195_groupi_n_9736;
  wire csa_tree_add_190_195_groupi_n_9737, csa_tree_add_190_195_groupi_n_9738, csa_tree_add_190_195_groupi_n_9739, csa_tree_add_190_195_groupi_n_9740, csa_tree_add_190_195_groupi_n_9741, csa_tree_add_190_195_groupi_n_9742, csa_tree_add_190_195_groupi_n_9743, csa_tree_add_190_195_groupi_n_9744;
  wire csa_tree_add_190_195_groupi_n_9745, csa_tree_add_190_195_groupi_n_9746, csa_tree_add_190_195_groupi_n_9747, csa_tree_add_190_195_groupi_n_9748, csa_tree_add_190_195_groupi_n_9749, csa_tree_add_190_195_groupi_n_9750, csa_tree_add_190_195_groupi_n_9751, csa_tree_add_190_195_groupi_n_9752;
  wire csa_tree_add_190_195_groupi_n_9753, csa_tree_add_190_195_groupi_n_9754, csa_tree_add_190_195_groupi_n_9755, csa_tree_add_190_195_groupi_n_9756, csa_tree_add_190_195_groupi_n_9757, csa_tree_add_190_195_groupi_n_9758, csa_tree_add_190_195_groupi_n_9759, csa_tree_add_190_195_groupi_n_9760;
  wire csa_tree_add_190_195_groupi_n_9761, csa_tree_add_190_195_groupi_n_9762, csa_tree_add_190_195_groupi_n_9763, csa_tree_add_190_195_groupi_n_9764, csa_tree_add_190_195_groupi_n_9765, csa_tree_add_190_195_groupi_n_9766, csa_tree_add_190_195_groupi_n_9767, csa_tree_add_190_195_groupi_n_9768;
  wire csa_tree_add_190_195_groupi_n_9769, csa_tree_add_190_195_groupi_n_9770, csa_tree_add_190_195_groupi_n_9771, csa_tree_add_190_195_groupi_n_9772, csa_tree_add_190_195_groupi_n_9773, csa_tree_add_190_195_groupi_n_9774, csa_tree_add_190_195_groupi_n_9775, csa_tree_add_190_195_groupi_n_9776;
  wire csa_tree_add_190_195_groupi_n_9777, csa_tree_add_190_195_groupi_n_9778, csa_tree_add_190_195_groupi_n_9779, csa_tree_add_190_195_groupi_n_9780, csa_tree_add_190_195_groupi_n_9781, csa_tree_add_190_195_groupi_n_9782, csa_tree_add_190_195_groupi_n_9783, csa_tree_add_190_195_groupi_n_9784;
  wire csa_tree_add_190_195_groupi_n_9785, csa_tree_add_190_195_groupi_n_9786, csa_tree_add_190_195_groupi_n_9787, csa_tree_add_190_195_groupi_n_9788, csa_tree_add_190_195_groupi_n_9789, csa_tree_add_190_195_groupi_n_9790, csa_tree_add_190_195_groupi_n_9791, csa_tree_add_190_195_groupi_n_9792;
  wire csa_tree_add_190_195_groupi_n_9793, csa_tree_add_190_195_groupi_n_9794, csa_tree_add_190_195_groupi_n_9795, csa_tree_add_190_195_groupi_n_9796, csa_tree_add_190_195_groupi_n_9797, csa_tree_add_190_195_groupi_n_9798, csa_tree_add_190_195_groupi_n_9799, csa_tree_add_190_195_groupi_n_9800;
  wire csa_tree_add_190_195_groupi_n_9801, csa_tree_add_190_195_groupi_n_9802, csa_tree_add_190_195_groupi_n_9803, csa_tree_add_190_195_groupi_n_9804, csa_tree_add_190_195_groupi_n_9805, csa_tree_add_190_195_groupi_n_9806, csa_tree_add_190_195_groupi_n_9807, csa_tree_add_190_195_groupi_n_9808;
  wire csa_tree_add_190_195_groupi_n_9809, csa_tree_add_190_195_groupi_n_9810, csa_tree_add_190_195_groupi_n_9811, csa_tree_add_190_195_groupi_n_9812, csa_tree_add_190_195_groupi_n_9813, csa_tree_add_190_195_groupi_n_9814, csa_tree_add_190_195_groupi_n_9815, csa_tree_add_190_195_groupi_n_9816;
  wire csa_tree_add_190_195_groupi_n_9817, csa_tree_add_190_195_groupi_n_9818, csa_tree_add_190_195_groupi_n_9819, csa_tree_add_190_195_groupi_n_9820, csa_tree_add_190_195_groupi_n_9821, csa_tree_add_190_195_groupi_n_9822, csa_tree_add_190_195_groupi_n_9823, csa_tree_add_190_195_groupi_n_9824;
  wire csa_tree_add_190_195_groupi_n_9825, csa_tree_add_190_195_groupi_n_9826, csa_tree_add_190_195_groupi_n_9827, csa_tree_add_190_195_groupi_n_9828, csa_tree_add_190_195_groupi_n_9829, csa_tree_add_190_195_groupi_n_9830, csa_tree_add_190_195_groupi_n_9831, csa_tree_add_190_195_groupi_n_9832;
  wire csa_tree_add_190_195_groupi_n_9833, csa_tree_add_190_195_groupi_n_9834, csa_tree_add_190_195_groupi_n_9835, csa_tree_add_190_195_groupi_n_9836, csa_tree_add_190_195_groupi_n_9837, csa_tree_add_190_195_groupi_n_9838, csa_tree_add_190_195_groupi_n_9839, csa_tree_add_190_195_groupi_n_9840;
  wire csa_tree_add_190_195_groupi_n_9841, csa_tree_add_190_195_groupi_n_9842, csa_tree_add_190_195_groupi_n_9843, csa_tree_add_190_195_groupi_n_9844, csa_tree_add_190_195_groupi_n_9845, csa_tree_add_190_195_groupi_n_9846, csa_tree_add_190_195_groupi_n_9847, csa_tree_add_190_195_groupi_n_9848;
  wire csa_tree_add_190_195_groupi_n_9849, csa_tree_add_190_195_groupi_n_9850, csa_tree_add_190_195_groupi_n_9851, csa_tree_add_190_195_groupi_n_9852, csa_tree_add_190_195_groupi_n_9853, csa_tree_add_190_195_groupi_n_9854, csa_tree_add_190_195_groupi_n_9855, csa_tree_add_190_195_groupi_n_9856;
  wire csa_tree_add_190_195_groupi_n_9857, csa_tree_add_190_195_groupi_n_9858, csa_tree_add_190_195_groupi_n_9859, csa_tree_add_190_195_groupi_n_9860, csa_tree_add_190_195_groupi_n_9861, csa_tree_add_190_195_groupi_n_9862, csa_tree_add_190_195_groupi_n_9863, csa_tree_add_190_195_groupi_n_9864;
  wire csa_tree_add_190_195_groupi_n_9865, csa_tree_add_190_195_groupi_n_9866, csa_tree_add_190_195_groupi_n_9867, csa_tree_add_190_195_groupi_n_9868, csa_tree_add_190_195_groupi_n_9869, csa_tree_add_190_195_groupi_n_9870, csa_tree_add_190_195_groupi_n_9871, csa_tree_add_190_195_groupi_n_9872;
  wire csa_tree_add_190_195_groupi_n_9873, csa_tree_add_190_195_groupi_n_9874, csa_tree_add_190_195_groupi_n_9875, csa_tree_add_190_195_groupi_n_9876, csa_tree_add_190_195_groupi_n_9877, csa_tree_add_190_195_groupi_n_9878, csa_tree_add_190_195_groupi_n_9879, csa_tree_add_190_195_groupi_n_9880;
  wire csa_tree_add_190_195_groupi_n_9881, csa_tree_add_190_195_groupi_n_9882, csa_tree_add_190_195_groupi_n_9883, csa_tree_add_190_195_groupi_n_9884, csa_tree_add_190_195_groupi_n_9885, csa_tree_add_190_195_groupi_n_9886, csa_tree_add_190_195_groupi_n_9887, csa_tree_add_190_195_groupi_n_9888;
  wire csa_tree_add_190_195_groupi_n_9889, csa_tree_add_190_195_groupi_n_9890, csa_tree_add_190_195_groupi_n_9891, csa_tree_add_190_195_groupi_n_9892, csa_tree_add_190_195_groupi_n_9893, csa_tree_add_190_195_groupi_n_9894, csa_tree_add_190_195_groupi_n_9895, csa_tree_add_190_195_groupi_n_9896;
  wire csa_tree_add_190_195_groupi_n_9897, csa_tree_add_190_195_groupi_n_9898, csa_tree_add_190_195_groupi_n_9899, csa_tree_add_190_195_groupi_n_9900, csa_tree_add_190_195_groupi_n_9901, csa_tree_add_190_195_groupi_n_9902, csa_tree_add_190_195_groupi_n_9903, csa_tree_add_190_195_groupi_n_9904;
  wire csa_tree_add_190_195_groupi_n_9905, csa_tree_add_190_195_groupi_n_9906, csa_tree_add_190_195_groupi_n_9907, csa_tree_add_190_195_groupi_n_9908, csa_tree_add_190_195_groupi_n_9909, csa_tree_add_190_195_groupi_n_9910, csa_tree_add_190_195_groupi_n_9911, csa_tree_add_190_195_groupi_n_9912;
  wire csa_tree_add_190_195_groupi_n_9913, csa_tree_add_190_195_groupi_n_9914, csa_tree_add_190_195_groupi_n_9915, csa_tree_add_190_195_groupi_n_9916, csa_tree_add_190_195_groupi_n_9917, csa_tree_add_190_195_groupi_n_9918, csa_tree_add_190_195_groupi_n_9919, csa_tree_add_190_195_groupi_n_9920;
  wire csa_tree_add_190_195_groupi_n_9921, csa_tree_add_190_195_groupi_n_9922, csa_tree_add_190_195_groupi_n_9923, csa_tree_add_190_195_groupi_n_9924, csa_tree_add_190_195_groupi_n_9925, csa_tree_add_190_195_groupi_n_9926, csa_tree_add_190_195_groupi_n_9927, csa_tree_add_190_195_groupi_n_9928;
  wire csa_tree_add_190_195_groupi_n_9929, csa_tree_add_190_195_groupi_n_9930, csa_tree_add_190_195_groupi_n_9931, csa_tree_add_190_195_groupi_n_9932, csa_tree_add_190_195_groupi_n_9933, csa_tree_add_190_195_groupi_n_9934, csa_tree_add_190_195_groupi_n_9935, csa_tree_add_190_195_groupi_n_9936;
  wire csa_tree_add_190_195_groupi_n_9937, csa_tree_add_190_195_groupi_n_9938, csa_tree_add_190_195_groupi_n_9939, csa_tree_add_190_195_groupi_n_9940, csa_tree_add_190_195_groupi_n_9941, csa_tree_add_190_195_groupi_n_9942, csa_tree_add_190_195_groupi_n_9943, csa_tree_add_190_195_groupi_n_9944;
  wire csa_tree_add_190_195_groupi_n_9945, csa_tree_add_190_195_groupi_n_9946, csa_tree_add_190_195_groupi_n_9947, csa_tree_add_190_195_groupi_n_9948, csa_tree_add_190_195_groupi_n_9949, csa_tree_add_190_195_groupi_n_9950, csa_tree_add_190_195_groupi_n_9951, csa_tree_add_190_195_groupi_n_9952;
  wire csa_tree_add_190_195_groupi_n_9953, csa_tree_add_190_195_groupi_n_9954, csa_tree_add_190_195_groupi_n_9955, csa_tree_add_190_195_groupi_n_9956, csa_tree_add_190_195_groupi_n_9957, csa_tree_add_190_195_groupi_n_9958, csa_tree_add_190_195_groupi_n_9959, csa_tree_add_190_195_groupi_n_9960;
  wire csa_tree_add_190_195_groupi_n_9961, csa_tree_add_190_195_groupi_n_9962, csa_tree_add_190_195_groupi_n_9963, csa_tree_add_190_195_groupi_n_9964, csa_tree_add_190_195_groupi_n_9965, csa_tree_add_190_195_groupi_n_9966, csa_tree_add_190_195_groupi_n_9967, csa_tree_add_190_195_groupi_n_9968;
  wire csa_tree_add_190_195_groupi_n_9969, csa_tree_add_190_195_groupi_n_9970, csa_tree_add_190_195_groupi_n_9971, csa_tree_add_190_195_groupi_n_9972, csa_tree_add_190_195_groupi_n_9973, csa_tree_add_190_195_groupi_n_9974, csa_tree_add_190_195_groupi_n_9975, csa_tree_add_190_195_groupi_n_9976;
  wire csa_tree_add_190_195_groupi_n_9977, csa_tree_add_190_195_groupi_n_9978, csa_tree_add_190_195_groupi_n_9979, csa_tree_add_190_195_groupi_n_9980, csa_tree_add_190_195_groupi_n_9981, csa_tree_add_190_195_groupi_n_9982, csa_tree_add_190_195_groupi_n_9983, csa_tree_add_190_195_groupi_n_9984;
  wire csa_tree_add_190_195_groupi_n_9985, csa_tree_add_190_195_groupi_n_9986, csa_tree_add_190_195_groupi_n_9987, csa_tree_add_190_195_groupi_n_9988, csa_tree_add_190_195_groupi_n_9989, csa_tree_add_190_195_groupi_n_9990, csa_tree_add_190_195_groupi_n_9991, csa_tree_add_190_195_groupi_n_9992;
  wire csa_tree_add_190_195_groupi_n_9993, csa_tree_add_190_195_groupi_n_9994, csa_tree_add_190_195_groupi_n_9995, csa_tree_add_190_195_groupi_n_9996, csa_tree_add_190_195_groupi_n_9997, csa_tree_add_190_195_groupi_n_9998, csa_tree_add_190_195_groupi_n_9999, csa_tree_add_190_195_groupi_n_10000;
  wire csa_tree_add_190_195_groupi_n_10001, csa_tree_add_190_195_groupi_n_10002, csa_tree_add_190_195_groupi_n_10003, csa_tree_add_190_195_groupi_n_10004, csa_tree_add_190_195_groupi_n_10005, csa_tree_add_190_195_groupi_n_10006, csa_tree_add_190_195_groupi_n_10007, csa_tree_add_190_195_groupi_n_10008;
  wire csa_tree_add_190_195_groupi_n_10009, csa_tree_add_190_195_groupi_n_10010, csa_tree_add_190_195_groupi_n_10011, csa_tree_add_190_195_groupi_n_10012, csa_tree_add_190_195_groupi_n_10013, csa_tree_add_190_195_groupi_n_10014, csa_tree_add_190_195_groupi_n_10015, csa_tree_add_190_195_groupi_n_10016;
  wire csa_tree_add_190_195_groupi_n_10017, csa_tree_add_190_195_groupi_n_10018, csa_tree_add_190_195_groupi_n_10019, csa_tree_add_190_195_groupi_n_10020, csa_tree_add_190_195_groupi_n_10021, csa_tree_add_190_195_groupi_n_10022, csa_tree_add_190_195_groupi_n_10023, csa_tree_add_190_195_groupi_n_10024;
  wire csa_tree_add_190_195_groupi_n_10025, csa_tree_add_190_195_groupi_n_10026, csa_tree_add_190_195_groupi_n_10027, csa_tree_add_190_195_groupi_n_10028, csa_tree_add_190_195_groupi_n_10029, csa_tree_add_190_195_groupi_n_10030, csa_tree_add_190_195_groupi_n_10031, csa_tree_add_190_195_groupi_n_10032;
  wire csa_tree_add_190_195_groupi_n_10033, csa_tree_add_190_195_groupi_n_10034, csa_tree_add_190_195_groupi_n_10035, csa_tree_add_190_195_groupi_n_10036, csa_tree_add_190_195_groupi_n_10037, csa_tree_add_190_195_groupi_n_10038, csa_tree_add_190_195_groupi_n_10039, csa_tree_add_190_195_groupi_n_10040;
  wire csa_tree_add_190_195_groupi_n_10041, csa_tree_add_190_195_groupi_n_10042, csa_tree_add_190_195_groupi_n_10043, csa_tree_add_190_195_groupi_n_10044, csa_tree_add_190_195_groupi_n_10045, csa_tree_add_190_195_groupi_n_10046, csa_tree_add_190_195_groupi_n_10047, csa_tree_add_190_195_groupi_n_10048;
  wire csa_tree_add_190_195_groupi_n_10049, csa_tree_add_190_195_groupi_n_10050, csa_tree_add_190_195_groupi_n_10051, csa_tree_add_190_195_groupi_n_10052, csa_tree_add_190_195_groupi_n_10053, csa_tree_add_190_195_groupi_n_10054, csa_tree_add_190_195_groupi_n_10055, csa_tree_add_190_195_groupi_n_10056;
  wire csa_tree_add_190_195_groupi_n_10057, csa_tree_add_190_195_groupi_n_10058, csa_tree_add_190_195_groupi_n_10059, csa_tree_add_190_195_groupi_n_10060, csa_tree_add_190_195_groupi_n_10061, csa_tree_add_190_195_groupi_n_10062, csa_tree_add_190_195_groupi_n_10063, csa_tree_add_190_195_groupi_n_10064;
  wire csa_tree_add_190_195_groupi_n_10065, csa_tree_add_190_195_groupi_n_10066, csa_tree_add_190_195_groupi_n_10067, csa_tree_add_190_195_groupi_n_10068, csa_tree_add_190_195_groupi_n_10069, csa_tree_add_190_195_groupi_n_10070, csa_tree_add_190_195_groupi_n_10071, csa_tree_add_190_195_groupi_n_10072;
  wire csa_tree_add_190_195_groupi_n_10073, csa_tree_add_190_195_groupi_n_10074, csa_tree_add_190_195_groupi_n_10075, csa_tree_add_190_195_groupi_n_10076, csa_tree_add_190_195_groupi_n_10077, csa_tree_add_190_195_groupi_n_10078, csa_tree_add_190_195_groupi_n_10079, csa_tree_add_190_195_groupi_n_10080;
  wire csa_tree_add_190_195_groupi_n_10081, csa_tree_add_190_195_groupi_n_10082, csa_tree_add_190_195_groupi_n_10083, csa_tree_add_190_195_groupi_n_10084, csa_tree_add_190_195_groupi_n_10085, csa_tree_add_190_195_groupi_n_10086, csa_tree_add_190_195_groupi_n_10087, csa_tree_add_190_195_groupi_n_10088;
  wire csa_tree_add_190_195_groupi_n_10089, csa_tree_add_190_195_groupi_n_10090, csa_tree_add_190_195_groupi_n_10091, csa_tree_add_190_195_groupi_n_10092, csa_tree_add_190_195_groupi_n_10093, csa_tree_add_190_195_groupi_n_10094, csa_tree_add_190_195_groupi_n_10095, csa_tree_add_190_195_groupi_n_10096;
  wire csa_tree_add_190_195_groupi_n_10097, csa_tree_add_190_195_groupi_n_10098, csa_tree_add_190_195_groupi_n_10099, csa_tree_add_190_195_groupi_n_10100, csa_tree_add_190_195_groupi_n_10101, csa_tree_add_190_195_groupi_n_10102, csa_tree_add_190_195_groupi_n_10103, csa_tree_add_190_195_groupi_n_10104;
  wire csa_tree_add_190_195_groupi_n_10105, csa_tree_add_190_195_groupi_n_10106, csa_tree_add_190_195_groupi_n_10107, csa_tree_add_190_195_groupi_n_10108, csa_tree_add_190_195_groupi_n_10109, csa_tree_add_190_195_groupi_n_10110, csa_tree_add_190_195_groupi_n_10111, csa_tree_add_190_195_groupi_n_10112;
  wire csa_tree_add_190_195_groupi_n_10113, csa_tree_add_190_195_groupi_n_10114, csa_tree_add_190_195_groupi_n_10115, csa_tree_add_190_195_groupi_n_10117, csa_tree_add_190_195_groupi_n_10118, csa_tree_add_190_195_groupi_n_10119, csa_tree_add_190_195_groupi_n_10120, csa_tree_add_190_195_groupi_n_10121;
  wire csa_tree_add_190_195_groupi_n_10122, csa_tree_add_190_195_groupi_n_10123, csa_tree_add_190_195_groupi_n_10124, csa_tree_add_190_195_groupi_n_10125, csa_tree_add_190_195_groupi_n_10126, csa_tree_add_190_195_groupi_n_10127, csa_tree_add_190_195_groupi_n_10128, csa_tree_add_190_195_groupi_n_10129;
  wire csa_tree_add_190_195_groupi_n_10130, csa_tree_add_190_195_groupi_n_10131, csa_tree_add_190_195_groupi_n_10132, csa_tree_add_190_195_groupi_n_10133, csa_tree_add_190_195_groupi_n_10134, csa_tree_add_190_195_groupi_n_10135, csa_tree_add_190_195_groupi_n_10136, csa_tree_add_190_195_groupi_n_10137;
  wire csa_tree_add_190_195_groupi_n_10138, csa_tree_add_190_195_groupi_n_10139, csa_tree_add_190_195_groupi_n_10140, csa_tree_add_190_195_groupi_n_10141, csa_tree_add_190_195_groupi_n_10142, csa_tree_add_190_195_groupi_n_10143, csa_tree_add_190_195_groupi_n_10144, csa_tree_add_190_195_groupi_n_10145;
  wire csa_tree_add_190_195_groupi_n_10146, csa_tree_add_190_195_groupi_n_10147, csa_tree_add_190_195_groupi_n_10148, csa_tree_add_190_195_groupi_n_10149, csa_tree_add_190_195_groupi_n_10150, csa_tree_add_190_195_groupi_n_10151, csa_tree_add_190_195_groupi_n_10152, csa_tree_add_190_195_groupi_n_10153;
  wire csa_tree_add_190_195_groupi_n_10154, csa_tree_add_190_195_groupi_n_10155, csa_tree_add_190_195_groupi_n_10156, csa_tree_add_190_195_groupi_n_10157, csa_tree_add_190_195_groupi_n_10158, csa_tree_add_190_195_groupi_n_10159, csa_tree_add_190_195_groupi_n_10160, csa_tree_add_190_195_groupi_n_10161;
  wire csa_tree_add_190_195_groupi_n_10162, csa_tree_add_190_195_groupi_n_10163, csa_tree_add_190_195_groupi_n_10164, csa_tree_add_190_195_groupi_n_10165, csa_tree_add_190_195_groupi_n_10166, csa_tree_add_190_195_groupi_n_10167, csa_tree_add_190_195_groupi_n_10168, csa_tree_add_190_195_groupi_n_10169;
  wire csa_tree_add_190_195_groupi_n_10170, csa_tree_add_190_195_groupi_n_10171, csa_tree_add_190_195_groupi_n_10172, csa_tree_add_190_195_groupi_n_10173, csa_tree_add_190_195_groupi_n_10174, csa_tree_add_190_195_groupi_n_10175, csa_tree_add_190_195_groupi_n_10176, csa_tree_add_190_195_groupi_n_10177;
  wire csa_tree_add_190_195_groupi_n_10178, csa_tree_add_190_195_groupi_n_10179, csa_tree_add_190_195_groupi_n_10180, csa_tree_add_190_195_groupi_n_10181, csa_tree_add_190_195_groupi_n_10182, csa_tree_add_190_195_groupi_n_10183, csa_tree_add_190_195_groupi_n_10184, csa_tree_add_190_195_groupi_n_10185;
  wire csa_tree_add_190_195_groupi_n_10186, csa_tree_add_190_195_groupi_n_10187, csa_tree_add_190_195_groupi_n_10188, csa_tree_add_190_195_groupi_n_10189, csa_tree_add_190_195_groupi_n_10190, csa_tree_add_190_195_groupi_n_10191, csa_tree_add_190_195_groupi_n_10192, csa_tree_add_190_195_groupi_n_10193;
  wire csa_tree_add_190_195_groupi_n_10194, csa_tree_add_190_195_groupi_n_10195, csa_tree_add_190_195_groupi_n_10196, csa_tree_add_190_195_groupi_n_10197, csa_tree_add_190_195_groupi_n_10198, csa_tree_add_190_195_groupi_n_10199, csa_tree_add_190_195_groupi_n_10200, csa_tree_add_190_195_groupi_n_10201;
  wire csa_tree_add_190_195_groupi_n_10202, csa_tree_add_190_195_groupi_n_10203, csa_tree_add_190_195_groupi_n_10204, csa_tree_add_190_195_groupi_n_10205, csa_tree_add_190_195_groupi_n_10206, csa_tree_add_190_195_groupi_n_10207, csa_tree_add_190_195_groupi_n_10208, csa_tree_add_190_195_groupi_n_10209;
  wire csa_tree_add_190_195_groupi_n_10210, csa_tree_add_190_195_groupi_n_10211, csa_tree_add_190_195_groupi_n_10212, csa_tree_add_190_195_groupi_n_10213, csa_tree_add_190_195_groupi_n_10214, csa_tree_add_190_195_groupi_n_10215, csa_tree_add_190_195_groupi_n_10216, csa_tree_add_190_195_groupi_n_10217;
  wire csa_tree_add_190_195_groupi_n_10218, csa_tree_add_190_195_groupi_n_10219, csa_tree_add_190_195_groupi_n_10220, csa_tree_add_190_195_groupi_n_10221, csa_tree_add_190_195_groupi_n_10222, csa_tree_add_190_195_groupi_n_10223, csa_tree_add_190_195_groupi_n_10224, csa_tree_add_190_195_groupi_n_10225;
  wire csa_tree_add_190_195_groupi_n_10226, csa_tree_add_190_195_groupi_n_10227, csa_tree_add_190_195_groupi_n_10228, csa_tree_add_190_195_groupi_n_10229, csa_tree_add_190_195_groupi_n_10230, csa_tree_add_190_195_groupi_n_10231, csa_tree_add_190_195_groupi_n_10232, csa_tree_add_190_195_groupi_n_10233;
  wire csa_tree_add_190_195_groupi_n_10234, csa_tree_add_190_195_groupi_n_10235, csa_tree_add_190_195_groupi_n_10236, csa_tree_add_190_195_groupi_n_10237, csa_tree_add_190_195_groupi_n_10238, csa_tree_add_190_195_groupi_n_10239, csa_tree_add_190_195_groupi_n_10240, csa_tree_add_190_195_groupi_n_10241;
  wire csa_tree_add_190_195_groupi_n_10242, csa_tree_add_190_195_groupi_n_10243, csa_tree_add_190_195_groupi_n_10244, csa_tree_add_190_195_groupi_n_10245, csa_tree_add_190_195_groupi_n_10246, csa_tree_add_190_195_groupi_n_10247, csa_tree_add_190_195_groupi_n_10248, csa_tree_add_190_195_groupi_n_10249;
  wire csa_tree_add_190_195_groupi_n_10250, csa_tree_add_190_195_groupi_n_10251, csa_tree_add_190_195_groupi_n_10252, csa_tree_add_190_195_groupi_n_10253, csa_tree_add_190_195_groupi_n_10254, csa_tree_add_190_195_groupi_n_10255, csa_tree_add_190_195_groupi_n_10256, csa_tree_add_190_195_groupi_n_10257;
  wire csa_tree_add_190_195_groupi_n_10258, csa_tree_add_190_195_groupi_n_10259, csa_tree_add_190_195_groupi_n_10260, csa_tree_add_190_195_groupi_n_10261, csa_tree_add_190_195_groupi_n_10262, csa_tree_add_190_195_groupi_n_10263, csa_tree_add_190_195_groupi_n_10264, csa_tree_add_190_195_groupi_n_10265;
  wire csa_tree_add_190_195_groupi_n_10266, csa_tree_add_190_195_groupi_n_10267, csa_tree_add_190_195_groupi_n_10268, csa_tree_add_190_195_groupi_n_10269, csa_tree_add_190_195_groupi_n_10270, csa_tree_add_190_195_groupi_n_10271, csa_tree_add_190_195_groupi_n_10272, csa_tree_add_190_195_groupi_n_10273;
  wire csa_tree_add_190_195_groupi_n_10274, csa_tree_add_190_195_groupi_n_10275, csa_tree_add_190_195_groupi_n_10276, csa_tree_add_190_195_groupi_n_10277, csa_tree_add_190_195_groupi_n_10278, csa_tree_add_190_195_groupi_n_10279, csa_tree_add_190_195_groupi_n_10280, csa_tree_add_190_195_groupi_n_10281;
  wire csa_tree_add_190_195_groupi_n_10282, csa_tree_add_190_195_groupi_n_10283, csa_tree_add_190_195_groupi_n_10284, csa_tree_add_190_195_groupi_n_10285, csa_tree_add_190_195_groupi_n_10286, csa_tree_add_190_195_groupi_n_10287, csa_tree_add_190_195_groupi_n_10288, csa_tree_add_190_195_groupi_n_10289;
  wire csa_tree_add_190_195_groupi_n_10290, csa_tree_add_190_195_groupi_n_10291, csa_tree_add_190_195_groupi_n_10292, csa_tree_add_190_195_groupi_n_10293, csa_tree_add_190_195_groupi_n_10294, csa_tree_add_190_195_groupi_n_10295, csa_tree_add_190_195_groupi_n_10296, csa_tree_add_190_195_groupi_n_10297;
  wire csa_tree_add_190_195_groupi_n_10298, csa_tree_add_190_195_groupi_n_10299, csa_tree_add_190_195_groupi_n_10300, csa_tree_add_190_195_groupi_n_10301, csa_tree_add_190_195_groupi_n_10302, csa_tree_add_190_195_groupi_n_10303, csa_tree_add_190_195_groupi_n_10304, csa_tree_add_190_195_groupi_n_10305;
  wire csa_tree_add_190_195_groupi_n_10306, csa_tree_add_190_195_groupi_n_10307, csa_tree_add_190_195_groupi_n_10308, csa_tree_add_190_195_groupi_n_10309, csa_tree_add_190_195_groupi_n_10310, csa_tree_add_190_195_groupi_n_10311, csa_tree_add_190_195_groupi_n_10312, csa_tree_add_190_195_groupi_n_10313;
  wire csa_tree_add_190_195_groupi_n_10314, csa_tree_add_190_195_groupi_n_10315, csa_tree_add_190_195_groupi_n_10316, csa_tree_add_190_195_groupi_n_10317, csa_tree_add_190_195_groupi_n_10318, csa_tree_add_190_195_groupi_n_10319, csa_tree_add_190_195_groupi_n_10320, csa_tree_add_190_195_groupi_n_10321;
  wire csa_tree_add_190_195_groupi_n_10322, csa_tree_add_190_195_groupi_n_10323, csa_tree_add_190_195_groupi_n_10324, csa_tree_add_190_195_groupi_n_10325, csa_tree_add_190_195_groupi_n_10326, csa_tree_add_190_195_groupi_n_10327, csa_tree_add_190_195_groupi_n_10328, csa_tree_add_190_195_groupi_n_10329;
  wire csa_tree_add_190_195_groupi_n_10330, csa_tree_add_190_195_groupi_n_10331, csa_tree_add_190_195_groupi_n_10332, csa_tree_add_190_195_groupi_n_10333, csa_tree_add_190_195_groupi_n_10334, csa_tree_add_190_195_groupi_n_10335, csa_tree_add_190_195_groupi_n_10336, csa_tree_add_190_195_groupi_n_10337;
  wire csa_tree_add_190_195_groupi_n_10338, csa_tree_add_190_195_groupi_n_10339, csa_tree_add_190_195_groupi_n_10340, csa_tree_add_190_195_groupi_n_10341, csa_tree_add_190_195_groupi_n_10342, csa_tree_add_190_195_groupi_n_10343, csa_tree_add_190_195_groupi_n_10344, csa_tree_add_190_195_groupi_n_10345;
  wire csa_tree_add_190_195_groupi_n_10346, csa_tree_add_190_195_groupi_n_10347, csa_tree_add_190_195_groupi_n_10348, csa_tree_add_190_195_groupi_n_10349, csa_tree_add_190_195_groupi_n_10350, csa_tree_add_190_195_groupi_n_10351, csa_tree_add_190_195_groupi_n_10352, csa_tree_add_190_195_groupi_n_10353;
  wire csa_tree_add_190_195_groupi_n_10354, csa_tree_add_190_195_groupi_n_10355, csa_tree_add_190_195_groupi_n_10356, csa_tree_add_190_195_groupi_n_10357, csa_tree_add_190_195_groupi_n_10358, csa_tree_add_190_195_groupi_n_10359, csa_tree_add_190_195_groupi_n_10360, csa_tree_add_190_195_groupi_n_10361;
  wire csa_tree_add_190_195_groupi_n_10362, csa_tree_add_190_195_groupi_n_10363, csa_tree_add_190_195_groupi_n_10364, csa_tree_add_190_195_groupi_n_10365, csa_tree_add_190_195_groupi_n_10366, csa_tree_add_190_195_groupi_n_10367, csa_tree_add_190_195_groupi_n_10368, csa_tree_add_190_195_groupi_n_10369;
  wire csa_tree_add_190_195_groupi_n_10370, csa_tree_add_190_195_groupi_n_10371, csa_tree_add_190_195_groupi_n_10372, csa_tree_add_190_195_groupi_n_10373, csa_tree_add_190_195_groupi_n_10374, csa_tree_add_190_195_groupi_n_10375, csa_tree_add_190_195_groupi_n_10376, csa_tree_add_190_195_groupi_n_10377;
  wire csa_tree_add_190_195_groupi_n_10378, csa_tree_add_190_195_groupi_n_10379, csa_tree_add_190_195_groupi_n_10380, csa_tree_add_190_195_groupi_n_10381, csa_tree_add_190_195_groupi_n_10382, csa_tree_add_190_195_groupi_n_10383, csa_tree_add_190_195_groupi_n_10384, csa_tree_add_190_195_groupi_n_10385;
  wire csa_tree_add_190_195_groupi_n_10386, csa_tree_add_190_195_groupi_n_10387, csa_tree_add_190_195_groupi_n_10388, csa_tree_add_190_195_groupi_n_10389, csa_tree_add_190_195_groupi_n_10390, csa_tree_add_190_195_groupi_n_10391, csa_tree_add_190_195_groupi_n_10392, csa_tree_add_190_195_groupi_n_10393;
  wire csa_tree_add_190_195_groupi_n_10394, csa_tree_add_190_195_groupi_n_10395, csa_tree_add_190_195_groupi_n_10396, csa_tree_add_190_195_groupi_n_10397, csa_tree_add_190_195_groupi_n_10398, csa_tree_add_190_195_groupi_n_10399, csa_tree_add_190_195_groupi_n_10400, csa_tree_add_190_195_groupi_n_10401;
  wire csa_tree_add_190_195_groupi_n_10402, csa_tree_add_190_195_groupi_n_10403, csa_tree_add_190_195_groupi_n_10404, csa_tree_add_190_195_groupi_n_10405, csa_tree_add_190_195_groupi_n_10406, csa_tree_add_190_195_groupi_n_10407, csa_tree_add_190_195_groupi_n_10408, csa_tree_add_190_195_groupi_n_10409;
  wire csa_tree_add_190_195_groupi_n_10410, csa_tree_add_190_195_groupi_n_10411, csa_tree_add_190_195_groupi_n_10412, csa_tree_add_190_195_groupi_n_10413, csa_tree_add_190_195_groupi_n_10414, csa_tree_add_190_195_groupi_n_10415, csa_tree_add_190_195_groupi_n_10416, csa_tree_add_190_195_groupi_n_10417;
  wire csa_tree_add_190_195_groupi_n_10418, csa_tree_add_190_195_groupi_n_10419, csa_tree_add_190_195_groupi_n_10420, csa_tree_add_190_195_groupi_n_10421, csa_tree_add_190_195_groupi_n_10422, csa_tree_add_190_195_groupi_n_10423, csa_tree_add_190_195_groupi_n_10424, csa_tree_add_190_195_groupi_n_10425;
  wire csa_tree_add_190_195_groupi_n_10426, csa_tree_add_190_195_groupi_n_10427, csa_tree_add_190_195_groupi_n_10428, csa_tree_add_190_195_groupi_n_10429, csa_tree_add_190_195_groupi_n_10430, csa_tree_add_190_195_groupi_n_10431, csa_tree_add_190_195_groupi_n_10432, csa_tree_add_190_195_groupi_n_10433;
  wire csa_tree_add_190_195_groupi_n_10434, csa_tree_add_190_195_groupi_n_10435, csa_tree_add_190_195_groupi_n_10436, csa_tree_add_190_195_groupi_n_10437, csa_tree_add_190_195_groupi_n_10438, csa_tree_add_190_195_groupi_n_10439, csa_tree_add_190_195_groupi_n_10440, csa_tree_add_190_195_groupi_n_10441;
  wire csa_tree_add_190_195_groupi_n_10442, csa_tree_add_190_195_groupi_n_10443, csa_tree_add_190_195_groupi_n_10444, csa_tree_add_190_195_groupi_n_10445, csa_tree_add_190_195_groupi_n_10446, csa_tree_add_190_195_groupi_n_10447, csa_tree_add_190_195_groupi_n_10448, csa_tree_add_190_195_groupi_n_10449;
  wire csa_tree_add_190_195_groupi_n_10450, csa_tree_add_190_195_groupi_n_10451, csa_tree_add_190_195_groupi_n_10452, csa_tree_add_190_195_groupi_n_10453, csa_tree_add_190_195_groupi_n_10454, csa_tree_add_190_195_groupi_n_10455, csa_tree_add_190_195_groupi_n_10456, csa_tree_add_190_195_groupi_n_10457;
  wire csa_tree_add_190_195_groupi_n_10458, csa_tree_add_190_195_groupi_n_10459, csa_tree_add_190_195_groupi_n_10460, csa_tree_add_190_195_groupi_n_10461, csa_tree_add_190_195_groupi_n_10462, csa_tree_add_190_195_groupi_n_10463, csa_tree_add_190_195_groupi_n_10464, csa_tree_add_190_195_groupi_n_10465;
  wire csa_tree_add_190_195_groupi_n_10466, csa_tree_add_190_195_groupi_n_10467, csa_tree_add_190_195_groupi_n_10468, csa_tree_add_190_195_groupi_n_10469, csa_tree_add_190_195_groupi_n_10470, csa_tree_add_190_195_groupi_n_10471, csa_tree_add_190_195_groupi_n_10472, csa_tree_add_190_195_groupi_n_10473;
  wire csa_tree_add_190_195_groupi_n_10474, csa_tree_add_190_195_groupi_n_10475, csa_tree_add_190_195_groupi_n_10476, csa_tree_add_190_195_groupi_n_10477, csa_tree_add_190_195_groupi_n_10478, csa_tree_add_190_195_groupi_n_10479, csa_tree_add_190_195_groupi_n_10480, csa_tree_add_190_195_groupi_n_10481;
  wire csa_tree_add_190_195_groupi_n_10482, csa_tree_add_190_195_groupi_n_10483, csa_tree_add_190_195_groupi_n_10484, csa_tree_add_190_195_groupi_n_10485, csa_tree_add_190_195_groupi_n_10486, csa_tree_add_190_195_groupi_n_10487, csa_tree_add_190_195_groupi_n_10488, csa_tree_add_190_195_groupi_n_10489;
  wire csa_tree_add_190_195_groupi_n_10490, csa_tree_add_190_195_groupi_n_10491, csa_tree_add_190_195_groupi_n_10492, csa_tree_add_190_195_groupi_n_10493, csa_tree_add_190_195_groupi_n_10494, csa_tree_add_190_195_groupi_n_10495, csa_tree_add_190_195_groupi_n_10496, csa_tree_add_190_195_groupi_n_10497;
  wire csa_tree_add_190_195_groupi_n_10498, csa_tree_add_190_195_groupi_n_10499, csa_tree_add_190_195_groupi_n_10500, csa_tree_add_190_195_groupi_n_10501, csa_tree_add_190_195_groupi_n_10502, csa_tree_add_190_195_groupi_n_10503, csa_tree_add_190_195_groupi_n_10504, csa_tree_add_190_195_groupi_n_10505;
  wire csa_tree_add_190_195_groupi_n_10506, csa_tree_add_190_195_groupi_n_10507, csa_tree_add_190_195_groupi_n_10508, csa_tree_add_190_195_groupi_n_10509, csa_tree_add_190_195_groupi_n_10510, csa_tree_add_190_195_groupi_n_10511, csa_tree_add_190_195_groupi_n_10512, csa_tree_add_190_195_groupi_n_10513;
  wire csa_tree_add_190_195_groupi_n_10514, csa_tree_add_190_195_groupi_n_10515, csa_tree_add_190_195_groupi_n_10516, csa_tree_add_190_195_groupi_n_10517, csa_tree_add_190_195_groupi_n_10518, csa_tree_add_190_195_groupi_n_10519, csa_tree_add_190_195_groupi_n_10520, csa_tree_add_190_195_groupi_n_10521;
  wire csa_tree_add_190_195_groupi_n_10522, csa_tree_add_190_195_groupi_n_10523, csa_tree_add_190_195_groupi_n_10524, csa_tree_add_190_195_groupi_n_10525, csa_tree_add_190_195_groupi_n_10526, csa_tree_add_190_195_groupi_n_10527, csa_tree_add_190_195_groupi_n_10528, csa_tree_add_190_195_groupi_n_10529;
  wire csa_tree_add_190_195_groupi_n_10530, csa_tree_add_190_195_groupi_n_10531, csa_tree_add_190_195_groupi_n_10532, csa_tree_add_190_195_groupi_n_10533, csa_tree_add_190_195_groupi_n_10534, csa_tree_add_190_195_groupi_n_10535, csa_tree_add_190_195_groupi_n_10536, csa_tree_add_190_195_groupi_n_10537;
  wire csa_tree_add_190_195_groupi_n_10538, csa_tree_add_190_195_groupi_n_10539, csa_tree_add_190_195_groupi_n_10540, csa_tree_add_190_195_groupi_n_10541, csa_tree_add_190_195_groupi_n_10542, csa_tree_add_190_195_groupi_n_10543, csa_tree_add_190_195_groupi_n_10544, csa_tree_add_190_195_groupi_n_10545;
  wire csa_tree_add_190_195_groupi_n_10546, csa_tree_add_190_195_groupi_n_10547, csa_tree_add_190_195_groupi_n_10548, csa_tree_add_190_195_groupi_n_10549, csa_tree_add_190_195_groupi_n_10550, csa_tree_add_190_195_groupi_n_10551, csa_tree_add_190_195_groupi_n_10552, csa_tree_add_190_195_groupi_n_10553;
  wire csa_tree_add_190_195_groupi_n_10554, csa_tree_add_190_195_groupi_n_10555, csa_tree_add_190_195_groupi_n_10556, csa_tree_add_190_195_groupi_n_10557, csa_tree_add_190_195_groupi_n_10558, csa_tree_add_190_195_groupi_n_10559, csa_tree_add_190_195_groupi_n_10560, csa_tree_add_190_195_groupi_n_10561;
  wire csa_tree_add_190_195_groupi_n_10562, csa_tree_add_190_195_groupi_n_10563, csa_tree_add_190_195_groupi_n_10564, csa_tree_add_190_195_groupi_n_10565, csa_tree_add_190_195_groupi_n_10566, csa_tree_add_190_195_groupi_n_10567, csa_tree_add_190_195_groupi_n_10568, csa_tree_add_190_195_groupi_n_10569;
  wire csa_tree_add_190_195_groupi_n_10570, csa_tree_add_190_195_groupi_n_10571, csa_tree_add_190_195_groupi_n_10572, csa_tree_add_190_195_groupi_n_10573, csa_tree_add_190_195_groupi_n_10574, csa_tree_add_190_195_groupi_n_10575, csa_tree_add_190_195_groupi_n_10576, csa_tree_add_190_195_groupi_n_10577;
  wire csa_tree_add_190_195_groupi_n_10578, csa_tree_add_190_195_groupi_n_10579, csa_tree_add_190_195_groupi_n_10580, csa_tree_add_190_195_groupi_n_10581, csa_tree_add_190_195_groupi_n_10582, csa_tree_add_190_195_groupi_n_10583, csa_tree_add_190_195_groupi_n_10584, csa_tree_add_190_195_groupi_n_10585;
  wire csa_tree_add_190_195_groupi_n_10586, csa_tree_add_190_195_groupi_n_10587, csa_tree_add_190_195_groupi_n_10588, csa_tree_add_190_195_groupi_n_10589, csa_tree_add_190_195_groupi_n_10590, csa_tree_add_190_195_groupi_n_10591, csa_tree_add_190_195_groupi_n_10592, csa_tree_add_190_195_groupi_n_10593;
  wire csa_tree_add_190_195_groupi_n_10594, csa_tree_add_190_195_groupi_n_10595, csa_tree_add_190_195_groupi_n_10596, csa_tree_add_190_195_groupi_n_10597, csa_tree_add_190_195_groupi_n_10598, csa_tree_add_190_195_groupi_n_10599, csa_tree_add_190_195_groupi_n_10600, csa_tree_add_190_195_groupi_n_10601;
  wire csa_tree_add_190_195_groupi_n_10602, csa_tree_add_190_195_groupi_n_10603, csa_tree_add_190_195_groupi_n_10604, csa_tree_add_190_195_groupi_n_10605, csa_tree_add_190_195_groupi_n_10606, csa_tree_add_190_195_groupi_n_10607, csa_tree_add_190_195_groupi_n_10608, csa_tree_add_190_195_groupi_n_10609;
  wire csa_tree_add_190_195_groupi_n_10610, csa_tree_add_190_195_groupi_n_10611, csa_tree_add_190_195_groupi_n_10612, csa_tree_add_190_195_groupi_n_10613, csa_tree_add_190_195_groupi_n_10614, csa_tree_add_190_195_groupi_n_10615, csa_tree_add_190_195_groupi_n_10616, csa_tree_add_190_195_groupi_n_10617;
  wire csa_tree_add_190_195_groupi_n_10618, csa_tree_add_190_195_groupi_n_10619, csa_tree_add_190_195_groupi_n_10620, csa_tree_add_190_195_groupi_n_10621, csa_tree_add_190_195_groupi_n_10622, csa_tree_add_190_195_groupi_n_10623, csa_tree_add_190_195_groupi_n_10624, csa_tree_add_190_195_groupi_n_10625;
  wire csa_tree_add_190_195_groupi_n_10626, csa_tree_add_190_195_groupi_n_10627, csa_tree_add_190_195_groupi_n_10628, csa_tree_add_190_195_groupi_n_10629, csa_tree_add_190_195_groupi_n_10630, csa_tree_add_190_195_groupi_n_10631, csa_tree_add_190_195_groupi_n_10632, csa_tree_add_190_195_groupi_n_10633;
  wire csa_tree_add_190_195_groupi_n_10634, csa_tree_add_190_195_groupi_n_10635, csa_tree_add_190_195_groupi_n_10636, csa_tree_add_190_195_groupi_n_10637, csa_tree_add_190_195_groupi_n_10638, csa_tree_add_190_195_groupi_n_10639, csa_tree_add_190_195_groupi_n_10640, csa_tree_add_190_195_groupi_n_10641;
  wire csa_tree_add_190_195_groupi_n_10642, csa_tree_add_190_195_groupi_n_10643, csa_tree_add_190_195_groupi_n_10644, csa_tree_add_190_195_groupi_n_10645, csa_tree_add_190_195_groupi_n_10646, csa_tree_add_190_195_groupi_n_10647, csa_tree_add_190_195_groupi_n_10648, csa_tree_add_190_195_groupi_n_10649;
  wire csa_tree_add_190_195_groupi_n_10650, csa_tree_add_190_195_groupi_n_10651, csa_tree_add_190_195_groupi_n_10652, csa_tree_add_190_195_groupi_n_10653, csa_tree_add_190_195_groupi_n_10654, csa_tree_add_190_195_groupi_n_10655, csa_tree_add_190_195_groupi_n_10656, csa_tree_add_190_195_groupi_n_10657;
  wire csa_tree_add_190_195_groupi_n_10658, csa_tree_add_190_195_groupi_n_10659, csa_tree_add_190_195_groupi_n_10660, csa_tree_add_190_195_groupi_n_10661, csa_tree_add_190_195_groupi_n_10662, csa_tree_add_190_195_groupi_n_10663, csa_tree_add_190_195_groupi_n_10664, csa_tree_add_190_195_groupi_n_10665;
  wire csa_tree_add_190_195_groupi_n_10666, csa_tree_add_190_195_groupi_n_10667, csa_tree_add_190_195_groupi_n_10668, csa_tree_add_190_195_groupi_n_10669, csa_tree_add_190_195_groupi_n_10670, csa_tree_add_190_195_groupi_n_10671, csa_tree_add_190_195_groupi_n_10672, csa_tree_add_190_195_groupi_n_10673;
  wire csa_tree_add_190_195_groupi_n_10674, csa_tree_add_190_195_groupi_n_10675, csa_tree_add_190_195_groupi_n_10676, csa_tree_add_190_195_groupi_n_10677, csa_tree_add_190_195_groupi_n_10678, csa_tree_add_190_195_groupi_n_10679, csa_tree_add_190_195_groupi_n_10680, csa_tree_add_190_195_groupi_n_10681;
  wire csa_tree_add_190_195_groupi_n_10682, csa_tree_add_190_195_groupi_n_10683, csa_tree_add_190_195_groupi_n_10684, csa_tree_add_190_195_groupi_n_10685, csa_tree_add_190_195_groupi_n_10686, csa_tree_add_190_195_groupi_n_10687, csa_tree_add_190_195_groupi_n_10688, csa_tree_add_190_195_groupi_n_10689;
  wire csa_tree_add_190_195_groupi_n_10690, csa_tree_add_190_195_groupi_n_10691, csa_tree_add_190_195_groupi_n_10692, csa_tree_add_190_195_groupi_n_10693, csa_tree_add_190_195_groupi_n_10694, csa_tree_add_190_195_groupi_n_10695, csa_tree_add_190_195_groupi_n_10696, csa_tree_add_190_195_groupi_n_10697;
  wire csa_tree_add_190_195_groupi_n_10698, csa_tree_add_190_195_groupi_n_10699, csa_tree_add_190_195_groupi_n_10700, csa_tree_add_190_195_groupi_n_10701, csa_tree_add_190_195_groupi_n_10702, csa_tree_add_190_195_groupi_n_10703, csa_tree_add_190_195_groupi_n_10704, csa_tree_add_190_195_groupi_n_10705;
  wire csa_tree_add_190_195_groupi_n_10706, csa_tree_add_190_195_groupi_n_10707, csa_tree_add_190_195_groupi_n_10708, csa_tree_add_190_195_groupi_n_10709, csa_tree_add_190_195_groupi_n_10710, csa_tree_add_190_195_groupi_n_10711, csa_tree_add_190_195_groupi_n_10712, csa_tree_add_190_195_groupi_n_10713;
  wire csa_tree_add_190_195_groupi_n_10714, csa_tree_add_190_195_groupi_n_10715, csa_tree_add_190_195_groupi_n_10716, csa_tree_add_190_195_groupi_n_10717, csa_tree_add_190_195_groupi_n_10718, csa_tree_add_190_195_groupi_n_10719, csa_tree_add_190_195_groupi_n_10720, csa_tree_add_190_195_groupi_n_10721;
  wire csa_tree_add_190_195_groupi_n_10722, csa_tree_add_190_195_groupi_n_10723, csa_tree_add_190_195_groupi_n_10724, csa_tree_add_190_195_groupi_n_10725, csa_tree_add_190_195_groupi_n_10726, csa_tree_add_190_195_groupi_n_10727, csa_tree_add_190_195_groupi_n_10728, csa_tree_add_190_195_groupi_n_10729;
  wire csa_tree_add_190_195_groupi_n_10730, csa_tree_add_190_195_groupi_n_10731, csa_tree_add_190_195_groupi_n_10732, csa_tree_add_190_195_groupi_n_10733, csa_tree_add_190_195_groupi_n_10734, csa_tree_add_190_195_groupi_n_10735, csa_tree_add_190_195_groupi_n_10736, csa_tree_add_190_195_groupi_n_10737;
  wire csa_tree_add_190_195_groupi_n_10738, csa_tree_add_190_195_groupi_n_10739, csa_tree_add_190_195_groupi_n_10740, csa_tree_add_190_195_groupi_n_10741, csa_tree_add_190_195_groupi_n_10742, csa_tree_add_190_195_groupi_n_10743, csa_tree_add_190_195_groupi_n_10744, csa_tree_add_190_195_groupi_n_10745;
  wire csa_tree_add_190_195_groupi_n_10746, csa_tree_add_190_195_groupi_n_10747, csa_tree_add_190_195_groupi_n_10748, csa_tree_add_190_195_groupi_n_10749, csa_tree_add_190_195_groupi_n_10750, csa_tree_add_190_195_groupi_n_10751, csa_tree_add_190_195_groupi_n_10752, csa_tree_add_190_195_groupi_n_10753;
  wire csa_tree_add_190_195_groupi_n_10754, csa_tree_add_190_195_groupi_n_10755, csa_tree_add_190_195_groupi_n_10756, csa_tree_add_190_195_groupi_n_10757, csa_tree_add_190_195_groupi_n_10758, csa_tree_add_190_195_groupi_n_10759, csa_tree_add_190_195_groupi_n_10760, csa_tree_add_190_195_groupi_n_10761;
  wire csa_tree_add_190_195_groupi_n_10762, csa_tree_add_190_195_groupi_n_10763, csa_tree_add_190_195_groupi_n_10764, csa_tree_add_190_195_groupi_n_10765, csa_tree_add_190_195_groupi_n_10766, csa_tree_add_190_195_groupi_n_10767, csa_tree_add_190_195_groupi_n_10768, csa_tree_add_190_195_groupi_n_10769;
  wire csa_tree_add_190_195_groupi_n_10770, csa_tree_add_190_195_groupi_n_10771, csa_tree_add_190_195_groupi_n_10772, csa_tree_add_190_195_groupi_n_10773, csa_tree_add_190_195_groupi_n_10774, csa_tree_add_190_195_groupi_n_10775, csa_tree_add_190_195_groupi_n_10776, csa_tree_add_190_195_groupi_n_10777;
  wire csa_tree_add_190_195_groupi_n_10778, csa_tree_add_190_195_groupi_n_10779, csa_tree_add_190_195_groupi_n_10780, csa_tree_add_190_195_groupi_n_10781, csa_tree_add_190_195_groupi_n_10782, csa_tree_add_190_195_groupi_n_10783, csa_tree_add_190_195_groupi_n_10784, csa_tree_add_190_195_groupi_n_10785;
  wire csa_tree_add_190_195_groupi_n_10786, csa_tree_add_190_195_groupi_n_10787, csa_tree_add_190_195_groupi_n_10788, csa_tree_add_190_195_groupi_n_10789, csa_tree_add_190_195_groupi_n_10790, csa_tree_add_190_195_groupi_n_10791, csa_tree_add_190_195_groupi_n_10792, csa_tree_add_190_195_groupi_n_10793;
  wire csa_tree_add_190_195_groupi_n_10794, csa_tree_add_190_195_groupi_n_10795, csa_tree_add_190_195_groupi_n_10796, csa_tree_add_190_195_groupi_n_10797, csa_tree_add_190_195_groupi_n_10798, csa_tree_add_190_195_groupi_n_10799, csa_tree_add_190_195_groupi_n_10800, csa_tree_add_190_195_groupi_n_10801;
  wire csa_tree_add_190_195_groupi_n_10802, csa_tree_add_190_195_groupi_n_10803, csa_tree_add_190_195_groupi_n_10804, csa_tree_add_190_195_groupi_n_10805, csa_tree_add_190_195_groupi_n_10806, csa_tree_add_190_195_groupi_n_10807, csa_tree_add_190_195_groupi_n_10808, csa_tree_add_190_195_groupi_n_10809;
  wire csa_tree_add_190_195_groupi_n_10810, csa_tree_add_190_195_groupi_n_10811, csa_tree_add_190_195_groupi_n_10812, csa_tree_add_190_195_groupi_n_10813, csa_tree_add_190_195_groupi_n_10814, csa_tree_add_190_195_groupi_n_10815, csa_tree_add_190_195_groupi_n_10816, csa_tree_add_190_195_groupi_n_10817;
  wire csa_tree_add_190_195_groupi_n_10818, csa_tree_add_190_195_groupi_n_10819, csa_tree_add_190_195_groupi_n_10820, csa_tree_add_190_195_groupi_n_10821, csa_tree_add_190_195_groupi_n_10822, csa_tree_add_190_195_groupi_n_10823, csa_tree_add_190_195_groupi_n_10824, csa_tree_add_190_195_groupi_n_10825;
  wire csa_tree_add_190_195_groupi_n_10826, csa_tree_add_190_195_groupi_n_10827, csa_tree_add_190_195_groupi_n_10828, csa_tree_add_190_195_groupi_n_10829, csa_tree_add_190_195_groupi_n_10830, csa_tree_add_190_195_groupi_n_10831, csa_tree_add_190_195_groupi_n_10832, csa_tree_add_190_195_groupi_n_10833;
  wire csa_tree_add_190_195_groupi_n_10834, csa_tree_add_190_195_groupi_n_10835, csa_tree_add_190_195_groupi_n_10836, csa_tree_add_190_195_groupi_n_10837, csa_tree_add_190_195_groupi_n_10838, csa_tree_add_190_195_groupi_n_10839, csa_tree_add_190_195_groupi_n_10840, csa_tree_add_190_195_groupi_n_10841;
  wire csa_tree_add_190_195_groupi_n_10842, csa_tree_add_190_195_groupi_n_10843, csa_tree_add_190_195_groupi_n_10844, csa_tree_add_190_195_groupi_n_10845, csa_tree_add_190_195_groupi_n_10846, csa_tree_add_190_195_groupi_n_10847, csa_tree_add_190_195_groupi_n_10848, csa_tree_add_190_195_groupi_n_10849;
  wire csa_tree_add_190_195_groupi_n_10850, csa_tree_add_190_195_groupi_n_10851, csa_tree_add_190_195_groupi_n_10852, csa_tree_add_190_195_groupi_n_10853, csa_tree_add_190_195_groupi_n_10854, csa_tree_add_190_195_groupi_n_10855, csa_tree_add_190_195_groupi_n_10856, csa_tree_add_190_195_groupi_n_10857;
  wire csa_tree_add_190_195_groupi_n_10858, csa_tree_add_190_195_groupi_n_10859, csa_tree_add_190_195_groupi_n_10860, csa_tree_add_190_195_groupi_n_10861, csa_tree_add_190_195_groupi_n_10862, csa_tree_add_190_195_groupi_n_10863, csa_tree_add_190_195_groupi_n_10864, csa_tree_add_190_195_groupi_n_10865;
  wire csa_tree_add_190_195_groupi_n_10866, csa_tree_add_190_195_groupi_n_10867, csa_tree_add_190_195_groupi_n_10868, csa_tree_add_190_195_groupi_n_10869, csa_tree_add_190_195_groupi_n_10870, csa_tree_add_190_195_groupi_n_10871, csa_tree_add_190_195_groupi_n_10872, csa_tree_add_190_195_groupi_n_10873;
  wire csa_tree_add_190_195_groupi_n_10874, csa_tree_add_190_195_groupi_n_10875, csa_tree_add_190_195_groupi_n_10876, csa_tree_add_190_195_groupi_n_10877, csa_tree_add_190_195_groupi_n_10878, csa_tree_add_190_195_groupi_n_10879, csa_tree_add_190_195_groupi_n_10880, csa_tree_add_190_195_groupi_n_10881;
  wire csa_tree_add_190_195_groupi_n_10882, csa_tree_add_190_195_groupi_n_10883, csa_tree_add_190_195_groupi_n_10884, csa_tree_add_190_195_groupi_n_10885, csa_tree_add_190_195_groupi_n_10886, csa_tree_add_190_195_groupi_n_10887, csa_tree_add_190_195_groupi_n_10888, csa_tree_add_190_195_groupi_n_10889;
  wire csa_tree_add_190_195_groupi_n_10890, csa_tree_add_190_195_groupi_n_10891, csa_tree_add_190_195_groupi_n_10892, csa_tree_add_190_195_groupi_n_10893, csa_tree_add_190_195_groupi_n_10894, csa_tree_add_190_195_groupi_n_10895, csa_tree_add_190_195_groupi_n_10896, csa_tree_add_190_195_groupi_n_10897;
  wire csa_tree_add_190_195_groupi_n_10898, csa_tree_add_190_195_groupi_n_10899, csa_tree_add_190_195_groupi_n_10900, csa_tree_add_190_195_groupi_n_10901, csa_tree_add_190_195_groupi_n_10902, csa_tree_add_190_195_groupi_n_10903, csa_tree_add_190_195_groupi_n_10904, csa_tree_add_190_195_groupi_n_10905;
  wire csa_tree_add_190_195_groupi_n_10906, csa_tree_add_190_195_groupi_n_10907, csa_tree_add_190_195_groupi_n_10908, csa_tree_add_190_195_groupi_n_10909, csa_tree_add_190_195_groupi_n_10910, csa_tree_add_190_195_groupi_n_10911, csa_tree_add_190_195_groupi_n_10912, csa_tree_add_190_195_groupi_n_10913;
  wire csa_tree_add_190_195_groupi_n_10914, csa_tree_add_190_195_groupi_n_10915, csa_tree_add_190_195_groupi_n_10916, csa_tree_add_190_195_groupi_n_10917, csa_tree_add_190_195_groupi_n_10918, csa_tree_add_190_195_groupi_n_10919, csa_tree_add_190_195_groupi_n_10920, csa_tree_add_190_195_groupi_n_10921;
  wire csa_tree_add_190_195_groupi_n_10922, csa_tree_add_190_195_groupi_n_10923, csa_tree_add_190_195_groupi_n_10924, csa_tree_add_190_195_groupi_n_10925, csa_tree_add_190_195_groupi_n_10926, csa_tree_add_190_195_groupi_n_10927, csa_tree_add_190_195_groupi_n_10928, csa_tree_add_190_195_groupi_n_10929;
  wire csa_tree_add_190_195_groupi_n_10930, csa_tree_add_190_195_groupi_n_10931, csa_tree_add_190_195_groupi_n_10932, csa_tree_add_190_195_groupi_n_10933, csa_tree_add_190_195_groupi_n_10934, csa_tree_add_190_195_groupi_n_10935, csa_tree_add_190_195_groupi_n_10936, csa_tree_add_190_195_groupi_n_10937;
  wire csa_tree_add_190_195_groupi_n_10938, csa_tree_add_190_195_groupi_n_10939, csa_tree_add_190_195_groupi_n_10940, csa_tree_add_190_195_groupi_n_10941, csa_tree_add_190_195_groupi_n_10942, csa_tree_add_190_195_groupi_n_10943, csa_tree_add_190_195_groupi_n_10944, csa_tree_add_190_195_groupi_n_10945;
  wire csa_tree_add_190_195_groupi_n_10946, csa_tree_add_190_195_groupi_n_10947, csa_tree_add_190_195_groupi_n_10948, csa_tree_add_190_195_groupi_n_10949, csa_tree_add_190_195_groupi_n_10950, csa_tree_add_190_195_groupi_n_10951, csa_tree_add_190_195_groupi_n_10952, csa_tree_add_190_195_groupi_n_10953;
  wire csa_tree_add_190_195_groupi_n_10954, csa_tree_add_190_195_groupi_n_10955, csa_tree_add_190_195_groupi_n_10956, csa_tree_add_190_195_groupi_n_10957, csa_tree_add_190_195_groupi_n_10958, csa_tree_add_190_195_groupi_n_10959, csa_tree_add_190_195_groupi_n_10960, csa_tree_add_190_195_groupi_n_10961;
  wire csa_tree_add_190_195_groupi_n_10962, csa_tree_add_190_195_groupi_n_10963, csa_tree_add_190_195_groupi_n_10964, csa_tree_add_190_195_groupi_n_10965, csa_tree_add_190_195_groupi_n_10966, csa_tree_add_190_195_groupi_n_10967, csa_tree_add_190_195_groupi_n_10968, csa_tree_add_190_195_groupi_n_10969;
  wire csa_tree_add_190_195_groupi_n_10970, csa_tree_add_190_195_groupi_n_10971, csa_tree_add_190_195_groupi_n_10972, csa_tree_add_190_195_groupi_n_10973, csa_tree_add_190_195_groupi_n_10974, csa_tree_add_190_195_groupi_n_10975, csa_tree_add_190_195_groupi_n_10976, csa_tree_add_190_195_groupi_n_10977;
  wire csa_tree_add_190_195_groupi_n_10978, csa_tree_add_190_195_groupi_n_10979, csa_tree_add_190_195_groupi_n_10980, csa_tree_add_190_195_groupi_n_10981, csa_tree_add_190_195_groupi_n_10982, csa_tree_add_190_195_groupi_n_10983, csa_tree_add_190_195_groupi_n_10984, csa_tree_add_190_195_groupi_n_10985;
  wire csa_tree_add_190_195_groupi_n_10986, csa_tree_add_190_195_groupi_n_10987, csa_tree_add_190_195_groupi_n_10988, csa_tree_add_190_195_groupi_n_10989, csa_tree_add_190_195_groupi_n_10990, csa_tree_add_190_195_groupi_n_10991, csa_tree_add_190_195_groupi_n_10992, csa_tree_add_190_195_groupi_n_10993;
  wire csa_tree_add_190_195_groupi_n_10994, csa_tree_add_190_195_groupi_n_10995, csa_tree_add_190_195_groupi_n_10996, csa_tree_add_190_195_groupi_n_10997, csa_tree_add_190_195_groupi_n_10998, csa_tree_add_190_195_groupi_n_10999, csa_tree_add_190_195_groupi_n_11000, csa_tree_add_190_195_groupi_n_11001;
  wire csa_tree_add_190_195_groupi_n_11002, csa_tree_add_190_195_groupi_n_11004, csa_tree_add_190_195_groupi_n_11005, csa_tree_add_190_195_groupi_n_11006, csa_tree_add_190_195_groupi_n_11007, csa_tree_add_190_195_groupi_n_11008, csa_tree_add_190_195_groupi_n_11009, csa_tree_add_190_195_groupi_n_11010;
  wire csa_tree_add_190_195_groupi_n_11011, csa_tree_add_190_195_groupi_n_11012, csa_tree_add_190_195_groupi_n_11013, csa_tree_add_190_195_groupi_n_11014, csa_tree_add_190_195_groupi_n_11015, csa_tree_add_190_195_groupi_n_11016, csa_tree_add_190_195_groupi_n_11017, csa_tree_add_190_195_groupi_n_11018;
  wire csa_tree_add_190_195_groupi_n_11019, csa_tree_add_190_195_groupi_n_11020, csa_tree_add_190_195_groupi_n_11021, csa_tree_add_190_195_groupi_n_11022, csa_tree_add_190_195_groupi_n_11023, csa_tree_add_190_195_groupi_n_11024, csa_tree_add_190_195_groupi_n_11025, csa_tree_add_190_195_groupi_n_11026;
  wire csa_tree_add_190_195_groupi_n_11027, csa_tree_add_190_195_groupi_n_11028, csa_tree_add_190_195_groupi_n_11029, csa_tree_add_190_195_groupi_n_11030, csa_tree_add_190_195_groupi_n_11031, csa_tree_add_190_195_groupi_n_11032, csa_tree_add_190_195_groupi_n_11033, csa_tree_add_190_195_groupi_n_11034;
  wire csa_tree_add_190_195_groupi_n_11035, csa_tree_add_190_195_groupi_n_11036, csa_tree_add_190_195_groupi_n_11037, csa_tree_add_190_195_groupi_n_11038, csa_tree_add_190_195_groupi_n_11039, csa_tree_add_190_195_groupi_n_11040, csa_tree_add_190_195_groupi_n_11041, csa_tree_add_190_195_groupi_n_11042;
  wire csa_tree_add_190_195_groupi_n_11043, csa_tree_add_190_195_groupi_n_11044, csa_tree_add_190_195_groupi_n_11045, csa_tree_add_190_195_groupi_n_11046, csa_tree_add_190_195_groupi_n_11047, csa_tree_add_190_195_groupi_n_11048, csa_tree_add_190_195_groupi_n_11049, csa_tree_add_190_195_groupi_n_11050;
  wire csa_tree_add_190_195_groupi_n_11051, csa_tree_add_190_195_groupi_n_11052, csa_tree_add_190_195_groupi_n_11053, csa_tree_add_190_195_groupi_n_11054, csa_tree_add_190_195_groupi_n_11055, csa_tree_add_190_195_groupi_n_11056, csa_tree_add_190_195_groupi_n_11057, csa_tree_add_190_195_groupi_n_11058;
  wire csa_tree_add_190_195_groupi_n_11059, csa_tree_add_190_195_groupi_n_11060, csa_tree_add_190_195_groupi_n_11061, csa_tree_add_190_195_groupi_n_11062, csa_tree_add_190_195_groupi_n_11063, csa_tree_add_190_195_groupi_n_11064, csa_tree_add_190_195_groupi_n_11065, csa_tree_add_190_195_groupi_n_11066;
  wire csa_tree_add_190_195_groupi_n_11067, csa_tree_add_190_195_groupi_n_11068, csa_tree_add_190_195_groupi_n_11069, csa_tree_add_190_195_groupi_n_11070, csa_tree_add_190_195_groupi_n_11071, csa_tree_add_190_195_groupi_n_11072, csa_tree_add_190_195_groupi_n_11073, csa_tree_add_190_195_groupi_n_11074;
  wire csa_tree_add_190_195_groupi_n_11075, csa_tree_add_190_195_groupi_n_11076, csa_tree_add_190_195_groupi_n_11077, csa_tree_add_190_195_groupi_n_11078, csa_tree_add_190_195_groupi_n_11079, csa_tree_add_190_195_groupi_n_11080, csa_tree_add_190_195_groupi_n_11081, csa_tree_add_190_195_groupi_n_11082;
  wire csa_tree_add_190_195_groupi_n_11083, csa_tree_add_190_195_groupi_n_11084, csa_tree_add_190_195_groupi_n_11085, csa_tree_add_190_195_groupi_n_11086, csa_tree_add_190_195_groupi_n_11087, csa_tree_add_190_195_groupi_n_11088, csa_tree_add_190_195_groupi_n_11089, csa_tree_add_190_195_groupi_n_11090;
  wire csa_tree_add_190_195_groupi_n_11091, csa_tree_add_190_195_groupi_n_11092, csa_tree_add_190_195_groupi_n_11093, csa_tree_add_190_195_groupi_n_11094, csa_tree_add_190_195_groupi_n_11095, csa_tree_add_190_195_groupi_n_11096, csa_tree_add_190_195_groupi_n_11097, csa_tree_add_190_195_groupi_n_11098;
  wire csa_tree_add_190_195_groupi_n_11099, csa_tree_add_190_195_groupi_n_11100, csa_tree_add_190_195_groupi_n_11101, csa_tree_add_190_195_groupi_n_11102, csa_tree_add_190_195_groupi_n_11103, csa_tree_add_190_195_groupi_n_11104, csa_tree_add_190_195_groupi_n_11105, csa_tree_add_190_195_groupi_n_11106;
  wire csa_tree_add_190_195_groupi_n_11107, csa_tree_add_190_195_groupi_n_11108, csa_tree_add_190_195_groupi_n_11109, csa_tree_add_190_195_groupi_n_11110, csa_tree_add_190_195_groupi_n_11111, csa_tree_add_190_195_groupi_n_11112, csa_tree_add_190_195_groupi_n_11113, csa_tree_add_190_195_groupi_n_11114;
  wire csa_tree_add_190_195_groupi_n_11115, csa_tree_add_190_195_groupi_n_11116, csa_tree_add_190_195_groupi_n_11117, csa_tree_add_190_195_groupi_n_11118, csa_tree_add_190_195_groupi_n_11119, csa_tree_add_190_195_groupi_n_11120, csa_tree_add_190_195_groupi_n_11121, csa_tree_add_190_195_groupi_n_11122;
  wire csa_tree_add_190_195_groupi_n_11123, csa_tree_add_190_195_groupi_n_11124, csa_tree_add_190_195_groupi_n_11125, csa_tree_add_190_195_groupi_n_11126, csa_tree_add_190_195_groupi_n_11127, csa_tree_add_190_195_groupi_n_11128, csa_tree_add_190_195_groupi_n_11129, csa_tree_add_190_195_groupi_n_11130;
  wire csa_tree_add_190_195_groupi_n_11131, csa_tree_add_190_195_groupi_n_11132, csa_tree_add_190_195_groupi_n_11133, csa_tree_add_190_195_groupi_n_11134, csa_tree_add_190_195_groupi_n_11135, csa_tree_add_190_195_groupi_n_11136, csa_tree_add_190_195_groupi_n_11137, csa_tree_add_190_195_groupi_n_11138;
  wire csa_tree_add_190_195_groupi_n_11139, csa_tree_add_190_195_groupi_n_11140, csa_tree_add_190_195_groupi_n_11141, csa_tree_add_190_195_groupi_n_11142, csa_tree_add_190_195_groupi_n_11143, csa_tree_add_190_195_groupi_n_11144, csa_tree_add_190_195_groupi_n_11145, csa_tree_add_190_195_groupi_n_11146;
  wire csa_tree_add_190_195_groupi_n_11147, csa_tree_add_190_195_groupi_n_11148, csa_tree_add_190_195_groupi_n_11149, csa_tree_add_190_195_groupi_n_11150, csa_tree_add_190_195_groupi_n_11151, csa_tree_add_190_195_groupi_n_11152, csa_tree_add_190_195_groupi_n_11153, csa_tree_add_190_195_groupi_n_11154;
  wire csa_tree_add_190_195_groupi_n_11155, csa_tree_add_190_195_groupi_n_11156, csa_tree_add_190_195_groupi_n_11157, csa_tree_add_190_195_groupi_n_11158, csa_tree_add_190_195_groupi_n_11159, csa_tree_add_190_195_groupi_n_11160, csa_tree_add_190_195_groupi_n_11161, csa_tree_add_190_195_groupi_n_11162;
  wire csa_tree_add_190_195_groupi_n_11163, csa_tree_add_190_195_groupi_n_11164, csa_tree_add_190_195_groupi_n_11165, csa_tree_add_190_195_groupi_n_11166, csa_tree_add_190_195_groupi_n_11167, csa_tree_add_190_195_groupi_n_11168, csa_tree_add_190_195_groupi_n_11169, csa_tree_add_190_195_groupi_n_11170;
  wire csa_tree_add_190_195_groupi_n_11171, csa_tree_add_190_195_groupi_n_11172, csa_tree_add_190_195_groupi_n_11173, csa_tree_add_190_195_groupi_n_11174, csa_tree_add_190_195_groupi_n_11175, csa_tree_add_190_195_groupi_n_11176, csa_tree_add_190_195_groupi_n_11177, csa_tree_add_190_195_groupi_n_11178;
  wire csa_tree_add_190_195_groupi_n_11179, csa_tree_add_190_195_groupi_n_11180, csa_tree_add_190_195_groupi_n_11181, csa_tree_add_190_195_groupi_n_11182, csa_tree_add_190_195_groupi_n_11183, csa_tree_add_190_195_groupi_n_11184, csa_tree_add_190_195_groupi_n_11185, csa_tree_add_190_195_groupi_n_11186;
  wire csa_tree_add_190_195_groupi_n_11187, csa_tree_add_190_195_groupi_n_11188, csa_tree_add_190_195_groupi_n_11189, csa_tree_add_190_195_groupi_n_11190, csa_tree_add_190_195_groupi_n_11191, csa_tree_add_190_195_groupi_n_11192, csa_tree_add_190_195_groupi_n_11193, csa_tree_add_190_195_groupi_n_11194;
  wire csa_tree_add_190_195_groupi_n_11195, csa_tree_add_190_195_groupi_n_11196, csa_tree_add_190_195_groupi_n_11197, csa_tree_add_190_195_groupi_n_11198, csa_tree_add_190_195_groupi_n_11199, csa_tree_add_190_195_groupi_n_11200, csa_tree_add_190_195_groupi_n_11201, csa_tree_add_190_195_groupi_n_11202;
  wire csa_tree_add_190_195_groupi_n_11203, csa_tree_add_190_195_groupi_n_11204, csa_tree_add_190_195_groupi_n_11205, csa_tree_add_190_195_groupi_n_11206, csa_tree_add_190_195_groupi_n_11207, csa_tree_add_190_195_groupi_n_11208, csa_tree_add_190_195_groupi_n_11209, csa_tree_add_190_195_groupi_n_11210;
  wire csa_tree_add_190_195_groupi_n_11211, csa_tree_add_190_195_groupi_n_11212, csa_tree_add_190_195_groupi_n_11213, csa_tree_add_190_195_groupi_n_11214, csa_tree_add_190_195_groupi_n_11215, csa_tree_add_190_195_groupi_n_11216, csa_tree_add_190_195_groupi_n_11217, csa_tree_add_190_195_groupi_n_11218;
  wire csa_tree_add_190_195_groupi_n_11219, csa_tree_add_190_195_groupi_n_11220, csa_tree_add_190_195_groupi_n_11221, csa_tree_add_190_195_groupi_n_11222, csa_tree_add_190_195_groupi_n_11223, csa_tree_add_190_195_groupi_n_11224, csa_tree_add_190_195_groupi_n_11225, csa_tree_add_190_195_groupi_n_11226;
  wire csa_tree_add_190_195_groupi_n_11227, csa_tree_add_190_195_groupi_n_11228, csa_tree_add_190_195_groupi_n_11229, csa_tree_add_190_195_groupi_n_11230, csa_tree_add_190_195_groupi_n_11231, csa_tree_add_190_195_groupi_n_11232, csa_tree_add_190_195_groupi_n_11233, csa_tree_add_190_195_groupi_n_11234;
  wire csa_tree_add_190_195_groupi_n_11235, csa_tree_add_190_195_groupi_n_11236, csa_tree_add_190_195_groupi_n_11237, csa_tree_add_190_195_groupi_n_11238, csa_tree_add_190_195_groupi_n_11239, csa_tree_add_190_195_groupi_n_11240, csa_tree_add_190_195_groupi_n_11241, csa_tree_add_190_195_groupi_n_11242;
  wire csa_tree_add_190_195_groupi_n_11243, csa_tree_add_190_195_groupi_n_11244, csa_tree_add_190_195_groupi_n_11245, csa_tree_add_190_195_groupi_n_11246, csa_tree_add_190_195_groupi_n_11247, csa_tree_add_190_195_groupi_n_11248, csa_tree_add_190_195_groupi_n_11249, csa_tree_add_190_195_groupi_n_11250;
  wire csa_tree_add_190_195_groupi_n_11251, csa_tree_add_190_195_groupi_n_11252, csa_tree_add_190_195_groupi_n_11253, csa_tree_add_190_195_groupi_n_11254, csa_tree_add_190_195_groupi_n_11255, csa_tree_add_190_195_groupi_n_11256, csa_tree_add_190_195_groupi_n_11257, csa_tree_add_190_195_groupi_n_11258;
  wire csa_tree_add_190_195_groupi_n_11259, csa_tree_add_190_195_groupi_n_11260, csa_tree_add_190_195_groupi_n_11261, csa_tree_add_190_195_groupi_n_11262, csa_tree_add_190_195_groupi_n_11263, csa_tree_add_190_195_groupi_n_11264, csa_tree_add_190_195_groupi_n_11265, csa_tree_add_190_195_groupi_n_11266;
  wire csa_tree_add_190_195_groupi_n_11267, csa_tree_add_190_195_groupi_n_11268, csa_tree_add_190_195_groupi_n_11269, csa_tree_add_190_195_groupi_n_11270, csa_tree_add_190_195_groupi_n_11271, csa_tree_add_190_195_groupi_n_11272, csa_tree_add_190_195_groupi_n_11273, csa_tree_add_190_195_groupi_n_11274;
  wire csa_tree_add_190_195_groupi_n_11275, csa_tree_add_190_195_groupi_n_11276, csa_tree_add_190_195_groupi_n_11277, csa_tree_add_190_195_groupi_n_11278, csa_tree_add_190_195_groupi_n_11279, csa_tree_add_190_195_groupi_n_11280, csa_tree_add_190_195_groupi_n_11281, csa_tree_add_190_195_groupi_n_11282;
  wire csa_tree_add_190_195_groupi_n_11283, csa_tree_add_190_195_groupi_n_11284, csa_tree_add_190_195_groupi_n_11285, csa_tree_add_190_195_groupi_n_11286, csa_tree_add_190_195_groupi_n_11287, csa_tree_add_190_195_groupi_n_11288, csa_tree_add_190_195_groupi_n_11289, csa_tree_add_190_195_groupi_n_11290;
  wire csa_tree_add_190_195_groupi_n_11291, csa_tree_add_190_195_groupi_n_11292, csa_tree_add_190_195_groupi_n_11293, csa_tree_add_190_195_groupi_n_11294, csa_tree_add_190_195_groupi_n_11295, csa_tree_add_190_195_groupi_n_11296, csa_tree_add_190_195_groupi_n_11297, csa_tree_add_190_195_groupi_n_11298;
  wire csa_tree_add_190_195_groupi_n_11299, csa_tree_add_190_195_groupi_n_11300, csa_tree_add_190_195_groupi_n_11301, csa_tree_add_190_195_groupi_n_11302, csa_tree_add_190_195_groupi_n_11303, csa_tree_add_190_195_groupi_n_11304, csa_tree_add_190_195_groupi_n_11305, csa_tree_add_190_195_groupi_n_11306;
  wire csa_tree_add_190_195_groupi_n_11307, csa_tree_add_190_195_groupi_n_11308, csa_tree_add_190_195_groupi_n_11309, csa_tree_add_190_195_groupi_n_11310, csa_tree_add_190_195_groupi_n_11311, csa_tree_add_190_195_groupi_n_11312, csa_tree_add_190_195_groupi_n_11313, csa_tree_add_190_195_groupi_n_11314;
  wire csa_tree_add_190_195_groupi_n_11315, csa_tree_add_190_195_groupi_n_11316, csa_tree_add_190_195_groupi_n_11317, csa_tree_add_190_195_groupi_n_11318, csa_tree_add_190_195_groupi_n_11319, csa_tree_add_190_195_groupi_n_11320, csa_tree_add_190_195_groupi_n_11321, csa_tree_add_190_195_groupi_n_11322;
  wire csa_tree_add_190_195_groupi_n_11323, csa_tree_add_190_195_groupi_n_11324, csa_tree_add_190_195_groupi_n_11325, csa_tree_add_190_195_groupi_n_11326, csa_tree_add_190_195_groupi_n_11327, csa_tree_add_190_195_groupi_n_11328, csa_tree_add_190_195_groupi_n_11329, csa_tree_add_190_195_groupi_n_11330;
  wire csa_tree_add_190_195_groupi_n_11331, csa_tree_add_190_195_groupi_n_11332, csa_tree_add_190_195_groupi_n_11333, csa_tree_add_190_195_groupi_n_11334, csa_tree_add_190_195_groupi_n_11335, csa_tree_add_190_195_groupi_n_11336, csa_tree_add_190_195_groupi_n_11337, csa_tree_add_190_195_groupi_n_11338;
  wire csa_tree_add_190_195_groupi_n_11339, csa_tree_add_190_195_groupi_n_11340, csa_tree_add_190_195_groupi_n_11341, csa_tree_add_190_195_groupi_n_11342, csa_tree_add_190_195_groupi_n_11343, csa_tree_add_190_195_groupi_n_11344, csa_tree_add_190_195_groupi_n_11345, csa_tree_add_190_195_groupi_n_11346;
  wire csa_tree_add_190_195_groupi_n_11347, csa_tree_add_190_195_groupi_n_11348, csa_tree_add_190_195_groupi_n_11349, csa_tree_add_190_195_groupi_n_11350, csa_tree_add_190_195_groupi_n_11351, csa_tree_add_190_195_groupi_n_11352, csa_tree_add_190_195_groupi_n_11353, csa_tree_add_190_195_groupi_n_11354;
  wire csa_tree_add_190_195_groupi_n_11355, csa_tree_add_190_195_groupi_n_11356, csa_tree_add_190_195_groupi_n_11357, csa_tree_add_190_195_groupi_n_11358, csa_tree_add_190_195_groupi_n_11359, csa_tree_add_190_195_groupi_n_11360, csa_tree_add_190_195_groupi_n_11361, csa_tree_add_190_195_groupi_n_11362;
  wire csa_tree_add_190_195_groupi_n_11363, csa_tree_add_190_195_groupi_n_11364, csa_tree_add_190_195_groupi_n_11365, csa_tree_add_190_195_groupi_n_11366, csa_tree_add_190_195_groupi_n_11367, csa_tree_add_190_195_groupi_n_11368, csa_tree_add_190_195_groupi_n_11369, csa_tree_add_190_195_groupi_n_11370;
  wire csa_tree_add_190_195_groupi_n_11371, csa_tree_add_190_195_groupi_n_11372, csa_tree_add_190_195_groupi_n_11373, csa_tree_add_190_195_groupi_n_11374, csa_tree_add_190_195_groupi_n_11375, csa_tree_add_190_195_groupi_n_11376, csa_tree_add_190_195_groupi_n_11377, csa_tree_add_190_195_groupi_n_11378;
  wire csa_tree_add_190_195_groupi_n_11379, csa_tree_add_190_195_groupi_n_11380, csa_tree_add_190_195_groupi_n_11381, csa_tree_add_190_195_groupi_n_11382, csa_tree_add_190_195_groupi_n_11383, csa_tree_add_190_195_groupi_n_11384, csa_tree_add_190_195_groupi_n_11385, csa_tree_add_190_195_groupi_n_11386;
  wire csa_tree_add_190_195_groupi_n_11387, csa_tree_add_190_195_groupi_n_11388, csa_tree_add_190_195_groupi_n_11389, csa_tree_add_190_195_groupi_n_11390, csa_tree_add_190_195_groupi_n_11391, csa_tree_add_190_195_groupi_n_11392, csa_tree_add_190_195_groupi_n_11393, csa_tree_add_190_195_groupi_n_11394;
  wire csa_tree_add_190_195_groupi_n_11395, csa_tree_add_190_195_groupi_n_11396, csa_tree_add_190_195_groupi_n_11397, csa_tree_add_190_195_groupi_n_11398, csa_tree_add_190_195_groupi_n_11399, csa_tree_add_190_195_groupi_n_11400, csa_tree_add_190_195_groupi_n_11401, csa_tree_add_190_195_groupi_n_11402;
  wire csa_tree_add_190_195_groupi_n_11403, csa_tree_add_190_195_groupi_n_11404, csa_tree_add_190_195_groupi_n_11405, csa_tree_add_190_195_groupi_n_11406, csa_tree_add_190_195_groupi_n_11407, csa_tree_add_190_195_groupi_n_11408, csa_tree_add_190_195_groupi_n_11409, csa_tree_add_190_195_groupi_n_11410;
  wire csa_tree_add_190_195_groupi_n_11411, csa_tree_add_190_195_groupi_n_11412, csa_tree_add_190_195_groupi_n_11413, csa_tree_add_190_195_groupi_n_11414, csa_tree_add_190_195_groupi_n_11415, csa_tree_add_190_195_groupi_n_11416, csa_tree_add_190_195_groupi_n_11417, csa_tree_add_190_195_groupi_n_11418;
  wire csa_tree_add_190_195_groupi_n_11419, csa_tree_add_190_195_groupi_n_11420, csa_tree_add_190_195_groupi_n_11421, csa_tree_add_190_195_groupi_n_11422, csa_tree_add_190_195_groupi_n_11423, csa_tree_add_190_195_groupi_n_11424, csa_tree_add_190_195_groupi_n_11425, csa_tree_add_190_195_groupi_n_11426;
  wire csa_tree_add_190_195_groupi_n_11427, csa_tree_add_190_195_groupi_n_11428, csa_tree_add_190_195_groupi_n_11429, csa_tree_add_190_195_groupi_n_11430, csa_tree_add_190_195_groupi_n_11431, csa_tree_add_190_195_groupi_n_11432, csa_tree_add_190_195_groupi_n_11433, csa_tree_add_190_195_groupi_n_11434;
  wire csa_tree_add_190_195_groupi_n_11435, csa_tree_add_190_195_groupi_n_11436, csa_tree_add_190_195_groupi_n_11437, csa_tree_add_190_195_groupi_n_11438, csa_tree_add_190_195_groupi_n_11439, csa_tree_add_190_195_groupi_n_11440, csa_tree_add_190_195_groupi_n_11441, csa_tree_add_190_195_groupi_n_11442;
  wire csa_tree_add_190_195_groupi_n_11443, csa_tree_add_190_195_groupi_n_11444, csa_tree_add_190_195_groupi_n_11445, csa_tree_add_190_195_groupi_n_11446, csa_tree_add_190_195_groupi_n_11447, csa_tree_add_190_195_groupi_n_11448, csa_tree_add_190_195_groupi_n_11449, csa_tree_add_190_195_groupi_n_11450;
  wire csa_tree_add_190_195_groupi_n_11451, csa_tree_add_190_195_groupi_n_11452, csa_tree_add_190_195_groupi_n_11453, csa_tree_add_190_195_groupi_n_11454, csa_tree_add_190_195_groupi_n_11455, csa_tree_add_190_195_groupi_n_11456, csa_tree_add_190_195_groupi_n_11457, csa_tree_add_190_195_groupi_n_11458;
  wire csa_tree_add_190_195_groupi_n_11459, csa_tree_add_190_195_groupi_n_11460, csa_tree_add_190_195_groupi_n_11461, csa_tree_add_190_195_groupi_n_11462, csa_tree_add_190_195_groupi_n_11463, csa_tree_add_190_195_groupi_n_11464, csa_tree_add_190_195_groupi_n_11465, csa_tree_add_190_195_groupi_n_11466;
  wire csa_tree_add_190_195_groupi_n_11467, csa_tree_add_190_195_groupi_n_11468, csa_tree_add_190_195_groupi_n_11469, csa_tree_add_190_195_groupi_n_11470, csa_tree_add_190_195_groupi_n_11471, csa_tree_add_190_195_groupi_n_11472, csa_tree_add_190_195_groupi_n_11473, csa_tree_add_190_195_groupi_n_11474;
  wire csa_tree_add_190_195_groupi_n_11475, csa_tree_add_190_195_groupi_n_11476, csa_tree_add_190_195_groupi_n_11477, csa_tree_add_190_195_groupi_n_11478, csa_tree_add_190_195_groupi_n_11479, csa_tree_add_190_195_groupi_n_11480, csa_tree_add_190_195_groupi_n_11481, csa_tree_add_190_195_groupi_n_11482;
  wire csa_tree_add_190_195_groupi_n_11483, csa_tree_add_190_195_groupi_n_11484, csa_tree_add_190_195_groupi_n_11485, csa_tree_add_190_195_groupi_n_11486, csa_tree_add_190_195_groupi_n_11487, csa_tree_add_190_195_groupi_n_11488, csa_tree_add_190_195_groupi_n_11489, csa_tree_add_190_195_groupi_n_11490;
  wire csa_tree_add_190_195_groupi_n_11491, csa_tree_add_190_195_groupi_n_11492, csa_tree_add_190_195_groupi_n_11493, csa_tree_add_190_195_groupi_n_11494, csa_tree_add_190_195_groupi_n_11495, csa_tree_add_190_195_groupi_n_11496, csa_tree_add_190_195_groupi_n_11497, csa_tree_add_190_195_groupi_n_11498;
  wire csa_tree_add_190_195_groupi_n_11499, csa_tree_add_190_195_groupi_n_11500, csa_tree_add_190_195_groupi_n_11501, csa_tree_add_190_195_groupi_n_11502, csa_tree_add_190_195_groupi_n_11503, csa_tree_add_190_195_groupi_n_11504, csa_tree_add_190_195_groupi_n_11505, csa_tree_add_190_195_groupi_n_11506;
  wire csa_tree_add_190_195_groupi_n_11507, csa_tree_add_190_195_groupi_n_11508, csa_tree_add_190_195_groupi_n_11509, csa_tree_add_190_195_groupi_n_11510, csa_tree_add_190_195_groupi_n_11511, csa_tree_add_190_195_groupi_n_11512, csa_tree_add_190_195_groupi_n_11513, csa_tree_add_190_195_groupi_n_11514;
  wire csa_tree_add_190_195_groupi_n_11515, csa_tree_add_190_195_groupi_n_11516, csa_tree_add_190_195_groupi_n_11517, csa_tree_add_190_195_groupi_n_11518, csa_tree_add_190_195_groupi_n_11519, csa_tree_add_190_195_groupi_n_11520, csa_tree_add_190_195_groupi_n_11521, csa_tree_add_190_195_groupi_n_11522;
  wire csa_tree_add_190_195_groupi_n_11523, csa_tree_add_190_195_groupi_n_11524, csa_tree_add_190_195_groupi_n_11525, csa_tree_add_190_195_groupi_n_11526, csa_tree_add_190_195_groupi_n_11527, csa_tree_add_190_195_groupi_n_11528, csa_tree_add_190_195_groupi_n_11529, csa_tree_add_190_195_groupi_n_11530;
  wire csa_tree_add_190_195_groupi_n_11531, csa_tree_add_190_195_groupi_n_11532, csa_tree_add_190_195_groupi_n_11533, csa_tree_add_190_195_groupi_n_11534, csa_tree_add_190_195_groupi_n_11535, csa_tree_add_190_195_groupi_n_11536, csa_tree_add_190_195_groupi_n_11537, csa_tree_add_190_195_groupi_n_11538;
  wire csa_tree_add_190_195_groupi_n_11539, csa_tree_add_190_195_groupi_n_11540, csa_tree_add_190_195_groupi_n_11541, csa_tree_add_190_195_groupi_n_11542, csa_tree_add_190_195_groupi_n_11543, csa_tree_add_190_195_groupi_n_11544, csa_tree_add_190_195_groupi_n_11545, csa_tree_add_190_195_groupi_n_11546;
  wire csa_tree_add_190_195_groupi_n_11547, csa_tree_add_190_195_groupi_n_11548, csa_tree_add_190_195_groupi_n_11549, csa_tree_add_190_195_groupi_n_11550, csa_tree_add_190_195_groupi_n_11551, csa_tree_add_190_195_groupi_n_11552, csa_tree_add_190_195_groupi_n_11553, csa_tree_add_190_195_groupi_n_11554;
  wire csa_tree_add_190_195_groupi_n_11555, csa_tree_add_190_195_groupi_n_11556, csa_tree_add_190_195_groupi_n_11557, csa_tree_add_190_195_groupi_n_11558, csa_tree_add_190_195_groupi_n_11559, csa_tree_add_190_195_groupi_n_11560, csa_tree_add_190_195_groupi_n_11561, csa_tree_add_190_195_groupi_n_11562;
  wire csa_tree_add_190_195_groupi_n_11563, csa_tree_add_190_195_groupi_n_11564, csa_tree_add_190_195_groupi_n_11565, csa_tree_add_190_195_groupi_n_11566, csa_tree_add_190_195_groupi_n_11567, csa_tree_add_190_195_groupi_n_11568, csa_tree_add_190_195_groupi_n_11569, csa_tree_add_190_195_groupi_n_11570;
  wire csa_tree_add_190_195_groupi_n_11571, csa_tree_add_190_195_groupi_n_11572, csa_tree_add_190_195_groupi_n_11573, csa_tree_add_190_195_groupi_n_11574, csa_tree_add_190_195_groupi_n_11575, csa_tree_add_190_195_groupi_n_11576, csa_tree_add_190_195_groupi_n_11577, csa_tree_add_190_195_groupi_n_11578;
  wire csa_tree_add_190_195_groupi_n_11579, csa_tree_add_190_195_groupi_n_11580, csa_tree_add_190_195_groupi_n_11581, csa_tree_add_190_195_groupi_n_11582, csa_tree_add_190_195_groupi_n_11583, csa_tree_add_190_195_groupi_n_11584, csa_tree_add_190_195_groupi_n_11585, csa_tree_add_190_195_groupi_n_11586;
  wire csa_tree_add_190_195_groupi_n_11587, csa_tree_add_190_195_groupi_n_11588, csa_tree_add_190_195_groupi_n_11589, csa_tree_add_190_195_groupi_n_11590, csa_tree_add_190_195_groupi_n_11591, csa_tree_add_190_195_groupi_n_11592, csa_tree_add_190_195_groupi_n_11593, csa_tree_add_190_195_groupi_n_11594;
  wire csa_tree_add_190_195_groupi_n_11595, csa_tree_add_190_195_groupi_n_11596, csa_tree_add_190_195_groupi_n_11597, csa_tree_add_190_195_groupi_n_11598, csa_tree_add_190_195_groupi_n_11599, csa_tree_add_190_195_groupi_n_11600, csa_tree_add_190_195_groupi_n_11601, csa_tree_add_190_195_groupi_n_11602;
  wire csa_tree_add_190_195_groupi_n_11603, csa_tree_add_190_195_groupi_n_11604, csa_tree_add_190_195_groupi_n_11605, csa_tree_add_190_195_groupi_n_11606, csa_tree_add_190_195_groupi_n_11607, csa_tree_add_190_195_groupi_n_11608, csa_tree_add_190_195_groupi_n_11609, csa_tree_add_190_195_groupi_n_11610;
  wire csa_tree_add_190_195_groupi_n_11611, csa_tree_add_190_195_groupi_n_11612, csa_tree_add_190_195_groupi_n_11613, csa_tree_add_190_195_groupi_n_11614, csa_tree_add_190_195_groupi_n_11615, csa_tree_add_190_195_groupi_n_11616, csa_tree_add_190_195_groupi_n_11617, csa_tree_add_190_195_groupi_n_11618;
  wire csa_tree_add_190_195_groupi_n_11619, csa_tree_add_190_195_groupi_n_11620, csa_tree_add_190_195_groupi_n_11621, csa_tree_add_190_195_groupi_n_11622, csa_tree_add_190_195_groupi_n_11623, csa_tree_add_190_195_groupi_n_11624, csa_tree_add_190_195_groupi_n_11625, csa_tree_add_190_195_groupi_n_11626;
  wire csa_tree_add_190_195_groupi_n_11627, csa_tree_add_190_195_groupi_n_11628, csa_tree_add_190_195_groupi_n_11630, csa_tree_add_190_195_groupi_n_11631, csa_tree_add_190_195_groupi_n_11632, csa_tree_add_190_195_groupi_n_11633, csa_tree_add_190_195_groupi_n_11634, csa_tree_add_190_195_groupi_n_11635;
  wire csa_tree_add_190_195_groupi_n_11636, csa_tree_add_190_195_groupi_n_11637, csa_tree_add_190_195_groupi_n_11638, csa_tree_add_190_195_groupi_n_11639, csa_tree_add_190_195_groupi_n_11640, csa_tree_add_190_195_groupi_n_11641, csa_tree_add_190_195_groupi_n_11642, csa_tree_add_190_195_groupi_n_11643;
  wire csa_tree_add_190_195_groupi_n_11644, csa_tree_add_190_195_groupi_n_11645, csa_tree_add_190_195_groupi_n_11646, csa_tree_add_190_195_groupi_n_11647, csa_tree_add_190_195_groupi_n_11648, csa_tree_add_190_195_groupi_n_11649, csa_tree_add_190_195_groupi_n_11650, csa_tree_add_190_195_groupi_n_11651;
  wire csa_tree_add_190_195_groupi_n_11652, csa_tree_add_190_195_groupi_n_11653, csa_tree_add_190_195_groupi_n_11654, csa_tree_add_190_195_groupi_n_11655, csa_tree_add_190_195_groupi_n_11656, csa_tree_add_190_195_groupi_n_11657, csa_tree_add_190_195_groupi_n_11658, csa_tree_add_190_195_groupi_n_11659;
  wire csa_tree_add_190_195_groupi_n_11660, csa_tree_add_190_195_groupi_n_11661, csa_tree_add_190_195_groupi_n_11662, csa_tree_add_190_195_groupi_n_11663, csa_tree_add_190_195_groupi_n_11664, csa_tree_add_190_195_groupi_n_11665, csa_tree_add_190_195_groupi_n_11666, csa_tree_add_190_195_groupi_n_11667;
  wire csa_tree_add_190_195_groupi_n_11668, csa_tree_add_190_195_groupi_n_11669, csa_tree_add_190_195_groupi_n_11670, csa_tree_add_190_195_groupi_n_11671, csa_tree_add_190_195_groupi_n_11672, csa_tree_add_190_195_groupi_n_11673, csa_tree_add_190_195_groupi_n_11674, csa_tree_add_190_195_groupi_n_11675;
  wire csa_tree_add_190_195_groupi_n_11676, csa_tree_add_190_195_groupi_n_11677, csa_tree_add_190_195_groupi_n_11678, csa_tree_add_190_195_groupi_n_11679, csa_tree_add_190_195_groupi_n_11680, csa_tree_add_190_195_groupi_n_11681, csa_tree_add_190_195_groupi_n_11682, csa_tree_add_190_195_groupi_n_11683;
  wire csa_tree_add_190_195_groupi_n_11684, csa_tree_add_190_195_groupi_n_11685, csa_tree_add_190_195_groupi_n_11686, csa_tree_add_190_195_groupi_n_11687, csa_tree_add_190_195_groupi_n_11688, csa_tree_add_190_195_groupi_n_11689, csa_tree_add_190_195_groupi_n_11690, csa_tree_add_190_195_groupi_n_11691;
  wire csa_tree_add_190_195_groupi_n_11692, csa_tree_add_190_195_groupi_n_11693, csa_tree_add_190_195_groupi_n_11694, csa_tree_add_190_195_groupi_n_11695, csa_tree_add_190_195_groupi_n_11696, csa_tree_add_190_195_groupi_n_11697, csa_tree_add_190_195_groupi_n_11698, csa_tree_add_190_195_groupi_n_11699;
  wire csa_tree_add_190_195_groupi_n_11700, csa_tree_add_190_195_groupi_n_11701, csa_tree_add_190_195_groupi_n_11702, csa_tree_add_190_195_groupi_n_11703, csa_tree_add_190_195_groupi_n_11704, csa_tree_add_190_195_groupi_n_11705, csa_tree_add_190_195_groupi_n_11706, csa_tree_add_190_195_groupi_n_11707;
  wire csa_tree_add_190_195_groupi_n_11708, csa_tree_add_190_195_groupi_n_11709, csa_tree_add_190_195_groupi_n_11710, csa_tree_add_190_195_groupi_n_11711, csa_tree_add_190_195_groupi_n_11712, csa_tree_add_190_195_groupi_n_11713, csa_tree_add_190_195_groupi_n_11714, csa_tree_add_190_195_groupi_n_11715;
  wire csa_tree_add_190_195_groupi_n_11716, csa_tree_add_190_195_groupi_n_11717, csa_tree_add_190_195_groupi_n_11718, csa_tree_add_190_195_groupi_n_11719, csa_tree_add_190_195_groupi_n_11720, csa_tree_add_190_195_groupi_n_11721, csa_tree_add_190_195_groupi_n_11722, csa_tree_add_190_195_groupi_n_11723;
  wire csa_tree_add_190_195_groupi_n_11724, csa_tree_add_190_195_groupi_n_11725, csa_tree_add_190_195_groupi_n_11726, csa_tree_add_190_195_groupi_n_11727, csa_tree_add_190_195_groupi_n_11728, csa_tree_add_190_195_groupi_n_11729, csa_tree_add_190_195_groupi_n_11730, csa_tree_add_190_195_groupi_n_11731;
  wire csa_tree_add_190_195_groupi_n_11732, csa_tree_add_190_195_groupi_n_11733, csa_tree_add_190_195_groupi_n_11734, csa_tree_add_190_195_groupi_n_11735, csa_tree_add_190_195_groupi_n_11736, csa_tree_add_190_195_groupi_n_11737, csa_tree_add_190_195_groupi_n_11738, csa_tree_add_190_195_groupi_n_11739;
  wire csa_tree_add_190_195_groupi_n_11740, csa_tree_add_190_195_groupi_n_11741, csa_tree_add_190_195_groupi_n_11742, csa_tree_add_190_195_groupi_n_11743, csa_tree_add_190_195_groupi_n_11744, csa_tree_add_190_195_groupi_n_11745, csa_tree_add_190_195_groupi_n_11746, csa_tree_add_190_195_groupi_n_11747;
  wire csa_tree_add_190_195_groupi_n_11748, csa_tree_add_190_195_groupi_n_11749, csa_tree_add_190_195_groupi_n_11750, csa_tree_add_190_195_groupi_n_11751, csa_tree_add_190_195_groupi_n_11752, csa_tree_add_190_195_groupi_n_11753, csa_tree_add_190_195_groupi_n_11754, csa_tree_add_190_195_groupi_n_11755;
  wire csa_tree_add_190_195_groupi_n_11756, csa_tree_add_190_195_groupi_n_11757, csa_tree_add_190_195_groupi_n_11758, csa_tree_add_190_195_groupi_n_11759, csa_tree_add_190_195_groupi_n_11760, csa_tree_add_190_195_groupi_n_11761, csa_tree_add_190_195_groupi_n_11762, csa_tree_add_190_195_groupi_n_11763;
  wire csa_tree_add_190_195_groupi_n_11764, csa_tree_add_190_195_groupi_n_11765, csa_tree_add_190_195_groupi_n_11766, csa_tree_add_190_195_groupi_n_11767, csa_tree_add_190_195_groupi_n_11768, csa_tree_add_190_195_groupi_n_11769, csa_tree_add_190_195_groupi_n_11770, csa_tree_add_190_195_groupi_n_11771;
  wire csa_tree_add_190_195_groupi_n_11772, csa_tree_add_190_195_groupi_n_11773, csa_tree_add_190_195_groupi_n_11774, csa_tree_add_190_195_groupi_n_11775, csa_tree_add_190_195_groupi_n_11776, csa_tree_add_190_195_groupi_n_11777, csa_tree_add_190_195_groupi_n_11778, csa_tree_add_190_195_groupi_n_11779;
  wire csa_tree_add_190_195_groupi_n_11780, csa_tree_add_190_195_groupi_n_11781, csa_tree_add_190_195_groupi_n_11782, csa_tree_add_190_195_groupi_n_11783, csa_tree_add_190_195_groupi_n_11784, csa_tree_add_190_195_groupi_n_11785, csa_tree_add_190_195_groupi_n_11786, csa_tree_add_190_195_groupi_n_11787;
  wire csa_tree_add_190_195_groupi_n_11788, csa_tree_add_190_195_groupi_n_11789, csa_tree_add_190_195_groupi_n_11790, csa_tree_add_190_195_groupi_n_11791, csa_tree_add_190_195_groupi_n_11792, csa_tree_add_190_195_groupi_n_11793, csa_tree_add_190_195_groupi_n_11794, csa_tree_add_190_195_groupi_n_11795;
  wire csa_tree_add_190_195_groupi_n_11796, csa_tree_add_190_195_groupi_n_11797, csa_tree_add_190_195_groupi_n_11798, csa_tree_add_190_195_groupi_n_11799, csa_tree_add_190_195_groupi_n_11800, csa_tree_add_190_195_groupi_n_11801, csa_tree_add_190_195_groupi_n_11802, csa_tree_add_190_195_groupi_n_11803;
  wire csa_tree_add_190_195_groupi_n_11804, csa_tree_add_190_195_groupi_n_11805, csa_tree_add_190_195_groupi_n_11806, csa_tree_add_190_195_groupi_n_11807, csa_tree_add_190_195_groupi_n_11808, csa_tree_add_190_195_groupi_n_11809, csa_tree_add_190_195_groupi_n_11810, csa_tree_add_190_195_groupi_n_11811;
  wire csa_tree_add_190_195_groupi_n_11812, csa_tree_add_190_195_groupi_n_11813, csa_tree_add_190_195_groupi_n_11814, csa_tree_add_190_195_groupi_n_11815, csa_tree_add_190_195_groupi_n_11816, csa_tree_add_190_195_groupi_n_11817, csa_tree_add_190_195_groupi_n_11818, csa_tree_add_190_195_groupi_n_11819;
  wire csa_tree_add_190_195_groupi_n_11820, csa_tree_add_190_195_groupi_n_11821, csa_tree_add_190_195_groupi_n_11822, csa_tree_add_190_195_groupi_n_11823, csa_tree_add_190_195_groupi_n_11824, csa_tree_add_190_195_groupi_n_11825, csa_tree_add_190_195_groupi_n_11826, csa_tree_add_190_195_groupi_n_11827;
  wire csa_tree_add_190_195_groupi_n_11828, csa_tree_add_190_195_groupi_n_11829, csa_tree_add_190_195_groupi_n_11830, csa_tree_add_190_195_groupi_n_11831, csa_tree_add_190_195_groupi_n_11832, csa_tree_add_190_195_groupi_n_11833, csa_tree_add_190_195_groupi_n_11834, csa_tree_add_190_195_groupi_n_11835;
  wire csa_tree_add_190_195_groupi_n_11836, csa_tree_add_190_195_groupi_n_11837, csa_tree_add_190_195_groupi_n_11838, csa_tree_add_190_195_groupi_n_11839, csa_tree_add_190_195_groupi_n_11840, csa_tree_add_190_195_groupi_n_11841, csa_tree_add_190_195_groupi_n_11842, csa_tree_add_190_195_groupi_n_11843;
  wire csa_tree_add_190_195_groupi_n_11844, csa_tree_add_190_195_groupi_n_11845, csa_tree_add_190_195_groupi_n_11846, csa_tree_add_190_195_groupi_n_11847, csa_tree_add_190_195_groupi_n_11848, csa_tree_add_190_195_groupi_n_11849, csa_tree_add_190_195_groupi_n_11850, csa_tree_add_190_195_groupi_n_11851;
  wire csa_tree_add_190_195_groupi_n_11852, csa_tree_add_190_195_groupi_n_11853, csa_tree_add_190_195_groupi_n_11854, csa_tree_add_190_195_groupi_n_11855, csa_tree_add_190_195_groupi_n_11856, csa_tree_add_190_195_groupi_n_11857, csa_tree_add_190_195_groupi_n_11858, csa_tree_add_190_195_groupi_n_11859;
  wire csa_tree_add_190_195_groupi_n_11860, csa_tree_add_190_195_groupi_n_11861, csa_tree_add_190_195_groupi_n_11862, csa_tree_add_190_195_groupi_n_11863, csa_tree_add_190_195_groupi_n_11864, csa_tree_add_190_195_groupi_n_11865, csa_tree_add_190_195_groupi_n_11866, csa_tree_add_190_195_groupi_n_11867;
  wire csa_tree_add_190_195_groupi_n_11868, csa_tree_add_190_195_groupi_n_11869, csa_tree_add_190_195_groupi_n_11870, csa_tree_add_190_195_groupi_n_11871, csa_tree_add_190_195_groupi_n_11872, csa_tree_add_190_195_groupi_n_11873, csa_tree_add_190_195_groupi_n_11874, csa_tree_add_190_195_groupi_n_11875;
  wire csa_tree_add_190_195_groupi_n_11876, csa_tree_add_190_195_groupi_n_11877, csa_tree_add_190_195_groupi_n_11878, csa_tree_add_190_195_groupi_n_11879, csa_tree_add_190_195_groupi_n_11880, csa_tree_add_190_195_groupi_n_11881, csa_tree_add_190_195_groupi_n_11882, csa_tree_add_190_195_groupi_n_11883;
  wire csa_tree_add_190_195_groupi_n_11884, csa_tree_add_190_195_groupi_n_11885, csa_tree_add_190_195_groupi_n_11886, csa_tree_add_190_195_groupi_n_11887, csa_tree_add_190_195_groupi_n_11888, csa_tree_add_190_195_groupi_n_11889, csa_tree_add_190_195_groupi_n_11890, csa_tree_add_190_195_groupi_n_11891;
  wire csa_tree_add_190_195_groupi_n_11892, csa_tree_add_190_195_groupi_n_11893, csa_tree_add_190_195_groupi_n_11894, csa_tree_add_190_195_groupi_n_11895, csa_tree_add_190_195_groupi_n_11896, csa_tree_add_190_195_groupi_n_11897, csa_tree_add_190_195_groupi_n_11898, csa_tree_add_190_195_groupi_n_11899;
  wire csa_tree_add_190_195_groupi_n_11900, csa_tree_add_190_195_groupi_n_11901, csa_tree_add_190_195_groupi_n_11902, csa_tree_add_190_195_groupi_n_11903, csa_tree_add_190_195_groupi_n_11904, csa_tree_add_190_195_groupi_n_11905, csa_tree_add_190_195_groupi_n_11906, csa_tree_add_190_195_groupi_n_11907;
  wire csa_tree_add_190_195_groupi_n_11908, csa_tree_add_190_195_groupi_n_11909, csa_tree_add_190_195_groupi_n_11910, csa_tree_add_190_195_groupi_n_11911, csa_tree_add_190_195_groupi_n_11912, csa_tree_add_190_195_groupi_n_11913, csa_tree_add_190_195_groupi_n_11914, csa_tree_add_190_195_groupi_n_11915;
  wire csa_tree_add_190_195_groupi_n_11916, csa_tree_add_190_195_groupi_n_11917, csa_tree_add_190_195_groupi_n_11918, csa_tree_add_190_195_groupi_n_11919, csa_tree_add_190_195_groupi_n_11920, csa_tree_add_190_195_groupi_n_11921, csa_tree_add_190_195_groupi_n_11922, csa_tree_add_190_195_groupi_n_11923;
  wire csa_tree_add_190_195_groupi_n_11924, csa_tree_add_190_195_groupi_n_11925, csa_tree_add_190_195_groupi_n_11926, csa_tree_add_190_195_groupi_n_11927, csa_tree_add_190_195_groupi_n_11928, csa_tree_add_190_195_groupi_n_11929, csa_tree_add_190_195_groupi_n_11930, csa_tree_add_190_195_groupi_n_11931;
  wire csa_tree_add_190_195_groupi_n_11932, csa_tree_add_190_195_groupi_n_11934, csa_tree_add_190_195_groupi_n_11935, csa_tree_add_190_195_groupi_n_11936, csa_tree_add_190_195_groupi_n_11937, csa_tree_add_190_195_groupi_n_11938, csa_tree_add_190_195_groupi_n_11939, csa_tree_add_190_195_groupi_n_11940;
  wire csa_tree_add_190_195_groupi_n_11941, csa_tree_add_190_195_groupi_n_11942, csa_tree_add_190_195_groupi_n_11943, csa_tree_add_190_195_groupi_n_11944, csa_tree_add_190_195_groupi_n_11945, csa_tree_add_190_195_groupi_n_11946, csa_tree_add_190_195_groupi_n_11947, csa_tree_add_190_195_groupi_n_11948;
  wire csa_tree_add_190_195_groupi_n_11949, csa_tree_add_190_195_groupi_n_11950, csa_tree_add_190_195_groupi_n_11951, csa_tree_add_190_195_groupi_n_11952, csa_tree_add_190_195_groupi_n_11953, csa_tree_add_190_195_groupi_n_11954, csa_tree_add_190_195_groupi_n_11955, csa_tree_add_190_195_groupi_n_11956;
  wire csa_tree_add_190_195_groupi_n_11957, csa_tree_add_190_195_groupi_n_11958, csa_tree_add_190_195_groupi_n_11959, csa_tree_add_190_195_groupi_n_11960, csa_tree_add_190_195_groupi_n_11961, csa_tree_add_190_195_groupi_n_11962, csa_tree_add_190_195_groupi_n_11963, csa_tree_add_190_195_groupi_n_11964;
  wire csa_tree_add_190_195_groupi_n_11965, csa_tree_add_190_195_groupi_n_11966, csa_tree_add_190_195_groupi_n_11967, csa_tree_add_190_195_groupi_n_11968, csa_tree_add_190_195_groupi_n_11969, csa_tree_add_190_195_groupi_n_11970, csa_tree_add_190_195_groupi_n_11971, csa_tree_add_190_195_groupi_n_11972;
  wire csa_tree_add_190_195_groupi_n_11973, csa_tree_add_190_195_groupi_n_11974, csa_tree_add_190_195_groupi_n_11975, csa_tree_add_190_195_groupi_n_11976, csa_tree_add_190_195_groupi_n_11977, csa_tree_add_190_195_groupi_n_11978, csa_tree_add_190_195_groupi_n_11979, csa_tree_add_190_195_groupi_n_11980;
  wire csa_tree_add_190_195_groupi_n_11981, csa_tree_add_190_195_groupi_n_11982, csa_tree_add_190_195_groupi_n_11983, csa_tree_add_190_195_groupi_n_11984, csa_tree_add_190_195_groupi_n_11985, csa_tree_add_190_195_groupi_n_11986, csa_tree_add_190_195_groupi_n_11987, csa_tree_add_190_195_groupi_n_11988;
  wire csa_tree_add_190_195_groupi_n_11989, csa_tree_add_190_195_groupi_n_11990, csa_tree_add_190_195_groupi_n_11991, csa_tree_add_190_195_groupi_n_11992, csa_tree_add_190_195_groupi_n_11993, csa_tree_add_190_195_groupi_n_11994, csa_tree_add_190_195_groupi_n_11995, csa_tree_add_190_195_groupi_n_11996;
  wire csa_tree_add_190_195_groupi_n_11997, csa_tree_add_190_195_groupi_n_11998, csa_tree_add_190_195_groupi_n_11999, csa_tree_add_190_195_groupi_n_12000, csa_tree_add_190_195_groupi_n_12001, csa_tree_add_190_195_groupi_n_12002, csa_tree_add_190_195_groupi_n_12003, csa_tree_add_190_195_groupi_n_12004;
  wire csa_tree_add_190_195_groupi_n_12005, csa_tree_add_190_195_groupi_n_12006, csa_tree_add_190_195_groupi_n_12007, csa_tree_add_190_195_groupi_n_12008, csa_tree_add_190_195_groupi_n_12009, csa_tree_add_190_195_groupi_n_12010, csa_tree_add_190_195_groupi_n_12011, csa_tree_add_190_195_groupi_n_12012;
  wire csa_tree_add_190_195_groupi_n_12013, csa_tree_add_190_195_groupi_n_12014, csa_tree_add_190_195_groupi_n_12015, csa_tree_add_190_195_groupi_n_12016, csa_tree_add_190_195_groupi_n_12017, csa_tree_add_190_195_groupi_n_12018, csa_tree_add_190_195_groupi_n_12019, csa_tree_add_190_195_groupi_n_12020;
  wire csa_tree_add_190_195_groupi_n_12021, csa_tree_add_190_195_groupi_n_12022, csa_tree_add_190_195_groupi_n_12023, csa_tree_add_190_195_groupi_n_12024, csa_tree_add_190_195_groupi_n_12025, csa_tree_add_190_195_groupi_n_12026, csa_tree_add_190_195_groupi_n_12027, csa_tree_add_190_195_groupi_n_12028;
  wire csa_tree_add_190_195_groupi_n_12029, csa_tree_add_190_195_groupi_n_12030, csa_tree_add_190_195_groupi_n_12031, csa_tree_add_190_195_groupi_n_12032, csa_tree_add_190_195_groupi_n_12033, csa_tree_add_190_195_groupi_n_12034, csa_tree_add_190_195_groupi_n_12035, csa_tree_add_190_195_groupi_n_12036;
  wire csa_tree_add_190_195_groupi_n_12037, csa_tree_add_190_195_groupi_n_12038, csa_tree_add_190_195_groupi_n_12039, csa_tree_add_190_195_groupi_n_12040, csa_tree_add_190_195_groupi_n_12041, csa_tree_add_190_195_groupi_n_12042, csa_tree_add_190_195_groupi_n_12043, csa_tree_add_190_195_groupi_n_12044;
  wire csa_tree_add_190_195_groupi_n_12045, csa_tree_add_190_195_groupi_n_12046, csa_tree_add_190_195_groupi_n_12047, csa_tree_add_190_195_groupi_n_12048, csa_tree_add_190_195_groupi_n_12049, csa_tree_add_190_195_groupi_n_12050, csa_tree_add_190_195_groupi_n_12051, csa_tree_add_190_195_groupi_n_12052;
  wire csa_tree_add_190_195_groupi_n_12053, csa_tree_add_190_195_groupi_n_12054, csa_tree_add_190_195_groupi_n_12055, csa_tree_add_190_195_groupi_n_12056, csa_tree_add_190_195_groupi_n_12057, csa_tree_add_190_195_groupi_n_12058, csa_tree_add_190_195_groupi_n_12059, csa_tree_add_190_195_groupi_n_12060;
  wire csa_tree_add_190_195_groupi_n_12061, csa_tree_add_190_195_groupi_n_12062, csa_tree_add_190_195_groupi_n_12063, csa_tree_add_190_195_groupi_n_12064, csa_tree_add_190_195_groupi_n_12065, csa_tree_add_190_195_groupi_n_12066, csa_tree_add_190_195_groupi_n_12067, csa_tree_add_190_195_groupi_n_12068;
  wire csa_tree_add_190_195_groupi_n_12069, csa_tree_add_190_195_groupi_n_12070, csa_tree_add_190_195_groupi_n_12071, csa_tree_add_190_195_groupi_n_12072, csa_tree_add_190_195_groupi_n_12073, csa_tree_add_190_195_groupi_n_12074, csa_tree_add_190_195_groupi_n_12075, csa_tree_add_190_195_groupi_n_12076;
  wire csa_tree_add_190_195_groupi_n_12077, csa_tree_add_190_195_groupi_n_12078, csa_tree_add_190_195_groupi_n_12079, csa_tree_add_190_195_groupi_n_12080, csa_tree_add_190_195_groupi_n_12081, csa_tree_add_190_195_groupi_n_12082, csa_tree_add_190_195_groupi_n_12083, csa_tree_add_190_195_groupi_n_12084;
  wire csa_tree_add_190_195_groupi_n_12085, csa_tree_add_190_195_groupi_n_12086, csa_tree_add_190_195_groupi_n_12087, csa_tree_add_190_195_groupi_n_12088, csa_tree_add_190_195_groupi_n_12089, csa_tree_add_190_195_groupi_n_12090, csa_tree_add_190_195_groupi_n_12091, csa_tree_add_190_195_groupi_n_12092;
  wire csa_tree_add_190_195_groupi_n_12093, csa_tree_add_190_195_groupi_n_12094, csa_tree_add_190_195_groupi_n_12095, csa_tree_add_190_195_groupi_n_12096, csa_tree_add_190_195_groupi_n_12097, csa_tree_add_190_195_groupi_n_12098, csa_tree_add_190_195_groupi_n_12099, csa_tree_add_190_195_groupi_n_12100;
  wire csa_tree_add_190_195_groupi_n_12101, csa_tree_add_190_195_groupi_n_12102, csa_tree_add_190_195_groupi_n_12103, csa_tree_add_190_195_groupi_n_12104, csa_tree_add_190_195_groupi_n_12105, csa_tree_add_190_195_groupi_n_12106, csa_tree_add_190_195_groupi_n_12107, csa_tree_add_190_195_groupi_n_12108;
  wire csa_tree_add_190_195_groupi_n_12109, csa_tree_add_190_195_groupi_n_12110, csa_tree_add_190_195_groupi_n_12111, csa_tree_add_190_195_groupi_n_12112, csa_tree_add_190_195_groupi_n_12113, csa_tree_add_190_195_groupi_n_12114, csa_tree_add_190_195_groupi_n_12115, csa_tree_add_190_195_groupi_n_12116;
  wire csa_tree_add_190_195_groupi_n_12117, csa_tree_add_190_195_groupi_n_12118, csa_tree_add_190_195_groupi_n_12119, csa_tree_add_190_195_groupi_n_12120, csa_tree_add_190_195_groupi_n_12121, csa_tree_add_190_195_groupi_n_12122, csa_tree_add_190_195_groupi_n_12123, csa_tree_add_190_195_groupi_n_12124;
  wire csa_tree_add_190_195_groupi_n_12125, csa_tree_add_190_195_groupi_n_12126, csa_tree_add_190_195_groupi_n_12127, csa_tree_add_190_195_groupi_n_12128, csa_tree_add_190_195_groupi_n_12129, csa_tree_add_190_195_groupi_n_12130, csa_tree_add_190_195_groupi_n_12131, csa_tree_add_190_195_groupi_n_12132;
  wire csa_tree_add_190_195_groupi_n_12133, csa_tree_add_190_195_groupi_n_12134, csa_tree_add_190_195_groupi_n_12135, csa_tree_add_190_195_groupi_n_12136, csa_tree_add_190_195_groupi_n_12137, csa_tree_add_190_195_groupi_n_12138, csa_tree_add_190_195_groupi_n_12139, csa_tree_add_190_195_groupi_n_12140;
  wire csa_tree_add_190_195_groupi_n_12141, csa_tree_add_190_195_groupi_n_12142, csa_tree_add_190_195_groupi_n_12143, csa_tree_add_190_195_groupi_n_12144, csa_tree_add_190_195_groupi_n_12145, csa_tree_add_190_195_groupi_n_12146, csa_tree_add_190_195_groupi_n_12147, csa_tree_add_190_195_groupi_n_12148;
  wire csa_tree_add_190_195_groupi_n_12149, csa_tree_add_190_195_groupi_n_12150, csa_tree_add_190_195_groupi_n_12151, csa_tree_add_190_195_groupi_n_12152, csa_tree_add_190_195_groupi_n_12153, csa_tree_add_190_195_groupi_n_12154, csa_tree_add_190_195_groupi_n_12155, csa_tree_add_190_195_groupi_n_12156;
  wire csa_tree_add_190_195_groupi_n_12157, csa_tree_add_190_195_groupi_n_12158, csa_tree_add_190_195_groupi_n_12159, csa_tree_add_190_195_groupi_n_12160, csa_tree_add_190_195_groupi_n_12161, csa_tree_add_190_195_groupi_n_12162, csa_tree_add_190_195_groupi_n_12163, csa_tree_add_190_195_groupi_n_12164;
  wire csa_tree_add_190_195_groupi_n_12165, csa_tree_add_190_195_groupi_n_12166, csa_tree_add_190_195_groupi_n_12167, csa_tree_add_190_195_groupi_n_12168, csa_tree_add_190_195_groupi_n_12169, csa_tree_add_190_195_groupi_n_12170, csa_tree_add_190_195_groupi_n_12171, csa_tree_add_190_195_groupi_n_12172;
  wire csa_tree_add_190_195_groupi_n_12173, csa_tree_add_190_195_groupi_n_12174, csa_tree_add_190_195_groupi_n_12175, csa_tree_add_190_195_groupi_n_12176, csa_tree_add_190_195_groupi_n_12177, csa_tree_add_190_195_groupi_n_12179, csa_tree_add_190_195_groupi_n_12180, csa_tree_add_190_195_groupi_n_12181;
  wire csa_tree_add_190_195_groupi_n_12182, csa_tree_add_190_195_groupi_n_12183, csa_tree_add_190_195_groupi_n_12184, csa_tree_add_190_195_groupi_n_12185, csa_tree_add_190_195_groupi_n_12186, csa_tree_add_190_195_groupi_n_12187, csa_tree_add_190_195_groupi_n_12188, csa_tree_add_190_195_groupi_n_12189;
  wire csa_tree_add_190_195_groupi_n_12190, csa_tree_add_190_195_groupi_n_12191, csa_tree_add_190_195_groupi_n_12192, csa_tree_add_190_195_groupi_n_12193, csa_tree_add_190_195_groupi_n_12194, csa_tree_add_190_195_groupi_n_12195, csa_tree_add_190_195_groupi_n_12196, csa_tree_add_190_195_groupi_n_12197;
  wire csa_tree_add_190_195_groupi_n_12198, csa_tree_add_190_195_groupi_n_12199, csa_tree_add_190_195_groupi_n_12200, csa_tree_add_190_195_groupi_n_12201, csa_tree_add_190_195_groupi_n_12202, csa_tree_add_190_195_groupi_n_12203, csa_tree_add_190_195_groupi_n_12204, csa_tree_add_190_195_groupi_n_12205;
  wire csa_tree_add_190_195_groupi_n_12206, csa_tree_add_190_195_groupi_n_12207, csa_tree_add_190_195_groupi_n_12208, csa_tree_add_190_195_groupi_n_12209, csa_tree_add_190_195_groupi_n_12210, csa_tree_add_190_195_groupi_n_12211, csa_tree_add_190_195_groupi_n_12212, csa_tree_add_190_195_groupi_n_12213;
  wire csa_tree_add_190_195_groupi_n_12214, csa_tree_add_190_195_groupi_n_12215, csa_tree_add_190_195_groupi_n_12216, csa_tree_add_190_195_groupi_n_12217, csa_tree_add_190_195_groupi_n_12218, csa_tree_add_190_195_groupi_n_12219, csa_tree_add_190_195_groupi_n_12220, csa_tree_add_190_195_groupi_n_12221;
  wire csa_tree_add_190_195_groupi_n_12222, csa_tree_add_190_195_groupi_n_12223, csa_tree_add_190_195_groupi_n_12224, csa_tree_add_190_195_groupi_n_12225, csa_tree_add_190_195_groupi_n_12226, csa_tree_add_190_195_groupi_n_12227, csa_tree_add_190_195_groupi_n_12228, csa_tree_add_190_195_groupi_n_12229;
  wire csa_tree_add_190_195_groupi_n_12230, csa_tree_add_190_195_groupi_n_12232, csa_tree_add_190_195_groupi_n_12233, csa_tree_add_190_195_groupi_n_12234, csa_tree_add_190_195_groupi_n_12235, csa_tree_add_190_195_groupi_n_12236, csa_tree_add_190_195_groupi_n_12237, csa_tree_add_190_195_groupi_n_12238;
  wire csa_tree_add_190_195_groupi_n_12239, csa_tree_add_190_195_groupi_n_12240, csa_tree_add_190_195_groupi_n_12241, csa_tree_add_190_195_groupi_n_12242, csa_tree_add_190_195_groupi_n_12243, csa_tree_add_190_195_groupi_n_12244, csa_tree_add_190_195_groupi_n_12245, csa_tree_add_190_195_groupi_n_12246;
  wire csa_tree_add_190_195_groupi_n_12247, csa_tree_add_190_195_groupi_n_12248, csa_tree_add_190_195_groupi_n_12249, csa_tree_add_190_195_groupi_n_12250, csa_tree_add_190_195_groupi_n_12251, csa_tree_add_190_195_groupi_n_12252, csa_tree_add_190_195_groupi_n_12253, csa_tree_add_190_195_groupi_n_12254;
  wire csa_tree_add_190_195_groupi_n_12255, csa_tree_add_190_195_groupi_n_12256, csa_tree_add_190_195_groupi_n_12257, csa_tree_add_190_195_groupi_n_12258, csa_tree_add_190_195_groupi_n_12259, csa_tree_add_190_195_groupi_n_12260, csa_tree_add_190_195_groupi_n_12261, csa_tree_add_190_195_groupi_n_12262;
  wire csa_tree_add_190_195_groupi_n_12263, csa_tree_add_190_195_groupi_n_12264, csa_tree_add_190_195_groupi_n_12265, csa_tree_add_190_195_groupi_n_12266, csa_tree_add_190_195_groupi_n_12267, csa_tree_add_190_195_groupi_n_12268, csa_tree_add_190_195_groupi_n_12269, csa_tree_add_190_195_groupi_n_12270;
  wire csa_tree_add_190_195_groupi_n_12271, csa_tree_add_190_195_groupi_n_12272, csa_tree_add_190_195_groupi_n_12273, csa_tree_add_190_195_groupi_n_12274, csa_tree_add_190_195_groupi_n_12275, csa_tree_add_190_195_groupi_n_12276, csa_tree_add_190_195_groupi_n_12277, csa_tree_add_190_195_groupi_n_12278;
  wire csa_tree_add_190_195_groupi_n_12279, csa_tree_add_190_195_groupi_n_12280, csa_tree_add_190_195_groupi_n_12281, csa_tree_add_190_195_groupi_n_12282, csa_tree_add_190_195_groupi_n_12283, csa_tree_add_190_195_groupi_n_12284, csa_tree_add_190_195_groupi_n_12285, csa_tree_add_190_195_groupi_n_12286;
  wire csa_tree_add_190_195_groupi_n_12287, csa_tree_add_190_195_groupi_n_12288, csa_tree_add_190_195_groupi_n_12289, csa_tree_add_190_195_groupi_n_12290, csa_tree_add_190_195_groupi_n_12291, csa_tree_add_190_195_groupi_n_12292, csa_tree_add_190_195_groupi_n_12293, csa_tree_add_190_195_groupi_n_12294;
  wire csa_tree_add_190_195_groupi_n_12295, csa_tree_add_190_195_groupi_n_12296, csa_tree_add_190_195_groupi_n_12297, csa_tree_add_190_195_groupi_n_12298, csa_tree_add_190_195_groupi_n_12299, csa_tree_add_190_195_groupi_n_12300, csa_tree_add_190_195_groupi_n_12301, csa_tree_add_190_195_groupi_n_12302;
  wire csa_tree_add_190_195_groupi_n_12303, csa_tree_add_190_195_groupi_n_12304, csa_tree_add_190_195_groupi_n_12305, csa_tree_add_190_195_groupi_n_12306, csa_tree_add_190_195_groupi_n_12307, csa_tree_add_190_195_groupi_n_12308, csa_tree_add_190_195_groupi_n_12309, csa_tree_add_190_195_groupi_n_12310;
  wire csa_tree_add_190_195_groupi_n_12311, csa_tree_add_190_195_groupi_n_12312, csa_tree_add_190_195_groupi_n_12313, csa_tree_add_190_195_groupi_n_12314, csa_tree_add_190_195_groupi_n_12315, csa_tree_add_190_195_groupi_n_12316, csa_tree_add_190_195_groupi_n_12317, csa_tree_add_190_195_groupi_n_12318;
  wire csa_tree_add_190_195_groupi_n_12319, csa_tree_add_190_195_groupi_n_12320, csa_tree_add_190_195_groupi_n_12321, csa_tree_add_190_195_groupi_n_12322, csa_tree_add_190_195_groupi_n_12323, csa_tree_add_190_195_groupi_n_12324, csa_tree_add_190_195_groupi_n_12325, csa_tree_add_190_195_groupi_n_12326;
  wire csa_tree_add_190_195_groupi_n_12327, csa_tree_add_190_195_groupi_n_12328, csa_tree_add_190_195_groupi_n_12329, csa_tree_add_190_195_groupi_n_12330, csa_tree_add_190_195_groupi_n_12331, csa_tree_add_190_195_groupi_n_12332, csa_tree_add_190_195_groupi_n_12333, csa_tree_add_190_195_groupi_n_12334;
  wire csa_tree_add_190_195_groupi_n_12335, csa_tree_add_190_195_groupi_n_12336, csa_tree_add_190_195_groupi_n_12337, csa_tree_add_190_195_groupi_n_12338, csa_tree_add_190_195_groupi_n_12339, csa_tree_add_190_195_groupi_n_12340, csa_tree_add_190_195_groupi_n_12341, csa_tree_add_190_195_groupi_n_12342;
  wire csa_tree_add_190_195_groupi_n_12343, csa_tree_add_190_195_groupi_n_12344, csa_tree_add_190_195_groupi_n_12345, csa_tree_add_190_195_groupi_n_12346, csa_tree_add_190_195_groupi_n_12347, csa_tree_add_190_195_groupi_n_12348, csa_tree_add_190_195_groupi_n_12349, csa_tree_add_190_195_groupi_n_12350;
  wire csa_tree_add_190_195_groupi_n_12351, csa_tree_add_190_195_groupi_n_12352, csa_tree_add_190_195_groupi_n_12353, csa_tree_add_190_195_groupi_n_12354, csa_tree_add_190_195_groupi_n_12355, csa_tree_add_190_195_groupi_n_12356, csa_tree_add_190_195_groupi_n_12357, csa_tree_add_190_195_groupi_n_12358;
  wire csa_tree_add_190_195_groupi_n_12359, csa_tree_add_190_195_groupi_n_12360, csa_tree_add_190_195_groupi_n_12361, csa_tree_add_190_195_groupi_n_12362, csa_tree_add_190_195_groupi_n_12363, csa_tree_add_190_195_groupi_n_12364, csa_tree_add_190_195_groupi_n_12365, csa_tree_add_190_195_groupi_n_12366;
  wire csa_tree_add_190_195_groupi_n_12367, csa_tree_add_190_195_groupi_n_12368, csa_tree_add_190_195_groupi_n_12369, csa_tree_add_190_195_groupi_n_12370, csa_tree_add_190_195_groupi_n_12371, csa_tree_add_190_195_groupi_n_12372, csa_tree_add_190_195_groupi_n_12373, csa_tree_add_190_195_groupi_n_12374;
  wire csa_tree_add_190_195_groupi_n_12375, csa_tree_add_190_195_groupi_n_12376, csa_tree_add_190_195_groupi_n_12377, csa_tree_add_190_195_groupi_n_12378, csa_tree_add_190_195_groupi_n_12379, csa_tree_add_190_195_groupi_n_12380, csa_tree_add_190_195_groupi_n_12382, csa_tree_add_190_195_groupi_n_12383;
  wire csa_tree_add_190_195_groupi_n_12384, csa_tree_add_190_195_groupi_n_12385, csa_tree_add_190_195_groupi_n_12386, csa_tree_add_190_195_groupi_n_12387, csa_tree_add_190_195_groupi_n_12388, csa_tree_add_190_195_groupi_n_12389, csa_tree_add_190_195_groupi_n_12390, csa_tree_add_190_195_groupi_n_12391;
  wire csa_tree_add_190_195_groupi_n_12392, csa_tree_add_190_195_groupi_n_12393, csa_tree_add_190_195_groupi_n_12394, csa_tree_add_190_195_groupi_n_12395, csa_tree_add_190_195_groupi_n_12396, csa_tree_add_190_195_groupi_n_12397, csa_tree_add_190_195_groupi_n_12398, csa_tree_add_190_195_groupi_n_12399;
  wire csa_tree_add_190_195_groupi_n_12400, csa_tree_add_190_195_groupi_n_12401, csa_tree_add_190_195_groupi_n_12402, csa_tree_add_190_195_groupi_n_12403, csa_tree_add_190_195_groupi_n_12404, csa_tree_add_190_195_groupi_n_12405, csa_tree_add_190_195_groupi_n_12406, csa_tree_add_190_195_groupi_n_12407;
  wire csa_tree_add_190_195_groupi_n_12408, csa_tree_add_190_195_groupi_n_12409, csa_tree_add_190_195_groupi_n_12410, csa_tree_add_190_195_groupi_n_12411, csa_tree_add_190_195_groupi_n_12412, csa_tree_add_190_195_groupi_n_12413, csa_tree_add_190_195_groupi_n_12414, csa_tree_add_190_195_groupi_n_12415;
  wire csa_tree_add_190_195_groupi_n_12416, csa_tree_add_190_195_groupi_n_12417, csa_tree_add_190_195_groupi_n_12418, csa_tree_add_190_195_groupi_n_12419, csa_tree_add_190_195_groupi_n_12420, csa_tree_add_190_195_groupi_n_12421, csa_tree_add_190_195_groupi_n_12422, csa_tree_add_190_195_groupi_n_12423;
  wire csa_tree_add_190_195_groupi_n_12424, csa_tree_add_190_195_groupi_n_12425, csa_tree_add_190_195_groupi_n_12426, csa_tree_add_190_195_groupi_n_12427, csa_tree_add_190_195_groupi_n_12428, csa_tree_add_190_195_groupi_n_12429, csa_tree_add_190_195_groupi_n_12430, csa_tree_add_190_195_groupi_n_12431;
  wire csa_tree_add_190_195_groupi_n_12432, csa_tree_add_190_195_groupi_n_12433, csa_tree_add_190_195_groupi_n_12434, csa_tree_add_190_195_groupi_n_12435, csa_tree_add_190_195_groupi_n_12436, csa_tree_add_190_195_groupi_n_12437, csa_tree_add_190_195_groupi_n_12438, csa_tree_add_190_195_groupi_n_12439;
  wire csa_tree_add_190_195_groupi_n_12440, csa_tree_add_190_195_groupi_n_12441, csa_tree_add_190_195_groupi_n_12442, csa_tree_add_190_195_groupi_n_12443, csa_tree_add_190_195_groupi_n_12444, csa_tree_add_190_195_groupi_n_12445, csa_tree_add_190_195_groupi_n_12446, csa_tree_add_190_195_groupi_n_12447;
  wire csa_tree_add_190_195_groupi_n_12448, csa_tree_add_190_195_groupi_n_12449, csa_tree_add_190_195_groupi_n_12450, csa_tree_add_190_195_groupi_n_12451, csa_tree_add_190_195_groupi_n_12452, csa_tree_add_190_195_groupi_n_12453, csa_tree_add_190_195_groupi_n_12454, csa_tree_add_190_195_groupi_n_12455;
  wire csa_tree_add_190_195_groupi_n_12456, csa_tree_add_190_195_groupi_n_12457, csa_tree_add_190_195_groupi_n_12458, csa_tree_add_190_195_groupi_n_12459, csa_tree_add_190_195_groupi_n_12460, csa_tree_add_190_195_groupi_n_12461, csa_tree_add_190_195_groupi_n_12462, csa_tree_add_190_195_groupi_n_12463;
  wire csa_tree_add_190_195_groupi_n_12464, csa_tree_add_190_195_groupi_n_12465, csa_tree_add_190_195_groupi_n_12466, csa_tree_add_190_195_groupi_n_12467, csa_tree_add_190_195_groupi_n_12468, csa_tree_add_190_195_groupi_n_12469, csa_tree_add_190_195_groupi_n_12470, csa_tree_add_190_195_groupi_n_12471;
  wire csa_tree_add_190_195_groupi_n_12472, csa_tree_add_190_195_groupi_n_12473, csa_tree_add_190_195_groupi_n_12474, csa_tree_add_190_195_groupi_n_12475, csa_tree_add_190_195_groupi_n_12476, csa_tree_add_190_195_groupi_n_12477, csa_tree_add_190_195_groupi_n_12478, csa_tree_add_190_195_groupi_n_12479;
  wire csa_tree_add_190_195_groupi_n_12480, csa_tree_add_190_195_groupi_n_12481, csa_tree_add_190_195_groupi_n_12482, csa_tree_add_190_195_groupi_n_12483, csa_tree_add_190_195_groupi_n_12484, csa_tree_add_190_195_groupi_n_12485, csa_tree_add_190_195_groupi_n_12486, csa_tree_add_190_195_groupi_n_12487;
  wire csa_tree_add_190_195_groupi_n_12488, csa_tree_add_190_195_groupi_n_12489, csa_tree_add_190_195_groupi_n_12490, csa_tree_add_190_195_groupi_n_12491, csa_tree_add_190_195_groupi_n_12492, csa_tree_add_190_195_groupi_n_12493, csa_tree_add_190_195_groupi_n_12494, csa_tree_add_190_195_groupi_n_12495;
  wire csa_tree_add_190_195_groupi_n_12496, csa_tree_add_190_195_groupi_n_12497, csa_tree_add_190_195_groupi_n_12498, csa_tree_add_190_195_groupi_n_12499, csa_tree_add_190_195_groupi_n_12500, csa_tree_add_190_195_groupi_n_12501, csa_tree_add_190_195_groupi_n_12502, csa_tree_add_190_195_groupi_n_12503;
  wire csa_tree_add_190_195_groupi_n_12504, csa_tree_add_190_195_groupi_n_12505, csa_tree_add_190_195_groupi_n_12506, csa_tree_add_190_195_groupi_n_12507, csa_tree_add_190_195_groupi_n_12508, csa_tree_add_190_195_groupi_n_12509, csa_tree_add_190_195_groupi_n_12510, csa_tree_add_190_195_groupi_n_12511;
  wire csa_tree_add_190_195_groupi_n_12512, csa_tree_add_190_195_groupi_n_12513, csa_tree_add_190_195_groupi_n_12514, csa_tree_add_190_195_groupi_n_12515, csa_tree_add_190_195_groupi_n_12516, csa_tree_add_190_195_groupi_n_12517, csa_tree_add_190_195_groupi_n_12518, csa_tree_add_190_195_groupi_n_12519;
  wire csa_tree_add_190_195_groupi_n_12520, csa_tree_add_190_195_groupi_n_12521, csa_tree_add_190_195_groupi_n_12522, csa_tree_add_190_195_groupi_n_12523, csa_tree_add_190_195_groupi_n_12524, csa_tree_add_190_195_groupi_n_12525, csa_tree_add_190_195_groupi_n_12526, csa_tree_add_190_195_groupi_n_12527;
  wire csa_tree_add_190_195_groupi_n_12528, csa_tree_add_190_195_groupi_n_12529, csa_tree_add_190_195_groupi_n_12530, csa_tree_add_190_195_groupi_n_12531, csa_tree_add_190_195_groupi_n_12532, csa_tree_add_190_195_groupi_n_12533, csa_tree_add_190_195_groupi_n_12534, csa_tree_add_190_195_groupi_n_12535;
  wire csa_tree_add_190_195_groupi_n_12536, csa_tree_add_190_195_groupi_n_12537, csa_tree_add_190_195_groupi_n_12538, csa_tree_add_190_195_groupi_n_12539, csa_tree_add_190_195_groupi_n_12540, csa_tree_add_190_195_groupi_n_12541, csa_tree_add_190_195_groupi_n_12542, csa_tree_add_190_195_groupi_n_12543;
  wire csa_tree_add_190_195_groupi_n_12544, csa_tree_add_190_195_groupi_n_12545, csa_tree_add_190_195_groupi_n_12546, csa_tree_add_190_195_groupi_n_12547, csa_tree_add_190_195_groupi_n_12548, csa_tree_add_190_195_groupi_n_12549, csa_tree_add_190_195_groupi_n_12550, csa_tree_add_190_195_groupi_n_12551;
  wire csa_tree_add_190_195_groupi_n_12552, csa_tree_add_190_195_groupi_n_12553, csa_tree_add_190_195_groupi_n_12555, csa_tree_add_190_195_groupi_n_12556, csa_tree_add_190_195_groupi_n_12557, csa_tree_add_190_195_groupi_n_12558, csa_tree_add_190_195_groupi_n_12559, csa_tree_add_190_195_groupi_n_12560;
  wire csa_tree_add_190_195_groupi_n_12561, csa_tree_add_190_195_groupi_n_12562, csa_tree_add_190_195_groupi_n_12563, csa_tree_add_190_195_groupi_n_12564, csa_tree_add_190_195_groupi_n_12565, csa_tree_add_190_195_groupi_n_12566, csa_tree_add_190_195_groupi_n_12567, csa_tree_add_190_195_groupi_n_12568;
  wire csa_tree_add_190_195_groupi_n_12569, csa_tree_add_190_195_groupi_n_12570, csa_tree_add_190_195_groupi_n_12571, csa_tree_add_190_195_groupi_n_12572, csa_tree_add_190_195_groupi_n_12573, csa_tree_add_190_195_groupi_n_12574, csa_tree_add_190_195_groupi_n_12575, csa_tree_add_190_195_groupi_n_12576;
  wire csa_tree_add_190_195_groupi_n_12578, csa_tree_add_190_195_groupi_n_12579, csa_tree_add_190_195_groupi_n_12580, csa_tree_add_190_195_groupi_n_12581, csa_tree_add_190_195_groupi_n_12582, csa_tree_add_190_195_groupi_n_12583, csa_tree_add_190_195_groupi_n_12585, csa_tree_add_190_195_groupi_n_12586;
  wire csa_tree_add_190_195_groupi_n_12587, csa_tree_add_190_195_groupi_n_12588, csa_tree_add_190_195_groupi_n_12589, csa_tree_add_190_195_groupi_n_12590, csa_tree_add_190_195_groupi_n_12591, csa_tree_add_190_195_groupi_n_12592, csa_tree_add_190_195_groupi_n_12593, csa_tree_add_190_195_groupi_n_12594;
  wire csa_tree_add_190_195_groupi_n_12595, csa_tree_add_190_195_groupi_n_12596, csa_tree_add_190_195_groupi_n_12597, csa_tree_add_190_195_groupi_n_12598, csa_tree_add_190_195_groupi_n_12599, csa_tree_add_190_195_groupi_n_12600, csa_tree_add_190_195_groupi_n_12601, csa_tree_add_190_195_groupi_n_12602;
  wire csa_tree_add_190_195_groupi_n_12603, csa_tree_add_190_195_groupi_n_12604, csa_tree_add_190_195_groupi_n_12605, csa_tree_add_190_195_groupi_n_12606, csa_tree_add_190_195_groupi_n_12607, csa_tree_add_190_195_groupi_n_12608, csa_tree_add_190_195_groupi_n_12609, csa_tree_add_190_195_groupi_n_12610;
  wire inc_add_191_21_n_1, inc_add_191_21_n_2, inc_add_191_21_n_5, inc_add_191_21_n_6, inc_add_191_21_n_7, inc_add_191_21_n_8, inc_add_191_21_n_9, inc_add_191_21_n_10;
  wire inc_add_191_21_n_11, inc_add_191_21_n_12, inc_add_191_21_n_13, inc_add_191_21_n_14, inc_add_191_21_n_15, inc_add_191_21_n_16, inc_add_191_21_n_17, inc_add_191_21_n_18;
  wire inc_add_191_21_n_19, inc_add_191_21_n_20, inc_add_191_21_n_21, inc_add_191_21_n_22, inc_add_191_21_n_23, inc_add_191_21_n_24, inc_add_191_21_n_25, inc_add_191_21_n_26;
  wire inc_add_191_21_n_27, inc_add_191_21_n_28, inc_add_191_21_n_29, inc_add_191_21_n_30, inc_add_191_21_n_31, inc_add_191_21_n_32, inc_add_191_21_n_33, inc_add_191_21_n_34;
  wire inc_add_191_21_n_36, inc_add_191_21_n_37, inc_add_191_21_n_38, inc_add_191_21_n_39, inc_add_191_21_n_40, inc_add_191_21_n_42, inc_add_191_21_n_43, inc_add_191_21_n_46;
  wire inc_add_191_21_n_47, inc_add_191_21_n_49, inc_add_191_21_n_50, inc_add_191_21_n_51, inc_add_191_21_n_52, inc_add_191_21_n_53, inc_add_191_21_n_55, inc_add_191_21_n_56;
  wire inc_add_191_21_n_57, inc_add_191_21_n_61, inc_add_191_21_n_62, inc_add_191_21_n_66, n_1, n_2, n_3, n_4;
  wire n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12;
  wire n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20;
  wire n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
  wire n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340;
  wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
  wire n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356;
  wire n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364;
  wire n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  wire n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  or add_128_19_g341__2398(n_34 ,add_128_19_n_29 ,add_128_19_n_92);
  xnor add_128_19_g342__5107(n_33 ,add_128_19_n_91 ,add_128_19_n_39);
  nor add_128_19_g343__6260(add_128_19_n_92 ,add_128_19_n_15 ,add_128_19_n_91);
  or add_128_19_g344__4319(add_128_19_n_91 ,add_128_19_n_24 ,add_128_19_n_89);
  xnor add_128_19_g345__8428(n_32 ,add_128_19_n_88 ,add_128_19_n_38);
  and add_128_19_g346__5526(add_128_19_n_89 ,add_128_19_n_9 ,add_128_19_n_88);
  or add_128_19_g347__6783(add_128_19_n_88 ,add_128_19_n_20 ,add_128_19_n_86);
  xnor add_128_19_g348__3680(n_31 ,add_128_19_n_85 ,add_128_19_n_37);
  and add_128_19_g349__1617(add_128_19_n_86 ,add_128_19_n_16 ,add_128_19_n_85);
  or add_128_19_g350__2802(add_128_19_n_85 ,add_128_19_n_10 ,add_128_19_n_83);
  xnor add_128_19_g351__1705(n_30 ,add_128_19_n_82 ,add_128_19_n_36);
  and add_128_19_g352__5122(add_128_19_n_83 ,add_128_19_n_12 ,add_128_19_n_82);
  or add_128_19_g353__8246(add_128_19_n_82 ,add_128_19_n_8 ,add_128_19_n_80);
  xnor add_128_19_g354__7098(n_29 ,add_128_19_n_79 ,add_128_19_n_35);
  and add_128_19_g355__6131(add_128_19_n_80 ,add_128_19_n_22 ,add_128_19_n_79);
  or add_128_19_g356__1881(add_128_19_n_79 ,add_128_19_n_32 ,add_128_19_n_77);
  xnor add_128_19_g357__5115(n_28 ,add_128_19_n_76 ,add_128_19_n_42);
  and add_128_19_g358__7482(add_128_19_n_77 ,add_128_19_n_2 ,add_128_19_n_76);
  or add_128_19_g359__4733(add_128_19_n_76 ,add_128_19_n_21 ,add_128_19_n_74);
  xnor add_128_19_g360__6161(n_27 ,add_128_19_n_73 ,add_128_19_n_48);
  and add_128_19_g361__9315(add_128_19_n_74 ,add_128_19_n_19 ,add_128_19_n_73);
  or add_128_19_g362__9945(add_128_19_n_73 ,add_128_19_n_28 ,add_128_19_n_71);
  xnor add_128_19_g363__2883(n_26 ,add_128_19_n_70 ,add_128_19_n_47);
  and add_128_19_g364__2346(add_128_19_n_71 ,add_128_19_n_11 ,add_128_19_n_70);
  or add_128_19_g365__1666(add_128_19_n_70 ,add_128_19_n_17 ,add_128_19_n_68);
  xnor add_128_19_g366__7410(n_25 ,add_128_19_n_67 ,add_128_19_n_46);
  and add_128_19_g367__6417(add_128_19_n_68 ,add_128_19_n_25 ,add_128_19_n_67);
  or add_128_19_g368__5477(add_128_19_n_67 ,add_128_19_n_6 ,add_128_19_n_65);
  xnor add_128_19_g369__2398(n_24 ,add_128_19_n_64 ,add_128_19_n_45);
  and add_128_19_g370__5107(add_128_19_n_65 ,add_128_19_n_18 ,add_128_19_n_64);
  or add_128_19_g371__6260(add_128_19_n_64 ,add_128_19_n_3 ,add_128_19_n_62);
  xnor add_128_19_g372__4319(n_23 ,add_128_19_n_61 ,add_128_19_n_44);
  and add_128_19_g373__8428(add_128_19_n_62 ,add_128_19_n_30 ,add_128_19_n_61);
  or add_128_19_g374__5526(add_128_19_n_61 ,add_128_19_n_31 ,add_128_19_n_59);
  xnor add_128_19_g375__6783(n_22 ,add_128_19_n_58 ,add_128_19_n_43);
  and add_128_19_g376__3680(add_128_19_n_59 ,add_128_19_n_26 ,add_128_19_n_58);
  or add_128_19_g377__1617(add_128_19_n_58 ,add_128_19_n_27 ,add_128_19_n_56);
  xnor add_128_19_g378__2802(n_21 ,add_128_19_n_55 ,add_128_19_n_34);
  and add_128_19_g379__1705(add_128_19_n_56 ,add_128_19_n_7 ,add_128_19_n_55);
  or add_128_19_g380__5122(add_128_19_n_55 ,add_128_19_n_5 ,add_128_19_n_53);
  xnor add_128_19_g381__8246(n_20 ,add_128_19_n_51 ,add_128_19_n_41);
  and add_128_19_g382__7098(add_128_19_n_53 ,add_128_19_n_23 ,add_128_19_n_51);
  xor add_128_19_g383__6131(n_19 ,add_128_19_n_33 ,add_128_19_n_40);
  or add_128_19_g384__1881(add_128_19_n_51 ,add_128_19_n_4 ,add_128_19_n_49);
  and add_128_19_g385__5115(n_18 ,add_128_19_n_33 ,add_128_19_n_13);
  nor add_128_19_g386__7482(add_128_19_n_49 ,add_128_19_n_33 ,add_128_19_n_14);
  xnor add_128_19_g387__4733(add_128_19_n_48 ,in1[9] ,in2[9]);
  xnor add_128_19_g388__6161(add_128_19_n_47 ,in1[8] ,in2[8]);
  xnor add_128_19_g389__9315(add_128_19_n_46 ,in1[7] ,in2[7]);
  xnor add_128_19_g390__9945(add_128_19_n_45 ,in1[6] ,in2[6]);
  xnor add_128_19_g391__2883(add_128_19_n_44 ,in1[5] ,in2[5]);
  xnor add_128_19_g392__2346(add_128_19_n_43 ,in1[4] ,in2[4]);
  xnor add_128_19_g393__1666(add_128_19_n_42 ,in1[10] ,in2[10]);
  xnor add_128_19_g394__7410(add_128_19_n_41 ,in1[2] ,in2[2]);
  xnor add_128_19_g395__6417(add_128_19_n_40 ,in1[1] ,in2[1]);
  xnor add_128_19_g396__5477(add_128_19_n_39 ,in1[15] ,in2[15]);
  xnor add_128_19_g397__2398(add_128_19_n_38 ,in1[14] ,in2[14]);
  xnor add_128_19_g398__5107(add_128_19_n_37 ,in1[13] ,in2[13]);
  xnor add_128_19_g399__6260(add_128_19_n_36 ,in1[12] ,in2[12]);
  xnor add_128_19_g400__4319(add_128_19_n_35 ,in1[11] ,in2[11]);
  xnor add_128_19_g401__8428(add_128_19_n_34 ,in1[3] ,in2[3]);
  and add_128_19_g402__5526(add_128_19_n_32 ,in1[10] ,in2[10]);
  and add_128_19_g403__6783(add_128_19_n_31 ,in1[4] ,in2[4]);
  or add_128_19_g404__3680(add_128_19_n_30 ,in1[5] ,in2[5]);
  and add_128_19_g405__1617(add_128_19_n_29 ,in1[15] ,in2[15]);
  and add_128_19_g406__2802(add_128_19_n_28 ,in1[8] ,in2[8]);
  and add_128_19_g407__1705(add_128_19_n_27 ,in1[3] ,in2[3]);
  or add_128_19_g408__5122(add_128_19_n_26 ,in1[4] ,in2[4]);
  or add_128_19_g409__8246(add_128_19_n_25 ,in1[7] ,in2[7]);
  and add_128_19_g410__7098(add_128_19_n_24 ,in1[14] ,in2[14]);
  or add_128_19_g411__6131(add_128_19_n_23 ,in1[2] ,in2[2]);
  or add_128_19_g412__1881(add_128_19_n_22 ,in1[11] ,in2[11]);
  and add_128_19_g413__5115(add_128_19_n_21 ,in1[9] ,in2[9]);
  and add_128_19_g414__7482(add_128_19_n_20 ,in1[13] ,in2[13]);
  or add_128_19_g415__4733(add_128_19_n_19 ,in1[9] ,in2[9]);
  or add_128_19_g416__6161(add_128_19_n_18 ,in1[6] ,in2[6]);
  or add_128_19_g417__9315(add_128_19_n_33 ,add_128_19_n_1 ,add_128_19_n_0);
  and add_128_19_g418__9945(add_128_19_n_17 ,in1[7] ,in2[7]);
  or add_128_19_g419__2883(add_128_19_n_16 ,in1[13] ,in2[13]);
  nor add_128_19_g420__2346(add_128_19_n_15 ,in1[15] ,in2[15]);
  nor add_128_19_g421__1666(add_128_19_n_14 ,in1[1] ,in2[1]);
  or add_128_19_g422__7410(add_128_19_n_13 ,in1[0] ,in2[0]);
  or add_128_19_g423__6417(add_128_19_n_12 ,in1[12] ,in2[12]);
  or add_128_19_g424__5477(add_128_19_n_11 ,in1[8] ,in2[8]);
  and add_128_19_g425__2398(add_128_19_n_10 ,in1[12] ,in2[12]);
  or add_128_19_g426__5107(add_128_19_n_9 ,in1[14] ,in2[14]);
  and add_128_19_g427__6260(add_128_19_n_8 ,in1[11] ,in2[11]);
  or add_128_19_g428__4319(add_128_19_n_7 ,in1[3] ,in2[3]);
  and add_128_19_g429__8428(add_128_19_n_6 ,in1[6] ,in2[6]);
  and add_128_19_g430__5526(add_128_19_n_5 ,in1[2] ,in2[2]);
  and add_128_19_g431__6783(add_128_19_n_4 ,in1[1] ,in2[1]);
  and add_128_19_g432__3680(add_128_19_n_3 ,in1[5] ,in2[5]);
  or add_128_19_g433__1617(add_128_19_n_2 ,in1[10] ,in2[10]);
  not add_128_19_g434(add_128_19_n_1 ,in1[0]);
  not add_128_19_g435(add_128_19_n_0 ,in2[0]);
  or add_130_19_g341__2802(n_17 ,add_130_19_n_29 ,add_130_19_n_92);
  xnor add_130_19_g342__1705(n_16 ,add_130_19_n_91 ,add_130_19_n_39);
  nor add_130_19_g343__5122(add_130_19_n_92 ,add_130_19_n_15 ,add_130_19_n_91);
  or add_130_19_g344__8246(add_130_19_n_91 ,add_130_19_n_24 ,add_130_19_n_89);
  xnor add_130_19_g345__7098(n_15 ,add_130_19_n_88 ,add_130_19_n_38);
  and add_130_19_g346__6131(add_130_19_n_89 ,add_130_19_n_9 ,add_130_19_n_88);
  or add_130_19_g347__1881(add_130_19_n_88 ,add_130_19_n_20 ,add_130_19_n_86);
  xnor add_130_19_g348__5115(n_14 ,add_130_19_n_85 ,add_130_19_n_37);
  and add_130_19_g349__7482(add_130_19_n_86 ,add_130_19_n_16 ,add_130_19_n_85);
  or add_130_19_g350__4733(add_130_19_n_85 ,add_130_19_n_10 ,add_130_19_n_83);
  xnor add_130_19_g351__6161(n_13 ,add_130_19_n_82 ,add_130_19_n_36);
  and add_130_19_g352__9315(add_130_19_n_83 ,add_130_19_n_12 ,add_130_19_n_82);
  or add_130_19_g353__9945(add_130_19_n_82 ,add_130_19_n_8 ,add_130_19_n_80);
  xnor add_130_19_g354__2883(n_12 ,add_130_19_n_79 ,add_130_19_n_35);
  and add_130_19_g355__2346(add_130_19_n_80 ,add_130_19_n_22 ,add_130_19_n_79);
  or add_130_19_g356__1666(add_130_19_n_79 ,add_130_19_n_32 ,add_130_19_n_77);
  xnor add_130_19_g357__7410(n_11 ,add_130_19_n_76 ,add_130_19_n_42);
  and add_130_19_g358__6417(add_130_19_n_77 ,add_130_19_n_2 ,add_130_19_n_76);
  or add_130_19_g359__5477(add_130_19_n_76 ,add_130_19_n_21 ,add_130_19_n_74);
  xnor add_130_19_g360__2398(n_10 ,add_130_19_n_73 ,add_130_19_n_48);
  and add_130_19_g361__5107(add_130_19_n_74 ,add_130_19_n_19 ,add_130_19_n_73);
  or add_130_19_g362__6260(add_130_19_n_73 ,add_130_19_n_28 ,add_130_19_n_71);
  xnor add_130_19_g363__4319(n_9 ,add_130_19_n_70 ,add_130_19_n_47);
  and add_130_19_g364__8428(add_130_19_n_71 ,add_130_19_n_11 ,add_130_19_n_70);
  or add_130_19_g365__5526(add_130_19_n_70 ,add_130_19_n_17 ,add_130_19_n_68);
  xnor add_130_19_g366__6783(n_8 ,add_130_19_n_67 ,add_130_19_n_46);
  and add_130_19_g367__3680(add_130_19_n_68 ,add_130_19_n_25 ,add_130_19_n_67);
  or add_130_19_g368__1617(add_130_19_n_67 ,add_130_19_n_6 ,add_130_19_n_65);
  xnor add_130_19_g369__2802(n_7 ,add_130_19_n_64 ,add_130_19_n_45);
  and add_130_19_g370__1705(add_130_19_n_65 ,add_130_19_n_18 ,add_130_19_n_64);
  or add_130_19_g371__5122(add_130_19_n_64 ,add_130_19_n_3 ,add_130_19_n_62);
  xnor add_130_19_g372__8246(n_6 ,add_130_19_n_61 ,add_130_19_n_44);
  and add_130_19_g373__7098(add_130_19_n_62 ,add_130_19_n_30 ,add_130_19_n_61);
  or add_130_19_g374__6131(add_130_19_n_61 ,add_130_19_n_31 ,add_130_19_n_59);
  xnor add_130_19_g375__1881(n_5 ,add_130_19_n_58 ,add_130_19_n_43);
  and add_130_19_g376__5115(add_130_19_n_59 ,add_130_19_n_26 ,add_130_19_n_58);
  or add_130_19_g377__7482(add_130_19_n_58 ,add_130_19_n_27 ,add_130_19_n_56);
  xnor add_130_19_g378__4733(n_4 ,add_130_19_n_55 ,add_130_19_n_34);
  and add_130_19_g379__6161(add_130_19_n_56 ,add_130_19_n_7 ,add_130_19_n_55);
  or add_130_19_g380__9315(add_130_19_n_55 ,add_130_19_n_5 ,add_130_19_n_53);
  xnor add_130_19_g381__9945(n_3 ,add_130_19_n_51 ,add_130_19_n_41);
  and add_130_19_g382__2883(add_130_19_n_53 ,add_130_19_n_23 ,add_130_19_n_51);
  xor add_130_19_g383__2346(n_2 ,add_130_19_n_33 ,add_130_19_n_40);
  or add_130_19_g384__1666(add_130_19_n_51 ,add_130_19_n_4 ,add_130_19_n_49);
  and add_130_19_g385__7410(n_1 ,add_130_19_n_33 ,add_130_19_n_13);
  nor add_130_19_g386__6417(add_130_19_n_49 ,add_130_19_n_33 ,add_130_19_n_14);
  xnor add_130_19_g387__5477(add_130_19_n_48 ,in3[9] ,in4[9]);
  xnor add_130_19_g388__2398(add_130_19_n_47 ,in3[8] ,in4[8]);
  xnor add_130_19_g389__5107(add_130_19_n_46 ,in3[7] ,in4[7]);
  xnor add_130_19_g390__6260(add_130_19_n_45 ,in3[6] ,in4[6]);
  xnor add_130_19_g391__4319(add_130_19_n_44 ,in3[5] ,in4[5]);
  xnor add_130_19_g392__8428(add_130_19_n_43 ,in3[4] ,in4[4]);
  xnor add_130_19_g393__5526(add_130_19_n_42 ,in3[10] ,in4[10]);
  xnor add_130_19_g394__6783(add_130_19_n_41 ,in3[2] ,in4[2]);
  xnor add_130_19_g395__3680(add_130_19_n_40 ,in3[1] ,in4[1]);
  xnor add_130_19_g396__1617(add_130_19_n_39 ,in3[15] ,in4[15]);
  xnor add_130_19_g397__2802(add_130_19_n_38 ,in3[14] ,in4[14]);
  xnor add_130_19_g398__1705(add_130_19_n_37 ,in3[13] ,in4[13]);
  xnor add_130_19_g399__5122(add_130_19_n_36 ,in3[12] ,in4[12]);
  xnor add_130_19_g400__8246(add_130_19_n_35 ,in3[11] ,in4[11]);
  xnor add_130_19_g401__7098(add_130_19_n_34 ,in3[3] ,in4[3]);
  and add_130_19_g402__6131(add_130_19_n_32 ,in3[10] ,in4[10]);
  and add_130_19_g403__1881(add_130_19_n_31 ,in3[4] ,in4[4]);
  or add_130_19_g404__5115(add_130_19_n_30 ,in3[5] ,in4[5]);
  and add_130_19_g405__7482(add_130_19_n_29 ,in3[15] ,in4[15]);
  and add_130_19_g406__4733(add_130_19_n_28 ,in3[8] ,in4[8]);
  and add_130_19_g407__6161(add_130_19_n_27 ,in3[3] ,in4[3]);
  or add_130_19_g408__9315(add_130_19_n_26 ,in3[4] ,in4[4]);
  or add_130_19_g409__9945(add_130_19_n_25 ,in3[7] ,in4[7]);
  and add_130_19_g410__2883(add_130_19_n_24 ,in3[14] ,in4[14]);
  or add_130_19_g411__2346(add_130_19_n_23 ,in3[2] ,in4[2]);
  or add_130_19_g412__1666(add_130_19_n_22 ,in3[11] ,in4[11]);
  and add_130_19_g413__7410(add_130_19_n_21 ,in3[9] ,in4[9]);
  and add_130_19_g414__6417(add_130_19_n_20 ,in3[13] ,in4[13]);
  or add_130_19_g415__5477(add_130_19_n_19 ,in3[9] ,in4[9]);
  or add_130_19_g416__2398(add_130_19_n_18 ,in3[6] ,in4[6]);
  or add_130_19_g417__5107(add_130_19_n_33 ,add_130_19_n_1 ,add_130_19_n_0);
  and add_130_19_g418__6260(add_130_19_n_17 ,in3[7] ,in4[7]);
  or add_130_19_g419__4319(add_130_19_n_16 ,in3[13] ,in4[13]);
  nor add_130_19_g420__8428(add_130_19_n_15 ,in3[15] ,in4[15]);
  nor add_130_19_g421__5526(add_130_19_n_14 ,in3[1] ,in4[1]);
  or add_130_19_g422__6783(add_130_19_n_13 ,in3[0] ,in4[0]);
  or add_130_19_g423__3680(add_130_19_n_12 ,in3[12] ,in4[12]);
  or add_130_19_g424__1617(add_130_19_n_11 ,in3[8] ,in4[8]);
  and add_130_19_g425__2802(add_130_19_n_10 ,in3[12] ,in4[12]);
  or add_130_19_g426__1705(add_130_19_n_9 ,in3[14] ,in4[14]);
  and add_130_19_g427__5122(add_130_19_n_8 ,in3[11] ,in4[11]);
  or add_130_19_g428__8246(add_130_19_n_7 ,in3[3] ,in4[3]);
  and add_130_19_g429__7098(add_130_19_n_6 ,in3[6] ,in4[6]);
  and add_130_19_g430__6131(add_130_19_n_5 ,in3[2] ,in4[2]);
  and add_130_19_g431__1881(add_130_19_n_4 ,in3[1] ,in4[1]);
  and add_130_19_g432__5115(add_130_19_n_3 ,in3[5] ,in4[5]);
  or add_130_19_g433__7482(add_130_19_n_2 ,in3[10] ,in4[10]);
  not add_130_19_g434(add_130_19_n_1 ,in3[0]);
  not add_130_19_g435(add_130_19_n_0 ,in4[0]);
  or add_132_19_g341__4733(n_51 ,add_132_19_n_29 ,add_132_19_n_92);
  xnor add_132_19_g342__6161(n_50 ,add_132_19_n_91 ,add_132_19_n_39);
  nor add_132_19_g343__9315(add_132_19_n_92 ,add_132_19_n_15 ,add_132_19_n_91);
  or add_132_19_g344__9945(add_132_19_n_91 ,add_132_19_n_24 ,add_132_19_n_89);
  xnor add_132_19_g345__2883(n_49 ,add_132_19_n_88 ,add_132_19_n_38);
  and add_132_19_g346__2346(add_132_19_n_89 ,add_132_19_n_9 ,add_132_19_n_88);
  or add_132_19_g347__1666(add_132_19_n_88 ,add_132_19_n_20 ,add_132_19_n_86);
  xnor add_132_19_g348__7410(n_48 ,add_132_19_n_85 ,add_132_19_n_37);
  and add_132_19_g349__6417(add_132_19_n_86 ,add_132_19_n_16 ,add_132_19_n_85);
  or add_132_19_g350__5477(add_132_19_n_85 ,add_132_19_n_10 ,add_132_19_n_83);
  xnor add_132_19_g351__2398(n_47 ,add_132_19_n_82 ,add_132_19_n_36);
  and add_132_19_g352__5107(add_132_19_n_83 ,add_132_19_n_12 ,add_132_19_n_82);
  or add_132_19_g353__6260(add_132_19_n_82 ,add_132_19_n_8 ,add_132_19_n_80);
  xnor add_132_19_g354__4319(n_46 ,add_132_19_n_79 ,add_132_19_n_35);
  and add_132_19_g355__8428(add_132_19_n_80 ,add_132_19_n_22 ,add_132_19_n_79);
  or add_132_19_g356__5526(add_132_19_n_79 ,add_132_19_n_32 ,add_132_19_n_77);
  xnor add_132_19_g357__6783(n_45 ,add_132_19_n_76 ,add_132_19_n_42);
  and add_132_19_g358__3680(add_132_19_n_77 ,add_132_19_n_2 ,add_132_19_n_76);
  or add_132_19_g359__1617(add_132_19_n_76 ,add_132_19_n_21 ,add_132_19_n_74);
  xnor add_132_19_g360__2802(n_44 ,add_132_19_n_73 ,add_132_19_n_48);
  and add_132_19_g361__1705(add_132_19_n_74 ,add_132_19_n_19 ,add_132_19_n_73);
  or add_132_19_g362__5122(add_132_19_n_73 ,add_132_19_n_28 ,add_132_19_n_71);
  xnor add_132_19_g363__8246(n_43 ,add_132_19_n_70 ,add_132_19_n_47);
  and add_132_19_g364__7098(add_132_19_n_71 ,add_132_19_n_11 ,add_132_19_n_70);
  or add_132_19_g365__6131(add_132_19_n_70 ,add_132_19_n_17 ,add_132_19_n_68);
  xnor add_132_19_g366__1881(n_42 ,add_132_19_n_67 ,add_132_19_n_46);
  and add_132_19_g367__5115(add_132_19_n_68 ,add_132_19_n_25 ,add_132_19_n_67);
  or add_132_19_g368__7482(add_132_19_n_67 ,add_132_19_n_6 ,add_132_19_n_65);
  xnor add_132_19_g369__4733(n_41 ,add_132_19_n_64 ,add_132_19_n_45);
  and add_132_19_g370__6161(add_132_19_n_65 ,add_132_19_n_18 ,add_132_19_n_64);
  or add_132_19_g371__9315(add_132_19_n_64 ,add_132_19_n_3 ,add_132_19_n_62);
  xnor add_132_19_g372__9945(n_40 ,add_132_19_n_61 ,add_132_19_n_44);
  and add_132_19_g373__2883(add_132_19_n_62 ,add_132_19_n_30 ,add_132_19_n_61);
  or add_132_19_g374__2346(add_132_19_n_61 ,add_132_19_n_31 ,add_132_19_n_59);
  xnor add_132_19_g375__1666(n_39 ,add_132_19_n_58 ,add_132_19_n_43);
  and add_132_19_g376__7410(add_132_19_n_59 ,add_132_19_n_26 ,add_132_19_n_58);
  or add_132_19_g377__6417(add_132_19_n_58 ,add_132_19_n_27 ,add_132_19_n_56);
  xnor add_132_19_g378__5477(n_38 ,add_132_19_n_55 ,add_132_19_n_34);
  and add_132_19_g379__2398(add_132_19_n_56 ,add_132_19_n_7 ,add_132_19_n_55);
  or add_132_19_g380__5107(add_132_19_n_55 ,add_132_19_n_5 ,add_132_19_n_53);
  xnor add_132_19_g381__6260(n_37 ,add_132_19_n_51 ,add_132_19_n_41);
  and add_132_19_g382__4319(add_132_19_n_53 ,add_132_19_n_23 ,add_132_19_n_51);
  xor add_132_19_g383__8428(n_36 ,add_132_19_n_33 ,add_132_19_n_40);
  or add_132_19_g384__5526(add_132_19_n_51 ,add_132_19_n_4 ,add_132_19_n_49);
  and add_132_19_g385__6783(n_35 ,add_132_19_n_33 ,add_132_19_n_13);
  nor add_132_19_g386__3680(add_132_19_n_49 ,add_132_19_n_33 ,add_132_19_n_14);
  xnor add_132_19_g387__1617(add_132_19_n_48 ,in5[9] ,in6[9]);
  xnor add_132_19_g388__2802(add_132_19_n_47 ,in5[8] ,in6[8]);
  xnor add_132_19_g389__1705(add_132_19_n_46 ,in5[7] ,in6[7]);
  xnor add_132_19_g390__5122(add_132_19_n_45 ,in5[6] ,in6[6]);
  xnor add_132_19_g391__8246(add_132_19_n_44 ,in5[5] ,in6[5]);
  xnor add_132_19_g392__7098(add_132_19_n_43 ,in5[4] ,in6[4]);
  xnor add_132_19_g393__6131(add_132_19_n_42 ,in5[10] ,in6[10]);
  xnor add_132_19_g394__1881(add_132_19_n_41 ,in5[2] ,in6[2]);
  xnor add_132_19_g395__5115(add_132_19_n_40 ,in5[1] ,in6[1]);
  xnor add_132_19_g396__7482(add_132_19_n_39 ,in5[15] ,in6[15]);
  xnor add_132_19_g397__4733(add_132_19_n_38 ,in5[14] ,in6[14]);
  xnor add_132_19_g398__6161(add_132_19_n_37 ,in5[13] ,in6[13]);
  xnor add_132_19_g399__9315(add_132_19_n_36 ,in5[12] ,in6[12]);
  xnor add_132_19_g400__9945(add_132_19_n_35 ,in5[11] ,in6[11]);
  xnor add_132_19_g401__2883(add_132_19_n_34 ,in5[3] ,in6[3]);
  and add_132_19_g402__2346(add_132_19_n_32 ,in5[10] ,in6[10]);
  and add_132_19_g403__1666(add_132_19_n_31 ,in5[4] ,in6[4]);
  or add_132_19_g404__7410(add_132_19_n_30 ,in5[5] ,in6[5]);
  and add_132_19_g405__6417(add_132_19_n_29 ,in5[15] ,in6[15]);
  and add_132_19_g406__5477(add_132_19_n_28 ,in5[8] ,in6[8]);
  and add_132_19_g407__2398(add_132_19_n_27 ,in5[3] ,in6[3]);
  or add_132_19_g408__5107(add_132_19_n_26 ,in5[4] ,in6[4]);
  or add_132_19_g409__6260(add_132_19_n_25 ,in5[7] ,in6[7]);
  and add_132_19_g410__4319(add_132_19_n_24 ,in5[14] ,in6[14]);
  or add_132_19_g411__8428(add_132_19_n_23 ,in5[2] ,in6[2]);
  or add_132_19_g412__5526(add_132_19_n_22 ,in5[11] ,in6[11]);
  and add_132_19_g413__6783(add_132_19_n_21 ,in5[9] ,in6[9]);
  and add_132_19_g414__3680(add_132_19_n_20 ,in5[13] ,in6[13]);
  or add_132_19_g415__1617(add_132_19_n_19 ,in5[9] ,in6[9]);
  or add_132_19_g416__2802(add_132_19_n_18 ,in5[6] ,in6[6]);
  or add_132_19_g417__1705(add_132_19_n_33 ,add_132_19_n_1 ,add_132_19_n_0);
  and add_132_19_g418__5122(add_132_19_n_17 ,in5[7] ,in6[7]);
  or add_132_19_g419__8246(add_132_19_n_16 ,in5[13] ,in6[13]);
  nor add_132_19_g420__7098(add_132_19_n_15 ,in5[15] ,in6[15]);
  nor add_132_19_g421__6131(add_132_19_n_14 ,in5[1] ,in6[1]);
  or add_132_19_g422__1881(add_132_19_n_13 ,in5[0] ,in6[0]);
  or add_132_19_g423__5115(add_132_19_n_12 ,in5[12] ,in6[12]);
  or add_132_19_g424__7482(add_132_19_n_11 ,in5[8] ,in6[8]);
  and add_132_19_g425__4733(add_132_19_n_10 ,in5[12] ,in6[12]);
  or add_132_19_g426__6161(add_132_19_n_9 ,in5[14] ,in6[14]);
  and add_132_19_g427__9315(add_132_19_n_8 ,in5[11] ,in6[11]);
  or add_132_19_g428__9945(add_132_19_n_7 ,in5[3] ,in6[3]);
  and add_132_19_g429__2883(add_132_19_n_6 ,in5[6] ,in6[6]);
  and add_132_19_g430__2346(add_132_19_n_5 ,in5[2] ,in6[2]);
  and add_132_19_g431__1666(add_132_19_n_4 ,in5[1] ,in6[1]);
  and add_132_19_g432__7410(add_132_19_n_3 ,in5[5] ,in6[5]);
  or add_132_19_g433__6417(add_132_19_n_2 ,in5[10] ,in6[10]);
  not add_132_19_g434(add_132_19_n_1 ,in5[0]);
  not add_132_19_g435(add_132_19_n_0 ,in6[0]);
  or add_134_19_g341__5477(n_68 ,add_134_19_n_29 ,add_134_19_n_92);
  xnor add_134_19_g342__2398(n_67 ,add_134_19_n_91 ,add_134_19_n_39);
  nor add_134_19_g343__5107(add_134_19_n_92 ,add_134_19_n_15 ,add_134_19_n_91);
  or add_134_19_g344__6260(add_134_19_n_91 ,add_134_19_n_24 ,add_134_19_n_89);
  xnor add_134_19_g345__4319(n_66 ,add_134_19_n_88 ,add_134_19_n_38);
  and add_134_19_g346__8428(add_134_19_n_89 ,add_134_19_n_9 ,add_134_19_n_88);
  or add_134_19_g347__5526(add_134_19_n_88 ,add_134_19_n_20 ,add_134_19_n_86);
  xnor add_134_19_g348__6783(n_65 ,add_134_19_n_85 ,add_134_19_n_37);
  and add_134_19_g349__3680(add_134_19_n_86 ,add_134_19_n_16 ,add_134_19_n_85);
  or add_134_19_g350__1617(add_134_19_n_85 ,add_134_19_n_10 ,add_134_19_n_83);
  xnor add_134_19_g351__2802(n_64 ,add_134_19_n_82 ,add_134_19_n_36);
  and add_134_19_g352__1705(add_134_19_n_83 ,add_134_19_n_12 ,add_134_19_n_82);
  or add_134_19_g353__5122(add_134_19_n_82 ,add_134_19_n_8 ,add_134_19_n_80);
  xnor add_134_19_g354__8246(n_63 ,add_134_19_n_79 ,add_134_19_n_35);
  and add_134_19_g355__7098(add_134_19_n_80 ,add_134_19_n_22 ,add_134_19_n_79);
  or add_134_19_g356__6131(add_134_19_n_79 ,add_134_19_n_32 ,add_134_19_n_77);
  xnor add_134_19_g357__1881(n_62 ,add_134_19_n_76 ,add_134_19_n_42);
  and add_134_19_g358__5115(add_134_19_n_77 ,add_134_19_n_2 ,add_134_19_n_76);
  or add_134_19_g359__7482(add_134_19_n_76 ,add_134_19_n_21 ,add_134_19_n_74);
  xnor add_134_19_g360__4733(n_61 ,add_134_19_n_73 ,add_134_19_n_48);
  and add_134_19_g361__6161(add_134_19_n_74 ,add_134_19_n_19 ,add_134_19_n_73);
  or add_134_19_g362__9315(add_134_19_n_73 ,add_134_19_n_28 ,add_134_19_n_71);
  xnor add_134_19_g363__9945(n_60 ,add_134_19_n_70 ,add_134_19_n_47);
  and add_134_19_g364__2883(add_134_19_n_71 ,add_134_19_n_11 ,add_134_19_n_70);
  or add_134_19_g365__2346(add_134_19_n_70 ,add_134_19_n_17 ,add_134_19_n_68);
  xnor add_134_19_g366__1666(n_59 ,add_134_19_n_67 ,add_134_19_n_46);
  and add_134_19_g367__7410(add_134_19_n_68 ,add_134_19_n_25 ,add_134_19_n_67);
  or add_134_19_g368__6417(add_134_19_n_67 ,add_134_19_n_6 ,add_134_19_n_65);
  xnor add_134_19_g369__5477(n_58 ,add_134_19_n_64 ,add_134_19_n_45);
  and add_134_19_g370__2398(add_134_19_n_65 ,add_134_19_n_18 ,add_134_19_n_64);
  or add_134_19_g371__5107(add_134_19_n_64 ,add_134_19_n_3 ,add_134_19_n_62);
  xnor add_134_19_g372__6260(n_57 ,add_134_19_n_61 ,add_134_19_n_44);
  and add_134_19_g373__4319(add_134_19_n_62 ,add_134_19_n_30 ,add_134_19_n_61);
  or add_134_19_g374__8428(add_134_19_n_61 ,add_134_19_n_31 ,add_134_19_n_59);
  xnor add_134_19_g375__5526(n_56 ,add_134_19_n_58 ,add_134_19_n_43);
  and add_134_19_g376__6783(add_134_19_n_59 ,add_134_19_n_26 ,add_134_19_n_58);
  or add_134_19_g377__3680(add_134_19_n_58 ,add_134_19_n_27 ,add_134_19_n_56);
  xnor add_134_19_g378__1617(n_55 ,add_134_19_n_55 ,add_134_19_n_34);
  and add_134_19_g379__2802(add_134_19_n_56 ,add_134_19_n_7 ,add_134_19_n_55);
  or add_134_19_g380__1705(add_134_19_n_55 ,add_134_19_n_5 ,add_134_19_n_53);
  xnor add_134_19_g381__5122(n_54 ,add_134_19_n_51 ,add_134_19_n_41);
  and add_134_19_g382__8246(add_134_19_n_53 ,add_134_19_n_23 ,add_134_19_n_51);
  xor add_134_19_g383__7098(n_53 ,add_134_19_n_33 ,add_134_19_n_40);
  or add_134_19_g384__6131(add_134_19_n_51 ,add_134_19_n_4 ,add_134_19_n_49);
  and add_134_19_g385__1881(n_52 ,add_134_19_n_33 ,add_134_19_n_13);
  nor add_134_19_g386__5115(add_134_19_n_49 ,add_134_19_n_33 ,add_134_19_n_14);
  xnor add_134_19_g387__7482(add_134_19_n_48 ,in7[9] ,in8[9]);
  xnor add_134_19_g388__4733(add_134_19_n_47 ,in7[8] ,in8[8]);
  xnor add_134_19_g389__6161(add_134_19_n_46 ,in7[7] ,in8[7]);
  xnor add_134_19_g390__9315(add_134_19_n_45 ,in7[6] ,in8[6]);
  xnor add_134_19_g391__9945(add_134_19_n_44 ,in7[5] ,in8[5]);
  xnor add_134_19_g392__2883(add_134_19_n_43 ,in7[4] ,in8[4]);
  xnor add_134_19_g393__2346(add_134_19_n_42 ,in7[10] ,in8[10]);
  xnor add_134_19_g394__1666(add_134_19_n_41 ,in7[2] ,in8[2]);
  xnor add_134_19_g395__7410(add_134_19_n_40 ,in7[1] ,in8[1]);
  xnor add_134_19_g396__6417(add_134_19_n_39 ,in7[15] ,in8[15]);
  xnor add_134_19_g397__5477(add_134_19_n_38 ,in7[14] ,in8[14]);
  xnor add_134_19_g398__2398(add_134_19_n_37 ,in7[13] ,in8[13]);
  xnor add_134_19_g399__5107(add_134_19_n_36 ,in7[12] ,in8[12]);
  xnor add_134_19_g400__6260(add_134_19_n_35 ,in7[11] ,in8[11]);
  xnor add_134_19_g401__4319(add_134_19_n_34 ,in7[3] ,in8[3]);
  and add_134_19_g402__8428(add_134_19_n_32 ,in7[10] ,in8[10]);
  and add_134_19_g403__5526(add_134_19_n_31 ,in7[4] ,in8[4]);
  or add_134_19_g404__6783(add_134_19_n_30 ,in7[5] ,in8[5]);
  and add_134_19_g405__3680(add_134_19_n_29 ,in7[15] ,in8[15]);
  and add_134_19_g406__1617(add_134_19_n_28 ,in7[8] ,in8[8]);
  and add_134_19_g407__2802(add_134_19_n_27 ,in7[3] ,in8[3]);
  or add_134_19_g408__1705(add_134_19_n_26 ,in7[4] ,in8[4]);
  or add_134_19_g409__5122(add_134_19_n_25 ,in7[7] ,in8[7]);
  and add_134_19_g410__8246(add_134_19_n_24 ,in7[14] ,in8[14]);
  or add_134_19_g411__7098(add_134_19_n_23 ,in7[2] ,in8[2]);
  or add_134_19_g412__6131(add_134_19_n_22 ,in7[11] ,in8[11]);
  and add_134_19_g413__1881(add_134_19_n_21 ,in7[9] ,in8[9]);
  and add_134_19_g414__5115(add_134_19_n_20 ,in7[13] ,in8[13]);
  or add_134_19_g415__7482(add_134_19_n_19 ,in7[9] ,in8[9]);
  or add_134_19_g416__4733(add_134_19_n_18 ,in7[6] ,in8[6]);
  or add_134_19_g417__6161(add_134_19_n_33 ,add_134_19_n_1 ,add_134_19_n_0);
  and add_134_19_g418__9315(add_134_19_n_17 ,in7[7] ,in8[7]);
  or add_134_19_g419__9945(add_134_19_n_16 ,in7[13] ,in8[13]);
  nor add_134_19_g420__2883(add_134_19_n_15 ,in7[15] ,in8[15]);
  nor add_134_19_g421__2346(add_134_19_n_14 ,in7[1] ,in8[1]);
  or add_134_19_g422__1666(add_134_19_n_13 ,in7[0] ,in8[0]);
  or add_134_19_g423__7410(add_134_19_n_12 ,in7[12] ,in8[12]);
  or add_134_19_g424__6417(add_134_19_n_11 ,in7[8] ,in8[8]);
  and add_134_19_g425__5477(add_134_19_n_10 ,in7[12] ,in8[12]);
  or add_134_19_g426__2398(add_134_19_n_9 ,in7[14] ,in8[14]);
  and add_134_19_g427__5107(add_134_19_n_8 ,in7[11] ,in8[11]);
  or add_134_19_g428__6260(add_134_19_n_7 ,in7[3] ,in8[3]);
  and add_134_19_g429__4319(add_134_19_n_6 ,in7[6] ,in8[6]);
  and add_134_19_g430__8428(add_134_19_n_5 ,in7[2] ,in8[2]);
  and add_134_19_g431__5526(add_134_19_n_4 ,in7[1] ,in8[1]);
  and add_134_19_g432__6783(add_134_19_n_3 ,in7[5] ,in8[5]);
  or add_134_19_g433__3680(add_134_19_n_2 ,in7[10] ,in8[10]);
  not add_134_19_g434(add_134_19_n_1 ,in7[0]);
  not add_134_19_g435(add_134_19_n_0 ,in8[0]);
  or add_136_19_g341__1617(n_85 ,add_136_19_n_29 ,add_136_19_n_92);
  xnor add_136_19_g342__2802(n_84 ,add_136_19_n_91 ,add_136_19_n_39);
  nor add_136_19_g343__1705(add_136_19_n_92 ,add_136_19_n_15 ,add_136_19_n_91);
  or add_136_19_g344__5122(add_136_19_n_91 ,add_136_19_n_24 ,add_136_19_n_89);
  xnor add_136_19_g345__8246(n_83 ,add_136_19_n_88 ,add_136_19_n_38);
  and add_136_19_g346__7098(add_136_19_n_89 ,add_136_19_n_9 ,add_136_19_n_88);
  or add_136_19_g347__6131(add_136_19_n_88 ,add_136_19_n_20 ,add_136_19_n_86);
  xnor add_136_19_g348__1881(n_82 ,add_136_19_n_85 ,add_136_19_n_37);
  and add_136_19_g349__5115(add_136_19_n_86 ,add_136_19_n_16 ,add_136_19_n_85);
  or add_136_19_g350__7482(add_136_19_n_85 ,add_136_19_n_10 ,add_136_19_n_83);
  xnor add_136_19_g351__4733(n_81 ,add_136_19_n_82 ,add_136_19_n_36);
  and add_136_19_g352__6161(add_136_19_n_83 ,add_136_19_n_12 ,add_136_19_n_82);
  or add_136_19_g353__9315(add_136_19_n_82 ,add_136_19_n_8 ,add_136_19_n_80);
  xnor add_136_19_g354__9945(n_80 ,add_136_19_n_79 ,add_136_19_n_35);
  and add_136_19_g355__2883(add_136_19_n_80 ,add_136_19_n_22 ,add_136_19_n_79);
  or add_136_19_g356__2346(add_136_19_n_79 ,add_136_19_n_32 ,add_136_19_n_77);
  xnor add_136_19_g357__1666(n_79 ,add_136_19_n_76 ,add_136_19_n_42);
  and add_136_19_g358__7410(add_136_19_n_77 ,add_136_19_n_2 ,add_136_19_n_76);
  or add_136_19_g359__6417(add_136_19_n_76 ,add_136_19_n_21 ,add_136_19_n_74);
  xnor add_136_19_g360__5477(n_78 ,add_136_19_n_73 ,add_136_19_n_48);
  and add_136_19_g361__2398(add_136_19_n_74 ,add_136_19_n_19 ,add_136_19_n_73);
  or add_136_19_g362__5107(add_136_19_n_73 ,add_136_19_n_28 ,add_136_19_n_71);
  xnor add_136_19_g363__6260(n_77 ,add_136_19_n_70 ,add_136_19_n_47);
  and add_136_19_g364__4319(add_136_19_n_71 ,add_136_19_n_11 ,add_136_19_n_70);
  or add_136_19_g365__8428(add_136_19_n_70 ,add_136_19_n_17 ,add_136_19_n_68);
  xnor add_136_19_g366__5526(n_76 ,add_136_19_n_67 ,add_136_19_n_46);
  and add_136_19_g367__6783(add_136_19_n_68 ,add_136_19_n_25 ,add_136_19_n_67);
  or add_136_19_g368__3680(add_136_19_n_67 ,add_136_19_n_6 ,add_136_19_n_65);
  xnor add_136_19_g369__1617(n_75 ,add_136_19_n_64 ,add_136_19_n_45);
  and add_136_19_g370__2802(add_136_19_n_65 ,add_136_19_n_18 ,add_136_19_n_64);
  or add_136_19_g371__1705(add_136_19_n_64 ,add_136_19_n_3 ,add_136_19_n_62);
  xnor add_136_19_g372__5122(n_74 ,add_136_19_n_61 ,add_136_19_n_44);
  and add_136_19_g373__8246(add_136_19_n_62 ,add_136_19_n_30 ,add_136_19_n_61);
  or add_136_19_g374__7098(add_136_19_n_61 ,add_136_19_n_31 ,add_136_19_n_59);
  xnor add_136_19_g375__6131(n_73 ,add_136_19_n_58 ,add_136_19_n_43);
  and add_136_19_g376__1881(add_136_19_n_59 ,add_136_19_n_26 ,add_136_19_n_58);
  or add_136_19_g377__5115(add_136_19_n_58 ,add_136_19_n_27 ,add_136_19_n_56);
  xnor add_136_19_g378__7482(n_72 ,add_136_19_n_55 ,add_136_19_n_34);
  and add_136_19_g379__4733(add_136_19_n_56 ,add_136_19_n_7 ,add_136_19_n_55);
  or add_136_19_g380__6161(add_136_19_n_55 ,add_136_19_n_5 ,add_136_19_n_53);
  xnor add_136_19_g381__9315(n_71 ,add_136_19_n_51 ,add_136_19_n_41);
  and add_136_19_g382__9945(add_136_19_n_53 ,add_136_19_n_23 ,add_136_19_n_51);
  xor add_136_19_g383__2883(n_70 ,add_136_19_n_33 ,add_136_19_n_40);
  or add_136_19_g384__2346(add_136_19_n_51 ,add_136_19_n_4 ,add_136_19_n_49);
  and add_136_19_g385__1666(n_69 ,add_136_19_n_33 ,add_136_19_n_13);
  nor add_136_19_g386__7410(add_136_19_n_49 ,add_136_19_n_33 ,add_136_19_n_14);
  xnor add_136_19_g387__6417(add_136_19_n_48 ,in9[9] ,in10[9]);
  xnor add_136_19_g388__5477(add_136_19_n_47 ,in9[8] ,in10[8]);
  xnor add_136_19_g389__2398(add_136_19_n_46 ,in9[7] ,in10[7]);
  xnor add_136_19_g390__5107(add_136_19_n_45 ,in9[6] ,in10[6]);
  xnor add_136_19_g391__6260(add_136_19_n_44 ,in9[5] ,in10[5]);
  xnor add_136_19_g392__4319(add_136_19_n_43 ,in9[4] ,in10[4]);
  xnor add_136_19_g393__8428(add_136_19_n_42 ,in9[10] ,in10[10]);
  xnor add_136_19_g394__5526(add_136_19_n_41 ,in9[2] ,in10[2]);
  xnor add_136_19_g395__6783(add_136_19_n_40 ,in9[1] ,in10[1]);
  xnor add_136_19_g396__3680(add_136_19_n_39 ,in9[15] ,in10[15]);
  xnor add_136_19_g397__1617(add_136_19_n_38 ,in9[14] ,in10[14]);
  xnor add_136_19_g398__2802(add_136_19_n_37 ,in9[13] ,in10[13]);
  xnor add_136_19_g399__1705(add_136_19_n_36 ,in9[12] ,in10[12]);
  xnor add_136_19_g400__5122(add_136_19_n_35 ,in9[11] ,in10[11]);
  xnor add_136_19_g401__8246(add_136_19_n_34 ,in9[3] ,in10[3]);
  and add_136_19_g402__7098(add_136_19_n_32 ,in9[10] ,in10[10]);
  and add_136_19_g403__6131(add_136_19_n_31 ,in9[4] ,in10[4]);
  or add_136_19_g404__1881(add_136_19_n_30 ,in9[5] ,in10[5]);
  and add_136_19_g405__5115(add_136_19_n_29 ,in9[15] ,in10[15]);
  and add_136_19_g406__7482(add_136_19_n_28 ,in9[8] ,in10[8]);
  and add_136_19_g407__4733(add_136_19_n_27 ,in9[3] ,in10[3]);
  or add_136_19_g408__6161(add_136_19_n_26 ,in9[4] ,in10[4]);
  or add_136_19_g409__9315(add_136_19_n_25 ,in9[7] ,in10[7]);
  and add_136_19_g410__9945(add_136_19_n_24 ,in9[14] ,in10[14]);
  or add_136_19_g411__2883(add_136_19_n_23 ,in9[2] ,in10[2]);
  or add_136_19_g412__2346(add_136_19_n_22 ,in9[11] ,in10[11]);
  and add_136_19_g413__1666(add_136_19_n_21 ,in9[9] ,in10[9]);
  and add_136_19_g414__7410(add_136_19_n_20 ,in9[13] ,in10[13]);
  or add_136_19_g415__6417(add_136_19_n_19 ,in9[9] ,in10[9]);
  or add_136_19_g416__5477(add_136_19_n_18 ,in9[6] ,in10[6]);
  or add_136_19_g417__2398(add_136_19_n_33 ,add_136_19_n_1 ,add_136_19_n_0);
  and add_136_19_g418__5107(add_136_19_n_17 ,in9[7] ,in10[7]);
  or add_136_19_g419__6260(add_136_19_n_16 ,in9[13] ,in10[13]);
  nor add_136_19_g420__4319(add_136_19_n_15 ,in9[15] ,in10[15]);
  nor add_136_19_g421__8428(add_136_19_n_14 ,in9[1] ,in10[1]);
  or add_136_19_g422__5526(add_136_19_n_13 ,in9[0] ,in10[0]);
  or add_136_19_g423__6783(add_136_19_n_12 ,in9[12] ,in10[12]);
  or add_136_19_g424__3680(add_136_19_n_11 ,in9[8] ,in10[8]);
  and add_136_19_g425__1617(add_136_19_n_10 ,in9[12] ,in10[12]);
  or add_136_19_g426__2802(add_136_19_n_9 ,in9[14] ,in10[14]);
  and add_136_19_g427__1705(add_136_19_n_8 ,in9[11] ,in10[11]);
  or add_136_19_g428__5122(add_136_19_n_7 ,in9[3] ,in10[3]);
  and add_136_19_g429__8246(add_136_19_n_6 ,in9[6] ,in10[6]);
  and add_136_19_g430__7098(add_136_19_n_5 ,in9[2] ,in10[2]);
  and add_136_19_g431__6131(add_136_19_n_4 ,in9[1] ,in10[1]);
  and add_136_19_g432__1881(add_136_19_n_3 ,in9[5] ,in10[5]);
  or add_136_19_g433__5115(add_136_19_n_2 ,in9[10] ,in10[10]);
  not add_136_19_g434(add_136_19_n_1 ,in9[0]);
  not add_136_19_g435(add_136_19_n_0 ,in10[0]);
  or add_138_20_g341__7482(n_102 ,add_138_20_n_29 ,add_138_20_n_92);
  xnor add_138_20_g342__4733(n_101 ,add_138_20_n_91 ,add_138_20_n_39);
  nor add_138_20_g343__6161(add_138_20_n_92 ,add_138_20_n_15 ,add_138_20_n_91);
  or add_138_20_g344__9315(add_138_20_n_91 ,add_138_20_n_24 ,add_138_20_n_89);
  xnor add_138_20_g345__9945(n_100 ,add_138_20_n_88 ,add_138_20_n_38);
  and add_138_20_g346__2883(add_138_20_n_89 ,add_138_20_n_9 ,add_138_20_n_88);
  or add_138_20_g347__2346(add_138_20_n_88 ,add_138_20_n_20 ,add_138_20_n_86);
  xnor add_138_20_g348__1666(n_99 ,add_138_20_n_85 ,add_138_20_n_37);
  and add_138_20_g349__7410(add_138_20_n_86 ,add_138_20_n_16 ,add_138_20_n_85);
  or add_138_20_g350__6417(add_138_20_n_85 ,add_138_20_n_10 ,add_138_20_n_83);
  xnor add_138_20_g351__5477(n_98 ,add_138_20_n_82 ,add_138_20_n_36);
  and add_138_20_g352__2398(add_138_20_n_83 ,add_138_20_n_12 ,add_138_20_n_82);
  or add_138_20_g353__5107(add_138_20_n_82 ,add_138_20_n_8 ,add_138_20_n_80);
  xnor add_138_20_g354__6260(n_97 ,add_138_20_n_79 ,add_138_20_n_35);
  and add_138_20_g355__4319(add_138_20_n_80 ,add_138_20_n_22 ,add_138_20_n_79);
  or add_138_20_g356__8428(add_138_20_n_79 ,add_138_20_n_32 ,add_138_20_n_77);
  xnor add_138_20_g357__5526(n_96 ,add_138_20_n_76 ,add_138_20_n_42);
  and add_138_20_g358__6783(add_138_20_n_77 ,add_138_20_n_2 ,add_138_20_n_76);
  or add_138_20_g359__3680(add_138_20_n_76 ,add_138_20_n_21 ,add_138_20_n_74);
  xnor add_138_20_g360__1617(n_95 ,add_138_20_n_73 ,add_138_20_n_48);
  and add_138_20_g361__2802(add_138_20_n_74 ,add_138_20_n_19 ,add_138_20_n_73);
  or add_138_20_g362__1705(add_138_20_n_73 ,add_138_20_n_28 ,add_138_20_n_71);
  xnor add_138_20_g363__5122(n_94 ,add_138_20_n_70 ,add_138_20_n_47);
  and add_138_20_g364__8246(add_138_20_n_71 ,add_138_20_n_11 ,add_138_20_n_70);
  or add_138_20_g365__7098(add_138_20_n_70 ,add_138_20_n_17 ,add_138_20_n_68);
  xnor add_138_20_g366__6131(n_93 ,add_138_20_n_67 ,add_138_20_n_46);
  and add_138_20_g367__1881(add_138_20_n_68 ,add_138_20_n_25 ,add_138_20_n_67);
  or add_138_20_g368__5115(add_138_20_n_67 ,add_138_20_n_6 ,add_138_20_n_65);
  xnor add_138_20_g369__7482(n_92 ,add_138_20_n_64 ,add_138_20_n_45);
  and add_138_20_g370__4733(add_138_20_n_65 ,add_138_20_n_18 ,add_138_20_n_64);
  or add_138_20_g371__6161(add_138_20_n_64 ,add_138_20_n_3 ,add_138_20_n_62);
  xnor add_138_20_g372__9315(n_91 ,add_138_20_n_61 ,add_138_20_n_44);
  and add_138_20_g373__9945(add_138_20_n_62 ,add_138_20_n_30 ,add_138_20_n_61);
  or add_138_20_g374__2883(add_138_20_n_61 ,add_138_20_n_31 ,add_138_20_n_59);
  xnor add_138_20_g375__2346(n_90 ,add_138_20_n_58 ,add_138_20_n_43);
  and add_138_20_g376__1666(add_138_20_n_59 ,add_138_20_n_26 ,add_138_20_n_58);
  or add_138_20_g377__7410(add_138_20_n_58 ,add_138_20_n_27 ,add_138_20_n_56);
  xnor add_138_20_g378__6417(n_89 ,add_138_20_n_55 ,add_138_20_n_34);
  and add_138_20_g379__5477(add_138_20_n_56 ,add_138_20_n_7 ,add_138_20_n_55);
  or add_138_20_g380__2398(add_138_20_n_55 ,add_138_20_n_5 ,add_138_20_n_53);
  xnor add_138_20_g381__5107(n_88 ,add_138_20_n_51 ,add_138_20_n_41);
  and add_138_20_g382__6260(add_138_20_n_53 ,add_138_20_n_23 ,add_138_20_n_51);
  xor add_138_20_g383__4319(n_87 ,add_138_20_n_33 ,add_138_20_n_40);
  or add_138_20_g384__8428(add_138_20_n_51 ,add_138_20_n_4 ,add_138_20_n_49);
  and add_138_20_g385__5526(n_86 ,add_138_20_n_33 ,add_138_20_n_13);
  nor add_138_20_g386__6783(add_138_20_n_49 ,add_138_20_n_33 ,add_138_20_n_14);
  xnor add_138_20_g387__3680(add_138_20_n_48 ,in11[9] ,in12[9]);
  xnor add_138_20_g388__1617(add_138_20_n_47 ,in11[8] ,in12[8]);
  xnor add_138_20_g389__2802(add_138_20_n_46 ,in11[7] ,in12[7]);
  xnor add_138_20_g390__1705(add_138_20_n_45 ,in11[6] ,in12[6]);
  xnor add_138_20_g391__5122(add_138_20_n_44 ,in11[5] ,in12[5]);
  xnor add_138_20_g392__8246(add_138_20_n_43 ,in11[4] ,in12[4]);
  xnor add_138_20_g393__7098(add_138_20_n_42 ,in11[10] ,in12[10]);
  xnor add_138_20_g394__6131(add_138_20_n_41 ,in11[2] ,in12[2]);
  xnor add_138_20_g395__1881(add_138_20_n_40 ,in11[1] ,in12[1]);
  xnor add_138_20_g396__5115(add_138_20_n_39 ,in11[15] ,in12[15]);
  xnor add_138_20_g397__7482(add_138_20_n_38 ,in11[14] ,in12[14]);
  xnor add_138_20_g398__4733(add_138_20_n_37 ,in11[13] ,in12[13]);
  xnor add_138_20_g399__6161(add_138_20_n_36 ,in11[12] ,in12[12]);
  xnor add_138_20_g400__9315(add_138_20_n_35 ,in11[11] ,in12[11]);
  xnor add_138_20_g401__9945(add_138_20_n_34 ,in11[3] ,in12[3]);
  and add_138_20_g402__2883(add_138_20_n_32 ,in11[10] ,in12[10]);
  and add_138_20_g403__2346(add_138_20_n_31 ,in11[4] ,in12[4]);
  or add_138_20_g404__1666(add_138_20_n_30 ,in11[5] ,in12[5]);
  and add_138_20_g405__7410(add_138_20_n_29 ,in11[15] ,in12[15]);
  and add_138_20_g406__6417(add_138_20_n_28 ,in11[8] ,in12[8]);
  and add_138_20_g407__5477(add_138_20_n_27 ,in11[3] ,in12[3]);
  or add_138_20_g408__2398(add_138_20_n_26 ,in11[4] ,in12[4]);
  or add_138_20_g409__5107(add_138_20_n_25 ,in11[7] ,in12[7]);
  and add_138_20_g410__6260(add_138_20_n_24 ,in11[14] ,in12[14]);
  or add_138_20_g411__4319(add_138_20_n_23 ,in11[2] ,in12[2]);
  or add_138_20_g412__8428(add_138_20_n_22 ,in11[11] ,in12[11]);
  and add_138_20_g413__5526(add_138_20_n_21 ,in11[9] ,in12[9]);
  and add_138_20_g414__6783(add_138_20_n_20 ,in11[13] ,in12[13]);
  or add_138_20_g415__3680(add_138_20_n_19 ,in11[9] ,in12[9]);
  or add_138_20_g416__1617(add_138_20_n_18 ,in11[6] ,in12[6]);
  or add_138_20_g417__2802(add_138_20_n_33 ,add_138_20_n_1 ,add_138_20_n_0);
  and add_138_20_g418__1705(add_138_20_n_17 ,in11[7] ,in12[7]);
  or add_138_20_g419__5122(add_138_20_n_16 ,in11[13] ,in12[13]);
  nor add_138_20_g420__8246(add_138_20_n_15 ,in11[15] ,in12[15]);
  nor add_138_20_g421__7098(add_138_20_n_14 ,in11[1] ,in12[1]);
  or add_138_20_g422__6131(add_138_20_n_13 ,in11[0] ,in12[0]);
  or add_138_20_g423__1881(add_138_20_n_12 ,in11[12] ,in12[12]);
  or add_138_20_g424__5115(add_138_20_n_11 ,in11[8] ,in12[8]);
  and add_138_20_g425__7482(add_138_20_n_10 ,in11[12] ,in12[12]);
  or add_138_20_g426__4733(add_138_20_n_9 ,in11[14] ,in12[14]);
  and add_138_20_g427__6161(add_138_20_n_8 ,in11[11] ,in12[11]);
  or add_138_20_g428__9315(add_138_20_n_7 ,in11[3] ,in12[3]);
  and add_138_20_g429__9945(add_138_20_n_6 ,in11[6] ,in12[6]);
  and add_138_20_g430__2883(add_138_20_n_5 ,in11[2] ,in12[2]);
  and add_138_20_g431__2346(add_138_20_n_4 ,in11[1] ,in12[1]);
  and add_138_20_g432__1666(add_138_20_n_3 ,in11[5] ,in12[5]);
  or add_138_20_g433__7410(add_138_20_n_2 ,in11[10] ,in12[10]);
  not add_138_20_g434(add_138_20_n_1 ,in11[0]);
  not add_138_20_g435(add_138_20_n_0 ,in12[0]);
  or add_140_21_g341__6417(n_119 ,add_140_21_n_29 ,add_140_21_n_92);
  xnor add_140_21_g342__5477(n_118 ,add_140_21_n_91 ,add_140_21_n_39);
  nor add_140_21_g343__2398(add_140_21_n_92 ,add_140_21_n_15 ,add_140_21_n_91);
  or add_140_21_g344__5107(add_140_21_n_91 ,add_140_21_n_24 ,add_140_21_n_89);
  xnor add_140_21_g345__6260(n_117 ,add_140_21_n_88 ,add_140_21_n_38);
  and add_140_21_g346__4319(add_140_21_n_89 ,add_140_21_n_9 ,add_140_21_n_88);
  or add_140_21_g347__8428(add_140_21_n_88 ,add_140_21_n_20 ,add_140_21_n_86);
  xnor add_140_21_g348__5526(n_116 ,add_140_21_n_85 ,add_140_21_n_37);
  and add_140_21_g349__6783(add_140_21_n_86 ,add_140_21_n_16 ,add_140_21_n_85);
  or add_140_21_g350__3680(add_140_21_n_85 ,add_140_21_n_10 ,add_140_21_n_83);
  xnor add_140_21_g351__1617(n_115 ,add_140_21_n_82 ,add_140_21_n_36);
  and add_140_21_g352__2802(add_140_21_n_83 ,add_140_21_n_12 ,add_140_21_n_82);
  or add_140_21_g353__1705(add_140_21_n_82 ,add_140_21_n_8 ,add_140_21_n_80);
  xnor add_140_21_g354__5122(n_114 ,add_140_21_n_79 ,add_140_21_n_35);
  and add_140_21_g355__8246(add_140_21_n_80 ,add_140_21_n_22 ,add_140_21_n_79);
  or add_140_21_g356__7098(add_140_21_n_79 ,add_140_21_n_32 ,add_140_21_n_77);
  xnor add_140_21_g357__6131(n_113 ,add_140_21_n_76 ,add_140_21_n_42);
  and add_140_21_g358__1881(add_140_21_n_77 ,add_140_21_n_2 ,add_140_21_n_76);
  or add_140_21_g359__5115(add_140_21_n_76 ,add_140_21_n_21 ,add_140_21_n_74);
  xnor add_140_21_g360__7482(n_112 ,add_140_21_n_73 ,add_140_21_n_48);
  and add_140_21_g361__4733(add_140_21_n_74 ,add_140_21_n_19 ,add_140_21_n_73);
  or add_140_21_g362__6161(add_140_21_n_73 ,add_140_21_n_28 ,add_140_21_n_71);
  xnor add_140_21_g363__9315(n_111 ,add_140_21_n_70 ,add_140_21_n_47);
  and add_140_21_g364__9945(add_140_21_n_71 ,add_140_21_n_11 ,add_140_21_n_70);
  or add_140_21_g365__2883(add_140_21_n_70 ,add_140_21_n_17 ,add_140_21_n_68);
  xnor add_140_21_g366__2346(n_110 ,add_140_21_n_67 ,add_140_21_n_46);
  and add_140_21_g367__1666(add_140_21_n_68 ,add_140_21_n_25 ,add_140_21_n_67);
  or add_140_21_g368__7410(add_140_21_n_67 ,add_140_21_n_6 ,add_140_21_n_65);
  xnor add_140_21_g369__6417(n_109 ,add_140_21_n_64 ,add_140_21_n_45);
  and add_140_21_g370__5477(add_140_21_n_65 ,add_140_21_n_18 ,add_140_21_n_64);
  or add_140_21_g371__2398(add_140_21_n_64 ,add_140_21_n_3 ,add_140_21_n_62);
  xnor add_140_21_g372__5107(n_108 ,add_140_21_n_61 ,add_140_21_n_44);
  and add_140_21_g373__6260(add_140_21_n_62 ,add_140_21_n_30 ,add_140_21_n_61);
  or add_140_21_g374__4319(add_140_21_n_61 ,add_140_21_n_31 ,add_140_21_n_59);
  xnor add_140_21_g375__8428(n_107 ,add_140_21_n_58 ,add_140_21_n_43);
  and add_140_21_g376__5526(add_140_21_n_59 ,add_140_21_n_26 ,add_140_21_n_58);
  or add_140_21_g377__6783(add_140_21_n_58 ,add_140_21_n_27 ,add_140_21_n_56);
  xnor add_140_21_g378__3680(n_106 ,add_140_21_n_55 ,add_140_21_n_34);
  and add_140_21_g379__1617(add_140_21_n_56 ,add_140_21_n_7 ,add_140_21_n_55);
  or add_140_21_g380__2802(add_140_21_n_55 ,add_140_21_n_5 ,add_140_21_n_53);
  xnor add_140_21_g381__1705(n_105 ,add_140_21_n_51 ,add_140_21_n_41);
  and add_140_21_g382__5122(add_140_21_n_53 ,add_140_21_n_23 ,add_140_21_n_51);
  xor add_140_21_g383__8246(n_104 ,add_140_21_n_33 ,add_140_21_n_40);
  or add_140_21_g384__7098(add_140_21_n_51 ,add_140_21_n_4 ,add_140_21_n_49);
  and add_140_21_g385__6131(n_103 ,add_140_21_n_33 ,add_140_21_n_13);
  nor add_140_21_g386__1881(add_140_21_n_49 ,add_140_21_n_33 ,add_140_21_n_14);
  xnor add_140_21_g387__5115(add_140_21_n_48 ,in13[9] ,in14[9]);
  xnor add_140_21_g388__7482(add_140_21_n_47 ,in13[8] ,in14[8]);
  xnor add_140_21_g389__4733(add_140_21_n_46 ,in13[7] ,in14[7]);
  xnor add_140_21_g390__6161(add_140_21_n_45 ,in13[6] ,in14[6]);
  xnor add_140_21_g391__9315(add_140_21_n_44 ,in13[5] ,in14[5]);
  xnor add_140_21_g392__9945(add_140_21_n_43 ,in13[4] ,in14[4]);
  xnor add_140_21_g393__2883(add_140_21_n_42 ,in13[10] ,in14[10]);
  xnor add_140_21_g394__2346(add_140_21_n_41 ,in13[2] ,in14[2]);
  xnor add_140_21_g395__1666(add_140_21_n_40 ,in13[1] ,in14[1]);
  xnor add_140_21_g396__7410(add_140_21_n_39 ,in13[15] ,in14[15]);
  xnor add_140_21_g397__6417(add_140_21_n_38 ,in13[14] ,in14[14]);
  xnor add_140_21_g398__5477(add_140_21_n_37 ,in13[13] ,in14[13]);
  xnor add_140_21_g399__2398(add_140_21_n_36 ,in13[12] ,in14[12]);
  xnor add_140_21_g400__5107(add_140_21_n_35 ,in13[11] ,in14[11]);
  xnor add_140_21_g401__6260(add_140_21_n_34 ,in13[3] ,in14[3]);
  and add_140_21_g402__4319(add_140_21_n_32 ,in13[10] ,in14[10]);
  and add_140_21_g403__8428(add_140_21_n_31 ,in13[4] ,in14[4]);
  or add_140_21_g404__5526(add_140_21_n_30 ,in13[5] ,in14[5]);
  and add_140_21_g405__6783(add_140_21_n_29 ,in13[15] ,in14[15]);
  and add_140_21_g406__3680(add_140_21_n_28 ,in13[8] ,in14[8]);
  and add_140_21_g407__1617(add_140_21_n_27 ,in13[3] ,in14[3]);
  or add_140_21_g408__2802(add_140_21_n_26 ,in13[4] ,in14[4]);
  or add_140_21_g409__1705(add_140_21_n_25 ,in13[7] ,in14[7]);
  and add_140_21_g410__5122(add_140_21_n_24 ,in13[14] ,in14[14]);
  or add_140_21_g411__8246(add_140_21_n_23 ,in13[2] ,in14[2]);
  or add_140_21_g412__7098(add_140_21_n_22 ,in13[11] ,in14[11]);
  and add_140_21_g413__6131(add_140_21_n_21 ,in13[9] ,in14[9]);
  and add_140_21_g414__1881(add_140_21_n_20 ,in13[13] ,in14[13]);
  or add_140_21_g415__5115(add_140_21_n_19 ,in13[9] ,in14[9]);
  or add_140_21_g416__7482(add_140_21_n_18 ,in13[6] ,in14[6]);
  or add_140_21_g417__4733(add_140_21_n_33 ,add_140_21_n_1 ,add_140_21_n_0);
  and add_140_21_g418__6161(add_140_21_n_17 ,in13[7] ,in14[7]);
  or add_140_21_g419__9315(add_140_21_n_16 ,in13[13] ,in14[13]);
  nor add_140_21_g420__9945(add_140_21_n_15 ,in13[15] ,in14[15]);
  nor add_140_21_g421__2883(add_140_21_n_14 ,in13[1] ,in14[1]);
  or add_140_21_g422__2346(add_140_21_n_13 ,in13[0] ,in14[0]);
  or add_140_21_g423__1666(add_140_21_n_12 ,in13[12] ,in14[12]);
  or add_140_21_g424__7410(add_140_21_n_11 ,in13[8] ,in14[8]);
  and add_140_21_g425__6417(add_140_21_n_10 ,in13[12] ,in14[12]);
  or add_140_21_g426__5477(add_140_21_n_9 ,in13[14] ,in14[14]);
  and add_140_21_g427__2398(add_140_21_n_8 ,in13[11] ,in14[11]);
  or add_140_21_g428__5107(add_140_21_n_7 ,in13[3] ,in14[3]);
  and add_140_21_g429__6260(add_140_21_n_6 ,in13[6] ,in14[6]);
  and add_140_21_g430__4319(add_140_21_n_5 ,in13[2] ,in14[2]);
  and add_140_21_g431__8428(add_140_21_n_4 ,in13[1] ,in14[1]);
  and add_140_21_g432__5526(add_140_21_n_3 ,in13[5] ,in14[5]);
  or add_140_21_g433__6783(add_140_21_n_2 ,in13[10] ,in14[10]);
  not add_140_21_g434(add_140_21_n_1 ,in13[0]);
  not add_140_21_g435(add_140_21_n_0 ,in14[0]);
  or add_142_21_g341__3680(n_136 ,add_142_21_n_29 ,add_142_21_n_92);
  xnor add_142_21_g342__1617(n_135 ,add_142_21_n_91 ,add_142_21_n_39);
  nor add_142_21_g343__2802(add_142_21_n_92 ,add_142_21_n_15 ,add_142_21_n_91);
  or add_142_21_g344__1705(add_142_21_n_91 ,add_142_21_n_24 ,add_142_21_n_89);
  xnor add_142_21_g345__5122(n_134 ,add_142_21_n_88 ,add_142_21_n_38);
  and add_142_21_g346__8246(add_142_21_n_89 ,add_142_21_n_9 ,add_142_21_n_88);
  or add_142_21_g347__7098(add_142_21_n_88 ,add_142_21_n_20 ,add_142_21_n_86);
  xnor add_142_21_g348__6131(n_133 ,add_142_21_n_85 ,add_142_21_n_37);
  and add_142_21_g349__1881(add_142_21_n_86 ,add_142_21_n_16 ,add_142_21_n_85);
  or add_142_21_g350__5115(add_142_21_n_85 ,add_142_21_n_10 ,add_142_21_n_83);
  xnor add_142_21_g351__7482(n_132 ,add_142_21_n_82 ,add_142_21_n_36);
  and add_142_21_g352__4733(add_142_21_n_83 ,add_142_21_n_12 ,add_142_21_n_82);
  or add_142_21_g353__6161(add_142_21_n_82 ,add_142_21_n_8 ,add_142_21_n_80);
  xnor add_142_21_g354__9315(n_131 ,add_142_21_n_79 ,add_142_21_n_35);
  and add_142_21_g355__9945(add_142_21_n_80 ,add_142_21_n_22 ,add_142_21_n_79);
  or add_142_21_g356__2883(add_142_21_n_79 ,add_142_21_n_32 ,add_142_21_n_77);
  xnor add_142_21_g357__2346(n_130 ,add_142_21_n_76 ,add_142_21_n_42);
  and add_142_21_g358__1666(add_142_21_n_77 ,add_142_21_n_2 ,add_142_21_n_76);
  or add_142_21_g359__7410(add_142_21_n_76 ,add_142_21_n_21 ,add_142_21_n_74);
  xnor add_142_21_g360__6417(n_129 ,add_142_21_n_73 ,add_142_21_n_48);
  and add_142_21_g361__5477(add_142_21_n_74 ,add_142_21_n_19 ,add_142_21_n_73);
  or add_142_21_g362__2398(add_142_21_n_73 ,add_142_21_n_28 ,add_142_21_n_71);
  xnor add_142_21_g363__5107(n_128 ,add_142_21_n_70 ,add_142_21_n_47);
  and add_142_21_g364__6260(add_142_21_n_71 ,add_142_21_n_11 ,add_142_21_n_70);
  or add_142_21_g365__4319(add_142_21_n_70 ,add_142_21_n_17 ,add_142_21_n_68);
  xnor add_142_21_g366__8428(n_127 ,add_142_21_n_67 ,add_142_21_n_46);
  and add_142_21_g367__5526(add_142_21_n_68 ,add_142_21_n_25 ,add_142_21_n_67);
  or add_142_21_g368__6783(add_142_21_n_67 ,add_142_21_n_6 ,add_142_21_n_65);
  xnor add_142_21_g369__3680(n_126 ,add_142_21_n_64 ,add_142_21_n_45);
  and add_142_21_g370__1617(add_142_21_n_65 ,add_142_21_n_18 ,add_142_21_n_64);
  or add_142_21_g371__2802(add_142_21_n_64 ,add_142_21_n_3 ,add_142_21_n_62);
  xnor add_142_21_g372__1705(n_125 ,add_142_21_n_61 ,add_142_21_n_44);
  and add_142_21_g373__5122(add_142_21_n_62 ,add_142_21_n_30 ,add_142_21_n_61);
  or add_142_21_g374__8246(add_142_21_n_61 ,add_142_21_n_31 ,add_142_21_n_59);
  xnor add_142_21_g375__7098(n_124 ,add_142_21_n_58 ,add_142_21_n_43);
  and add_142_21_g376__6131(add_142_21_n_59 ,add_142_21_n_26 ,add_142_21_n_58);
  or add_142_21_g377__1881(add_142_21_n_58 ,add_142_21_n_27 ,add_142_21_n_56);
  xnor add_142_21_g378__5115(n_123 ,add_142_21_n_55 ,add_142_21_n_34);
  and add_142_21_g379__7482(add_142_21_n_56 ,add_142_21_n_7 ,add_142_21_n_55);
  or add_142_21_g380__4733(add_142_21_n_55 ,add_142_21_n_5 ,add_142_21_n_53);
  xnor add_142_21_g381__6161(n_122 ,add_142_21_n_51 ,add_142_21_n_41);
  and add_142_21_g382__9315(add_142_21_n_53 ,add_142_21_n_23 ,add_142_21_n_51);
  xor add_142_21_g383__9945(n_121 ,add_142_21_n_33 ,add_142_21_n_40);
  or add_142_21_g384__2883(add_142_21_n_51 ,add_142_21_n_4 ,add_142_21_n_49);
  and add_142_21_g385__2346(n_120 ,add_142_21_n_33 ,add_142_21_n_13);
  nor add_142_21_g386__1666(add_142_21_n_49 ,add_142_21_n_33 ,add_142_21_n_14);
  xnor add_142_21_g387__7410(add_142_21_n_48 ,in15[9] ,in16[9]);
  xnor add_142_21_g388__6417(add_142_21_n_47 ,in15[8] ,in16[8]);
  xnor add_142_21_g389__5477(add_142_21_n_46 ,in15[7] ,in16[7]);
  xnor add_142_21_g390__2398(add_142_21_n_45 ,in15[6] ,in16[6]);
  xnor add_142_21_g391__5107(add_142_21_n_44 ,in15[5] ,in16[5]);
  xnor add_142_21_g392__6260(add_142_21_n_43 ,in15[4] ,in16[4]);
  xnor add_142_21_g393__4319(add_142_21_n_42 ,in15[10] ,in16[10]);
  xnor add_142_21_g394__8428(add_142_21_n_41 ,in15[2] ,in16[2]);
  xnor add_142_21_g395__5526(add_142_21_n_40 ,in15[1] ,in16[1]);
  xnor add_142_21_g396__6783(add_142_21_n_39 ,in15[15] ,in16[15]);
  xnor add_142_21_g397__3680(add_142_21_n_38 ,in15[14] ,in16[14]);
  xnor add_142_21_g398__1617(add_142_21_n_37 ,in15[13] ,in16[13]);
  xnor add_142_21_g399__2802(add_142_21_n_36 ,in15[12] ,in16[12]);
  xnor add_142_21_g400__1705(add_142_21_n_35 ,in15[11] ,in16[11]);
  xnor add_142_21_g401__5122(add_142_21_n_34 ,in15[3] ,in16[3]);
  and add_142_21_g402__8246(add_142_21_n_32 ,in15[10] ,in16[10]);
  and add_142_21_g403__7098(add_142_21_n_31 ,in15[4] ,in16[4]);
  or add_142_21_g404__6131(add_142_21_n_30 ,in15[5] ,in16[5]);
  and add_142_21_g405__1881(add_142_21_n_29 ,in15[15] ,in16[15]);
  and add_142_21_g406__5115(add_142_21_n_28 ,in15[8] ,in16[8]);
  and add_142_21_g407__7482(add_142_21_n_27 ,in15[3] ,in16[3]);
  or add_142_21_g408__4733(add_142_21_n_26 ,in15[4] ,in16[4]);
  or add_142_21_g409__6161(add_142_21_n_25 ,in15[7] ,in16[7]);
  and add_142_21_g410__9315(add_142_21_n_24 ,in15[14] ,in16[14]);
  or add_142_21_g411__9945(add_142_21_n_23 ,in15[2] ,in16[2]);
  or add_142_21_g412__2883(add_142_21_n_22 ,in15[11] ,in16[11]);
  and add_142_21_g413__2346(add_142_21_n_21 ,in15[9] ,in16[9]);
  and add_142_21_g414__1666(add_142_21_n_20 ,in15[13] ,in16[13]);
  or add_142_21_g415__7410(add_142_21_n_19 ,in15[9] ,in16[9]);
  or add_142_21_g416__6417(add_142_21_n_18 ,in15[6] ,in16[6]);
  or add_142_21_g417__5477(add_142_21_n_33 ,add_142_21_n_1 ,add_142_21_n_0);
  and add_142_21_g418__2398(add_142_21_n_17 ,in15[7] ,in16[7]);
  or add_142_21_g419__5107(add_142_21_n_16 ,in15[13] ,in16[13]);
  nor add_142_21_g420__6260(add_142_21_n_15 ,in15[15] ,in16[15]);
  nor add_142_21_g421__4319(add_142_21_n_14 ,in15[1] ,in16[1]);
  or add_142_21_g422__8428(add_142_21_n_13 ,in15[0] ,in16[0]);
  or add_142_21_g423__5526(add_142_21_n_12 ,in15[12] ,in16[12]);
  or add_142_21_g424__6783(add_142_21_n_11 ,in15[8] ,in16[8]);
  and add_142_21_g425__3680(add_142_21_n_10 ,in15[12] ,in16[12]);
  or add_142_21_g426__1617(add_142_21_n_9 ,in15[14] ,in16[14]);
  and add_142_21_g427__2802(add_142_21_n_8 ,in15[11] ,in16[11]);
  or add_142_21_g428__1705(add_142_21_n_7 ,in15[3] ,in16[3]);
  and add_142_21_g429__5122(add_142_21_n_6 ,in15[6] ,in16[6]);
  and add_142_21_g430__8246(add_142_21_n_5 ,in15[2] ,in16[2]);
  and add_142_21_g431__7098(add_142_21_n_4 ,in15[1] ,in16[1]);
  and add_142_21_g432__6131(add_142_21_n_3 ,in15[5] ,in16[5]);
  or add_142_21_g433__1881(add_142_21_n_2 ,in15[10] ,in16[10]);
  not add_142_21_g434(add_142_21_n_1 ,in15[0]);
  not add_142_21_g435(add_142_21_n_0 ,in16[0]);
  or add_144_21_g341__5115(n_153 ,add_144_21_n_29 ,add_144_21_n_92);
  xnor add_144_21_g342__7482(n_152 ,add_144_21_n_91 ,add_144_21_n_39);
  nor add_144_21_g343__4733(add_144_21_n_92 ,add_144_21_n_15 ,add_144_21_n_91);
  or add_144_21_g344__6161(add_144_21_n_91 ,add_144_21_n_24 ,add_144_21_n_89);
  xnor add_144_21_g345__9315(n_151 ,add_144_21_n_88 ,add_144_21_n_38);
  and add_144_21_g346__9945(add_144_21_n_89 ,add_144_21_n_9 ,add_144_21_n_88);
  or add_144_21_g347__2883(add_144_21_n_88 ,add_144_21_n_20 ,add_144_21_n_86);
  xnor add_144_21_g348__2346(n_150 ,add_144_21_n_85 ,add_144_21_n_37);
  and add_144_21_g349__1666(add_144_21_n_86 ,add_144_21_n_16 ,add_144_21_n_85);
  or add_144_21_g350__7410(add_144_21_n_85 ,add_144_21_n_10 ,add_144_21_n_83);
  xnor add_144_21_g351__6417(n_149 ,add_144_21_n_82 ,add_144_21_n_36);
  and add_144_21_g352__5477(add_144_21_n_83 ,add_144_21_n_12 ,add_144_21_n_82);
  or add_144_21_g353__2398(add_144_21_n_82 ,add_144_21_n_8 ,add_144_21_n_80);
  xnor add_144_21_g354__5107(n_148 ,add_144_21_n_79 ,add_144_21_n_35);
  and add_144_21_g355__6260(add_144_21_n_80 ,add_144_21_n_22 ,add_144_21_n_79);
  or add_144_21_g356__4319(add_144_21_n_79 ,add_144_21_n_32 ,add_144_21_n_77);
  xnor add_144_21_g357__8428(n_147 ,add_144_21_n_76 ,add_144_21_n_42);
  and add_144_21_g358__5526(add_144_21_n_77 ,add_144_21_n_2 ,add_144_21_n_76);
  or add_144_21_g359__6783(add_144_21_n_76 ,add_144_21_n_21 ,add_144_21_n_74);
  xnor add_144_21_g360__3680(n_146 ,add_144_21_n_73 ,add_144_21_n_48);
  and add_144_21_g361__1617(add_144_21_n_74 ,add_144_21_n_19 ,add_144_21_n_73);
  or add_144_21_g362__2802(add_144_21_n_73 ,add_144_21_n_28 ,add_144_21_n_71);
  xnor add_144_21_g363__1705(n_145 ,add_144_21_n_70 ,add_144_21_n_47);
  and add_144_21_g364__5122(add_144_21_n_71 ,add_144_21_n_11 ,add_144_21_n_70);
  or add_144_21_g365__8246(add_144_21_n_70 ,add_144_21_n_17 ,add_144_21_n_68);
  xnor add_144_21_g366__7098(n_144 ,add_144_21_n_67 ,add_144_21_n_46);
  and add_144_21_g367__6131(add_144_21_n_68 ,add_144_21_n_25 ,add_144_21_n_67);
  or add_144_21_g368__1881(add_144_21_n_67 ,add_144_21_n_6 ,add_144_21_n_65);
  xnor add_144_21_g369__5115(n_143 ,add_144_21_n_64 ,add_144_21_n_45);
  and add_144_21_g370__7482(add_144_21_n_65 ,add_144_21_n_18 ,add_144_21_n_64);
  or add_144_21_g371__4733(add_144_21_n_64 ,add_144_21_n_3 ,add_144_21_n_62);
  xnor add_144_21_g372__6161(n_142 ,add_144_21_n_61 ,add_144_21_n_44);
  and add_144_21_g373__9315(add_144_21_n_62 ,add_144_21_n_30 ,add_144_21_n_61);
  or add_144_21_g374__9945(add_144_21_n_61 ,add_144_21_n_31 ,add_144_21_n_59);
  xnor add_144_21_g375__2883(n_141 ,add_144_21_n_58 ,add_144_21_n_43);
  and add_144_21_g376__2346(add_144_21_n_59 ,add_144_21_n_26 ,add_144_21_n_58);
  or add_144_21_g377__1666(add_144_21_n_58 ,add_144_21_n_27 ,add_144_21_n_56);
  xnor add_144_21_g378__7410(n_140 ,add_144_21_n_55 ,add_144_21_n_34);
  and add_144_21_g379__6417(add_144_21_n_56 ,add_144_21_n_7 ,add_144_21_n_55);
  or add_144_21_g380__5477(add_144_21_n_55 ,add_144_21_n_5 ,add_144_21_n_53);
  xnor add_144_21_g381__2398(n_139 ,add_144_21_n_51 ,add_144_21_n_41);
  and add_144_21_g382__5107(add_144_21_n_53 ,add_144_21_n_23 ,add_144_21_n_51);
  xor add_144_21_g383__6260(n_138 ,add_144_21_n_33 ,add_144_21_n_40);
  or add_144_21_g384__4319(add_144_21_n_51 ,add_144_21_n_4 ,add_144_21_n_49);
  and add_144_21_g385__8428(n_137 ,add_144_21_n_33 ,add_144_21_n_13);
  nor add_144_21_g386__5526(add_144_21_n_49 ,add_144_21_n_33 ,add_144_21_n_14);
  xnor add_144_21_g387__6783(add_144_21_n_48 ,in17[9] ,in18[9]);
  xnor add_144_21_g388__3680(add_144_21_n_47 ,in17[8] ,in18[8]);
  xnor add_144_21_g389__1617(add_144_21_n_46 ,in17[7] ,in18[7]);
  xnor add_144_21_g390__2802(add_144_21_n_45 ,in17[6] ,in18[6]);
  xnor add_144_21_g391__1705(add_144_21_n_44 ,in17[5] ,in18[5]);
  xnor add_144_21_g392__5122(add_144_21_n_43 ,in17[4] ,in18[4]);
  xnor add_144_21_g393__8246(add_144_21_n_42 ,in17[10] ,in18[10]);
  xnor add_144_21_g394__7098(add_144_21_n_41 ,in17[2] ,in18[2]);
  xnor add_144_21_g395__6131(add_144_21_n_40 ,in17[1] ,in18[1]);
  xnor add_144_21_g396__1881(add_144_21_n_39 ,in17[15] ,in18[15]);
  xnor add_144_21_g397__5115(add_144_21_n_38 ,in17[14] ,in18[14]);
  xnor add_144_21_g398__7482(add_144_21_n_37 ,in17[13] ,in18[13]);
  xnor add_144_21_g399__4733(add_144_21_n_36 ,in17[12] ,in18[12]);
  xnor add_144_21_g400__6161(add_144_21_n_35 ,in17[11] ,in18[11]);
  xnor add_144_21_g401__9315(add_144_21_n_34 ,in17[3] ,in18[3]);
  and add_144_21_g402__9945(add_144_21_n_32 ,in17[10] ,in18[10]);
  and add_144_21_g403__2883(add_144_21_n_31 ,in17[4] ,in18[4]);
  or add_144_21_g404__2346(add_144_21_n_30 ,in17[5] ,in18[5]);
  and add_144_21_g405__1666(add_144_21_n_29 ,in17[15] ,in18[15]);
  and add_144_21_g406__7410(add_144_21_n_28 ,in17[8] ,in18[8]);
  and add_144_21_g407__6417(add_144_21_n_27 ,in17[3] ,in18[3]);
  or add_144_21_g408__5477(add_144_21_n_26 ,in17[4] ,in18[4]);
  or add_144_21_g409__2398(add_144_21_n_25 ,in17[7] ,in18[7]);
  and add_144_21_g410__5107(add_144_21_n_24 ,in17[14] ,in18[14]);
  or add_144_21_g411__6260(add_144_21_n_23 ,in17[2] ,in18[2]);
  or add_144_21_g412__4319(add_144_21_n_22 ,in17[11] ,in18[11]);
  and add_144_21_g413__8428(add_144_21_n_21 ,in17[9] ,in18[9]);
  and add_144_21_g414__5526(add_144_21_n_20 ,in17[13] ,in18[13]);
  or add_144_21_g415__6783(add_144_21_n_19 ,in17[9] ,in18[9]);
  or add_144_21_g416__3680(add_144_21_n_18 ,in17[6] ,in18[6]);
  or add_144_21_g417__1617(add_144_21_n_33 ,add_144_21_n_1 ,add_144_21_n_0);
  and add_144_21_g418__2802(add_144_21_n_17 ,in17[7] ,in18[7]);
  or add_144_21_g419__1705(add_144_21_n_16 ,in17[13] ,in18[13]);
  nor add_144_21_g420__5122(add_144_21_n_15 ,in17[15] ,in18[15]);
  nor add_144_21_g421__8246(add_144_21_n_14 ,in17[1] ,in18[1]);
  or add_144_21_g422__7098(add_144_21_n_13 ,in17[0] ,in18[0]);
  or add_144_21_g423__6131(add_144_21_n_12 ,in17[12] ,in18[12]);
  or add_144_21_g424__1881(add_144_21_n_11 ,in17[8] ,in18[8]);
  and add_144_21_g425__5115(add_144_21_n_10 ,in17[12] ,in18[12]);
  or add_144_21_g426__7482(add_144_21_n_9 ,in17[14] ,in18[14]);
  and add_144_21_g427__4733(add_144_21_n_8 ,in17[11] ,in18[11]);
  or add_144_21_g428__6161(add_144_21_n_7 ,in17[3] ,in18[3]);
  and add_144_21_g429__9315(add_144_21_n_6 ,in17[6] ,in18[6]);
  and add_144_21_g430__9945(add_144_21_n_5 ,in17[2] ,in18[2]);
  and add_144_21_g431__2883(add_144_21_n_4 ,in17[1] ,in18[1]);
  and add_144_21_g432__2346(add_144_21_n_3 ,in17[5] ,in18[5]);
  or add_144_21_g433__1666(add_144_21_n_2 ,in17[10] ,in18[10]);
  not add_144_21_g434(add_144_21_n_1 ,in17[0]);
  not add_144_21_g435(add_144_21_n_0 ,in18[0]);
  or add_146_21_g341__7410(n_170 ,add_146_21_n_29 ,add_146_21_n_92);
  xnor add_146_21_g342__6417(n_169 ,add_146_21_n_91 ,add_146_21_n_39);
  nor add_146_21_g343__5477(add_146_21_n_92 ,add_146_21_n_15 ,add_146_21_n_91);
  or add_146_21_g344__2398(add_146_21_n_91 ,add_146_21_n_24 ,add_146_21_n_89);
  xnor add_146_21_g345__5107(n_168 ,add_146_21_n_88 ,add_146_21_n_38);
  and add_146_21_g346__6260(add_146_21_n_89 ,add_146_21_n_9 ,add_146_21_n_88);
  or add_146_21_g347__4319(add_146_21_n_88 ,add_146_21_n_20 ,add_146_21_n_86);
  xnor add_146_21_g348__8428(n_167 ,add_146_21_n_85 ,add_146_21_n_37);
  and add_146_21_g349__5526(add_146_21_n_86 ,add_146_21_n_16 ,add_146_21_n_85);
  or add_146_21_g350__6783(add_146_21_n_85 ,add_146_21_n_10 ,add_146_21_n_83);
  xnor add_146_21_g351__3680(n_166 ,add_146_21_n_82 ,add_146_21_n_36);
  and add_146_21_g352__1617(add_146_21_n_83 ,add_146_21_n_12 ,add_146_21_n_82);
  or add_146_21_g353__2802(add_146_21_n_82 ,add_146_21_n_8 ,add_146_21_n_80);
  xnor add_146_21_g354__1705(n_165 ,add_146_21_n_79 ,add_146_21_n_35);
  and add_146_21_g355__5122(add_146_21_n_80 ,add_146_21_n_22 ,add_146_21_n_79);
  or add_146_21_g356__8246(add_146_21_n_79 ,add_146_21_n_32 ,add_146_21_n_77);
  xnor add_146_21_g357__7098(n_164 ,add_146_21_n_76 ,add_146_21_n_42);
  and add_146_21_g358__6131(add_146_21_n_77 ,add_146_21_n_2 ,add_146_21_n_76);
  or add_146_21_g359__1881(add_146_21_n_76 ,add_146_21_n_21 ,add_146_21_n_74);
  xnor add_146_21_g360__5115(n_163 ,add_146_21_n_73 ,add_146_21_n_48);
  and add_146_21_g361__7482(add_146_21_n_74 ,add_146_21_n_19 ,add_146_21_n_73);
  or add_146_21_g362__4733(add_146_21_n_73 ,add_146_21_n_28 ,add_146_21_n_71);
  xnor add_146_21_g363__6161(n_162 ,add_146_21_n_70 ,add_146_21_n_47);
  and add_146_21_g364__9315(add_146_21_n_71 ,add_146_21_n_11 ,add_146_21_n_70);
  or add_146_21_g365__9945(add_146_21_n_70 ,add_146_21_n_17 ,add_146_21_n_68);
  xnor add_146_21_g366__2883(n_161 ,add_146_21_n_67 ,add_146_21_n_46);
  and add_146_21_g367__2346(add_146_21_n_68 ,add_146_21_n_25 ,add_146_21_n_67);
  or add_146_21_g368__1666(add_146_21_n_67 ,add_146_21_n_6 ,add_146_21_n_65);
  xnor add_146_21_g369__7410(n_160 ,add_146_21_n_64 ,add_146_21_n_45);
  and add_146_21_g370__6417(add_146_21_n_65 ,add_146_21_n_18 ,add_146_21_n_64);
  or add_146_21_g371__5477(add_146_21_n_64 ,add_146_21_n_3 ,add_146_21_n_62);
  xnor add_146_21_g372__2398(n_159 ,add_146_21_n_61 ,add_146_21_n_44);
  and add_146_21_g373__5107(add_146_21_n_62 ,add_146_21_n_30 ,add_146_21_n_61);
  or add_146_21_g374__6260(add_146_21_n_61 ,add_146_21_n_31 ,add_146_21_n_59);
  xnor add_146_21_g375__4319(n_158 ,add_146_21_n_58 ,add_146_21_n_43);
  and add_146_21_g376__8428(add_146_21_n_59 ,add_146_21_n_26 ,add_146_21_n_58);
  or add_146_21_g377__5526(add_146_21_n_58 ,add_146_21_n_27 ,add_146_21_n_56);
  xnor add_146_21_g378__6783(n_157 ,add_146_21_n_55 ,add_146_21_n_34);
  and add_146_21_g379__3680(add_146_21_n_56 ,add_146_21_n_7 ,add_146_21_n_55);
  or add_146_21_g380__1617(add_146_21_n_55 ,add_146_21_n_5 ,add_146_21_n_53);
  xnor add_146_21_g381__2802(n_156 ,add_146_21_n_51 ,add_146_21_n_41);
  and add_146_21_g382__1705(add_146_21_n_53 ,add_146_21_n_23 ,add_146_21_n_51);
  xor add_146_21_g383__5122(n_155 ,add_146_21_n_33 ,add_146_21_n_40);
  or add_146_21_g384__8246(add_146_21_n_51 ,add_146_21_n_4 ,add_146_21_n_49);
  and add_146_21_g385__7098(n_154 ,add_146_21_n_33 ,add_146_21_n_13);
  nor add_146_21_g386__6131(add_146_21_n_49 ,add_146_21_n_33 ,add_146_21_n_14);
  xnor add_146_21_g387__1881(add_146_21_n_48 ,in19[9] ,in20[9]);
  xnor add_146_21_g388__5115(add_146_21_n_47 ,in19[8] ,in20[8]);
  xnor add_146_21_g389__7482(add_146_21_n_46 ,in19[7] ,in20[7]);
  xnor add_146_21_g390__4733(add_146_21_n_45 ,in19[6] ,in20[6]);
  xnor add_146_21_g391__6161(add_146_21_n_44 ,in19[5] ,in20[5]);
  xnor add_146_21_g392__9315(add_146_21_n_43 ,in19[4] ,in20[4]);
  xnor add_146_21_g393__9945(add_146_21_n_42 ,in19[10] ,in20[10]);
  xnor add_146_21_g394__2883(add_146_21_n_41 ,in19[2] ,in20[2]);
  xnor add_146_21_g395__2346(add_146_21_n_40 ,in19[1] ,in20[1]);
  xnor add_146_21_g396__1666(add_146_21_n_39 ,in19[15] ,in20[15]);
  xnor add_146_21_g397__7410(add_146_21_n_38 ,in19[14] ,in20[14]);
  xnor add_146_21_g398__6417(add_146_21_n_37 ,in19[13] ,in20[13]);
  xnor add_146_21_g399__5477(add_146_21_n_36 ,in19[12] ,in20[12]);
  xnor add_146_21_g400__2398(add_146_21_n_35 ,in19[11] ,in20[11]);
  xnor add_146_21_g401__5107(add_146_21_n_34 ,in19[3] ,in20[3]);
  and add_146_21_g402__6260(add_146_21_n_32 ,in19[10] ,in20[10]);
  and add_146_21_g403__4319(add_146_21_n_31 ,in19[4] ,in20[4]);
  or add_146_21_g404__8428(add_146_21_n_30 ,in19[5] ,in20[5]);
  and add_146_21_g405__5526(add_146_21_n_29 ,in19[15] ,in20[15]);
  and add_146_21_g406__6783(add_146_21_n_28 ,in19[8] ,in20[8]);
  and add_146_21_g407__3680(add_146_21_n_27 ,in19[3] ,in20[3]);
  or add_146_21_g408__1617(add_146_21_n_26 ,in19[4] ,in20[4]);
  or add_146_21_g409__2802(add_146_21_n_25 ,in19[7] ,in20[7]);
  and add_146_21_g410__1705(add_146_21_n_24 ,in19[14] ,in20[14]);
  or add_146_21_g411__5122(add_146_21_n_23 ,in19[2] ,in20[2]);
  or add_146_21_g412__8246(add_146_21_n_22 ,in19[11] ,in20[11]);
  and add_146_21_g413__7098(add_146_21_n_21 ,in19[9] ,in20[9]);
  and add_146_21_g414__6131(add_146_21_n_20 ,in19[13] ,in20[13]);
  or add_146_21_g415__1881(add_146_21_n_19 ,in19[9] ,in20[9]);
  or add_146_21_g416__5115(add_146_21_n_18 ,in19[6] ,in20[6]);
  or add_146_21_g417__7482(add_146_21_n_33 ,add_146_21_n_1 ,add_146_21_n_0);
  and add_146_21_g418__4733(add_146_21_n_17 ,in19[7] ,in20[7]);
  or add_146_21_g419__6161(add_146_21_n_16 ,in19[13] ,in20[13]);
  nor add_146_21_g420__9315(add_146_21_n_15 ,in19[15] ,in20[15]);
  nor add_146_21_g421__9945(add_146_21_n_14 ,in19[1] ,in20[1]);
  or add_146_21_g422__2883(add_146_21_n_13 ,in19[0] ,in20[0]);
  or add_146_21_g423__2346(add_146_21_n_12 ,in19[12] ,in20[12]);
  or add_146_21_g424__1666(add_146_21_n_11 ,in19[8] ,in20[8]);
  and add_146_21_g425__7410(add_146_21_n_10 ,in19[12] ,in20[12]);
  or add_146_21_g426__6417(add_146_21_n_9 ,in19[14] ,in20[14]);
  and add_146_21_g427__5477(add_146_21_n_8 ,in19[11] ,in20[11]);
  or add_146_21_g428__2398(add_146_21_n_7 ,in19[3] ,in20[3]);
  and add_146_21_g429__5107(add_146_21_n_6 ,in19[6] ,in20[6]);
  and add_146_21_g430__6260(add_146_21_n_5 ,in19[2] ,in20[2]);
  and add_146_21_g431__4319(add_146_21_n_4 ,in19[1] ,in20[1]);
  and add_146_21_g432__8428(add_146_21_n_3 ,in19[5] ,in20[5]);
  or add_146_21_g433__5526(add_146_21_n_2 ,in19[10] ,in20[10]);
  not add_146_21_g434(add_146_21_n_1 ,in19[0]);
  not add_146_21_g435(add_146_21_n_0 ,in20[0]);
  or add_148_21_g341__6783(n_187 ,add_148_21_n_29 ,add_148_21_n_92);
  xnor add_148_21_g342__3680(n_186 ,add_148_21_n_91 ,add_148_21_n_39);
  nor add_148_21_g343__1617(add_148_21_n_92 ,add_148_21_n_15 ,add_148_21_n_91);
  or add_148_21_g344__2802(add_148_21_n_91 ,add_148_21_n_24 ,add_148_21_n_89);
  xnor add_148_21_g345__1705(n_185 ,add_148_21_n_88 ,add_148_21_n_38);
  and add_148_21_g346__5122(add_148_21_n_89 ,add_148_21_n_9 ,add_148_21_n_88);
  or add_148_21_g347__8246(add_148_21_n_88 ,add_148_21_n_20 ,add_148_21_n_86);
  xnor add_148_21_g348__7098(n_184 ,add_148_21_n_85 ,add_148_21_n_37);
  and add_148_21_g349__6131(add_148_21_n_86 ,add_148_21_n_16 ,add_148_21_n_85);
  or add_148_21_g350__1881(add_148_21_n_85 ,add_148_21_n_10 ,add_148_21_n_83);
  xnor add_148_21_g351__5115(n_183 ,add_148_21_n_82 ,add_148_21_n_36);
  and add_148_21_g352__7482(add_148_21_n_83 ,add_148_21_n_12 ,add_148_21_n_82);
  or add_148_21_g353__4733(add_148_21_n_82 ,add_148_21_n_8 ,add_148_21_n_80);
  xnor add_148_21_g354__6161(n_182 ,add_148_21_n_79 ,add_148_21_n_35);
  and add_148_21_g355__9315(add_148_21_n_80 ,add_148_21_n_22 ,add_148_21_n_79);
  or add_148_21_g356__9945(add_148_21_n_79 ,add_148_21_n_32 ,add_148_21_n_77);
  xnor add_148_21_g357__2883(n_181 ,add_148_21_n_76 ,add_148_21_n_42);
  and add_148_21_g358__2346(add_148_21_n_77 ,add_148_21_n_2 ,add_148_21_n_76);
  or add_148_21_g359__1666(add_148_21_n_76 ,add_148_21_n_21 ,add_148_21_n_74);
  xnor add_148_21_g360__7410(n_180 ,add_148_21_n_73 ,add_148_21_n_48);
  and add_148_21_g361__6417(add_148_21_n_74 ,add_148_21_n_19 ,add_148_21_n_73);
  or add_148_21_g362__5477(add_148_21_n_73 ,add_148_21_n_28 ,add_148_21_n_71);
  xnor add_148_21_g363__2398(n_179 ,add_148_21_n_70 ,add_148_21_n_47);
  and add_148_21_g364__5107(add_148_21_n_71 ,add_148_21_n_11 ,add_148_21_n_70);
  or add_148_21_g365__6260(add_148_21_n_70 ,add_148_21_n_17 ,add_148_21_n_68);
  xnor add_148_21_g366__4319(n_178 ,add_148_21_n_67 ,add_148_21_n_46);
  and add_148_21_g367__8428(add_148_21_n_68 ,add_148_21_n_25 ,add_148_21_n_67);
  or add_148_21_g368__5526(add_148_21_n_67 ,add_148_21_n_6 ,add_148_21_n_65);
  xnor add_148_21_g369__6783(n_177 ,add_148_21_n_64 ,add_148_21_n_45);
  and add_148_21_g370__3680(add_148_21_n_65 ,add_148_21_n_18 ,add_148_21_n_64);
  or add_148_21_g371__1617(add_148_21_n_64 ,add_148_21_n_3 ,add_148_21_n_62);
  xnor add_148_21_g372__2802(n_176 ,add_148_21_n_61 ,add_148_21_n_44);
  and add_148_21_g373__1705(add_148_21_n_62 ,add_148_21_n_30 ,add_148_21_n_61);
  or add_148_21_g374__5122(add_148_21_n_61 ,add_148_21_n_31 ,add_148_21_n_59);
  xnor add_148_21_g375__8246(n_175 ,add_148_21_n_58 ,add_148_21_n_43);
  and add_148_21_g376__7098(add_148_21_n_59 ,add_148_21_n_26 ,add_148_21_n_58);
  or add_148_21_g377__6131(add_148_21_n_58 ,add_148_21_n_27 ,add_148_21_n_56);
  xnor add_148_21_g378__1881(n_174 ,add_148_21_n_55 ,add_148_21_n_34);
  and add_148_21_g379__5115(add_148_21_n_56 ,add_148_21_n_7 ,add_148_21_n_55);
  or add_148_21_g380__7482(add_148_21_n_55 ,add_148_21_n_5 ,add_148_21_n_53);
  xnor add_148_21_g381__4733(n_173 ,add_148_21_n_51 ,add_148_21_n_41);
  and add_148_21_g382__6161(add_148_21_n_53 ,add_148_21_n_23 ,add_148_21_n_51);
  xor add_148_21_g383__9315(n_172 ,add_148_21_n_33 ,add_148_21_n_40);
  or add_148_21_g384__9945(add_148_21_n_51 ,add_148_21_n_4 ,add_148_21_n_49);
  and add_148_21_g385__2883(n_171 ,add_148_21_n_33 ,add_148_21_n_13);
  nor add_148_21_g386__2346(add_148_21_n_49 ,add_148_21_n_33 ,add_148_21_n_14);
  xnor add_148_21_g387__1666(add_148_21_n_48 ,in21[9] ,in22[9]);
  xnor add_148_21_g388__7410(add_148_21_n_47 ,in21[8] ,in22[8]);
  xnor add_148_21_g389__6417(add_148_21_n_46 ,in21[7] ,in22[7]);
  xnor add_148_21_g390__5477(add_148_21_n_45 ,in21[6] ,in22[6]);
  xnor add_148_21_g391__2398(add_148_21_n_44 ,in21[5] ,in22[5]);
  xnor add_148_21_g392__5107(add_148_21_n_43 ,in21[4] ,in22[4]);
  xnor add_148_21_g393__6260(add_148_21_n_42 ,in21[10] ,in22[10]);
  xnor add_148_21_g394__4319(add_148_21_n_41 ,in21[2] ,in22[2]);
  xnor add_148_21_g395__8428(add_148_21_n_40 ,in21[1] ,in22[1]);
  xnor add_148_21_g396__5526(add_148_21_n_39 ,in21[15] ,in22[15]);
  xnor add_148_21_g397__6783(add_148_21_n_38 ,in21[14] ,in22[14]);
  xnor add_148_21_g398__3680(add_148_21_n_37 ,in21[13] ,in22[13]);
  xnor add_148_21_g399__1617(add_148_21_n_36 ,in21[12] ,in22[12]);
  xnor add_148_21_g400__2802(add_148_21_n_35 ,in21[11] ,in22[11]);
  xnor add_148_21_g401__1705(add_148_21_n_34 ,in21[3] ,in22[3]);
  and add_148_21_g402__5122(add_148_21_n_32 ,in21[10] ,in22[10]);
  and add_148_21_g403__8246(add_148_21_n_31 ,in21[4] ,in22[4]);
  or add_148_21_g404__7098(add_148_21_n_30 ,in21[5] ,in22[5]);
  and add_148_21_g405__6131(add_148_21_n_29 ,in21[15] ,in22[15]);
  and add_148_21_g406__1881(add_148_21_n_28 ,in21[8] ,in22[8]);
  and add_148_21_g407__5115(add_148_21_n_27 ,in21[3] ,in22[3]);
  or add_148_21_g408__7482(add_148_21_n_26 ,in21[4] ,in22[4]);
  or add_148_21_g409__4733(add_148_21_n_25 ,in21[7] ,in22[7]);
  and add_148_21_g410__6161(add_148_21_n_24 ,in21[14] ,in22[14]);
  or add_148_21_g411(add_148_21_n_23 ,in21[2] ,in22[2]);
  or add_148_21_g412(add_148_21_n_22 ,in21[11] ,in22[11]);
  and add_148_21_g413(add_148_21_n_21 ,in21[9] ,in22[9]);
  and add_148_21_g414(add_148_21_n_20 ,in21[13] ,in22[13]);
  or add_148_21_g415(add_148_21_n_19 ,in21[9] ,in22[9]);
  or add_148_21_g416(add_148_21_n_18 ,in21[6] ,in22[6]);
  or add_148_21_g417(add_148_21_n_33 ,add_148_21_n_1 ,add_148_21_n_0);
  and add_148_21_g418(add_148_21_n_17 ,in21[7] ,in22[7]);
  or add_148_21_g419(add_148_21_n_16 ,in21[13] ,in22[13]);
  nor add_148_21_g420(add_148_21_n_15 ,in21[15] ,in22[15]);
  nor add_148_21_g421(add_148_21_n_14 ,in21[1] ,in22[1]);
  or add_148_21_g422(add_148_21_n_13 ,in21[0] ,in22[0]);
  or add_148_21_g423(add_148_21_n_12 ,in21[12] ,in22[12]);
  or add_148_21_g424(add_148_21_n_11 ,in21[8] ,in22[8]);
  and add_148_21_g425(add_148_21_n_10 ,in21[12] ,in22[12]);
  or add_148_21_g426(add_148_21_n_9 ,in21[14] ,in22[14]);
  and add_148_21_g427(add_148_21_n_8 ,in21[11] ,in22[11]);
  or add_148_21_g428(add_148_21_n_7 ,in21[3] ,in22[3]);
  and add_148_21_g429(add_148_21_n_6 ,in21[6] ,in22[6]);
  and add_148_21_g430(add_148_21_n_5 ,in21[2] ,in22[2]);
  and add_148_21_g431(add_148_21_n_4 ,in21[1] ,in22[1]);
  and add_148_21_g432(add_148_21_n_3 ,in21[5] ,in22[5]);
  or add_148_21_g433(add_148_21_n_2 ,in21[10] ,in22[10]);
  not add_148_21_g434(add_148_21_n_1 ,in21[0]);
  not add_148_21_g435(add_148_21_n_0 ,in22[0]);
  or add_150_21_g341(n_204 ,add_150_21_n_29 ,add_150_21_n_92);
  xnor add_150_21_g342(n_203 ,add_150_21_n_91 ,add_150_21_n_39);
  nor add_150_21_g343(add_150_21_n_92 ,add_150_21_n_15 ,add_150_21_n_91);
  or add_150_21_g344(add_150_21_n_91 ,add_150_21_n_24 ,add_150_21_n_89);
  xnor add_150_21_g345(n_202 ,add_150_21_n_88 ,add_150_21_n_38);
  and add_150_21_g346(add_150_21_n_89 ,add_150_21_n_9 ,add_150_21_n_88);
  or add_150_21_g347(add_150_21_n_88 ,add_150_21_n_20 ,add_150_21_n_86);
  xnor add_150_21_g348(n_201 ,add_150_21_n_85 ,add_150_21_n_37);
  and add_150_21_g349(add_150_21_n_86 ,add_150_21_n_16 ,add_150_21_n_85);
  or add_150_21_g350(add_150_21_n_85 ,add_150_21_n_10 ,add_150_21_n_83);
  xnor add_150_21_g351(n_200 ,add_150_21_n_82 ,add_150_21_n_36);
  and add_150_21_g352(add_150_21_n_83 ,add_150_21_n_12 ,add_150_21_n_82);
  or add_150_21_g353(add_150_21_n_82 ,add_150_21_n_8 ,add_150_21_n_80);
  xnor add_150_21_g354(n_199 ,add_150_21_n_79 ,add_150_21_n_35);
  and add_150_21_g355(add_150_21_n_80 ,add_150_21_n_22 ,add_150_21_n_79);
  or add_150_21_g356(add_150_21_n_79 ,add_150_21_n_32 ,add_150_21_n_77);
  xnor add_150_21_g357(n_198 ,add_150_21_n_76 ,add_150_21_n_42);
  and add_150_21_g358(add_150_21_n_77 ,add_150_21_n_2 ,add_150_21_n_76);
  or add_150_21_g359(add_150_21_n_76 ,add_150_21_n_21 ,add_150_21_n_74);
  xnor add_150_21_g360(n_197 ,add_150_21_n_73 ,add_150_21_n_48);
  and add_150_21_g361(add_150_21_n_74 ,add_150_21_n_19 ,add_150_21_n_73);
  or add_150_21_g362(add_150_21_n_73 ,add_150_21_n_28 ,add_150_21_n_71);
  xnor add_150_21_g363(n_196 ,add_150_21_n_70 ,add_150_21_n_47);
  and add_150_21_g364(add_150_21_n_71 ,add_150_21_n_11 ,add_150_21_n_70);
  or add_150_21_g365(add_150_21_n_70 ,add_150_21_n_17 ,add_150_21_n_68);
  xnor add_150_21_g366(n_195 ,add_150_21_n_67 ,add_150_21_n_46);
  and add_150_21_g367(add_150_21_n_68 ,add_150_21_n_25 ,add_150_21_n_67);
  or add_150_21_g368(add_150_21_n_67 ,add_150_21_n_6 ,add_150_21_n_65);
  xnor add_150_21_g369(n_194 ,add_150_21_n_64 ,add_150_21_n_45);
  and add_150_21_g370(add_150_21_n_65 ,add_150_21_n_18 ,add_150_21_n_64);
  or add_150_21_g371(add_150_21_n_64 ,add_150_21_n_3 ,add_150_21_n_62);
  xnor add_150_21_g372(n_193 ,add_150_21_n_61 ,add_150_21_n_44);
  and add_150_21_g373(add_150_21_n_62 ,add_150_21_n_30 ,add_150_21_n_61);
  or add_150_21_g374(add_150_21_n_61 ,add_150_21_n_31 ,add_150_21_n_59);
  xnor add_150_21_g375(n_192 ,add_150_21_n_58 ,add_150_21_n_43);
  and add_150_21_g376(add_150_21_n_59 ,add_150_21_n_26 ,add_150_21_n_58);
  or add_150_21_g377(add_150_21_n_58 ,add_150_21_n_27 ,add_150_21_n_56);
  xnor add_150_21_g378(n_191 ,add_150_21_n_55 ,add_150_21_n_34);
  and add_150_21_g379(add_150_21_n_56 ,add_150_21_n_7 ,add_150_21_n_55);
  or add_150_21_g380(add_150_21_n_55 ,add_150_21_n_5 ,add_150_21_n_53);
  xnor add_150_21_g381(n_190 ,add_150_21_n_51 ,add_150_21_n_41);
  and add_150_21_g382(add_150_21_n_53 ,add_150_21_n_23 ,add_150_21_n_51);
  xor add_150_21_g383(n_189 ,add_150_21_n_33 ,add_150_21_n_40);
  or add_150_21_g384(add_150_21_n_51 ,add_150_21_n_4 ,add_150_21_n_49);
  and add_150_21_g385(n_188 ,add_150_21_n_33 ,add_150_21_n_13);
  nor add_150_21_g386(add_150_21_n_49 ,add_150_21_n_33 ,add_150_21_n_14);
  xnor add_150_21_g387(add_150_21_n_48 ,in23[9] ,in24[9]);
  xnor add_150_21_g388(add_150_21_n_47 ,in23[8] ,in24[8]);
  xnor add_150_21_g389(add_150_21_n_46 ,in23[7] ,in24[7]);
  xnor add_150_21_g390(add_150_21_n_45 ,in23[6] ,in24[6]);
  xnor add_150_21_g391(add_150_21_n_44 ,in23[5] ,in24[5]);
  xnor add_150_21_g392(add_150_21_n_43 ,in23[4] ,in24[4]);
  xnor add_150_21_g393(add_150_21_n_42 ,in23[10] ,in24[10]);
  xnor add_150_21_g394(add_150_21_n_41 ,in23[2] ,in24[2]);
  xnor add_150_21_g395(add_150_21_n_40 ,in23[1] ,in24[1]);
  xnor add_150_21_g396(add_150_21_n_39 ,in23[15] ,in24[15]);
  xnor add_150_21_g397(add_150_21_n_38 ,in23[14] ,in24[14]);
  xnor add_150_21_g398(add_150_21_n_37 ,in23[13] ,in24[13]);
  xnor add_150_21_g399(add_150_21_n_36 ,in23[12] ,in24[12]);
  xnor add_150_21_g400(add_150_21_n_35 ,in23[11] ,in24[11]);
  xnor add_150_21_g401(add_150_21_n_34 ,in23[3] ,in24[3]);
  and add_150_21_g402(add_150_21_n_32 ,in23[10] ,in24[10]);
  and add_150_21_g403(add_150_21_n_31 ,in23[4] ,in24[4]);
  or add_150_21_g404(add_150_21_n_30 ,in23[5] ,in24[5]);
  and add_150_21_g405(add_150_21_n_29 ,in23[15] ,in24[15]);
  and add_150_21_g406(add_150_21_n_28 ,in23[8] ,in24[8]);
  and add_150_21_g407(add_150_21_n_27 ,in23[3] ,in24[3]);
  or add_150_21_g408(add_150_21_n_26 ,in23[4] ,in24[4]);
  or add_150_21_g409(add_150_21_n_25 ,in23[7] ,in24[7]);
  and add_150_21_g410(add_150_21_n_24 ,in23[14] ,in24[14]);
  or add_150_21_g411(add_150_21_n_23 ,in23[2] ,in24[2]);
  or add_150_21_g412(add_150_21_n_22 ,in23[11] ,in24[11]);
  and add_150_21_g413(add_150_21_n_21 ,in23[9] ,in24[9]);
  and add_150_21_g414(add_150_21_n_20 ,in23[13] ,in24[13]);
  or add_150_21_g415(add_150_21_n_19 ,in23[9] ,in24[9]);
  or add_150_21_g416(add_150_21_n_18 ,in23[6] ,in24[6]);
  or add_150_21_g417(add_150_21_n_33 ,add_150_21_n_1 ,add_150_21_n_0);
  and add_150_21_g418(add_150_21_n_17 ,in23[7] ,in24[7]);
  or add_150_21_g419(add_150_21_n_16 ,in23[13] ,in24[13]);
  nor add_150_21_g420(add_150_21_n_15 ,in23[15] ,in24[15]);
  nor add_150_21_g421(add_150_21_n_14 ,in23[1] ,in24[1]);
  or add_150_21_g422(add_150_21_n_13 ,in23[0] ,in24[0]);
  or add_150_21_g423(add_150_21_n_12 ,in23[12] ,in24[12]);
  or add_150_21_g424(add_150_21_n_11 ,in23[8] ,in24[8]);
  and add_150_21_g425(add_150_21_n_10 ,in23[12] ,in24[12]);
  or add_150_21_g426(add_150_21_n_9 ,in23[14] ,in24[14]);
  and add_150_21_g427(add_150_21_n_8 ,in23[11] ,in24[11]);
  or add_150_21_g428(add_150_21_n_7 ,in23[3] ,in24[3]);
  and add_150_21_g429(add_150_21_n_6 ,in23[6] ,in24[6]);
  and add_150_21_g430(add_150_21_n_5 ,in23[2] ,in24[2]);
  and add_150_21_g431(add_150_21_n_4 ,in23[1] ,in24[1]);
  and add_150_21_g432(add_150_21_n_3 ,in23[5] ,in24[5]);
  or add_150_21_g433(add_150_21_n_2 ,in23[10] ,in24[10]);
  not add_150_21_g434(add_150_21_n_1 ,in23[0]);
  not add_150_21_g435(add_150_21_n_0 ,in24[0]);
  or add_152_21_g341(n_221 ,add_152_21_n_29 ,add_152_21_n_92);
  xnor add_152_21_g342(n_220 ,add_152_21_n_91 ,add_152_21_n_39);
  nor add_152_21_g343(add_152_21_n_92 ,add_152_21_n_15 ,add_152_21_n_91);
  or add_152_21_g344(add_152_21_n_91 ,add_152_21_n_24 ,add_152_21_n_89);
  xnor add_152_21_g345(n_219 ,add_152_21_n_88 ,add_152_21_n_38);
  and add_152_21_g346(add_152_21_n_89 ,add_152_21_n_9 ,add_152_21_n_88);
  or add_152_21_g347(add_152_21_n_88 ,add_152_21_n_20 ,add_152_21_n_86);
  xnor add_152_21_g348(n_218 ,add_152_21_n_85 ,add_152_21_n_37);
  and add_152_21_g349(add_152_21_n_86 ,add_152_21_n_16 ,add_152_21_n_85);
  or add_152_21_g350(add_152_21_n_85 ,add_152_21_n_10 ,add_152_21_n_83);
  xnor add_152_21_g351(n_217 ,add_152_21_n_82 ,add_152_21_n_36);
  and add_152_21_g352(add_152_21_n_83 ,add_152_21_n_12 ,add_152_21_n_82);
  or add_152_21_g353(add_152_21_n_82 ,add_152_21_n_8 ,add_152_21_n_80);
  xnor add_152_21_g354(n_216 ,add_152_21_n_79 ,add_152_21_n_35);
  and add_152_21_g355(add_152_21_n_80 ,add_152_21_n_22 ,add_152_21_n_79);
  or add_152_21_g356(add_152_21_n_79 ,add_152_21_n_32 ,add_152_21_n_77);
  xnor add_152_21_g357(n_215 ,add_152_21_n_76 ,add_152_21_n_42);
  and add_152_21_g358(add_152_21_n_77 ,add_152_21_n_2 ,add_152_21_n_76);
  or add_152_21_g359(add_152_21_n_76 ,add_152_21_n_21 ,add_152_21_n_74);
  xnor add_152_21_g360(n_214 ,add_152_21_n_73 ,add_152_21_n_48);
  and add_152_21_g361(add_152_21_n_74 ,add_152_21_n_19 ,add_152_21_n_73);
  or add_152_21_g362(add_152_21_n_73 ,add_152_21_n_28 ,add_152_21_n_71);
  xnor add_152_21_g363(n_213 ,add_152_21_n_70 ,add_152_21_n_47);
  and add_152_21_g364(add_152_21_n_71 ,add_152_21_n_11 ,add_152_21_n_70);
  or add_152_21_g365(add_152_21_n_70 ,add_152_21_n_17 ,add_152_21_n_68);
  xnor add_152_21_g366(n_212 ,add_152_21_n_67 ,add_152_21_n_46);
  and add_152_21_g367(add_152_21_n_68 ,add_152_21_n_25 ,add_152_21_n_67);
  or add_152_21_g368(add_152_21_n_67 ,add_152_21_n_6 ,add_152_21_n_65);
  xnor add_152_21_g369(n_211 ,add_152_21_n_64 ,add_152_21_n_45);
  and add_152_21_g370(add_152_21_n_65 ,add_152_21_n_18 ,add_152_21_n_64);
  or add_152_21_g371(add_152_21_n_64 ,add_152_21_n_3 ,add_152_21_n_62);
  xnor add_152_21_g372(n_210 ,add_152_21_n_61 ,add_152_21_n_44);
  and add_152_21_g373(add_152_21_n_62 ,add_152_21_n_30 ,add_152_21_n_61);
  or add_152_21_g374(add_152_21_n_61 ,add_152_21_n_31 ,add_152_21_n_59);
  xnor add_152_21_g375(n_209 ,add_152_21_n_58 ,add_152_21_n_43);
  and add_152_21_g376(add_152_21_n_59 ,add_152_21_n_26 ,add_152_21_n_58);
  or add_152_21_g377(add_152_21_n_58 ,add_152_21_n_27 ,add_152_21_n_56);
  xnor add_152_21_g378(n_208 ,add_152_21_n_55 ,add_152_21_n_34);
  and add_152_21_g379(add_152_21_n_56 ,add_152_21_n_7 ,add_152_21_n_55);
  or add_152_21_g380(add_152_21_n_55 ,add_152_21_n_5 ,add_152_21_n_53);
  xnor add_152_21_g381(n_207 ,add_152_21_n_51 ,add_152_21_n_41);
  and add_152_21_g382(add_152_21_n_53 ,add_152_21_n_23 ,add_152_21_n_51);
  xor add_152_21_g383(n_206 ,add_152_21_n_33 ,add_152_21_n_40);
  or add_152_21_g384(add_152_21_n_51 ,add_152_21_n_4 ,add_152_21_n_49);
  and add_152_21_g385(n_205 ,add_152_21_n_33 ,add_152_21_n_13);
  nor add_152_21_g386(add_152_21_n_49 ,add_152_21_n_33 ,add_152_21_n_14);
  xnor add_152_21_g387(add_152_21_n_48 ,in25[9] ,in26[9]);
  xnor add_152_21_g388(add_152_21_n_47 ,in25[8] ,in26[8]);
  xnor add_152_21_g389(add_152_21_n_46 ,in25[7] ,in26[7]);
  xnor add_152_21_g390(add_152_21_n_45 ,in25[6] ,in26[6]);
  xnor add_152_21_g391(add_152_21_n_44 ,in25[5] ,in26[5]);
  xnor add_152_21_g392(add_152_21_n_43 ,in25[4] ,in26[4]);
  xnor add_152_21_g393(add_152_21_n_42 ,in25[10] ,in26[10]);
  xnor add_152_21_g394(add_152_21_n_41 ,in25[2] ,in26[2]);
  xnor add_152_21_g395(add_152_21_n_40 ,in25[1] ,in26[1]);
  xnor add_152_21_g396(add_152_21_n_39 ,in25[15] ,in26[15]);
  xnor add_152_21_g397(add_152_21_n_38 ,in25[14] ,in26[14]);
  xnor add_152_21_g398(add_152_21_n_37 ,in25[13] ,in26[13]);
  xnor add_152_21_g399(add_152_21_n_36 ,in25[12] ,in26[12]);
  xnor add_152_21_g400(add_152_21_n_35 ,in25[11] ,in26[11]);
  xnor add_152_21_g401(add_152_21_n_34 ,in25[3] ,in26[3]);
  and add_152_21_g402(add_152_21_n_32 ,in25[10] ,in26[10]);
  and add_152_21_g403(add_152_21_n_31 ,in25[4] ,in26[4]);
  or add_152_21_g404(add_152_21_n_30 ,in25[5] ,in26[5]);
  and add_152_21_g405(add_152_21_n_29 ,in25[15] ,in26[15]);
  and add_152_21_g406(add_152_21_n_28 ,in25[8] ,in26[8]);
  and add_152_21_g407(add_152_21_n_27 ,in25[3] ,in26[3]);
  or add_152_21_g408(add_152_21_n_26 ,in25[4] ,in26[4]);
  or add_152_21_g409(add_152_21_n_25 ,in25[7] ,in26[7]);
  and add_152_21_g410(add_152_21_n_24 ,in25[14] ,in26[14]);
  or add_152_21_g411(add_152_21_n_23 ,in25[2] ,in26[2]);
  or add_152_21_g412(add_152_21_n_22 ,in25[11] ,in26[11]);
  and add_152_21_g413(add_152_21_n_21 ,in25[9] ,in26[9]);
  and add_152_21_g414(add_152_21_n_20 ,in25[13] ,in26[13]);
  or add_152_21_g415(add_152_21_n_19 ,in25[9] ,in26[9]);
  or add_152_21_g416(add_152_21_n_18 ,in25[6] ,in26[6]);
  or add_152_21_g417(add_152_21_n_33 ,add_152_21_n_1 ,add_152_21_n_0);
  and add_152_21_g418(add_152_21_n_17 ,in25[7] ,in26[7]);
  or add_152_21_g419(add_152_21_n_16 ,in25[13] ,in26[13]);
  nor add_152_21_g420(add_152_21_n_15 ,in25[15] ,in26[15]);
  nor add_152_21_g421(add_152_21_n_14 ,in25[1] ,in26[1]);
  or add_152_21_g422(add_152_21_n_13 ,in25[0] ,in26[0]);
  or add_152_21_g423(add_152_21_n_12 ,in25[12] ,in26[12]);
  or add_152_21_g424(add_152_21_n_11 ,in25[8] ,in26[8]);
  and add_152_21_g425(add_152_21_n_10 ,in25[12] ,in26[12]);
  or add_152_21_g426(add_152_21_n_9 ,in25[14] ,in26[14]);
  and add_152_21_g427(add_152_21_n_8 ,in25[11] ,in26[11]);
  or add_152_21_g428(add_152_21_n_7 ,in25[3] ,in26[3]);
  and add_152_21_g429(add_152_21_n_6 ,in25[6] ,in26[6]);
  and add_152_21_g430(add_152_21_n_5 ,in25[2] ,in26[2]);
  and add_152_21_g431(add_152_21_n_4 ,in25[1] ,in26[1]);
  and add_152_21_g432(add_152_21_n_3 ,in25[5] ,in26[5]);
  or add_152_21_g433(add_152_21_n_2 ,in25[10] ,in26[10]);
  not add_152_21_g434(add_152_21_n_1 ,in25[0]);
  not add_152_21_g435(add_152_21_n_0 ,in26[0]);
  or add_154_21_g341(n_238 ,add_154_21_n_29 ,add_154_21_n_92);
  xnor add_154_21_g342(n_237 ,add_154_21_n_91 ,add_154_21_n_39);
  nor add_154_21_g343(add_154_21_n_92 ,add_154_21_n_15 ,add_154_21_n_91);
  or add_154_21_g344(add_154_21_n_91 ,add_154_21_n_24 ,add_154_21_n_89);
  xnor add_154_21_g345(n_236 ,add_154_21_n_88 ,add_154_21_n_38);
  and add_154_21_g346(add_154_21_n_89 ,add_154_21_n_9 ,add_154_21_n_88);
  or add_154_21_g347(add_154_21_n_88 ,add_154_21_n_20 ,add_154_21_n_86);
  xnor add_154_21_g348(n_235 ,add_154_21_n_85 ,add_154_21_n_37);
  and add_154_21_g349(add_154_21_n_86 ,add_154_21_n_16 ,add_154_21_n_85);
  or add_154_21_g350(add_154_21_n_85 ,add_154_21_n_10 ,add_154_21_n_83);
  xnor add_154_21_g351(n_234 ,add_154_21_n_82 ,add_154_21_n_36);
  and add_154_21_g352(add_154_21_n_83 ,add_154_21_n_12 ,add_154_21_n_82);
  or add_154_21_g353(add_154_21_n_82 ,add_154_21_n_8 ,add_154_21_n_80);
  xnor add_154_21_g354(n_233 ,add_154_21_n_79 ,add_154_21_n_35);
  and add_154_21_g355(add_154_21_n_80 ,add_154_21_n_22 ,add_154_21_n_79);
  or add_154_21_g356(add_154_21_n_79 ,add_154_21_n_32 ,add_154_21_n_77);
  xnor add_154_21_g357(n_232 ,add_154_21_n_76 ,add_154_21_n_42);
  and add_154_21_g358(add_154_21_n_77 ,add_154_21_n_2 ,add_154_21_n_76);
  or add_154_21_g359(add_154_21_n_76 ,add_154_21_n_21 ,add_154_21_n_74);
  xnor add_154_21_g360(n_231 ,add_154_21_n_73 ,add_154_21_n_48);
  and add_154_21_g361(add_154_21_n_74 ,add_154_21_n_19 ,add_154_21_n_73);
  or add_154_21_g362(add_154_21_n_73 ,add_154_21_n_28 ,add_154_21_n_71);
  xnor add_154_21_g363(n_230 ,add_154_21_n_70 ,add_154_21_n_47);
  and add_154_21_g364(add_154_21_n_71 ,add_154_21_n_11 ,add_154_21_n_70);
  or add_154_21_g365(add_154_21_n_70 ,add_154_21_n_17 ,add_154_21_n_68);
  xnor add_154_21_g366(n_229 ,add_154_21_n_67 ,add_154_21_n_46);
  and add_154_21_g367(add_154_21_n_68 ,add_154_21_n_25 ,add_154_21_n_67);
  or add_154_21_g368(add_154_21_n_67 ,add_154_21_n_6 ,add_154_21_n_65);
  xnor add_154_21_g369(n_228 ,add_154_21_n_64 ,add_154_21_n_45);
  and add_154_21_g370(add_154_21_n_65 ,add_154_21_n_18 ,add_154_21_n_64);
  or add_154_21_g371(add_154_21_n_64 ,add_154_21_n_3 ,add_154_21_n_62);
  xnor add_154_21_g372(n_227 ,add_154_21_n_61 ,add_154_21_n_44);
  and add_154_21_g373(add_154_21_n_62 ,add_154_21_n_30 ,add_154_21_n_61);
  or add_154_21_g374(add_154_21_n_61 ,add_154_21_n_31 ,add_154_21_n_59);
  xnor add_154_21_g375(n_226 ,add_154_21_n_58 ,add_154_21_n_43);
  and add_154_21_g376(add_154_21_n_59 ,add_154_21_n_26 ,add_154_21_n_58);
  or add_154_21_g377(add_154_21_n_58 ,add_154_21_n_27 ,add_154_21_n_56);
  xnor add_154_21_g378(n_225 ,add_154_21_n_55 ,add_154_21_n_34);
  and add_154_21_g379(add_154_21_n_56 ,add_154_21_n_7 ,add_154_21_n_55);
  or add_154_21_g380(add_154_21_n_55 ,add_154_21_n_5 ,add_154_21_n_53);
  xnor add_154_21_g381(n_224 ,add_154_21_n_51 ,add_154_21_n_41);
  and add_154_21_g382(add_154_21_n_53 ,add_154_21_n_23 ,add_154_21_n_51);
  xor add_154_21_g383(n_223 ,add_154_21_n_33 ,add_154_21_n_40);
  or add_154_21_g384(add_154_21_n_51 ,add_154_21_n_4 ,add_154_21_n_49);
  and add_154_21_g385(n_222 ,add_154_21_n_33 ,add_154_21_n_13);
  nor add_154_21_g386(add_154_21_n_49 ,add_154_21_n_33 ,add_154_21_n_14);
  xnor add_154_21_g387(add_154_21_n_48 ,in27[9] ,in28[9]);
  xnor add_154_21_g388(add_154_21_n_47 ,in27[8] ,in28[8]);
  xnor add_154_21_g389(add_154_21_n_46 ,in27[7] ,in28[7]);
  xnor add_154_21_g390(add_154_21_n_45 ,in27[6] ,in28[6]);
  xnor add_154_21_g391(add_154_21_n_44 ,in27[5] ,in28[5]);
  xnor add_154_21_g392(add_154_21_n_43 ,in27[4] ,in28[4]);
  xnor add_154_21_g393(add_154_21_n_42 ,in27[10] ,in28[10]);
  xnor add_154_21_g394(add_154_21_n_41 ,in27[2] ,in28[2]);
  xnor add_154_21_g395(add_154_21_n_40 ,in27[1] ,in28[1]);
  xnor add_154_21_g396(add_154_21_n_39 ,in27[15] ,in28[15]);
  xnor add_154_21_g397(add_154_21_n_38 ,in27[14] ,in28[14]);
  xnor add_154_21_g398(add_154_21_n_37 ,in27[13] ,in28[13]);
  xnor add_154_21_g399(add_154_21_n_36 ,in27[12] ,in28[12]);
  xnor add_154_21_g400(add_154_21_n_35 ,in27[11] ,in28[11]);
  xnor add_154_21_g401(add_154_21_n_34 ,in27[3] ,in28[3]);
  and add_154_21_g402(add_154_21_n_32 ,in27[10] ,in28[10]);
  and add_154_21_g403(add_154_21_n_31 ,in27[4] ,in28[4]);
  or add_154_21_g404(add_154_21_n_30 ,in27[5] ,in28[5]);
  and add_154_21_g405(add_154_21_n_29 ,in27[15] ,in28[15]);
  and add_154_21_g406(add_154_21_n_28 ,in27[8] ,in28[8]);
  and add_154_21_g407(add_154_21_n_27 ,in27[3] ,in28[3]);
  or add_154_21_g408(add_154_21_n_26 ,in27[4] ,in28[4]);
  or add_154_21_g409(add_154_21_n_25 ,in27[7] ,in28[7]);
  and add_154_21_g410(add_154_21_n_24 ,in27[14] ,in28[14]);
  or add_154_21_g411(add_154_21_n_23 ,in27[2] ,in28[2]);
  or add_154_21_g412(add_154_21_n_22 ,in27[11] ,in28[11]);
  and add_154_21_g413(add_154_21_n_21 ,in27[9] ,in28[9]);
  and add_154_21_g414(add_154_21_n_20 ,in27[13] ,in28[13]);
  or add_154_21_g415(add_154_21_n_19 ,in27[9] ,in28[9]);
  or add_154_21_g416(add_154_21_n_18 ,in27[6] ,in28[6]);
  or add_154_21_g417(add_154_21_n_33 ,add_154_21_n_1 ,add_154_21_n_0);
  and add_154_21_g418(add_154_21_n_17 ,in27[7] ,in28[7]);
  or add_154_21_g419(add_154_21_n_16 ,in27[13] ,in28[13]);
  nor add_154_21_g420(add_154_21_n_15 ,in27[15] ,in28[15]);
  nor add_154_21_g421(add_154_21_n_14 ,in27[1] ,in28[1]);
  or add_154_21_g422(add_154_21_n_13 ,in27[0] ,in28[0]);
  or add_154_21_g423(add_154_21_n_12 ,in27[12] ,in28[12]);
  or add_154_21_g424(add_154_21_n_11 ,in27[8] ,in28[8]);
  and add_154_21_g425(add_154_21_n_10 ,in27[12] ,in28[12]);
  or add_154_21_g426(add_154_21_n_9 ,in27[14] ,in28[14]);
  and add_154_21_g427(add_154_21_n_8 ,in27[11] ,in28[11]);
  or add_154_21_g428(add_154_21_n_7 ,in27[3] ,in28[3]);
  and add_154_21_g429(add_154_21_n_6 ,in27[6] ,in28[6]);
  and add_154_21_g430(add_154_21_n_5 ,in27[2] ,in28[2]);
  and add_154_21_g431(add_154_21_n_4 ,in27[1] ,in28[1]);
  and add_154_21_g432(add_154_21_n_3 ,in27[5] ,in28[5]);
  or add_154_21_g433(add_154_21_n_2 ,in27[10] ,in28[10]);
  not add_154_21_g434(add_154_21_n_1 ,in27[0]);
  not add_154_21_g435(add_154_21_n_0 ,in28[0]);
  or add_156_21_g341(n_255 ,add_156_21_n_29 ,add_156_21_n_92);
  xnor add_156_21_g342(n_254 ,add_156_21_n_91 ,add_156_21_n_39);
  nor add_156_21_g343(add_156_21_n_92 ,add_156_21_n_15 ,add_156_21_n_91);
  or add_156_21_g344(add_156_21_n_91 ,add_156_21_n_24 ,add_156_21_n_89);
  xnor add_156_21_g345(n_253 ,add_156_21_n_88 ,add_156_21_n_38);
  and add_156_21_g346(add_156_21_n_89 ,add_156_21_n_9 ,add_156_21_n_88);
  or add_156_21_g347(add_156_21_n_88 ,add_156_21_n_20 ,add_156_21_n_86);
  xnor add_156_21_g348(n_252 ,add_156_21_n_85 ,add_156_21_n_37);
  and add_156_21_g349(add_156_21_n_86 ,add_156_21_n_16 ,add_156_21_n_85);
  or add_156_21_g350(add_156_21_n_85 ,add_156_21_n_10 ,add_156_21_n_83);
  xnor add_156_21_g351(n_251 ,add_156_21_n_82 ,add_156_21_n_36);
  and add_156_21_g352(add_156_21_n_83 ,add_156_21_n_12 ,add_156_21_n_82);
  or add_156_21_g353(add_156_21_n_82 ,add_156_21_n_8 ,add_156_21_n_80);
  xnor add_156_21_g354(n_250 ,add_156_21_n_79 ,add_156_21_n_35);
  and add_156_21_g355(add_156_21_n_80 ,add_156_21_n_22 ,add_156_21_n_79);
  or add_156_21_g356(add_156_21_n_79 ,add_156_21_n_32 ,add_156_21_n_77);
  xnor add_156_21_g357(n_249 ,add_156_21_n_76 ,add_156_21_n_42);
  and add_156_21_g358(add_156_21_n_77 ,add_156_21_n_2 ,add_156_21_n_76);
  or add_156_21_g359(add_156_21_n_76 ,add_156_21_n_21 ,add_156_21_n_74);
  xnor add_156_21_g360(n_248 ,add_156_21_n_73 ,add_156_21_n_48);
  and add_156_21_g361(add_156_21_n_74 ,add_156_21_n_19 ,add_156_21_n_73);
  or add_156_21_g362(add_156_21_n_73 ,add_156_21_n_28 ,add_156_21_n_71);
  xnor add_156_21_g363(n_247 ,add_156_21_n_70 ,add_156_21_n_47);
  and add_156_21_g364(add_156_21_n_71 ,add_156_21_n_11 ,add_156_21_n_70);
  or add_156_21_g365(add_156_21_n_70 ,add_156_21_n_17 ,add_156_21_n_68);
  xnor add_156_21_g366(n_246 ,add_156_21_n_67 ,add_156_21_n_46);
  and add_156_21_g367(add_156_21_n_68 ,add_156_21_n_25 ,add_156_21_n_67);
  or add_156_21_g368(add_156_21_n_67 ,add_156_21_n_6 ,add_156_21_n_65);
  xnor add_156_21_g369(n_245 ,add_156_21_n_64 ,add_156_21_n_45);
  and add_156_21_g370(add_156_21_n_65 ,add_156_21_n_18 ,add_156_21_n_64);
  or add_156_21_g371(add_156_21_n_64 ,add_156_21_n_3 ,add_156_21_n_62);
  xnor add_156_21_g372(n_244 ,add_156_21_n_61 ,add_156_21_n_44);
  and add_156_21_g373(add_156_21_n_62 ,add_156_21_n_30 ,add_156_21_n_61);
  or add_156_21_g374(add_156_21_n_61 ,add_156_21_n_31 ,add_156_21_n_59);
  xnor add_156_21_g375(n_243 ,add_156_21_n_58 ,add_156_21_n_43);
  and add_156_21_g376(add_156_21_n_59 ,add_156_21_n_26 ,add_156_21_n_58);
  or add_156_21_g377(add_156_21_n_58 ,add_156_21_n_27 ,add_156_21_n_56);
  xnor add_156_21_g378(n_242 ,add_156_21_n_55 ,add_156_21_n_34);
  and add_156_21_g379(add_156_21_n_56 ,add_156_21_n_7 ,add_156_21_n_55);
  or add_156_21_g380(add_156_21_n_55 ,add_156_21_n_5 ,add_156_21_n_53);
  xnor add_156_21_g381(n_241 ,add_156_21_n_51 ,add_156_21_n_41);
  and add_156_21_g382(add_156_21_n_53 ,add_156_21_n_23 ,add_156_21_n_51);
  xor add_156_21_g383(n_240 ,add_156_21_n_33 ,add_156_21_n_40);
  or add_156_21_g384(add_156_21_n_51 ,add_156_21_n_4 ,add_156_21_n_49);
  and add_156_21_g385(n_239 ,add_156_21_n_33 ,add_156_21_n_13);
  nor add_156_21_g386(add_156_21_n_49 ,add_156_21_n_33 ,add_156_21_n_14);
  xnor add_156_21_g387(add_156_21_n_48 ,in29[9] ,in30[9]);
  xnor add_156_21_g388(add_156_21_n_47 ,in29[8] ,in30[8]);
  xnor add_156_21_g389(add_156_21_n_46 ,in29[7] ,in30[7]);
  xnor add_156_21_g390(add_156_21_n_45 ,in29[6] ,in30[6]);
  xnor add_156_21_g391(add_156_21_n_44 ,in29[5] ,in30[5]);
  xnor add_156_21_g392(add_156_21_n_43 ,in29[4] ,in30[4]);
  xnor add_156_21_g393(add_156_21_n_42 ,in29[10] ,in30[10]);
  xnor add_156_21_g394(add_156_21_n_41 ,in29[2] ,in30[2]);
  xnor add_156_21_g395(add_156_21_n_40 ,in29[1] ,in30[1]);
  xnor add_156_21_g396(add_156_21_n_39 ,in29[15] ,in30[15]);
  xnor add_156_21_g397(add_156_21_n_38 ,in29[14] ,in30[14]);
  xnor add_156_21_g398(add_156_21_n_37 ,in29[13] ,in30[13]);
  xnor add_156_21_g399(add_156_21_n_36 ,in29[12] ,in30[12]);
  xnor add_156_21_g400(add_156_21_n_35 ,in29[11] ,in30[11]);
  xnor add_156_21_g401(add_156_21_n_34 ,in29[3] ,in30[3]);
  and add_156_21_g402(add_156_21_n_32 ,in29[10] ,in30[10]);
  and add_156_21_g403(add_156_21_n_31 ,in29[4] ,in30[4]);
  or add_156_21_g404(add_156_21_n_30 ,in29[5] ,in30[5]);
  and add_156_21_g405(add_156_21_n_29 ,in29[15] ,in30[15]);
  and add_156_21_g406(add_156_21_n_28 ,in29[8] ,in30[8]);
  and add_156_21_g407(add_156_21_n_27 ,in29[3] ,in30[3]);
  or add_156_21_g408(add_156_21_n_26 ,in29[4] ,in30[4]);
  or add_156_21_g409(add_156_21_n_25 ,in29[7] ,in30[7]);
  and add_156_21_g410(add_156_21_n_24 ,in29[14] ,in30[14]);
  or add_156_21_g411(add_156_21_n_23 ,in29[2] ,in30[2]);
  or add_156_21_g412(add_156_21_n_22 ,in29[11] ,in30[11]);
  and add_156_21_g413(add_156_21_n_21 ,in29[9] ,in30[9]);
  and add_156_21_g414(add_156_21_n_20 ,in29[13] ,in30[13]);
  or add_156_21_g415(add_156_21_n_19 ,in29[9] ,in30[9]);
  or add_156_21_g416(add_156_21_n_18 ,in29[6] ,in30[6]);
  or add_156_21_g417(add_156_21_n_33 ,add_156_21_n_1 ,add_156_21_n_0);
  and add_156_21_g418(add_156_21_n_17 ,in29[7] ,in30[7]);
  or add_156_21_g419(add_156_21_n_16 ,in29[13] ,in30[13]);
  nor add_156_21_g420(add_156_21_n_15 ,in29[15] ,in30[15]);
  nor add_156_21_g421(add_156_21_n_14 ,in29[1] ,in30[1]);
  or add_156_21_g422(add_156_21_n_13 ,in29[0] ,in30[0]);
  or add_156_21_g423(add_156_21_n_12 ,in29[12] ,in30[12]);
  or add_156_21_g424(add_156_21_n_11 ,in29[8] ,in30[8]);
  and add_156_21_g425(add_156_21_n_10 ,in29[12] ,in30[12]);
  or add_156_21_g426(add_156_21_n_9 ,in29[14] ,in30[14]);
  and add_156_21_g427(add_156_21_n_8 ,in29[11] ,in30[11]);
  or add_156_21_g428(add_156_21_n_7 ,in29[3] ,in30[3]);
  and add_156_21_g429(add_156_21_n_6 ,in29[6] ,in30[6]);
  and add_156_21_g430(add_156_21_n_5 ,in29[2] ,in30[2]);
  and add_156_21_g431(add_156_21_n_4 ,in29[1] ,in30[1]);
  and add_156_21_g432(add_156_21_n_3 ,in29[5] ,in30[5]);
  or add_156_21_g433(add_156_21_n_2 ,in29[10] ,in30[10]);
  not add_156_21_g434(add_156_21_n_1 ,in29[0]);
  not add_156_21_g435(add_156_21_n_0 ,in30[0]);
  or add_158_21_g341(n_272 ,add_158_21_n_29 ,add_158_21_n_92);
  xnor add_158_21_g342(n_271 ,add_158_21_n_91 ,add_158_21_n_39);
  nor add_158_21_g343(add_158_21_n_92 ,add_158_21_n_15 ,add_158_21_n_91);
  or add_158_21_g344(add_158_21_n_91 ,add_158_21_n_24 ,add_158_21_n_89);
  xnor add_158_21_g345(n_270 ,add_158_21_n_88 ,add_158_21_n_38);
  and add_158_21_g346(add_158_21_n_89 ,add_158_21_n_9 ,add_158_21_n_88);
  or add_158_21_g347(add_158_21_n_88 ,add_158_21_n_20 ,add_158_21_n_86);
  xnor add_158_21_g348(n_269 ,add_158_21_n_85 ,add_158_21_n_37);
  and add_158_21_g349(add_158_21_n_86 ,add_158_21_n_16 ,add_158_21_n_85);
  or add_158_21_g350(add_158_21_n_85 ,add_158_21_n_10 ,add_158_21_n_83);
  xnor add_158_21_g351(n_268 ,add_158_21_n_82 ,add_158_21_n_36);
  and add_158_21_g352(add_158_21_n_83 ,add_158_21_n_12 ,add_158_21_n_82);
  or add_158_21_g353(add_158_21_n_82 ,add_158_21_n_8 ,add_158_21_n_80);
  xnor add_158_21_g354(n_267 ,add_158_21_n_79 ,add_158_21_n_35);
  and add_158_21_g355(add_158_21_n_80 ,add_158_21_n_22 ,add_158_21_n_79);
  or add_158_21_g356(add_158_21_n_79 ,add_158_21_n_32 ,add_158_21_n_77);
  xnor add_158_21_g357(n_266 ,add_158_21_n_76 ,add_158_21_n_42);
  and add_158_21_g358(add_158_21_n_77 ,add_158_21_n_2 ,add_158_21_n_76);
  or add_158_21_g359(add_158_21_n_76 ,add_158_21_n_21 ,add_158_21_n_74);
  xnor add_158_21_g360(n_265 ,add_158_21_n_73 ,add_158_21_n_48);
  and add_158_21_g361(add_158_21_n_74 ,add_158_21_n_19 ,add_158_21_n_73);
  or add_158_21_g362(add_158_21_n_73 ,add_158_21_n_28 ,add_158_21_n_71);
  xnor add_158_21_g363(n_264 ,add_158_21_n_70 ,add_158_21_n_47);
  and add_158_21_g364(add_158_21_n_71 ,add_158_21_n_11 ,add_158_21_n_70);
  or add_158_21_g365(add_158_21_n_70 ,add_158_21_n_17 ,add_158_21_n_68);
  xnor add_158_21_g366(n_263 ,add_158_21_n_67 ,add_158_21_n_46);
  and add_158_21_g367(add_158_21_n_68 ,add_158_21_n_25 ,add_158_21_n_67);
  or add_158_21_g368(add_158_21_n_67 ,add_158_21_n_6 ,add_158_21_n_65);
  xnor add_158_21_g369(n_262 ,add_158_21_n_64 ,add_158_21_n_45);
  and add_158_21_g370(add_158_21_n_65 ,add_158_21_n_18 ,add_158_21_n_64);
  or add_158_21_g371(add_158_21_n_64 ,add_158_21_n_3 ,add_158_21_n_62);
  xnor add_158_21_g372(n_261 ,add_158_21_n_61 ,add_158_21_n_44);
  and add_158_21_g373(add_158_21_n_62 ,add_158_21_n_30 ,add_158_21_n_61);
  or add_158_21_g374(add_158_21_n_61 ,add_158_21_n_31 ,add_158_21_n_59);
  xnor add_158_21_g375(n_260 ,add_158_21_n_58 ,add_158_21_n_43);
  and add_158_21_g376(add_158_21_n_59 ,add_158_21_n_26 ,add_158_21_n_58);
  or add_158_21_g377(add_158_21_n_58 ,add_158_21_n_27 ,add_158_21_n_56);
  xnor add_158_21_g378(n_259 ,add_158_21_n_55 ,add_158_21_n_34);
  and add_158_21_g379(add_158_21_n_56 ,add_158_21_n_7 ,add_158_21_n_55);
  or add_158_21_g380(add_158_21_n_55 ,add_158_21_n_5 ,add_158_21_n_53);
  xnor add_158_21_g381(n_258 ,add_158_21_n_51 ,add_158_21_n_41);
  and add_158_21_g382(add_158_21_n_53 ,add_158_21_n_23 ,add_158_21_n_51);
  xor add_158_21_g383(n_257 ,add_158_21_n_33 ,add_158_21_n_40);
  or add_158_21_g384(add_158_21_n_51 ,add_158_21_n_4 ,add_158_21_n_49);
  and add_158_21_g385(n_256 ,add_158_21_n_33 ,add_158_21_n_13);
  nor add_158_21_g386(add_158_21_n_49 ,add_158_21_n_33 ,add_158_21_n_14);
  xnor add_158_21_g387(add_158_21_n_48 ,in31[9] ,in32[9]);
  xnor add_158_21_g388(add_158_21_n_47 ,in31[8] ,in32[8]);
  xnor add_158_21_g389(add_158_21_n_46 ,in31[7] ,in32[7]);
  xnor add_158_21_g390(add_158_21_n_45 ,in31[6] ,in32[6]);
  xnor add_158_21_g391(add_158_21_n_44 ,in31[5] ,in32[5]);
  xnor add_158_21_g392(add_158_21_n_43 ,in31[4] ,in32[4]);
  xnor add_158_21_g393(add_158_21_n_42 ,in31[10] ,in32[10]);
  xnor add_158_21_g394(add_158_21_n_41 ,in31[2] ,in32[2]);
  xnor add_158_21_g395(add_158_21_n_40 ,in31[1] ,in32[1]);
  xnor add_158_21_g396(add_158_21_n_39 ,in31[15] ,in32[15]);
  xnor add_158_21_g397(add_158_21_n_38 ,in31[14] ,in32[14]);
  xnor add_158_21_g398(add_158_21_n_37 ,in31[13] ,in32[13]);
  xnor add_158_21_g399(add_158_21_n_36 ,in31[12] ,in32[12]);
  xnor add_158_21_g400(add_158_21_n_35 ,in31[11] ,in32[11]);
  xnor add_158_21_g401(add_158_21_n_34 ,in31[3] ,in32[3]);
  and add_158_21_g402(add_158_21_n_32 ,in31[10] ,in32[10]);
  and add_158_21_g403(add_158_21_n_31 ,in31[4] ,in32[4]);
  or add_158_21_g404(add_158_21_n_30 ,in31[5] ,in32[5]);
  and add_158_21_g405(add_158_21_n_29 ,in31[15] ,in32[15]);
  and add_158_21_g406(add_158_21_n_28 ,in31[8] ,in32[8]);
  and add_158_21_g407(add_158_21_n_27 ,in31[3] ,in32[3]);
  or add_158_21_g408(add_158_21_n_26 ,in31[4] ,in32[4]);
  or add_158_21_g409(add_158_21_n_25 ,in31[7] ,in32[7]);
  and add_158_21_g410(add_158_21_n_24 ,in31[14] ,in32[14]);
  or add_158_21_g411(add_158_21_n_23 ,in31[2] ,in32[2]);
  or add_158_21_g412(add_158_21_n_22 ,in31[11] ,in32[11]);
  and add_158_21_g413(add_158_21_n_21 ,in31[9] ,in32[9]);
  and add_158_21_g414(add_158_21_n_20 ,in31[13] ,in32[13]);
  or add_158_21_g415(add_158_21_n_19 ,in31[9] ,in32[9]);
  or add_158_21_g416(add_158_21_n_18 ,in31[6] ,in32[6]);
  or add_158_21_g417(add_158_21_n_33 ,add_158_21_n_1 ,add_158_21_n_0);
  and add_158_21_g418(add_158_21_n_17 ,in31[7] ,in32[7]);
  or add_158_21_g419(add_158_21_n_16 ,in31[13] ,in32[13]);
  nor add_158_21_g420(add_158_21_n_15 ,in31[15] ,in32[15]);
  nor add_158_21_g421(add_158_21_n_14 ,in31[1] ,in32[1]);
  or add_158_21_g422(add_158_21_n_13 ,in31[0] ,in32[0]);
  or add_158_21_g423(add_158_21_n_12 ,in31[12] ,in32[12]);
  or add_158_21_g424(add_158_21_n_11 ,in31[8] ,in32[8]);
  and add_158_21_g425(add_158_21_n_10 ,in31[12] ,in32[12]);
  or add_158_21_g426(add_158_21_n_9 ,in31[14] ,in32[14]);
  and add_158_21_g427(add_158_21_n_8 ,in31[11] ,in32[11]);
  or add_158_21_g428(add_158_21_n_7 ,in31[3] ,in32[3]);
  and add_158_21_g429(add_158_21_n_6 ,in31[6] ,in32[6]);
  and add_158_21_g430(add_158_21_n_5 ,in31[2] ,in32[2]);
  and add_158_21_g431(add_158_21_n_4 ,in31[1] ,in32[1]);
  and add_158_21_g432(add_158_21_n_3 ,in31[5] ,in32[5]);
  or add_158_21_g433(add_158_21_n_2 ,in31[10] ,in32[10]);
  not add_158_21_g434(add_158_21_n_1 ,in31[0]);
  not add_158_21_g435(add_158_21_n_0 ,in32[0]);
  or add_160_21_g341(n_289 ,add_160_21_n_29 ,add_160_21_n_92);
  xnor add_160_21_g342(n_288 ,add_160_21_n_91 ,add_160_21_n_39);
  nor add_160_21_g343(add_160_21_n_92 ,add_160_21_n_15 ,add_160_21_n_91);
  or add_160_21_g344(add_160_21_n_91 ,add_160_21_n_24 ,add_160_21_n_89);
  xnor add_160_21_g345(n_287 ,add_160_21_n_88 ,add_160_21_n_38);
  and add_160_21_g346(add_160_21_n_89 ,add_160_21_n_9 ,add_160_21_n_88);
  or add_160_21_g347(add_160_21_n_88 ,add_160_21_n_20 ,add_160_21_n_86);
  xnor add_160_21_g348(n_286 ,add_160_21_n_85 ,add_160_21_n_37);
  and add_160_21_g349(add_160_21_n_86 ,add_160_21_n_16 ,add_160_21_n_85);
  or add_160_21_g350(add_160_21_n_85 ,add_160_21_n_10 ,add_160_21_n_83);
  xnor add_160_21_g351(n_285 ,add_160_21_n_82 ,add_160_21_n_36);
  and add_160_21_g352(add_160_21_n_83 ,add_160_21_n_12 ,add_160_21_n_82);
  or add_160_21_g353(add_160_21_n_82 ,add_160_21_n_8 ,add_160_21_n_80);
  xnor add_160_21_g354(n_284 ,add_160_21_n_79 ,add_160_21_n_35);
  and add_160_21_g355(add_160_21_n_80 ,add_160_21_n_22 ,add_160_21_n_79);
  or add_160_21_g356(add_160_21_n_79 ,add_160_21_n_32 ,add_160_21_n_77);
  xnor add_160_21_g357(n_283 ,add_160_21_n_76 ,add_160_21_n_42);
  and add_160_21_g358(add_160_21_n_77 ,add_160_21_n_2 ,add_160_21_n_76);
  or add_160_21_g359(add_160_21_n_76 ,add_160_21_n_21 ,add_160_21_n_74);
  xnor add_160_21_g360(n_282 ,add_160_21_n_73 ,add_160_21_n_48);
  and add_160_21_g361(add_160_21_n_74 ,add_160_21_n_19 ,add_160_21_n_73);
  or add_160_21_g362(add_160_21_n_73 ,add_160_21_n_28 ,add_160_21_n_71);
  xnor add_160_21_g363(n_281 ,add_160_21_n_70 ,add_160_21_n_47);
  and add_160_21_g364(add_160_21_n_71 ,add_160_21_n_11 ,add_160_21_n_70);
  or add_160_21_g365(add_160_21_n_70 ,add_160_21_n_17 ,add_160_21_n_68);
  xnor add_160_21_g366(n_280 ,add_160_21_n_67 ,add_160_21_n_46);
  and add_160_21_g367(add_160_21_n_68 ,add_160_21_n_25 ,add_160_21_n_67);
  or add_160_21_g368(add_160_21_n_67 ,add_160_21_n_6 ,add_160_21_n_65);
  xnor add_160_21_g369(n_279 ,add_160_21_n_64 ,add_160_21_n_45);
  and add_160_21_g370(add_160_21_n_65 ,add_160_21_n_18 ,add_160_21_n_64);
  or add_160_21_g371(add_160_21_n_64 ,add_160_21_n_3 ,add_160_21_n_62);
  xnor add_160_21_g372(n_278 ,add_160_21_n_61 ,add_160_21_n_44);
  and add_160_21_g373(add_160_21_n_62 ,add_160_21_n_30 ,add_160_21_n_61);
  or add_160_21_g374(add_160_21_n_61 ,add_160_21_n_31 ,add_160_21_n_59);
  xnor add_160_21_g375(n_277 ,add_160_21_n_58 ,add_160_21_n_43);
  and add_160_21_g376(add_160_21_n_59 ,add_160_21_n_26 ,add_160_21_n_58);
  or add_160_21_g377(add_160_21_n_58 ,add_160_21_n_27 ,add_160_21_n_56);
  xnor add_160_21_g378(n_276 ,add_160_21_n_55 ,add_160_21_n_34);
  and add_160_21_g379(add_160_21_n_56 ,add_160_21_n_7 ,add_160_21_n_55);
  or add_160_21_g380(add_160_21_n_55 ,add_160_21_n_5 ,add_160_21_n_53);
  xnor add_160_21_g381(n_275 ,add_160_21_n_51 ,add_160_21_n_41);
  and add_160_21_g382(add_160_21_n_53 ,add_160_21_n_23 ,add_160_21_n_51);
  xor add_160_21_g383(n_274 ,add_160_21_n_33 ,add_160_21_n_40);
  or add_160_21_g384(add_160_21_n_51 ,add_160_21_n_4 ,add_160_21_n_49);
  and add_160_21_g385(n_273 ,add_160_21_n_33 ,add_160_21_n_13);
  nor add_160_21_g386(add_160_21_n_49 ,add_160_21_n_33 ,add_160_21_n_14);
  xnor add_160_21_g387(add_160_21_n_48 ,in33[9] ,in34[9]);
  xnor add_160_21_g388(add_160_21_n_47 ,in33[8] ,in34[8]);
  xnor add_160_21_g389(add_160_21_n_46 ,in33[7] ,in34[7]);
  xnor add_160_21_g390(add_160_21_n_45 ,in33[6] ,in34[6]);
  xnor add_160_21_g391(add_160_21_n_44 ,in33[5] ,in34[5]);
  xnor add_160_21_g392(add_160_21_n_43 ,in33[4] ,in34[4]);
  xnor add_160_21_g393(add_160_21_n_42 ,in33[10] ,in34[10]);
  xnor add_160_21_g394(add_160_21_n_41 ,in33[2] ,in34[2]);
  xnor add_160_21_g395(add_160_21_n_40 ,in33[1] ,in34[1]);
  xnor add_160_21_g396(add_160_21_n_39 ,in33[15] ,in34[15]);
  xnor add_160_21_g397(add_160_21_n_38 ,in33[14] ,in34[14]);
  xnor add_160_21_g398(add_160_21_n_37 ,in33[13] ,in34[13]);
  xnor add_160_21_g399(add_160_21_n_36 ,in33[12] ,in34[12]);
  xnor add_160_21_g400(add_160_21_n_35 ,in33[11] ,in34[11]);
  xnor add_160_21_g401(add_160_21_n_34 ,in33[3] ,in34[3]);
  and add_160_21_g402(add_160_21_n_32 ,in33[10] ,in34[10]);
  and add_160_21_g403(add_160_21_n_31 ,in33[4] ,in34[4]);
  or add_160_21_g404(add_160_21_n_30 ,in33[5] ,in34[5]);
  and add_160_21_g405(add_160_21_n_29 ,in33[15] ,in34[15]);
  and add_160_21_g406(add_160_21_n_28 ,in33[8] ,in34[8]);
  and add_160_21_g407(add_160_21_n_27 ,in33[3] ,in34[3]);
  or add_160_21_g408(add_160_21_n_26 ,in33[4] ,in34[4]);
  or add_160_21_g409(add_160_21_n_25 ,in33[7] ,in34[7]);
  and add_160_21_g410(add_160_21_n_24 ,in33[14] ,in34[14]);
  or add_160_21_g411(add_160_21_n_23 ,in33[2] ,in34[2]);
  or add_160_21_g412(add_160_21_n_22 ,in33[11] ,in34[11]);
  and add_160_21_g413(add_160_21_n_21 ,in33[9] ,in34[9]);
  and add_160_21_g414(add_160_21_n_20 ,in33[13] ,in34[13]);
  or add_160_21_g415(add_160_21_n_19 ,in33[9] ,in34[9]);
  or add_160_21_g416(add_160_21_n_18 ,in33[6] ,in34[6]);
  or add_160_21_g417(add_160_21_n_33 ,add_160_21_n_1 ,add_160_21_n_0);
  and add_160_21_g418(add_160_21_n_17 ,in33[7] ,in34[7]);
  or add_160_21_g419(add_160_21_n_16 ,in33[13] ,in34[13]);
  nor add_160_21_g420(add_160_21_n_15 ,in33[15] ,in34[15]);
  nor add_160_21_g421(add_160_21_n_14 ,in33[1] ,in34[1]);
  or add_160_21_g422(add_160_21_n_13 ,in33[0] ,in34[0]);
  or add_160_21_g423(add_160_21_n_12 ,in33[12] ,in34[12]);
  or add_160_21_g424(add_160_21_n_11 ,in33[8] ,in34[8]);
  and add_160_21_g425(add_160_21_n_10 ,in33[12] ,in34[12]);
  or add_160_21_g426(add_160_21_n_9 ,in33[14] ,in34[14]);
  and add_160_21_g427(add_160_21_n_8 ,in33[11] ,in34[11]);
  or add_160_21_g428(add_160_21_n_7 ,in33[3] ,in34[3]);
  and add_160_21_g429(add_160_21_n_6 ,in33[6] ,in34[6]);
  and add_160_21_g430(add_160_21_n_5 ,in33[2] ,in34[2]);
  and add_160_21_g431(add_160_21_n_4 ,in33[1] ,in34[1]);
  and add_160_21_g432(add_160_21_n_3 ,in33[5] ,in34[5]);
  or add_160_21_g433(add_160_21_n_2 ,in33[10] ,in34[10]);
  not add_160_21_g434(add_160_21_n_1 ,in33[0]);
  not add_160_21_g435(add_160_21_n_0 ,in34[0]);
  or add_162_21_g341(n_306 ,add_162_21_n_29 ,add_162_21_n_92);
  xnor add_162_21_g342(n_305 ,add_162_21_n_91 ,add_162_21_n_39);
  nor add_162_21_g343(add_162_21_n_92 ,add_162_21_n_15 ,add_162_21_n_91);
  or add_162_21_g344(add_162_21_n_91 ,add_162_21_n_24 ,add_162_21_n_89);
  xnor add_162_21_g345(n_304 ,add_162_21_n_88 ,add_162_21_n_38);
  and add_162_21_g346(add_162_21_n_89 ,add_162_21_n_9 ,add_162_21_n_88);
  or add_162_21_g347(add_162_21_n_88 ,add_162_21_n_20 ,add_162_21_n_86);
  xnor add_162_21_g348(n_303 ,add_162_21_n_85 ,add_162_21_n_37);
  and add_162_21_g349(add_162_21_n_86 ,add_162_21_n_16 ,add_162_21_n_85);
  or add_162_21_g350(add_162_21_n_85 ,add_162_21_n_10 ,add_162_21_n_83);
  xnor add_162_21_g351(n_302 ,add_162_21_n_82 ,add_162_21_n_36);
  and add_162_21_g352(add_162_21_n_83 ,add_162_21_n_12 ,add_162_21_n_82);
  or add_162_21_g353(add_162_21_n_82 ,add_162_21_n_8 ,add_162_21_n_80);
  xnor add_162_21_g354(n_301 ,add_162_21_n_79 ,add_162_21_n_35);
  and add_162_21_g355(add_162_21_n_80 ,add_162_21_n_22 ,add_162_21_n_79);
  or add_162_21_g356(add_162_21_n_79 ,add_162_21_n_32 ,add_162_21_n_77);
  xnor add_162_21_g357(n_300 ,add_162_21_n_76 ,add_162_21_n_42);
  and add_162_21_g358(add_162_21_n_77 ,add_162_21_n_2 ,add_162_21_n_76);
  or add_162_21_g359(add_162_21_n_76 ,add_162_21_n_21 ,add_162_21_n_74);
  xnor add_162_21_g360(n_299 ,add_162_21_n_73 ,add_162_21_n_48);
  and add_162_21_g361(add_162_21_n_74 ,add_162_21_n_19 ,add_162_21_n_73);
  or add_162_21_g362(add_162_21_n_73 ,add_162_21_n_28 ,add_162_21_n_71);
  xnor add_162_21_g363(n_298 ,add_162_21_n_70 ,add_162_21_n_47);
  and add_162_21_g364(add_162_21_n_71 ,add_162_21_n_11 ,add_162_21_n_70);
  or add_162_21_g365(add_162_21_n_70 ,add_162_21_n_17 ,add_162_21_n_68);
  xnor add_162_21_g366(n_297 ,add_162_21_n_67 ,add_162_21_n_46);
  and add_162_21_g367(add_162_21_n_68 ,add_162_21_n_25 ,add_162_21_n_67);
  or add_162_21_g368(add_162_21_n_67 ,add_162_21_n_6 ,add_162_21_n_65);
  xnor add_162_21_g369(n_296 ,add_162_21_n_64 ,add_162_21_n_45);
  and add_162_21_g370(add_162_21_n_65 ,add_162_21_n_18 ,add_162_21_n_64);
  or add_162_21_g371(add_162_21_n_64 ,add_162_21_n_3 ,add_162_21_n_62);
  xnor add_162_21_g372(n_295 ,add_162_21_n_61 ,add_162_21_n_44);
  and add_162_21_g373(add_162_21_n_62 ,add_162_21_n_30 ,add_162_21_n_61);
  or add_162_21_g374(add_162_21_n_61 ,add_162_21_n_31 ,add_162_21_n_59);
  xnor add_162_21_g375(n_294 ,add_162_21_n_58 ,add_162_21_n_43);
  and add_162_21_g376(add_162_21_n_59 ,add_162_21_n_26 ,add_162_21_n_58);
  or add_162_21_g377(add_162_21_n_58 ,add_162_21_n_27 ,add_162_21_n_56);
  xnor add_162_21_g378(n_293 ,add_162_21_n_55 ,add_162_21_n_34);
  and add_162_21_g379(add_162_21_n_56 ,add_162_21_n_7 ,add_162_21_n_55);
  or add_162_21_g380(add_162_21_n_55 ,add_162_21_n_5 ,add_162_21_n_53);
  xnor add_162_21_g381(n_292 ,add_162_21_n_51 ,add_162_21_n_41);
  and add_162_21_g382(add_162_21_n_53 ,add_162_21_n_23 ,add_162_21_n_51);
  xor add_162_21_g383(n_291 ,add_162_21_n_33 ,add_162_21_n_40);
  or add_162_21_g384(add_162_21_n_51 ,add_162_21_n_4 ,add_162_21_n_49);
  and add_162_21_g385(n_290 ,add_162_21_n_33 ,add_162_21_n_13);
  nor add_162_21_g386(add_162_21_n_49 ,add_162_21_n_33 ,add_162_21_n_14);
  xnor add_162_21_g387(add_162_21_n_48 ,in35[9] ,in36[9]);
  xnor add_162_21_g388(add_162_21_n_47 ,in35[8] ,in36[8]);
  xnor add_162_21_g389(add_162_21_n_46 ,in35[7] ,in36[7]);
  xnor add_162_21_g390(add_162_21_n_45 ,in35[6] ,in36[6]);
  xnor add_162_21_g391(add_162_21_n_44 ,in35[5] ,in36[5]);
  xnor add_162_21_g392(add_162_21_n_43 ,in35[4] ,in36[4]);
  xnor add_162_21_g393(add_162_21_n_42 ,in35[10] ,in36[10]);
  xnor add_162_21_g394(add_162_21_n_41 ,in35[2] ,in36[2]);
  xnor add_162_21_g395(add_162_21_n_40 ,in35[1] ,in36[1]);
  xnor add_162_21_g396(add_162_21_n_39 ,in35[15] ,in36[15]);
  xnor add_162_21_g397(add_162_21_n_38 ,in35[14] ,in36[14]);
  xnor add_162_21_g398(add_162_21_n_37 ,in35[13] ,in36[13]);
  xnor add_162_21_g399(add_162_21_n_36 ,in35[12] ,in36[12]);
  xnor add_162_21_g400(add_162_21_n_35 ,in35[11] ,in36[11]);
  xnor add_162_21_g401(add_162_21_n_34 ,in35[3] ,in36[3]);
  and add_162_21_g402(add_162_21_n_32 ,in35[10] ,in36[10]);
  and add_162_21_g403(add_162_21_n_31 ,in35[4] ,in36[4]);
  or add_162_21_g404(add_162_21_n_30 ,in35[5] ,in36[5]);
  and add_162_21_g405(add_162_21_n_29 ,in35[15] ,in36[15]);
  and add_162_21_g406(add_162_21_n_28 ,in35[8] ,in36[8]);
  and add_162_21_g407(add_162_21_n_27 ,in35[3] ,in36[3]);
  or add_162_21_g408(add_162_21_n_26 ,in35[4] ,in36[4]);
  or add_162_21_g409(add_162_21_n_25 ,in35[7] ,in36[7]);
  and add_162_21_g410(add_162_21_n_24 ,in35[14] ,in36[14]);
  or add_162_21_g411(add_162_21_n_23 ,in35[2] ,in36[2]);
  or add_162_21_g412(add_162_21_n_22 ,in35[11] ,in36[11]);
  and add_162_21_g413(add_162_21_n_21 ,in35[9] ,in36[9]);
  and add_162_21_g414(add_162_21_n_20 ,in35[13] ,in36[13]);
  or add_162_21_g415(add_162_21_n_19 ,in35[9] ,in36[9]);
  or add_162_21_g416(add_162_21_n_18 ,in35[6] ,in36[6]);
  or add_162_21_g417(add_162_21_n_33 ,add_162_21_n_1 ,add_162_21_n_0);
  and add_162_21_g418(add_162_21_n_17 ,in35[7] ,in36[7]);
  or add_162_21_g419(add_162_21_n_16 ,in35[13] ,in36[13]);
  nor add_162_21_g420(add_162_21_n_15 ,in35[15] ,in36[15]);
  nor add_162_21_g421(add_162_21_n_14 ,in35[1] ,in36[1]);
  or add_162_21_g422(add_162_21_n_13 ,in35[0] ,in36[0]);
  or add_162_21_g423(add_162_21_n_12 ,in35[12] ,in36[12]);
  or add_162_21_g424(add_162_21_n_11 ,in35[8] ,in36[8]);
  and add_162_21_g425(add_162_21_n_10 ,in35[12] ,in36[12]);
  or add_162_21_g426(add_162_21_n_9 ,in35[14] ,in36[14]);
  and add_162_21_g427(add_162_21_n_8 ,in35[11] ,in36[11]);
  or add_162_21_g428(add_162_21_n_7 ,in35[3] ,in36[3]);
  and add_162_21_g429(add_162_21_n_6 ,in35[6] ,in36[6]);
  and add_162_21_g430(add_162_21_n_5 ,in35[2] ,in36[2]);
  and add_162_21_g431(add_162_21_n_4 ,in35[1] ,in36[1]);
  and add_162_21_g432(add_162_21_n_3 ,in35[5] ,in36[5]);
  or add_162_21_g433(add_162_21_n_2 ,in35[10] ,in36[10]);
  not add_162_21_g434(add_162_21_n_1 ,in35[0]);
  not add_162_21_g435(add_162_21_n_0 ,in36[0]);
  or add_164_21_g341(n_323 ,add_164_21_n_29 ,add_164_21_n_92);
  xnor add_164_21_g342(n_322 ,add_164_21_n_91 ,add_164_21_n_39);
  nor add_164_21_g343(add_164_21_n_92 ,add_164_21_n_15 ,add_164_21_n_91);
  or add_164_21_g344(add_164_21_n_91 ,add_164_21_n_24 ,add_164_21_n_89);
  xnor add_164_21_g345(n_321 ,add_164_21_n_88 ,add_164_21_n_38);
  and add_164_21_g346(add_164_21_n_89 ,add_164_21_n_9 ,add_164_21_n_88);
  or add_164_21_g347(add_164_21_n_88 ,add_164_21_n_20 ,add_164_21_n_86);
  xnor add_164_21_g348(n_320 ,add_164_21_n_85 ,add_164_21_n_37);
  and add_164_21_g349(add_164_21_n_86 ,add_164_21_n_16 ,add_164_21_n_85);
  or add_164_21_g350(add_164_21_n_85 ,add_164_21_n_10 ,add_164_21_n_83);
  xnor add_164_21_g351(n_319 ,add_164_21_n_82 ,add_164_21_n_36);
  and add_164_21_g352(add_164_21_n_83 ,add_164_21_n_12 ,add_164_21_n_82);
  or add_164_21_g353(add_164_21_n_82 ,add_164_21_n_8 ,add_164_21_n_80);
  xnor add_164_21_g354(n_318 ,add_164_21_n_79 ,add_164_21_n_35);
  and add_164_21_g355(add_164_21_n_80 ,add_164_21_n_22 ,add_164_21_n_79);
  or add_164_21_g356(add_164_21_n_79 ,add_164_21_n_32 ,add_164_21_n_77);
  xnor add_164_21_g357(n_317 ,add_164_21_n_76 ,add_164_21_n_42);
  and add_164_21_g358(add_164_21_n_77 ,add_164_21_n_2 ,add_164_21_n_76);
  or add_164_21_g359(add_164_21_n_76 ,add_164_21_n_21 ,add_164_21_n_74);
  xnor add_164_21_g360(n_316 ,add_164_21_n_73 ,add_164_21_n_48);
  and add_164_21_g361(add_164_21_n_74 ,add_164_21_n_19 ,add_164_21_n_73);
  or add_164_21_g362(add_164_21_n_73 ,add_164_21_n_28 ,add_164_21_n_71);
  xnor add_164_21_g363(n_315 ,add_164_21_n_70 ,add_164_21_n_47);
  and add_164_21_g364(add_164_21_n_71 ,add_164_21_n_11 ,add_164_21_n_70);
  or add_164_21_g365(add_164_21_n_70 ,add_164_21_n_17 ,add_164_21_n_68);
  xnor add_164_21_g366(n_314 ,add_164_21_n_67 ,add_164_21_n_46);
  and add_164_21_g367(add_164_21_n_68 ,add_164_21_n_25 ,add_164_21_n_67);
  or add_164_21_g368(add_164_21_n_67 ,add_164_21_n_6 ,add_164_21_n_65);
  xnor add_164_21_g369(n_313 ,add_164_21_n_64 ,add_164_21_n_45);
  and add_164_21_g370(add_164_21_n_65 ,add_164_21_n_18 ,add_164_21_n_64);
  or add_164_21_g371(add_164_21_n_64 ,add_164_21_n_3 ,add_164_21_n_62);
  xnor add_164_21_g372(n_312 ,add_164_21_n_61 ,add_164_21_n_44);
  and add_164_21_g373(add_164_21_n_62 ,add_164_21_n_30 ,add_164_21_n_61);
  or add_164_21_g374(add_164_21_n_61 ,add_164_21_n_31 ,add_164_21_n_59);
  xnor add_164_21_g375(n_311 ,add_164_21_n_58 ,add_164_21_n_43);
  and add_164_21_g376(add_164_21_n_59 ,add_164_21_n_26 ,add_164_21_n_58);
  or add_164_21_g377(add_164_21_n_58 ,add_164_21_n_27 ,add_164_21_n_56);
  xnor add_164_21_g378(n_310 ,add_164_21_n_55 ,add_164_21_n_34);
  and add_164_21_g379(add_164_21_n_56 ,add_164_21_n_7 ,add_164_21_n_55);
  or add_164_21_g380(add_164_21_n_55 ,add_164_21_n_5 ,add_164_21_n_53);
  xnor add_164_21_g381(n_309 ,add_164_21_n_51 ,add_164_21_n_41);
  and add_164_21_g382(add_164_21_n_53 ,add_164_21_n_23 ,add_164_21_n_51);
  xor add_164_21_g383(n_308 ,add_164_21_n_33 ,add_164_21_n_40);
  or add_164_21_g384(add_164_21_n_51 ,add_164_21_n_4 ,add_164_21_n_49);
  and add_164_21_g385(n_307 ,add_164_21_n_33 ,add_164_21_n_13);
  nor add_164_21_g386(add_164_21_n_49 ,add_164_21_n_33 ,add_164_21_n_14);
  xnor add_164_21_g387(add_164_21_n_48 ,in37[9] ,in38[9]);
  xnor add_164_21_g388(add_164_21_n_47 ,in37[8] ,in38[8]);
  xnor add_164_21_g389(add_164_21_n_46 ,in37[7] ,in38[7]);
  xnor add_164_21_g390(add_164_21_n_45 ,in37[6] ,in38[6]);
  xnor add_164_21_g391(add_164_21_n_44 ,in37[5] ,in38[5]);
  xnor add_164_21_g392(add_164_21_n_43 ,in37[4] ,in38[4]);
  xnor add_164_21_g393(add_164_21_n_42 ,in37[10] ,in38[10]);
  xnor add_164_21_g394(add_164_21_n_41 ,in37[2] ,in38[2]);
  xnor add_164_21_g395(add_164_21_n_40 ,in37[1] ,in38[1]);
  xnor add_164_21_g396(add_164_21_n_39 ,in37[15] ,in38[15]);
  xnor add_164_21_g397(add_164_21_n_38 ,in37[14] ,in38[14]);
  xnor add_164_21_g398(add_164_21_n_37 ,in37[13] ,in38[13]);
  xnor add_164_21_g399(add_164_21_n_36 ,in37[12] ,in38[12]);
  xnor add_164_21_g400(add_164_21_n_35 ,in37[11] ,in38[11]);
  xnor add_164_21_g401(add_164_21_n_34 ,in37[3] ,in38[3]);
  and add_164_21_g402(add_164_21_n_32 ,in37[10] ,in38[10]);
  and add_164_21_g403(add_164_21_n_31 ,in37[4] ,in38[4]);
  or add_164_21_g404(add_164_21_n_30 ,in37[5] ,in38[5]);
  and add_164_21_g405(add_164_21_n_29 ,in37[15] ,in38[15]);
  and add_164_21_g406(add_164_21_n_28 ,in37[8] ,in38[8]);
  and add_164_21_g407(add_164_21_n_27 ,in37[3] ,in38[3]);
  or add_164_21_g408(add_164_21_n_26 ,in37[4] ,in38[4]);
  or add_164_21_g409(add_164_21_n_25 ,in37[7] ,in38[7]);
  and add_164_21_g410(add_164_21_n_24 ,in37[14] ,in38[14]);
  or add_164_21_g411(add_164_21_n_23 ,in37[2] ,in38[2]);
  or add_164_21_g412(add_164_21_n_22 ,in37[11] ,in38[11]);
  and add_164_21_g413(add_164_21_n_21 ,in37[9] ,in38[9]);
  and add_164_21_g414(add_164_21_n_20 ,in37[13] ,in38[13]);
  or add_164_21_g415(add_164_21_n_19 ,in37[9] ,in38[9]);
  or add_164_21_g416(add_164_21_n_18 ,in37[6] ,in38[6]);
  or add_164_21_g417(add_164_21_n_33 ,add_164_21_n_1 ,add_164_21_n_0);
  and add_164_21_g418(add_164_21_n_17 ,in37[7] ,in38[7]);
  or add_164_21_g419(add_164_21_n_16 ,in37[13] ,in38[13]);
  nor add_164_21_g420(add_164_21_n_15 ,in37[15] ,in38[15]);
  nor add_164_21_g421(add_164_21_n_14 ,in37[1] ,in38[1]);
  or add_164_21_g422(add_164_21_n_13 ,in37[0] ,in38[0]);
  or add_164_21_g423(add_164_21_n_12 ,in37[12] ,in38[12]);
  or add_164_21_g424(add_164_21_n_11 ,in37[8] ,in38[8]);
  and add_164_21_g425(add_164_21_n_10 ,in37[12] ,in38[12]);
  or add_164_21_g426(add_164_21_n_9 ,in37[14] ,in38[14]);
  and add_164_21_g427(add_164_21_n_8 ,in37[11] ,in38[11]);
  or add_164_21_g428(add_164_21_n_7 ,in37[3] ,in38[3]);
  and add_164_21_g429(add_164_21_n_6 ,in37[6] ,in38[6]);
  and add_164_21_g430(add_164_21_n_5 ,in37[2] ,in38[2]);
  and add_164_21_g431(add_164_21_n_4 ,in37[1] ,in38[1]);
  and add_164_21_g432(add_164_21_n_3 ,in37[5] ,in38[5]);
  or add_164_21_g433(add_164_21_n_2 ,in37[10] ,in38[10]);
  not add_164_21_g434(add_164_21_n_1 ,in37[0]);
  not add_164_21_g435(add_164_21_n_0 ,in38[0]);
  or add_166_21_g341(n_340 ,add_166_21_n_29 ,add_166_21_n_92);
  xnor add_166_21_g342(n_339 ,add_166_21_n_91 ,add_166_21_n_39);
  nor add_166_21_g343(add_166_21_n_92 ,add_166_21_n_15 ,add_166_21_n_91);
  or add_166_21_g344(add_166_21_n_91 ,add_166_21_n_24 ,add_166_21_n_89);
  xnor add_166_21_g345(n_338 ,add_166_21_n_88 ,add_166_21_n_38);
  and add_166_21_g346(add_166_21_n_89 ,add_166_21_n_9 ,add_166_21_n_88);
  or add_166_21_g347(add_166_21_n_88 ,add_166_21_n_20 ,add_166_21_n_86);
  xnor add_166_21_g348(n_337 ,add_166_21_n_85 ,add_166_21_n_37);
  and add_166_21_g349(add_166_21_n_86 ,add_166_21_n_16 ,add_166_21_n_85);
  or add_166_21_g350(add_166_21_n_85 ,add_166_21_n_10 ,add_166_21_n_83);
  xnor add_166_21_g351(n_336 ,add_166_21_n_82 ,add_166_21_n_36);
  and add_166_21_g352(add_166_21_n_83 ,add_166_21_n_12 ,add_166_21_n_82);
  or add_166_21_g353(add_166_21_n_82 ,add_166_21_n_8 ,add_166_21_n_80);
  xnor add_166_21_g354(n_335 ,add_166_21_n_79 ,add_166_21_n_35);
  and add_166_21_g355(add_166_21_n_80 ,add_166_21_n_22 ,add_166_21_n_79);
  or add_166_21_g356(add_166_21_n_79 ,add_166_21_n_32 ,add_166_21_n_77);
  xnor add_166_21_g357(n_334 ,add_166_21_n_76 ,add_166_21_n_42);
  and add_166_21_g358(add_166_21_n_77 ,add_166_21_n_2 ,add_166_21_n_76);
  or add_166_21_g359(add_166_21_n_76 ,add_166_21_n_21 ,add_166_21_n_74);
  xnor add_166_21_g360(n_333 ,add_166_21_n_73 ,add_166_21_n_48);
  and add_166_21_g361(add_166_21_n_74 ,add_166_21_n_19 ,add_166_21_n_73);
  or add_166_21_g362(add_166_21_n_73 ,add_166_21_n_28 ,add_166_21_n_71);
  xnor add_166_21_g363(n_332 ,add_166_21_n_70 ,add_166_21_n_47);
  and add_166_21_g364(add_166_21_n_71 ,add_166_21_n_11 ,add_166_21_n_70);
  or add_166_21_g365(add_166_21_n_70 ,add_166_21_n_17 ,add_166_21_n_68);
  xnor add_166_21_g366(n_331 ,add_166_21_n_67 ,add_166_21_n_46);
  and add_166_21_g367(add_166_21_n_68 ,add_166_21_n_25 ,add_166_21_n_67);
  or add_166_21_g368(add_166_21_n_67 ,add_166_21_n_6 ,add_166_21_n_65);
  xnor add_166_21_g369(n_330 ,add_166_21_n_64 ,add_166_21_n_45);
  and add_166_21_g370(add_166_21_n_65 ,add_166_21_n_18 ,add_166_21_n_64);
  or add_166_21_g371(add_166_21_n_64 ,add_166_21_n_3 ,add_166_21_n_62);
  xnor add_166_21_g372(n_329 ,add_166_21_n_61 ,add_166_21_n_44);
  and add_166_21_g373(add_166_21_n_62 ,add_166_21_n_30 ,add_166_21_n_61);
  or add_166_21_g374(add_166_21_n_61 ,add_166_21_n_31 ,add_166_21_n_59);
  xnor add_166_21_g375(n_328 ,add_166_21_n_58 ,add_166_21_n_43);
  and add_166_21_g376(add_166_21_n_59 ,add_166_21_n_26 ,add_166_21_n_58);
  or add_166_21_g377(add_166_21_n_58 ,add_166_21_n_27 ,add_166_21_n_56);
  xnor add_166_21_g378(n_327 ,add_166_21_n_55 ,add_166_21_n_34);
  and add_166_21_g379(add_166_21_n_56 ,add_166_21_n_7 ,add_166_21_n_55);
  or add_166_21_g380(add_166_21_n_55 ,add_166_21_n_5 ,add_166_21_n_53);
  xnor add_166_21_g381(n_326 ,add_166_21_n_51 ,add_166_21_n_41);
  and add_166_21_g382(add_166_21_n_53 ,add_166_21_n_23 ,add_166_21_n_51);
  xor add_166_21_g383(n_325 ,add_166_21_n_33 ,add_166_21_n_40);
  or add_166_21_g384(add_166_21_n_51 ,add_166_21_n_4 ,add_166_21_n_49);
  and add_166_21_g385(n_324 ,add_166_21_n_33 ,add_166_21_n_13);
  nor add_166_21_g386(add_166_21_n_49 ,add_166_21_n_33 ,add_166_21_n_14);
  xnor add_166_21_g387(add_166_21_n_48 ,in39[9] ,in40[9]);
  xnor add_166_21_g388(add_166_21_n_47 ,in39[8] ,in40[8]);
  xnor add_166_21_g389(add_166_21_n_46 ,in39[7] ,in40[7]);
  xnor add_166_21_g390(add_166_21_n_45 ,in39[6] ,in40[6]);
  xnor add_166_21_g391(add_166_21_n_44 ,in39[5] ,in40[5]);
  xnor add_166_21_g392(add_166_21_n_43 ,in39[4] ,in40[4]);
  xnor add_166_21_g393(add_166_21_n_42 ,in39[10] ,in40[10]);
  xnor add_166_21_g394(add_166_21_n_41 ,in39[2] ,in40[2]);
  xnor add_166_21_g395(add_166_21_n_40 ,in39[1] ,in40[1]);
  xnor add_166_21_g396(add_166_21_n_39 ,in39[15] ,in40[15]);
  xnor add_166_21_g397(add_166_21_n_38 ,in39[14] ,in40[14]);
  xnor add_166_21_g398(add_166_21_n_37 ,in39[13] ,in40[13]);
  xnor add_166_21_g399(add_166_21_n_36 ,in39[12] ,in40[12]);
  xnor add_166_21_g400(add_166_21_n_35 ,in39[11] ,in40[11]);
  xnor add_166_21_g401(add_166_21_n_34 ,in39[3] ,in40[3]);
  and add_166_21_g402(add_166_21_n_32 ,in39[10] ,in40[10]);
  and add_166_21_g403(add_166_21_n_31 ,in39[4] ,in40[4]);
  or add_166_21_g404(add_166_21_n_30 ,in39[5] ,in40[5]);
  and add_166_21_g405(add_166_21_n_29 ,in39[15] ,in40[15]);
  and add_166_21_g406(add_166_21_n_28 ,in39[8] ,in40[8]);
  and add_166_21_g407(add_166_21_n_27 ,in39[3] ,in40[3]);
  or add_166_21_g408(add_166_21_n_26 ,in39[4] ,in40[4]);
  or add_166_21_g409(add_166_21_n_25 ,in39[7] ,in40[7]);
  and add_166_21_g410(add_166_21_n_24 ,in39[14] ,in40[14]);
  or add_166_21_g411(add_166_21_n_23 ,in39[2] ,in40[2]);
  or add_166_21_g412(add_166_21_n_22 ,in39[11] ,in40[11]);
  and add_166_21_g413(add_166_21_n_21 ,in39[9] ,in40[9]);
  and add_166_21_g414(add_166_21_n_20 ,in39[13] ,in40[13]);
  or add_166_21_g415(add_166_21_n_19 ,in39[9] ,in40[9]);
  or add_166_21_g416(add_166_21_n_18 ,in39[6] ,in40[6]);
  or add_166_21_g417(add_166_21_n_33 ,add_166_21_n_1 ,add_166_21_n_0);
  and add_166_21_g418(add_166_21_n_17 ,in39[7] ,in40[7]);
  or add_166_21_g419(add_166_21_n_16 ,in39[13] ,in40[13]);
  nor add_166_21_g420(add_166_21_n_15 ,in39[15] ,in40[15]);
  nor add_166_21_g421(add_166_21_n_14 ,in39[1] ,in40[1]);
  or add_166_21_g422(add_166_21_n_13 ,in39[0] ,in40[0]);
  or add_166_21_g423(add_166_21_n_12 ,in39[12] ,in40[12]);
  or add_166_21_g424(add_166_21_n_11 ,in39[8] ,in40[8]);
  and add_166_21_g425(add_166_21_n_10 ,in39[12] ,in40[12]);
  or add_166_21_g426(add_166_21_n_9 ,in39[14] ,in40[14]);
  and add_166_21_g427(add_166_21_n_8 ,in39[11] ,in40[11]);
  or add_166_21_g428(add_166_21_n_7 ,in39[3] ,in40[3]);
  and add_166_21_g429(add_166_21_n_6 ,in39[6] ,in40[6]);
  and add_166_21_g430(add_166_21_n_5 ,in39[2] ,in40[2]);
  and add_166_21_g431(add_166_21_n_4 ,in39[1] ,in40[1]);
  and add_166_21_g432(add_166_21_n_3 ,in39[5] ,in40[5]);
  or add_166_21_g433(add_166_21_n_2 ,in39[10] ,in40[10]);
  not add_166_21_g434(add_166_21_n_1 ,in39[0]);
  not add_166_21_g435(add_166_21_n_0 ,in40[0]);
  or add_168_21_g341(n_357 ,add_168_21_n_29 ,add_168_21_n_92);
  xnor add_168_21_g342(n_356 ,add_168_21_n_91 ,add_168_21_n_39);
  nor add_168_21_g343(add_168_21_n_92 ,add_168_21_n_15 ,add_168_21_n_91);
  or add_168_21_g344(add_168_21_n_91 ,add_168_21_n_24 ,add_168_21_n_89);
  xnor add_168_21_g345(n_355 ,add_168_21_n_88 ,add_168_21_n_38);
  and add_168_21_g346(add_168_21_n_89 ,add_168_21_n_9 ,add_168_21_n_88);
  or add_168_21_g347(add_168_21_n_88 ,add_168_21_n_20 ,add_168_21_n_86);
  xnor add_168_21_g348(n_354 ,add_168_21_n_85 ,add_168_21_n_37);
  and add_168_21_g349(add_168_21_n_86 ,add_168_21_n_16 ,add_168_21_n_85);
  or add_168_21_g350(add_168_21_n_85 ,add_168_21_n_10 ,add_168_21_n_83);
  xnor add_168_21_g351(n_353 ,add_168_21_n_82 ,add_168_21_n_36);
  and add_168_21_g352(add_168_21_n_83 ,add_168_21_n_12 ,add_168_21_n_82);
  or add_168_21_g353(add_168_21_n_82 ,add_168_21_n_8 ,add_168_21_n_80);
  xnor add_168_21_g354(n_352 ,add_168_21_n_79 ,add_168_21_n_35);
  and add_168_21_g355(add_168_21_n_80 ,add_168_21_n_22 ,add_168_21_n_79);
  or add_168_21_g356(add_168_21_n_79 ,add_168_21_n_32 ,add_168_21_n_77);
  xnor add_168_21_g357(n_351 ,add_168_21_n_76 ,add_168_21_n_42);
  and add_168_21_g358(add_168_21_n_77 ,add_168_21_n_2 ,add_168_21_n_76);
  or add_168_21_g359(add_168_21_n_76 ,add_168_21_n_21 ,add_168_21_n_74);
  xnor add_168_21_g360(n_350 ,add_168_21_n_73 ,add_168_21_n_48);
  and add_168_21_g361(add_168_21_n_74 ,add_168_21_n_19 ,add_168_21_n_73);
  or add_168_21_g362(add_168_21_n_73 ,add_168_21_n_28 ,add_168_21_n_71);
  xnor add_168_21_g363(n_349 ,add_168_21_n_70 ,add_168_21_n_47);
  and add_168_21_g364(add_168_21_n_71 ,add_168_21_n_11 ,add_168_21_n_70);
  or add_168_21_g365(add_168_21_n_70 ,add_168_21_n_17 ,add_168_21_n_68);
  xnor add_168_21_g366(n_348 ,add_168_21_n_67 ,add_168_21_n_46);
  and add_168_21_g367(add_168_21_n_68 ,add_168_21_n_25 ,add_168_21_n_67);
  or add_168_21_g368(add_168_21_n_67 ,add_168_21_n_6 ,add_168_21_n_65);
  xnor add_168_21_g369(n_347 ,add_168_21_n_64 ,add_168_21_n_45);
  and add_168_21_g370(add_168_21_n_65 ,add_168_21_n_18 ,add_168_21_n_64);
  or add_168_21_g371(add_168_21_n_64 ,add_168_21_n_3 ,add_168_21_n_62);
  xnor add_168_21_g372(n_346 ,add_168_21_n_61 ,add_168_21_n_44);
  and add_168_21_g373(add_168_21_n_62 ,add_168_21_n_30 ,add_168_21_n_61);
  or add_168_21_g374(add_168_21_n_61 ,add_168_21_n_31 ,add_168_21_n_59);
  xnor add_168_21_g375(n_345 ,add_168_21_n_58 ,add_168_21_n_43);
  and add_168_21_g376(add_168_21_n_59 ,add_168_21_n_26 ,add_168_21_n_58);
  or add_168_21_g377(add_168_21_n_58 ,add_168_21_n_27 ,add_168_21_n_56);
  xnor add_168_21_g378(n_344 ,add_168_21_n_55 ,add_168_21_n_34);
  and add_168_21_g379(add_168_21_n_56 ,add_168_21_n_7 ,add_168_21_n_55);
  or add_168_21_g380(add_168_21_n_55 ,add_168_21_n_5 ,add_168_21_n_53);
  xnor add_168_21_g381(n_343 ,add_168_21_n_51 ,add_168_21_n_41);
  and add_168_21_g382(add_168_21_n_53 ,add_168_21_n_23 ,add_168_21_n_51);
  xor add_168_21_g383(n_342 ,add_168_21_n_33 ,add_168_21_n_40);
  or add_168_21_g384(add_168_21_n_51 ,add_168_21_n_4 ,add_168_21_n_49);
  and add_168_21_g385(n_341 ,add_168_21_n_33 ,add_168_21_n_13);
  nor add_168_21_g386(add_168_21_n_49 ,add_168_21_n_33 ,add_168_21_n_14);
  xnor add_168_21_g387(add_168_21_n_48 ,in41[9] ,in42[9]);
  xnor add_168_21_g388(add_168_21_n_47 ,in41[8] ,in42[8]);
  xnor add_168_21_g389(add_168_21_n_46 ,in41[7] ,in42[7]);
  xnor add_168_21_g390(add_168_21_n_45 ,in41[6] ,in42[6]);
  xnor add_168_21_g391(add_168_21_n_44 ,in41[5] ,in42[5]);
  xnor add_168_21_g392(add_168_21_n_43 ,in41[4] ,in42[4]);
  xnor add_168_21_g393(add_168_21_n_42 ,in41[10] ,in42[10]);
  xnor add_168_21_g394(add_168_21_n_41 ,in41[2] ,in42[2]);
  xnor add_168_21_g395(add_168_21_n_40 ,in41[1] ,in42[1]);
  xnor add_168_21_g396(add_168_21_n_39 ,in41[15] ,in42[15]);
  xnor add_168_21_g397(add_168_21_n_38 ,in41[14] ,in42[14]);
  xnor add_168_21_g398(add_168_21_n_37 ,in41[13] ,in42[13]);
  xnor add_168_21_g399(add_168_21_n_36 ,in41[12] ,in42[12]);
  xnor add_168_21_g400(add_168_21_n_35 ,in41[11] ,in42[11]);
  xnor add_168_21_g401(add_168_21_n_34 ,in41[3] ,in42[3]);
  and add_168_21_g402(add_168_21_n_32 ,in41[10] ,in42[10]);
  and add_168_21_g403(add_168_21_n_31 ,in41[4] ,in42[4]);
  or add_168_21_g404(add_168_21_n_30 ,in41[5] ,in42[5]);
  and add_168_21_g405(add_168_21_n_29 ,in41[15] ,in42[15]);
  and add_168_21_g406(add_168_21_n_28 ,in41[8] ,in42[8]);
  and add_168_21_g407(add_168_21_n_27 ,in41[3] ,in42[3]);
  or add_168_21_g408(add_168_21_n_26 ,in41[4] ,in42[4]);
  or add_168_21_g409(add_168_21_n_25 ,in41[7] ,in42[7]);
  and add_168_21_g410(add_168_21_n_24 ,in41[14] ,in42[14]);
  or add_168_21_g411(add_168_21_n_23 ,in41[2] ,in42[2]);
  or add_168_21_g412(add_168_21_n_22 ,in41[11] ,in42[11]);
  and add_168_21_g413(add_168_21_n_21 ,in41[9] ,in42[9]);
  and add_168_21_g414(add_168_21_n_20 ,in41[13] ,in42[13]);
  or add_168_21_g415(add_168_21_n_19 ,in41[9] ,in42[9]);
  or add_168_21_g416(add_168_21_n_18 ,in41[6] ,in42[6]);
  or add_168_21_g417(add_168_21_n_33 ,add_168_21_n_1 ,add_168_21_n_0);
  and add_168_21_g418(add_168_21_n_17 ,in41[7] ,in42[7]);
  or add_168_21_g419(add_168_21_n_16 ,in41[13] ,in42[13]);
  nor add_168_21_g420(add_168_21_n_15 ,in41[15] ,in42[15]);
  nor add_168_21_g421(add_168_21_n_14 ,in41[1] ,in42[1]);
  or add_168_21_g422(add_168_21_n_13 ,in41[0] ,in42[0]);
  or add_168_21_g423(add_168_21_n_12 ,in41[12] ,in42[12]);
  or add_168_21_g424(add_168_21_n_11 ,in41[8] ,in42[8]);
  and add_168_21_g425(add_168_21_n_10 ,in41[12] ,in42[12]);
  or add_168_21_g426(add_168_21_n_9 ,in41[14] ,in42[14]);
  and add_168_21_g427(add_168_21_n_8 ,in41[11] ,in42[11]);
  or add_168_21_g428(add_168_21_n_7 ,in41[3] ,in42[3]);
  and add_168_21_g429(add_168_21_n_6 ,in41[6] ,in42[6]);
  and add_168_21_g430(add_168_21_n_5 ,in41[2] ,in42[2]);
  and add_168_21_g431(add_168_21_n_4 ,in41[1] ,in42[1]);
  and add_168_21_g432(add_168_21_n_3 ,in41[5] ,in42[5]);
  or add_168_21_g433(add_168_21_n_2 ,in41[10] ,in42[10]);
  not add_168_21_g434(add_168_21_n_1 ,in41[0]);
  not add_168_21_g435(add_168_21_n_0 ,in42[0]);
  or add_170_21_g341(n_374 ,add_170_21_n_29 ,add_170_21_n_92);
  xnor add_170_21_g342(n_373 ,add_170_21_n_91 ,add_170_21_n_39);
  nor add_170_21_g343(add_170_21_n_92 ,add_170_21_n_15 ,add_170_21_n_91);
  or add_170_21_g344(add_170_21_n_91 ,add_170_21_n_24 ,add_170_21_n_89);
  xnor add_170_21_g345(n_372 ,add_170_21_n_88 ,add_170_21_n_38);
  and add_170_21_g346(add_170_21_n_89 ,add_170_21_n_9 ,add_170_21_n_88);
  or add_170_21_g347(add_170_21_n_88 ,add_170_21_n_20 ,add_170_21_n_86);
  xnor add_170_21_g348(n_371 ,add_170_21_n_85 ,add_170_21_n_37);
  and add_170_21_g349(add_170_21_n_86 ,add_170_21_n_16 ,add_170_21_n_85);
  or add_170_21_g350(add_170_21_n_85 ,add_170_21_n_10 ,add_170_21_n_83);
  xnor add_170_21_g351(n_370 ,add_170_21_n_82 ,add_170_21_n_36);
  and add_170_21_g352(add_170_21_n_83 ,add_170_21_n_12 ,add_170_21_n_82);
  or add_170_21_g353(add_170_21_n_82 ,add_170_21_n_8 ,add_170_21_n_80);
  xnor add_170_21_g354(n_369 ,add_170_21_n_79 ,add_170_21_n_35);
  and add_170_21_g355(add_170_21_n_80 ,add_170_21_n_22 ,add_170_21_n_79);
  or add_170_21_g356(add_170_21_n_79 ,add_170_21_n_32 ,add_170_21_n_77);
  xnor add_170_21_g357(n_368 ,add_170_21_n_76 ,add_170_21_n_42);
  and add_170_21_g358(add_170_21_n_77 ,add_170_21_n_2 ,add_170_21_n_76);
  or add_170_21_g359(add_170_21_n_76 ,add_170_21_n_21 ,add_170_21_n_74);
  xnor add_170_21_g360(n_367 ,add_170_21_n_73 ,add_170_21_n_48);
  and add_170_21_g361(add_170_21_n_74 ,add_170_21_n_19 ,add_170_21_n_73);
  or add_170_21_g362(add_170_21_n_73 ,add_170_21_n_28 ,add_170_21_n_71);
  xnor add_170_21_g363(n_366 ,add_170_21_n_70 ,add_170_21_n_47);
  and add_170_21_g364(add_170_21_n_71 ,add_170_21_n_11 ,add_170_21_n_70);
  or add_170_21_g365(add_170_21_n_70 ,add_170_21_n_17 ,add_170_21_n_68);
  xnor add_170_21_g366(n_365 ,add_170_21_n_67 ,add_170_21_n_46);
  and add_170_21_g367(add_170_21_n_68 ,add_170_21_n_25 ,add_170_21_n_67);
  or add_170_21_g368(add_170_21_n_67 ,add_170_21_n_6 ,add_170_21_n_65);
  xnor add_170_21_g369(n_364 ,add_170_21_n_64 ,add_170_21_n_45);
  and add_170_21_g370(add_170_21_n_65 ,add_170_21_n_18 ,add_170_21_n_64);
  or add_170_21_g371(add_170_21_n_64 ,add_170_21_n_3 ,add_170_21_n_62);
  xnor add_170_21_g372(n_363 ,add_170_21_n_61 ,add_170_21_n_44);
  and add_170_21_g373(add_170_21_n_62 ,add_170_21_n_30 ,add_170_21_n_61);
  or add_170_21_g374(add_170_21_n_61 ,add_170_21_n_31 ,add_170_21_n_59);
  xnor add_170_21_g375(n_362 ,add_170_21_n_58 ,add_170_21_n_43);
  and add_170_21_g376(add_170_21_n_59 ,add_170_21_n_26 ,add_170_21_n_58);
  or add_170_21_g377(add_170_21_n_58 ,add_170_21_n_27 ,add_170_21_n_56);
  xnor add_170_21_g378(n_361 ,add_170_21_n_55 ,add_170_21_n_34);
  and add_170_21_g379(add_170_21_n_56 ,add_170_21_n_7 ,add_170_21_n_55);
  or add_170_21_g380(add_170_21_n_55 ,add_170_21_n_5 ,add_170_21_n_53);
  xnor add_170_21_g381(n_360 ,add_170_21_n_51 ,add_170_21_n_41);
  and add_170_21_g382(add_170_21_n_53 ,add_170_21_n_23 ,add_170_21_n_51);
  xor add_170_21_g383(n_359 ,add_170_21_n_33 ,add_170_21_n_40);
  or add_170_21_g384(add_170_21_n_51 ,add_170_21_n_4 ,add_170_21_n_49);
  and add_170_21_g385(n_358 ,add_170_21_n_33 ,add_170_21_n_13);
  nor add_170_21_g386(add_170_21_n_49 ,add_170_21_n_33 ,add_170_21_n_14);
  xnor add_170_21_g387(add_170_21_n_48 ,in43[9] ,in44[9]);
  xnor add_170_21_g388(add_170_21_n_47 ,in43[8] ,in44[8]);
  xnor add_170_21_g389(add_170_21_n_46 ,in43[7] ,in44[7]);
  xnor add_170_21_g390(add_170_21_n_45 ,in43[6] ,in44[6]);
  xnor add_170_21_g391(add_170_21_n_44 ,in43[5] ,in44[5]);
  xnor add_170_21_g392(add_170_21_n_43 ,in43[4] ,in44[4]);
  xnor add_170_21_g393(add_170_21_n_42 ,in43[10] ,in44[10]);
  xnor add_170_21_g394(add_170_21_n_41 ,in43[2] ,in44[2]);
  xnor add_170_21_g395(add_170_21_n_40 ,in43[1] ,in44[1]);
  xnor add_170_21_g396(add_170_21_n_39 ,in43[15] ,in44[15]);
  xnor add_170_21_g397(add_170_21_n_38 ,in43[14] ,in44[14]);
  xnor add_170_21_g398(add_170_21_n_37 ,in43[13] ,in44[13]);
  xnor add_170_21_g399(add_170_21_n_36 ,in43[12] ,in44[12]);
  xnor add_170_21_g400(add_170_21_n_35 ,in43[11] ,in44[11]);
  xnor add_170_21_g401(add_170_21_n_34 ,in43[3] ,in44[3]);
  and add_170_21_g402(add_170_21_n_32 ,in43[10] ,in44[10]);
  and add_170_21_g403(add_170_21_n_31 ,in43[4] ,in44[4]);
  or add_170_21_g404(add_170_21_n_30 ,in43[5] ,in44[5]);
  and add_170_21_g405(add_170_21_n_29 ,in43[15] ,in44[15]);
  and add_170_21_g406(add_170_21_n_28 ,in43[8] ,in44[8]);
  and add_170_21_g407(add_170_21_n_27 ,in43[3] ,in44[3]);
  or add_170_21_g408(add_170_21_n_26 ,in43[4] ,in44[4]);
  or add_170_21_g409(add_170_21_n_25 ,in43[7] ,in44[7]);
  and add_170_21_g410(add_170_21_n_24 ,in43[14] ,in44[14]);
  or add_170_21_g411(add_170_21_n_23 ,in43[2] ,in44[2]);
  or add_170_21_g412(add_170_21_n_22 ,in43[11] ,in44[11]);
  and add_170_21_g413(add_170_21_n_21 ,in43[9] ,in44[9]);
  and add_170_21_g414(add_170_21_n_20 ,in43[13] ,in44[13]);
  or add_170_21_g415(add_170_21_n_19 ,in43[9] ,in44[9]);
  or add_170_21_g416(add_170_21_n_18 ,in43[6] ,in44[6]);
  or add_170_21_g417(add_170_21_n_33 ,add_170_21_n_1 ,add_170_21_n_0);
  and add_170_21_g418(add_170_21_n_17 ,in43[7] ,in44[7]);
  or add_170_21_g419(add_170_21_n_16 ,in43[13] ,in44[13]);
  nor add_170_21_g420(add_170_21_n_15 ,in43[15] ,in44[15]);
  nor add_170_21_g421(add_170_21_n_14 ,in43[1] ,in44[1]);
  or add_170_21_g422(add_170_21_n_13 ,in43[0] ,in44[0]);
  or add_170_21_g423(add_170_21_n_12 ,in43[12] ,in44[12]);
  or add_170_21_g424(add_170_21_n_11 ,in43[8] ,in44[8]);
  and add_170_21_g425(add_170_21_n_10 ,in43[12] ,in44[12]);
  or add_170_21_g426(add_170_21_n_9 ,in43[14] ,in44[14]);
  and add_170_21_g427(add_170_21_n_8 ,in43[11] ,in44[11]);
  or add_170_21_g428(add_170_21_n_7 ,in43[3] ,in44[3]);
  and add_170_21_g429(add_170_21_n_6 ,in43[6] ,in44[6]);
  and add_170_21_g430(add_170_21_n_5 ,in43[2] ,in44[2]);
  and add_170_21_g431(add_170_21_n_4 ,in43[1] ,in44[1]);
  and add_170_21_g432(add_170_21_n_3 ,in43[5] ,in44[5]);
  or add_170_21_g433(add_170_21_n_2 ,in43[10] ,in44[10]);
  not add_170_21_g434(add_170_21_n_1 ,in43[0]);
  not add_170_21_g435(add_170_21_n_0 ,in44[0]);
  or add_172_21_g341(n_391 ,add_172_21_n_29 ,add_172_21_n_92);
  xnor add_172_21_g342(n_390 ,add_172_21_n_91 ,add_172_21_n_39);
  nor add_172_21_g343(add_172_21_n_92 ,add_172_21_n_15 ,add_172_21_n_91);
  or add_172_21_g344(add_172_21_n_91 ,add_172_21_n_24 ,add_172_21_n_89);
  xnor add_172_21_g345(n_389 ,add_172_21_n_88 ,add_172_21_n_38);
  and add_172_21_g346(add_172_21_n_89 ,add_172_21_n_9 ,add_172_21_n_88);
  or add_172_21_g347(add_172_21_n_88 ,add_172_21_n_20 ,add_172_21_n_86);
  xnor add_172_21_g348(n_388 ,add_172_21_n_85 ,add_172_21_n_37);
  and add_172_21_g349(add_172_21_n_86 ,add_172_21_n_16 ,add_172_21_n_85);
  or add_172_21_g350(add_172_21_n_85 ,add_172_21_n_10 ,add_172_21_n_83);
  xnor add_172_21_g351(n_387 ,add_172_21_n_82 ,add_172_21_n_36);
  and add_172_21_g352(add_172_21_n_83 ,add_172_21_n_12 ,add_172_21_n_82);
  or add_172_21_g353(add_172_21_n_82 ,add_172_21_n_8 ,add_172_21_n_80);
  xnor add_172_21_g354(n_386 ,add_172_21_n_79 ,add_172_21_n_35);
  and add_172_21_g355(add_172_21_n_80 ,add_172_21_n_22 ,add_172_21_n_79);
  or add_172_21_g356(add_172_21_n_79 ,add_172_21_n_32 ,add_172_21_n_77);
  xnor add_172_21_g357(n_385 ,add_172_21_n_76 ,add_172_21_n_42);
  and add_172_21_g358(add_172_21_n_77 ,add_172_21_n_2 ,add_172_21_n_76);
  or add_172_21_g359(add_172_21_n_76 ,add_172_21_n_21 ,add_172_21_n_74);
  xnor add_172_21_g360(n_384 ,add_172_21_n_73 ,add_172_21_n_48);
  and add_172_21_g361(add_172_21_n_74 ,add_172_21_n_19 ,add_172_21_n_73);
  or add_172_21_g362(add_172_21_n_73 ,add_172_21_n_28 ,add_172_21_n_71);
  xnor add_172_21_g363(n_383 ,add_172_21_n_70 ,add_172_21_n_47);
  and add_172_21_g364(add_172_21_n_71 ,add_172_21_n_11 ,add_172_21_n_70);
  or add_172_21_g365(add_172_21_n_70 ,add_172_21_n_17 ,add_172_21_n_68);
  xnor add_172_21_g366(n_382 ,add_172_21_n_67 ,add_172_21_n_46);
  and add_172_21_g367(add_172_21_n_68 ,add_172_21_n_25 ,add_172_21_n_67);
  or add_172_21_g368(add_172_21_n_67 ,add_172_21_n_6 ,add_172_21_n_65);
  xnor add_172_21_g369(n_381 ,add_172_21_n_64 ,add_172_21_n_45);
  and add_172_21_g370(add_172_21_n_65 ,add_172_21_n_18 ,add_172_21_n_64);
  or add_172_21_g371(add_172_21_n_64 ,add_172_21_n_3 ,add_172_21_n_62);
  xnor add_172_21_g372(n_380 ,add_172_21_n_61 ,add_172_21_n_44);
  and add_172_21_g373(add_172_21_n_62 ,add_172_21_n_30 ,add_172_21_n_61);
  or add_172_21_g374(add_172_21_n_61 ,add_172_21_n_31 ,add_172_21_n_59);
  xnor add_172_21_g375(n_379 ,add_172_21_n_58 ,add_172_21_n_43);
  and add_172_21_g376(add_172_21_n_59 ,add_172_21_n_26 ,add_172_21_n_58);
  or add_172_21_g377(add_172_21_n_58 ,add_172_21_n_27 ,add_172_21_n_56);
  xnor add_172_21_g378(n_378 ,add_172_21_n_55 ,add_172_21_n_34);
  and add_172_21_g379(add_172_21_n_56 ,add_172_21_n_7 ,add_172_21_n_55);
  or add_172_21_g380(add_172_21_n_55 ,add_172_21_n_5 ,add_172_21_n_53);
  xnor add_172_21_g381(n_377 ,add_172_21_n_51 ,add_172_21_n_41);
  and add_172_21_g382(add_172_21_n_53 ,add_172_21_n_23 ,add_172_21_n_51);
  xor add_172_21_g383(n_376 ,add_172_21_n_33 ,add_172_21_n_40);
  or add_172_21_g384(add_172_21_n_51 ,add_172_21_n_4 ,add_172_21_n_49);
  and add_172_21_g385(n_375 ,add_172_21_n_33 ,add_172_21_n_13);
  nor add_172_21_g386(add_172_21_n_49 ,add_172_21_n_33 ,add_172_21_n_14);
  xnor add_172_21_g387(add_172_21_n_48 ,in45[9] ,in46[9]);
  xnor add_172_21_g388(add_172_21_n_47 ,in45[8] ,in46[8]);
  xnor add_172_21_g389(add_172_21_n_46 ,in45[7] ,in46[7]);
  xnor add_172_21_g390(add_172_21_n_45 ,in45[6] ,in46[6]);
  xnor add_172_21_g391(add_172_21_n_44 ,in45[5] ,in46[5]);
  xnor add_172_21_g392(add_172_21_n_43 ,in45[4] ,in46[4]);
  xnor add_172_21_g393(add_172_21_n_42 ,in45[10] ,in46[10]);
  xnor add_172_21_g394(add_172_21_n_41 ,in45[2] ,in46[2]);
  xnor add_172_21_g395(add_172_21_n_40 ,in45[1] ,in46[1]);
  xnor add_172_21_g396(add_172_21_n_39 ,in45[15] ,in46[15]);
  xnor add_172_21_g397(add_172_21_n_38 ,in45[14] ,in46[14]);
  xnor add_172_21_g398(add_172_21_n_37 ,in45[13] ,in46[13]);
  xnor add_172_21_g399(add_172_21_n_36 ,in45[12] ,in46[12]);
  xnor add_172_21_g400(add_172_21_n_35 ,in45[11] ,in46[11]);
  xnor add_172_21_g401(add_172_21_n_34 ,in45[3] ,in46[3]);
  and add_172_21_g402(add_172_21_n_32 ,in45[10] ,in46[10]);
  and add_172_21_g403(add_172_21_n_31 ,in45[4] ,in46[4]);
  or add_172_21_g404(add_172_21_n_30 ,in45[5] ,in46[5]);
  and add_172_21_g405(add_172_21_n_29 ,in45[15] ,in46[15]);
  and add_172_21_g406(add_172_21_n_28 ,in45[8] ,in46[8]);
  and add_172_21_g407(add_172_21_n_27 ,in45[3] ,in46[3]);
  or add_172_21_g408(add_172_21_n_26 ,in45[4] ,in46[4]);
  or add_172_21_g409(add_172_21_n_25 ,in45[7] ,in46[7]);
  and add_172_21_g410(add_172_21_n_24 ,in45[14] ,in46[14]);
  or add_172_21_g411(add_172_21_n_23 ,in45[2] ,in46[2]);
  or add_172_21_g412(add_172_21_n_22 ,in45[11] ,in46[11]);
  and add_172_21_g413(add_172_21_n_21 ,in45[9] ,in46[9]);
  and add_172_21_g414(add_172_21_n_20 ,in45[13] ,in46[13]);
  or add_172_21_g415(add_172_21_n_19 ,in45[9] ,in46[9]);
  or add_172_21_g416(add_172_21_n_18 ,in45[6] ,in46[6]);
  or add_172_21_g417(add_172_21_n_33 ,add_172_21_n_1 ,add_172_21_n_0);
  and add_172_21_g418(add_172_21_n_17 ,in45[7] ,in46[7]);
  or add_172_21_g419(add_172_21_n_16 ,in45[13] ,in46[13]);
  nor add_172_21_g420(add_172_21_n_15 ,in45[15] ,in46[15]);
  nor add_172_21_g421(add_172_21_n_14 ,in45[1] ,in46[1]);
  or add_172_21_g422(add_172_21_n_13 ,in45[0] ,in46[0]);
  or add_172_21_g423(add_172_21_n_12 ,in45[12] ,in46[12]);
  or add_172_21_g424(add_172_21_n_11 ,in45[8] ,in46[8]);
  and add_172_21_g425(add_172_21_n_10 ,in45[12] ,in46[12]);
  or add_172_21_g426(add_172_21_n_9 ,in45[14] ,in46[14]);
  and add_172_21_g427(add_172_21_n_8 ,in45[11] ,in46[11]);
  or add_172_21_g428(add_172_21_n_7 ,in45[3] ,in46[3]);
  and add_172_21_g429(add_172_21_n_6 ,in45[6] ,in46[6]);
  and add_172_21_g430(add_172_21_n_5 ,in45[2] ,in46[2]);
  and add_172_21_g431(add_172_21_n_4 ,in45[1] ,in46[1]);
  and add_172_21_g432(add_172_21_n_3 ,in45[5] ,in46[5]);
  or add_172_21_g433(add_172_21_n_2 ,in45[10] ,in46[10]);
  not add_172_21_g434(add_172_21_n_1 ,in45[0]);
  not add_172_21_g435(add_172_21_n_0 ,in46[0]);
  or add_174_21_g341(n_408 ,add_174_21_n_29 ,add_174_21_n_92);
  xnor add_174_21_g342(n_407 ,add_174_21_n_91 ,add_174_21_n_39);
  nor add_174_21_g343(add_174_21_n_92 ,add_174_21_n_15 ,add_174_21_n_91);
  or add_174_21_g344(add_174_21_n_91 ,add_174_21_n_24 ,add_174_21_n_89);
  xnor add_174_21_g345(n_406 ,add_174_21_n_88 ,add_174_21_n_38);
  and add_174_21_g346(add_174_21_n_89 ,add_174_21_n_9 ,add_174_21_n_88);
  or add_174_21_g347(add_174_21_n_88 ,add_174_21_n_20 ,add_174_21_n_86);
  xnor add_174_21_g348(n_405 ,add_174_21_n_85 ,add_174_21_n_37);
  and add_174_21_g349(add_174_21_n_86 ,add_174_21_n_16 ,add_174_21_n_85);
  or add_174_21_g350(add_174_21_n_85 ,add_174_21_n_10 ,add_174_21_n_83);
  xnor add_174_21_g351(n_404 ,add_174_21_n_82 ,add_174_21_n_36);
  and add_174_21_g352(add_174_21_n_83 ,add_174_21_n_12 ,add_174_21_n_82);
  or add_174_21_g353(add_174_21_n_82 ,add_174_21_n_8 ,add_174_21_n_80);
  xnor add_174_21_g354(n_403 ,add_174_21_n_79 ,add_174_21_n_35);
  and add_174_21_g355(add_174_21_n_80 ,add_174_21_n_22 ,add_174_21_n_79);
  or add_174_21_g356(add_174_21_n_79 ,add_174_21_n_32 ,add_174_21_n_77);
  xnor add_174_21_g357(n_402 ,add_174_21_n_76 ,add_174_21_n_42);
  and add_174_21_g358(add_174_21_n_77 ,add_174_21_n_2 ,add_174_21_n_76);
  or add_174_21_g359(add_174_21_n_76 ,add_174_21_n_21 ,add_174_21_n_74);
  xnor add_174_21_g360(n_401 ,add_174_21_n_73 ,add_174_21_n_48);
  and add_174_21_g361(add_174_21_n_74 ,add_174_21_n_19 ,add_174_21_n_73);
  or add_174_21_g362(add_174_21_n_73 ,add_174_21_n_28 ,add_174_21_n_71);
  xnor add_174_21_g363(n_400 ,add_174_21_n_70 ,add_174_21_n_47);
  and add_174_21_g364(add_174_21_n_71 ,add_174_21_n_11 ,add_174_21_n_70);
  or add_174_21_g365(add_174_21_n_70 ,add_174_21_n_17 ,add_174_21_n_68);
  xnor add_174_21_g366(n_399 ,add_174_21_n_67 ,add_174_21_n_46);
  and add_174_21_g367(add_174_21_n_68 ,add_174_21_n_25 ,add_174_21_n_67);
  or add_174_21_g368(add_174_21_n_67 ,add_174_21_n_6 ,add_174_21_n_65);
  xnor add_174_21_g369(n_398 ,add_174_21_n_64 ,add_174_21_n_45);
  and add_174_21_g370(add_174_21_n_65 ,add_174_21_n_18 ,add_174_21_n_64);
  or add_174_21_g371(add_174_21_n_64 ,add_174_21_n_3 ,add_174_21_n_62);
  xnor add_174_21_g372(n_397 ,add_174_21_n_61 ,add_174_21_n_44);
  and add_174_21_g373(add_174_21_n_62 ,add_174_21_n_30 ,add_174_21_n_61);
  or add_174_21_g374(add_174_21_n_61 ,add_174_21_n_31 ,add_174_21_n_59);
  xnor add_174_21_g375(n_396 ,add_174_21_n_58 ,add_174_21_n_43);
  and add_174_21_g376(add_174_21_n_59 ,add_174_21_n_26 ,add_174_21_n_58);
  or add_174_21_g377(add_174_21_n_58 ,add_174_21_n_27 ,add_174_21_n_56);
  xnor add_174_21_g378(n_395 ,add_174_21_n_55 ,add_174_21_n_34);
  and add_174_21_g379(add_174_21_n_56 ,add_174_21_n_7 ,add_174_21_n_55);
  or add_174_21_g380(add_174_21_n_55 ,add_174_21_n_5 ,add_174_21_n_53);
  xnor add_174_21_g381(n_394 ,add_174_21_n_51 ,add_174_21_n_41);
  and add_174_21_g382(add_174_21_n_53 ,add_174_21_n_23 ,add_174_21_n_51);
  xor add_174_21_g383(n_393 ,add_174_21_n_33 ,add_174_21_n_40);
  or add_174_21_g384(add_174_21_n_51 ,add_174_21_n_4 ,add_174_21_n_49);
  and add_174_21_g385(n_392 ,add_174_21_n_33 ,add_174_21_n_13);
  nor add_174_21_g386(add_174_21_n_49 ,add_174_21_n_33 ,add_174_21_n_14);
  xnor add_174_21_g387(add_174_21_n_48 ,in47[9] ,in48[9]);
  xnor add_174_21_g388(add_174_21_n_47 ,in47[8] ,in48[8]);
  xnor add_174_21_g389(add_174_21_n_46 ,in47[7] ,in48[7]);
  xnor add_174_21_g390(add_174_21_n_45 ,in47[6] ,in48[6]);
  xnor add_174_21_g391(add_174_21_n_44 ,in47[5] ,in48[5]);
  xnor add_174_21_g392(add_174_21_n_43 ,in47[4] ,in48[4]);
  xnor add_174_21_g393(add_174_21_n_42 ,in47[10] ,in48[10]);
  xnor add_174_21_g394(add_174_21_n_41 ,in47[2] ,in48[2]);
  xnor add_174_21_g395(add_174_21_n_40 ,in47[1] ,in48[1]);
  xnor add_174_21_g396(add_174_21_n_39 ,in47[15] ,in48[15]);
  xnor add_174_21_g397(add_174_21_n_38 ,in47[14] ,in48[14]);
  xnor add_174_21_g398(add_174_21_n_37 ,in47[13] ,in48[13]);
  xnor add_174_21_g399(add_174_21_n_36 ,in47[12] ,in48[12]);
  xnor add_174_21_g400(add_174_21_n_35 ,in47[11] ,in48[11]);
  xnor add_174_21_g401(add_174_21_n_34 ,in47[3] ,in48[3]);
  and add_174_21_g402(add_174_21_n_32 ,in47[10] ,in48[10]);
  and add_174_21_g403(add_174_21_n_31 ,in47[4] ,in48[4]);
  or add_174_21_g404(add_174_21_n_30 ,in47[5] ,in48[5]);
  and add_174_21_g405(add_174_21_n_29 ,in47[15] ,in48[15]);
  and add_174_21_g406(add_174_21_n_28 ,in47[8] ,in48[8]);
  and add_174_21_g407(add_174_21_n_27 ,in47[3] ,in48[3]);
  or add_174_21_g408(add_174_21_n_26 ,in47[4] ,in48[4]);
  or add_174_21_g409(add_174_21_n_25 ,in47[7] ,in48[7]);
  and add_174_21_g410(add_174_21_n_24 ,in47[14] ,in48[14]);
  or add_174_21_g411(add_174_21_n_23 ,in47[2] ,in48[2]);
  or add_174_21_g412(add_174_21_n_22 ,in47[11] ,in48[11]);
  and add_174_21_g413(add_174_21_n_21 ,in47[9] ,in48[9]);
  and add_174_21_g414(add_174_21_n_20 ,in47[13] ,in48[13]);
  or add_174_21_g415(add_174_21_n_19 ,in47[9] ,in48[9]);
  or add_174_21_g416(add_174_21_n_18 ,in47[6] ,in48[6]);
  or add_174_21_g417(add_174_21_n_33 ,add_174_21_n_1 ,add_174_21_n_0);
  and add_174_21_g418(add_174_21_n_17 ,in47[7] ,in48[7]);
  or add_174_21_g419(add_174_21_n_16 ,in47[13] ,in48[13]);
  nor add_174_21_g420(add_174_21_n_15 ,in47[15] ,in48[15]);
  nor add_174_21_g421(add_174_21_n_14 ,in47[1] ,in48[1]);
  or add_174_21_g422(add_174_21_n_13 ,in47[0] ,in48[0]);
  or add_174_21_g423(add_174_21_n_12 ,in47[12] ,in48[12]);
  or add_174_21_g424(add_174_21_n_11 ,in47[8] ,in48[8]);
  and add_174_21_g425(add_174_21_n_10 ,in47[12] ,in48[12]);
  or add_174_21_g426(add_174_21_n_9 ,in47[14] ,in48[14]);
  and add_174_21_g427(add_174_21_n_8 ,in47[11] ,in48[11]);
  or add_174_21_g428(add_174_21_n_7 ,in47[3] ,in48[3]);
  and add_174_21_g429(add_174_21_n_6 ,in47[6] ,in48[6]);
  and add_174_21_g430(add_174_21_n_5 ,in47[2] ,in48[2]);
  and add_174_21_g431(add_174_21_n_4 ,in47[1] ,in48[1]);
  and add_174_21_g432(add_174_21_n_3 ,in47[5] ,in48[5]);
  or add_174_21_g433(add_174_21_n_2 ,in47[10] ,in48[10]);
  not add_174_21_g434(add_174_21_n_1 ,in47[0]);
  not add_174_21_g435(add_174_21_n_0 ,in48[0]);
  or add_176_21_g341(n_425 ,add_176_21_n_29 ,add_176_21_n_92);
  xnor add_176_21_g342(n_424 ,add_176_21_n_91 ,add_176_21_n_39);
  nor add_176_21_g343(add_176_21_n_92 ,add_176_21_n_15 ,add_176_21_n_91);
  or add_176_21_g344(add_176_21_n_91 ,add_176_21_n_24 ,add_176_21_n_89);
  xnor add_176_21_g345(n_423 ,add_176_21_n_88 ,add_176_21_n_38);
  and add_176_21_g346(add_176_21_n_89 ,add_176_21_n_9 ,add_176_21_n_88);
  or add_176_21_g347(add_176_21_n_88 ,add_176_21_n_20 ,add_176_21_n_86);
  xnor add_176_21_g348(n_422 ,add_176_21_n_85 ,add_176_21_n_37);
  and add_176_21_g349(add_176_21_n_86 ,add_176_21_n_16 ,add_176_21_n_85);
  or add_176_21_g350(add_176_21_n_85 ,add_176_21_n_10 ,add_176_21_n_83);
  xnor add_176_21_g351(n_421 ,add_176_21_n_82 ,add_176_21_n_36);
  and add_176_21_g352(add_176_21_n_83 ,add_176_21_n_12 ,add_176_21_n_82);
  or add_176_21_g353(add_176_21_n_82 ,add_176_21_n_8 ,add_176_21_n_80);
  xnor add_176_21_g354(n_420 ,add_176_21_n_79 ,add_176_21_n_35);
  and add_176_21_g355(add_176_21_n_80 ,add_176_21_n_22 ,add_176_21_n_79);
  or add_176_21_g356(add_176_21_n_79 ,add_176_21_n_32 ,add_176_21_n_77);
  xnor add_176_21_g357(n_419 ,add_176_21_n_76 ,add_176_21_n_42);
  and add_176_21_g358(add_176_21_n_77 ,add_176_21_n_2 ,add_176_21_n_76);
  or add_176_21_g359(add_176_21_n_76 ,add_176_21_n_21 ,add_176_21_n_74);
  xnor add_176_21_g360(n_418 ,add_176_21_n_73 ,add_176_21_n_48);
  and add_176_21_g361(add_176_21_n_74 ,add_176_21_n_19 ,add_176_21_n_73);
  or add_176_21_g362(add_176_21_n_73 ,add_176_21_n_28 ,add_176_21_n_71);
  xnor add_176_21_g363(n_417 ,add_176_21_n_70 ,add_176_21_n_47);
  and add_176_21_g364(add_176_21_n_71 ,add_176_21_n_11 ,add_176_21_n_70);
  or add_176_21_g365(add_176_21_n_70 ,add_176_21_n_17 ,add_176_21_n_68);
  xnor add_176_21_g366(n_416 ,add_176_21_n_67 ,add_176_21_n_46);
  and add_176_21_g367(add_176_21_n_68 ,add_176_21_n_25 ,add_176_21_n_67);
  or add_176_21_g368(add_176_21_n_67 ,add_176_21_n_6 ,add_176_21_n_65);
  xnor add_176_21_g369(n_415 ,add_176_21_n_64 ,add_176_21_n_45);
  and add_176_21_g370(add_176_21_n_65 ,add_176_21_n_18 ,add_176_21_n_64);
  or add_176_21_g371(add_176_21_n_64 ,add_176_21_n_3 ,add_176_21_n_62);
  xnor add_176_21_g372(n_414 ,add_176_21_n_61 ,add_176_21_n_44);
  and add_176_21_g373(add_176_21_n_62 ,add_176_21_n_30 ,add_176_21_n_61);
  or add_176_21_g374(add_176_21_n_61 ,add_176_21_n_31 ,add_176_21_n_59);
  xnor add_176_21_g375(n_413 ,add_176_21_n_58 ,add_176_21_n_43);
  and add_176_21_g376(add_176_21_n_59 ,add_176_21_n_26 ,add_176_21_n_58);
  or add_176_21_g377(add_176_21_n_58 ,add_176_21_n_27 ,add_176_21_n_56);
  xnor add_176_21_g378(n_412 ,add_176_21_n_55 ,add_176_21_n_34);
  and add_176_21_g379(add_176_21_n_56 ,add_176_21_n_7 ,add_176_21_n_55);
  or add_176_21_g380(add_176_21_n_55 ,add_176_21_n_5 ,add_176_21_n_53);
  xnor add_176_21_g381(n_411 ,add_176_21_n_51 ,add_176_21_n_41);
  and add_176_21_g382(add_176_21_n_53 ,add_176_21_n_23 ,add_176_21_n_51);
  xor add_176_21_g383(n_410 ,add_176_21_n_33 ,add_176_21_n_40);
  or add_176_21_g384(add_176_21_n_51 ,add_176_21_n_4 ,add_176_21_n_49);
  and add_176_21_g385(n_409 ,add_176_21_n_33 ,add_176_21_n_13);
  nor add_176_21_g386(add_176_21_n_49 ,add_176_21_n_33 ,add_176_21_n_14);
  xnor add_176_21_g387(add_176_21_n_48 ,in49[9] ,in50[9]);
  xnor add_176_21_g388(add_176_21_n_47 ,in49[8] ,in50[8]);
  xnor add_176_21_g389(add_176_21_n_46 ,in49[7] ,in50[7]);
  xnor add_176_21_g390(add_176_21_n_45 ,in49[6] ,in50[6]);
  xnor add_176_21_g391(add_176_21_n_44 ,in49[5] ,in50[5]);
  xnor add_176_21_g392(add_176_21_n_43 ,in49[4] ,in50[4]);
  xnor add_176_21_g393(add_176_21_n_42 ,in49[10] ,in50[10]);
  xnor add_176_21_g394(add_176_21_n_41 ,in49[2] ,in50[2]);
  xnor add_176_21_g395(add_176_21_n_40 ,in49[1] ,in50[1]);
  xnor add_176_21_g396(add_176_21_n_39 ,in49[15] ,in50[15]);
  xnor add_176_21_g397(add_176_21_n_38 ,in49[14] ,in50[14]);
  xnor add_176_21_g398(add_176_21_n_37 ,in49[13] ,in50[13]);
  xnor add_176_21_g399(add_176_21_n_36 ,in49[12] ,in50[12]);
  xnor add_176_21_g400(add_176_21_n_35 ,in49[11] ,in50[11]);
  xnor add_176_21_g401(add_176_21_n_34 ,in49[3] ,in50[3]);
  and add_176_21_g402(add_176_21_n_32 ,in49[10] ,in50[10]);
  and add_176_21_g403(add_176_21_n_31 ,in49[4] ,in50[4]);
  or add_176_21_g404(add_176_21_n_30 ,in49[5] ,in50[5]);
  and add_176_21_g405(add_176_21_n_29 ,in49[15] ,in50[15]);
  and add_176_21_g406(add_176_21_n_28 ,in49[8] ,in50[8]);
  and add_176_21_g407(add_176_21_n_27 ,in49[3] ,in50[3]);
  or add_176_21_g408(add_176_21_n_26 ,in49[4] ,in50[4]);
  or add_176_21_g409(add_176_21_n_25 ,in49[7] ,in50[7]);
  and add_176_21_g410(add_176_21_n_24 ,in49[14] ,in50[14]);
  or add_176_21_g411(add_176_21_n_23 ,in49[2] ,in50[2]);
  or add_176_21_g412(add_176_21_n_22 ,in49[11] ,in50[11]);
  and add_176_21_g413(add_176_21_n_21 ,in49[9] ,in50[9]);
  and add_176_21_g414(add_176_21_n_20 ,in49[13] ,in50[13]);
  or add_176_21_g415(add_176_21_n_19 ,in49[9] ,in50[9]);
  or add_176_21_g416(add_176_21_n_18 ,in49[6] ,in50[6]);
  or add_176_21_g417(add_176_21_n_33 ,add_176_21_n_1 ,add_176_21_n_0);
  and add_176_21_g418(add_176_21_n_17 ,in49[7] ,in50[7]);
  or add_176_21_g419(add_176_21_n_16 ,in49[13] ,in50[13]);
  nor add_176_21_g420(add_176_21_n_15 ,in49[15] ,in50[15]);
  nor add_176_21_g421(add_176_21_n_14 ,in49[1] ,in50[1]);
  or add_176_21_g422(add_176_21_n_13 ,in49[0] ,in50[0]);
  or add_176_21_g423(add_176_21_n_12 ,in49[12] ,in50[12]);
  or add_176_21_g424(add_176_21_n_11 ,in49[8] ,in50[8]);
  and add_176_21_g425(add_176_21_n_10 ,in49[12] ,in50[12]);
  or add_176_21_g426(add_176_21_n_9 ,in49[14] ,in50[14]);
  and add_176_21_g427(add_176_21_n_8 ,in49[11] ,in50[11]);
  or add_176_21_g428(add_176_21_n_7 ,in49[3] ,in50[3]);
  and add_176_21_g429(add_176_21_n_6 ,in49[6] ,in50[6]);
  and add_176_21_g430(add_176_21_n_5 ,in49[2] ,in50[2]);
  and add_176_21_g431(add_176_21_n_4 ,in49[1] ,in50[1]);
  and add_176_21_g432(add_176_21_n_3 ,in49[5] ,in50[5]);
  or add_176_21_g433(add_176_21_n_2 ,in49[10] ,in50[10]);
  not add_176_21_g434(add_176_21_n_1 ,in49[0]);
  not add_176_21_g435(add_176_21_n_0 ,in50[0]);
  or add_178_21_g341(n_442 ,add_178_21_n_29 ,add_178_21_n_92);
  xnor add_178_21_g342(n_441 ,add_178_21_n_91 ,add_178_21_n_39);
  nor add_178_21_g343(add_178_21_n_92 ,add_178_21_n_15 ,add_178_21_n_91);
  or add_178_21_g344(add_178_21_n_91 ,add_178_21_n_24 ,add_178_21_n_89);
  xnor add_178_21_g345(n_440 ,add_178_21_n_88 ,add_178_21_n_38);
  and add_178_21_g346(add_178_21_n_89 ,add_178_21_n_9 ,add_178_21_n_88);
  or add_178_21_g347(add_178_21_n_88 ,add_178_21_n_20 ,add_178_21_n_86);
  xnor add_178_21_g348(n_439 ,add_178_21_n_85 ,add_178_21_n_37);
  and add_178_21_g349(add_178_21_n_86 ,add_178_21_n_16 ,add_178_21_n_85);
  or add_178_21_g350(add_178_21_n_85 ,add_178_21_n_10 ,add_178_21_n_83);
  xnor add_178_21_g351(n_438 ,add_178_21_n_82 ,add_178_21_n_36);
  and add_178_21_g352(add_178_21_n_83 ,add_178_21_n_12 ,add_178_21_n_82);
  or add_178_21_g353(add_178_21_n_82 ,add_178_21_n_8 ,add_178_21_n_80);
  xnor add_178_21_g354(n_437 ,add_178_21_n_79 ,add_178_21_n_35);
  and add_178_21_g355(add_178_21_n_80 ,add_178_21_n_22 ,add_178_21_n_79);
  or add_178_21_g356(add_178_21_n_79 ,add_178_21_n_32 ,add_178_21_n_77);
  xnor add_178_21_g357(n_436 ,add_178_21_n_76 ,add_178_21_n_42);
  and add_178_21_g358(add_178_21_n_77 ,add_178_21_n_2 ,add_178_21_n_76);
  or add_178_21_g359(add_178_21_n_76 ,add_178_21_n_21 ,add_178_21_n_74);
  xnor add_178_21_g360(n_435 ,add_178_21_n_73 ,add_178_21_n_48);
  and add_178_21_g361(add_178_21_n_74 ,add_178_21_n_19 ,add_178_21_n_73);
  or add_178_21_g362(add_178_21_n_73 ,add_178_21_n_28 ,add_178_21_n_71);
  xnor add_178_21_g363(n_434 ,add_178_21_n_70 ,add_178_21_n_47);
  and add_178_21_g364(add_178_21_n_71 ,add_178_21_n_11 ,add_178_21_n_70);
  or add_178_21_g365(add_178_21_n_70 ,add_178_21_n_17 ,add_178_21_n_68);
  xnor add_178_21_g366(n_433 ,add_178_21_n_67 ,add_178_21_n_46);
  and add_178_21_g367(add_178_21_n_68 ,add_178_21_n_25 ,add_178_21_n_67);
  or add_178_21_g368(add_178_21_n_67 ,add_178_21_n_6 ,add_178_21_n_65);
  xnor add_178_21_g369(n_432 ,add_178_21_n_64 ,add_178_21_n_45);
  and add_178_21_g370(add_178_21_n_65 ,add_178_21_n_18 ,add_178_21_n_64);
  or add_178_21_g371(add_178_21_n_64 ,add_178_21_n_3 ,add_178_21_n_62);
  xnor add_178_21_g372(n_431 ,add_178_21_n_61 ,add_178_21_n_44);
  and add_178_21_g373(add_178_21_n_62 ,add_178_21_n_30 ,add_178_21_n_61);
  or add_178_21_g374(add_178_21_n_61 ,add_178_21_n_31 ,add_178_21_n_59);
  xnor add_178_21_g375(n_430 ,add_178_21_n_58 ,add_178_21_n_43);
  and add_178_21_g376(add_178_21_n_59 ,add_178_21_n_26 ,add_178_21_n_58);
  or add_178_21_g377(add_178_21_n_58 ,add_178_21_n_27 ,add_178_21_n_56);
  xnor add_178_21_g378(n_429 ,add_178_21_n_55 ,add_178_21_n_34);
  and add_178_21_g379(add_178_21_n_56 ,add_178_21_n_7 ,add_178_21_n_55);
  or add_178_21_g380(add_178_21_n_55 ,add_178_21_n_5 ,add_178_21_n_53);
  xnor add_178_21_g381(n_428 ,add_178_21_n_51 ,add_178_21_n_41);
  and add_178_21_g382(add_178_21_n_53 ,add_178_21_n_23 ,add_178_21_n_51);
  xor add_178_21_g383(n_427 ,add_178_21_n_33 ,add_178_21_n_40);
  or add_178_21_g384(add_178_21_n_51 ,add_178_21_n_4 ,add_178_21_n_49);
  and add_178_21_g385(n_426 ,add_178_21_n_33 ,add_178_21_n_13);
  nor add_178_21_g386(add_178_21_n_49 ,add_178_21_n_33 ,add_178_21_n_14);
  xnor add_178_21_g387(add_178_21_n_48 ,in51[9] ,in52[9]);
  xnor add_178_21_g388(add_178_21_n_47 ,in51[8] ,in52[8]);
  xnor add_178_21_g389(add_178_21_n_46 ,in51[7] ,in52[7]);
  xnor add_178_21_g390(add_178_21_n_45 ,in51[6] ,in52[6]);
  xnor add_178_21_g391(add_178_21_n_44 ,in51[5] ,in52[5]);
  xnor add_178_21_g392(add_178_21_n_43 ,in51[4] ,in52[4]);
  xnor add_178_21_g393(add_178_21_n_42 ,in51[10] ,in52[10]);
  xnor add_178_21_g394(add_178_21_n_41 ,in51[2] ,in52[2]);
  xnor add_178_21_g395(add_178_21_n_40 ,in51[1] ,in52[1]);
  xnor add_178_21_g396(add_178_21_n_39 ,in51[15] ,in52[15]);
  xnor add_178_21_g397(add_178_21_n_38 ,in51[14] ,in52[14]);
  xnor add_178_21_g398(add_178_21_n_37 ,in51[13] ,in52[13]);
  xnor add_178_21_g399(add_178_21_n_36 ,in51[12] ,in52[12]);
  xnor add_178_21_g400(add_178_21_n_35 ,in51[11] ,in52[11]);
  xnor add_178_21_g401(add_178_21_n_34 ,in51[3] ,in52[3]);
  and add_178_21_g402(add_178_21_n_32 ,in51[10] ,in52[10]);
  and add_178_21_g403(add_178_21_n_31 ,in51[4] ,in52[4]);
  or add_178_21_g404(add_178_21_n_30 ,in51[5] ,in52[5]);
  and add_178_21_g405(add_178_21_n_29 ,in51[15] ,in52[15]);
  and add_178_21_g406(add_178_21_n_28 ,in51[8] ,in52[8]);
  and add_178_21_g407(add_178_21_n_27 ,in51[3] ,in52[3]);
  or add_178_21_g408(add_178_21_n_26 ,in51[4] ,in52[4]);
  or add_178_21_g409(add_178_21_n_25 ,in51[7] ,in52[7]);
  and add_178_21_g410(add_178_21_n_24 ,in51[14] ,in52[14]);
  or add_178_21_g411(add_178_21_n_23 ,in51[2] ,in52[2]);
  or add_178_21_g412(add_178_21_n_22 ,in51[11] ,in52[11]);
  and add_178_21_g413(add_178_21_n_21 ,in51[9] ,in52[9]);
  and add_178_21_g414(add_178_21_n_20 ,in51[13] ,in52[13]);
  or add_178_21_g415(add_178_21_n_19 ,in51[9] ,in52[9]);
  or add_178_21_g416(add_178_21_n_18 ,in51[6] ,in52[6]);
  or add_178_21_g417(add_178_21_n_33 ,add_178_21_n_1 ,add_178_21_n_0);
  and add_178_21_g418(add_178_21_n_17 ,in51[7] ,in52[7]);
  or add_178_21_g419(add_178_21_n_16 ,in51[13] ,in52[13]);
  nor add_178_21_g420(add_178_21_n_15 ,in51[15] ,in52[15]);
  nor add_178_21_g421(add_178_21_n_14 ,in51[1] ,in52[1]);
  or add_178_21_g422(add_178_21_n_13 ,in51[0] ,in52[0]);
  or add_178_21_g423(add_178_21_n_12 ,in51[12] ,in52[12]);
  or add_178_21_g424(add_178_21_n_11 ,in51[8] ,in52[8]);
  and add_178_21_g425(add_178_21_n_10 ,in51[12] ,in52[12]);
  or add_178_21_g426(add_178_21_n_9 ,in51[14] ,in52[14]);
  and add_178_21_g427(add_178_21_n_8 ,in51[11] ,in52[11]);
  or add_178_21_g428(add_178_21_n_7 ,in51[3] ,in52[3]);
  and add_178_21_g429(add_178_21_n_6 ,in51[6] ,in52[6]);
  and add_178_21_g430(add_178_21_n_5 ,in51[2] ,in52[2]);
  and add_178_21_g431(add_178_21_n_4 ,in51[1] ,in52[1]);
  and add_178_21_g432(add_178_21_n_3 ,in51[5] ,in52[5]);
  or add_178_21_g433(add_178_21_n_2 ,in51[10] ,in52[10]);
  not add_178_21_g434(add_178_21_n_1 ,in51[0]);
  not add_178_21_g435(add_178_21_n_0 ,in52[0]);
  or add_180_21_g341(n_459 ,add_180_21_n_29 ,add_180_21_n_92);
  xnor add_180_21_g342(n_458 ,add_180_21_n_91 ,add_180_21_n_39);
  nor add_180_21_g343(add_180_21_n_92 ,add_180_21_n_15 ,add_180_21_n_91);
  or add_180_21_g344(add_180_21_n_91 ,add_180_21_n_24 ,add_180_21_n_89);
  xnor add_180_21_g345(n_457 ,add_180_21_n_88 ,add_180_21_n_38);
  and add_180_21_g346(add_180_21_n_89 ,add_180_21_n_9 ,add_180_21_n_88);
  or add_180_21_g347(add_180_21_n_88 ,add_180_21_n_20 ,add_180_21_n_86);
  xnor add_180_21_g348(n_456 ,add_180_21_n_85 ,add_180_21_n_37);
  and add_180_21_g349(add_180_21_n_86 ,add_180_21_n_16 ,add_180_21_n_85);
  or add_180_21_g350(add_180_21_n_85 ,add_180_21_n_10 ,add_180_21_n_83);
  xnor add_180_21_g351(n_455 ,add_180_21_n_82 ,add_180_21_n_36);
  and add_180_21_g352(add_180_21_n_83 ,add_180_21_n_12 ,add_180_21_n_82);
  or add_180_21_g353(add_180_21_n_82 ,add_180_21_n_8 ,add_180_21_n_80);
  xnor add_180_21_g354(n_454 ,add_180_21_n_79 ,add_180_21_n_35);
  and add_180_21_g355(add_180_21_n_80 ,add_180_21_n_22 ,add_180_21_n_79);
  or add_180_21_g356(add_180_21_n_79 ,add_180_21_n_32 ,add_180_21_n_77);
  xnor add_180_21_g357(n_453 ,add_180_21_n_76 ,add_180_21_n_42);
  and add_180_21_g358(add_180_21_n_77 ,add_180_21_n_2 ,add_180_21_n_76);
  or add_180_21_g359(add_180_21_n_76 ,add_180_21_n_21 ,add_180_21_n_74);
  xnor add_180_21_g360(n_452 ,add_180_21_n_73 ,add_180_21_n_48);
  and add_180_21_g361(add_180_21_n_74 ,add_180_21_n_19 ,add_180_21_n_73);
  or add_180_21_g362(add_180_21_n_73 ,add_180_21_n_28 ,add_180_21_n_71);
  xnor add_180_21_g363(n_451 ,add_180_21_n_70 ,add_180_21_n_47);
  and add_180_21_g364(add_180_21_n_71 ,add_180_21_n_11 ,add_180_21_n_70);
  or add_180_21_g365(add_180_21_n_70 ,add_180_21_n_17 ,add_180_21_n_68);
  xnor add_180_21_g366(n_450 ,add_180_21_n_67 ,add_180_21_n_46);
  and add_180_21_g367(add_180_21_n_68 ,add_180_21_n_25 ,add_180_21_n_67);
  or add_180_21_g368(add_180_21_n_67 ,add_180_21_n_6 ,add_180_21_n_65);
  xnor add_180_21_g369(n_449 ,add_180_21_n_64 ,add_180_21_n_45);
  and add_180_21_g370(add_180_21_n_65 ,add_180_21_n_18 ,add_180_21_n_64);
  or add_180_21_g371(add_180_21_n_64 ,add_180_21_n_3 ,add_180_21_n_62);
  xnor add_180_21_g372(n_448 ,add_180_21_n_61 ,add_180_21_n_44);
  and add_180_21_g373(add_180_21_n_62 ,add_180_21_n_30 ,add_180_21_n_61);
  or add_180_21_g374(add_180_21_n_61 ,add_180_21_n_31 ,add_180_21_n_59);
  xnor add_180_21_g375(n_447 ,add_180_21_n_58 ,add_180_21_n_43);
  and add_180_21_g376(add_180_21_n_59 ,add_180_21_n_26 ,add_180_21_n_58);
  or add_180_21_g377(add_180_21_n_58 ,add_180_21_n_27 ,add_180_21_n_56);
  xnor add_180_21_g378(n_446 ,add_180_21_n_55 ,add_180_21_n_34);
  and add_180_21_g379(add_180_21_n_56 ,add_180_21_n_7 ,add_180_21_n_55);
  or add_180_21_g380(add_180_21_n_55 ,add_180_21_n_5 ,add_180_21_n_53);
  xnor add_180_21_g381(n_445 ,add_180_21_n_51 ,add_180_21_n_41);
  and add_180_21_g382(add_180_21_n_53 ,add_180_21_n_23 ,add_180_21_n_51);
  xor add_180_21_g383(n_444 ,add_180_21_n_33 ,add_180_21_n_40);
  or add_180_21_g384(add_180_21_n_51 ,add_180_21_n_4 ,add_180_21_n_49);
  and add_180_21_g385(n_443 ,add_180_21_n_33 ,add_180_21_n_13);
  nor add_180_21_g386(add_180_21_n_49 ,add_180_21_n_33 ,add_180_21_n_14);
  xnor add_180_21_g387(add_180_21_n_48 ,in53[9] ,in54[9]);
  xnor add_180_21_g388(add_180_21_n_47 ,in53[8] ,in54[8]);
  xnor add_180_21_g389(add_180_21_n_46 ,in53[7] ,in54[7]);
  xnor add_180_21_g390(add_180_21_n_45 ,in53[6] ,in54[6]);
  xnor add_180_21_g391(add_180_21_n_44 ,in53[5] ,in54[5]);
  xnor add_180_21_g392(add_180_21_n_43 ,in53[4] ,in54[4]);
  xnor add_180_21_g393(add_180_21_n_42 ,in53[10] ,in54[10]);
  xnor add_180_21_g394(add_180_21_n_41 ,in53[2] ,in54[2]);
  xnor add_180_21_g395(add_180_21_n_40 ,in53[1] ,in54[1]);
  xnor add_180_21_g396(add_180_21_n_39 ,in53[15] ,in54[15]);
  xnor add_180_21_g397(add_180_21_n_38 ,in53[14] ,in54[14]);
  xnor add_180_21_g398(add_180_21_n_37 ,in53[13] ,in54[13]);
  xnor add_180_21_g399(add_180_21_n_36 ,in53[12] ,in54[12]);
  xnor add_180_21_g400(add_180_21_n_35 ,in53[11] ,in54[11]);
  xnor add_180_21_g401(add_180_21_n_34 ,in53[3] ,in54[3]);
  and add_180_21_g402(add_180_21_n_32 ,in53[10] ,in54[10]);
  and add_180_21_g403(add_180_21_n_31 ,in53[4] ,in54[4]);
  or add_180_21_g404(add_180_21_n_30 ,in53[5] ,in54[5]);
  and add_180_21_g405(add_180_21_n_29 ,in53[15] ,in54[15]);
  and add_180_21_g406(add_180_21_n_28 ,in53[8] ,in54[8]);
  and add_180_21_g407(add_180_21_n_27 ,in53[3] ,in54[3]);
  or add_180_21_g408(add_180_21_n_26 ,in53[4] ,in54[4]);
  or add_180_21_g409(add_180_21_n_25 ,in53[7] ,in54[7]);
  and add_180_21_g410(add_180_21_n_24 ,in53[14] ,in54[14]);
  or add_180_21_g411(add_180_21_n_23 ,in53[2] ,in54[2]);
  or add_180_21_g412(add_180_21_n_22 ,in53[11] ,in54[11]);
  and add_180_21_g413(add_180_21_n_21 ,in53[9] ,in54[9]);
  and add_180_21_g414(add_180_21_n_20 ,in53[13] ,in54[13]);
  or add_180_21_g415(add_180_21_n_19 ,in53[9] ,in54[9]);
  or add_180_21_g416(add_180_21_n_18 ,in53[6] ,in54[6]);
  or add_180_21_g417(add_180_21_n_33 ,add_180_21_n_1 ,add_180_21_n_0);
  and add_180_21_g418(add_180_21_n_17 ,in53[7] ,in54[7]);
  or add_180_21_g419(add_180_21_n_16 ,in53[13] ,in54[13]);
  nor add_180_21_g420(add_180_21_n_15 ,in53[15] ,in54[15]);
  nor add_180_21_g421(add_180_21_n_14 ,in53[1] ,in54[1]);
  or add_180_21_g422(add_180_21_n_13 ,in53[0] ,in54[0]);
  or add_180_21_g423(add_180_21_n_12 ,in53[12] ,in54[12]);
  or add_180_21_g424(add_180_21_n_11 ,in53[8] ,in54[8]);
  and add_180_21_g425(add_180_21_n_10 ,in53[12] ,in54[12]);
  or add_180_21_g426(add_180_21_n_9 ,in53[14] ,in54[14]);
  and add_180_21_g427(add_180_21_n_8 ,in53[11] ,in54[11]);
  or add_180_21_g428(add_180_21_n_7 ,in53[3] ,in54[3]);
  and add_180_21_g429(add_180_21_n_6 ,in53[6] ,in54[6]);
  and add_180_21_g430(add_180_21_n_5 ,in53[2] ,in54[2]);
  and add_180_21_g431(add_180_21_n_4 ,in53[1] ,in54[1]);
  and add_180_21_g432(add_180_21_n_3 ,in53[5] ,in54[5]);
  or add_180_21_g433(add_180_21_n_2 ,in53[10] ,in54[10]);
  not add_180_21_g434(add_180_21_n_1 ,in53[0]);
  not add_180_21_g435(add_180_21_n_0 ,in54[0]);
  xnor csa_tree_add_190_195_groupi_g36279(out1[28] ,csa_tree_add_190_195_groupi_n_12610 ,csa_tree_add_190_195_groupi_n_8314);
  or csa_tree_add_190_195_groupi_g36280(csa_tree_add_190_195_groupi_n_12610 ,csa_tree_add_190_195_groupi_n_11739 ,csa_tree_add_190_195_groupi_n_12608);
  xnor csa_tree_add_190_195_groupi_g36281(csa_tree_add_190_195_groupi_n_12609 ,csa_tree_add_190_195_groupi_n_12607 ,csa_tree_add_190_195_groupi_n_11843);
  nor csa_tree_add_190_195_groupi_g36282(csa_tree_add_190_195_groupi_n_12608 ,csa_tree_add_190_195_groupi_n_11791 ,csa_tree_add_190_195_groupi_n_12607);
  and csa_tree_add_190_195_groupi_g36283(csa_tree_add_190_195_groupi_n_12607 ,csa_tree_add_190_195_groupi_n_12318 ,csa_tree_add_190_195_groupi_n_12605);
  xnor csa_tree_add_190_195_groupi_g36284(csa_tree_add_190_195_groupi_n_12606 ,csa_tree_add_190_195_groupi_n_12604 ,csa_tree_add_190_195_groupi_n_12332);
  or csa_tree_add_190_195_groupi_g36285(csa_tree_add_190_195_groupi_n_12605 ,csa_tree_add_190_195_groupi_n_12604 ,csa_tree_add_190_195_groupi_n_12283);
  and csa_tree_add_190_195_groupi_g36286(csa_tree_add_190_195_groupi_n_12604 ,csa_tree_add_190_195_groupi_n_12363 ,csa_tree_add_190_195_groupi_n_12602);
  xnor csa_tree_add_190_195_groupi_g36287(csa_tree_add_190_195_groupi_n_12603 ,csa_tree_add_190_195_groupi_n_12601 ,csa_tree_add_190_195_groupi_n_12378);
  or csa_tree_add_190_195_groupi_g36288(csa_tree_add_190_195_groupi_n_12602 ,csa_tree_add_190_195_groupi_n_12354 ,csa_tree_add_190_195_groupi_n_12601);
  and csa_tree_add_190_195_groupi_g36289(csa_tree_add_190_195_groupi_n_12601 ,csa_tree_add_190_195_groupi_n_12468 ,csa_tree_add_190_195_groupi_n_12599);
  xnor csa_tree_add_190_195_groupi_g36290(csa_tree_add_190_195_groupi_n_12600 ,csa_tree_add_190_195_groupi_n_12598 ,csa_tree_add_190_195_groupi_n_12481);
  or csa_tree_add_190_195_groupi_g36291(csa_tree_add_190_195_groupi_n_12599 ,csa_tree_add_190_195_groupi_n_12467 ,csa_tree_add_190_195_groupi_n_12598);
  and csa_tree_add_190_195_groupi_g36292(csa_tree_add_190_195_groupi_n_12598 ,csa_tree_add_190_195_groupi_n_12492 ,csa_tree_add_190_195_groupi_n_12596);
  xnor csa_tree_add_190_195_groupi_g36293(csa_tree_add_190_195_groupi_n_12597 ,csa_tree_add_190_195_groupi_n_12595 ,csa_tree_add_190_195_groupi_n_180);
  or csa_tree_add_190_195_groupi_g36294(csa_tree_add_190_195_groupi_n_12596 ,csa_tree_add_190_195_groupi_n_12595 ,csa_tree_add_190_195_groupi_n_12484);
  and csa_tree_add_190_195_groupi_g36295(csa_tree_add_190_195_groupi_n_12595 ,csa_tree_add_190_195_groupi_n_12514 ,csa_tree_add_190_195_groupi_n_12593);
  xnor csa_tree_add_190_195_groupi_g36296(csa_tree_add_190_195_groupi_n_12594 ,csa_tree_add_190_195_groupi_n_12592 ,csa_tree_add_190_195_groupi_n_182);
  or csa_tree_add_190_195_groupi_g36297(csa_tree_add_190_195_groupi_n_12593 ,csa_tree_add_190_195_groupi_n_12592 ,csa_tree_add_190_195_groupi_n_12504);
  and csa_tree_add_190_195_groupi_g36298(csa_tree_add_190_195_groupi_n_12592 ,csa_tree_add_190_195_groupi_n_12537 ,csa_tree_add_190_195_groupi_n_12591);
  or csa_tree_add_190_195_groupi_g36300(csa_tree_add_190_195_groupi_n_12591 ,csa_tree_add_190_195_groupi_n_12590 ,csa_tree_add_190_195_groupi_n_12527);
  and csa_tree_add_190_195_groupi_g36302(csa_tree_add_190_195_groupi_n_12590 ,csa_tree_add_190_195_groupi_n_12588 ,csa_tree_add_190_195_groupi_n_12549);
  xnor csa_tree_add_190_195_groupi_g36303(csa_tree_add_190_195_groupi_n_12589 ,csa_tree_add_190_195_groupi_n_12587 ,csa_tree_add_190_195_groupi_n_12555);
  or csa_tree_add_190_195_groupi_g36304(csa_tree_add_190_195_groupi_n_12588 ,csa_tree_add_190_195_groupi_n_12587 ,csa_tree_add_190_195_groupi_n_12550);
  and csa_tree_add_190_195_groupi_g36305(csa_tree_add_190_195_groupi_n_12587 ,csa_tree_add_190_195_groupi_n_12586 ,csa_tree_add_190_195_groupi_n_12556);
  or csa_tree_add_190_195_groupi_g36307(csa_tree_add_190_195_groupi_n_12586 ,csa_tree_add_190_195_groupi_n_12557 ,csa_tree_add_190_195_groupi_n_12585);
  and csa_tree_add_190_195_groupi_g36309(csa_tree_add_190_195_groupi_n_12585 ,csa_tree_add_190_195_groupi_n_12559 ,csa_tree_add_190_195_groupi_n_12583);
  xnor csa_tree_add_190_195_groupi_g36310(out1[18] ,csa_tree_add_190_195_groupi_n_12581 ,csa_tree_add_190_195_groupi_n_12561);
  or csa_tree_add_190_195_groupi_g36311(csa_tree_add_190_195_groupi_n_12583 ,csa_tree_add_190_195_groupi_n_12558 ,csa_tree_add_190_195_groupi_n_12582);
  not csa_tree_add_190_195_groupi_g36312(csa_tree_add_190_195_groupi_n_12582 ,csa_tree_add_190_195_groupi_n_12581);
  or csa_tree_add_190_195_groupi_g36313(csa_tree_add_190_195_groupi_n_12581 ,csa_tree_add_190_195_groupi_n_12552 ,csa_tree_add_190_195_groupi_n_12579);
  xnor csa_tree_add_190_195_groupi_g36314(csa_tree_add_190_195_groupi_n_12580 ,csa_tree_add_190_195_groupi_n_12578 ,csa_tree_add_190_195_groupi_n_183);
  nor csa_tree_add_190_195_groupi_g36315(csa_tree_add_190_195_groupi_n_12579 ,csa_tree_add_190_195_groupi_n_12578 ,csa_tree_add_190_195_groupi_n_12553);
  and csa_tree_add_190_195_groupi_g36316(csa_tree_add_190_195_groupi_n_12578 ,csa_tree_add_190_195_groupi_n_12576 ,csa_tree_add_190_195_groupi_n_12528);
  xnor csa_tree_add_190_195_groupi_g36317(out1[16] ,csa_tree_add_190_195_groupi_n_12574 ,csa_tree_add_190_195_groupi_n_12543);
  or csa_tree_add_190_195_groupi_g36318(csa_tree_add_190_195_groupi_n_12576 ,csa_tree_add_190_195_groupi_n_12575 ,csa_tree_add_190_195_groupi_n_12539);
  not csa_tree_add_190_195_groupi_g36319(csa_tree_add_190_195_groupi_n_12575 ,csa_tree_add_190_195_groupi_n_12574);
  or csa_tree_add_190_195_groupi_g36320(csa_tree_add_190_195_groupi_n_12574 ,csa_tree_add_190_195_groupi_n_12535 ,csa_tree_add_190_195_groupi_n_12572);
  xnor csa_tree_add_190_195_groupi_g36321(csa_tree_add_190_195_groupi_n_12573 ,csa_tree_add_190_195_groupi_n_12571 ,csa_tree_add_190_195_groupi_n_12544);
  nor csa_tree_add_190_195_groupi_g36322(csa_tree_add_190_195_groupi_n_12572 ,csa_tree_add_190_195_groupi_n_12571 ,csa_tree_add_190_195_groupi_n_12534);
  and csa_tree_add_190_195_groupi_g36323(csa_tree_add_190_195_groupi_n_12571 ,csa_tree_add_190_195_groupi_n_12538 ,csa_tree_add_190_195_groupi_n_12569);
  xnor csa_tree_add_190_195_groupi_g36324(csa_tree_add_190_195_groupi_n_12570 ,csa_tree_add_190_195_groupi_n_12567 ,csa_tree_add_190_195_groupi_n_12541);
  or csa_tree_add_190_195_groupi_g36325(csa_tree_add_190_195_groupi_n_12569 ,csa_tree_add_190_195_groupi_n_12536 ,csa_tree_add_190_195_groupi_n_12568);
  not csa_tree_add_190_195_groupi_g36326(csa_tree_add_190_195_groupi_n_12568 ,csa_tree_add_190_195_groupi_n_12567);
  or csa_tree_add_190_195_groupi_g36327(csa_tree_add_190_195_groupi_n_12567 ,csa_tree_add_190_195_groupi_n_12515 ,csa_tree_add_190_195_groupi_n_12565);
  xnor csa_tree_add_190_195_groupi_g36328(csa_tree_add_190_195_groupi_n_12566 ,csa_tree_add_190_195_groupi_n_12564 ,csa_tree_add_190_195_groupi_n_12526);
  nor csa_tree_add_190_195_groupi_g36329(csa_tree_add_190_195_groupi_n_12565 ,csa_tree_add_190_195_groupi_n_12564 ,csa_tree_add_190_195_groupi_n_12505);
  and csa_tree_add_190_195_groupi_g36330(csa_tree_add_190_195_groupi_n_12564 ,csa_tree_add_190_195_groupi_n_12491 ,csa_tree_add_190_195_groupi_n_12563);
  or csa_tree_add_190_195_groupi_g36332(csa_tree_add_190_195_groupi_n_12563 ,csa_tree_add_190_195_groupi_n_12495 ,csa_tree_add_190_195_groupi_n_12560);
  xnor csa_tree_add_190_195_groupi_g36333(csa_tree_add_190_195_groupi_n_12562 ,csa_tree_add_190_195_groupi_n_12533 ,csa_tree_add_190_195_groupi_n_12548);
  xnor csa_tree_add_190_195_groupi_g36334(csa_tree_add_190_195_groupi_n_12561 ,csa_tree_add_190_195_groupi_n_12546 ,csa_tree_add_190_195_groupi_n_12519);
  and csa_tree_add_190_195_groupi_g36336(csa_tree_add_190_195_groupi_n_12560 ,csa_tree_add_190_195_groupi_n_12471 ,csa_tree_add_190_195_groupi_n_12551);
  or csa_tree_add_190_195_groupi_g36337(csa_tree_add_190_195_groupi_n_12559 ,csa_tree_add_190_195_groupi_n_12545 ,csa_tree_add_190_195_groupi_n_12518);
  nor csa_tree_add_190_195_groupi_g36338(csa_tree_add_190_195_groupi_n_12558 ,csa_tree_add_190_195_groupi_n_12546 ,csa_tree_add_190_195_groupi_n_12519);
  nor csa_tree_add_190_195_groupi_g36339(csa_tree_add_190_195_groupi_n_12557 ,csa_tree_add_190_195_groupi_n_12533 ,csa_tree_add_190_195_groupi_n_12548);
  or csa_tree_add_190_195_groupi_g36340(csa_tree_add_190_195_groupi_n_12556 ,csa_tree_add_190_195_groupi_n_12532 ,csa_tree_add_190_195_groupi_n_12547);
  xnor csa_tree_add_190_195_groupi_g36341(csa_tree_add_190_195_groupi_n_12555 ,csa_tree_add_190_195_groupi_n_12530 ,csa_tree_add_190_195_groupi_n_12521);
  xnor csa_tree_add_190_195_groupi_g36343(out1[11] ,csa_tree_add_190_195_groupi_n_12540 ,csa_tree_add_190_195_groupi_n_12480);
  and csa_tree_add_190_195_groupi_g36344(csa_tree_add_190_195_groupi_n_12553 ,csa_tree_add_190_195_groupi_n_12531 ,csa_tree_add_190_195_groupi_n_12525);
  nor csa_tree_add_190_195_groupi_g36345(csa_tree_add_190_195_groupi_n_12552 ,csa_tree_add_190_195_groupi_n_12531 ,csa_tree_add_190_195_groupi_n_12525);
  or csa_tree_add_190_195_groupi_g36346(csa_tree_add_190_195_groupi_n_12551 ,csa_tree_add_190_195_groupi_n_12540 ,csa_tree_add_190_195_groupi_n_12470);
  nor csa_tree_add_190_195_groupi_g36347(csa_tree_add_190_195_groupi_n_12550 ,csa_tree_add_190_195_groupi_n_12529 ,csa_tree_add_190_195_groupi_n_12521);
  or csa_tree_add_190_195_groupi_g36348(csa_tree_add_190_195_groupi_n_12549 ,csa_tree_add_190_195_groupi_n_12530 ,csa_tree_add_190_195_groupi_n_12520);
  not csa_tree_add_190_195_groupi_g36349(csa_tree_add_190_195_groupi_n_12548 ,csa_tree_add_190_195_groupi_n_12547);
  not csa_tree_add_190_195_groupi_g36350(csa_tree_add_190_195_groupi_n_12546 ,csa_tree_add_190_195_groupi_n_12545);
  xnor csa_tree_add_190_195_groupi_g36351(csa_tree_add_190_195_groupi_n_12544 ,csa_tree_add_190_195_groupi_n_12522 ,csa_tree_add_190_195_groupi_n_12510);
  xnor csa_tree_add_190_195_groupi_g36352(csa_tree_add_190_195_groupi_n_12543 ,csa_tree_add_190_195_groupi_n_12489 ,csa_tree_add_190_195_groupi_n_12507);
  xnor csa_tree_add_190_195_groupi_g36353(csa_tree_add_190_195_groupi_n_12542 ,csa_tree_add_190_195_groupi_n_12524 ,csa_tree_add_190_195_groupi_n_12513);
  xnor csa_tree_add_190_195_groupi_g36354(csa_tree_add_190_195_groupi_n_12541 ,csa_tree_add_190_195_groupi_n_12509 ,csa_tree_add_190_195_groupi_n_12476);
  xnor csa_tree_add_190_195_groupi_g36355(csa_tree_add_190_195_groupi_n_12547 ,csa_tree_add_190_195_groupi_n_12438 ,csa_tree_add_190_195_groupi_n_12501);
  xnor csa_tree_add_190_195_groupi_g36356(csa_tree_add_190_195_groupi_n_12545 ,csa_tree_add_190_195_groupi_n_12444 ,csa_tree_add_190_195_groupi_n_12502);
  nor csa_tree_add_190_195_groupi_g36357(csa_tree_add_190_195_groupi_n_12539 ,csa_tree_add_190_195_groupi_n_12489 ,csa_tree_add_190_195_groupi_n_12507);
  or csa_tree_add_190_195_groupi_g36358(csa_tree_add_190_195_groupi_n_12538 ,csa_tree_add_190_195_groupi_n_12508 ,csa_tree_add_190_195_groupi_n_12475);
  or csa_tree_add_190_195_groupi_g36359(csa_tree_add_190_195_groupi_n_12537 ,csa_tree_add_190_195_groupi_n_12523 ,csa_tree_add_190_195_groupi_n_12512);
  nor csa_tree_add_190_195_groupi_g36360(csa_tree_add_190_195_groupi_n_12536 ,csa_tree_add_190_195_groupi_n_12509 ,csa_tree_add_190_195_groupi_n_12476);
  nor csa_tree_add_190_195_groupi_g36361(csa_tree_add_190_195_groupi_n_12535 ,csa_tree_add_190_195_groupi_n_12522 ,csa_tree_add_190_195_groupi_n_12511);
  and csa_tree_add_190_195_groupi_g36362(csa_tree_add_190_195_groupi_n_12534 ,csa_tree_add_190_195_groupi_n_12522 ,csa_tree_add_190_195_groupi_n_12511);
  and csa_tree_add_190_195_groupi_g36363(csa_tree_add_190_195_groupi_n_12540 ,csa_tree_add_190_195_groupi_n_12419 ,csa_tree_add_190_195_groupi_n_12517);
  not csa_tree_add_190_195_groupi_g36364(csa_tree_add_190_195_groupi_n_12533 ,csa_tree_add_190_195_groupi_n_12532);
  not csa_tree_add_190_195_groupi_g36365(csa_tree_add_190_195_groupi_n_12530 ,csa_tree_add_190_195_groupi_n_12529);
  or csa_tree_add_190_195_groupi_g36366(csa_tree_add_190_195_groupi_n_12528 ,csa_tree_add_190_195_groupi_n_12488 ,csa_tree_add_190_195_groupi_n_12506);
  nor csa_tree_add_190_195_groupi_g36367(csa_tree_add_190_195_groupi_n_12527 ,csa_tree_add_190_195_groupi_n_12524 ,csa_tree_add_190_195_groupi_n_12513);
  xnor csa_tree_add_190_195_groupi_g36369(csa_tree_add_190_195_groupi_n_12526 ,csa_tree_add_190_195_groupi_n_12487 ,csa_tree_add_190_195_groupi_n_12477);
  and csa_tree_add_190_195_groupi_g36371(csa_tree_add_190_195_groupi_n_12532 ,csa_tree_add_190_195_groupi_n_12485 ,csa_tree_add_190_195_groupi_n_12516);
  xnor csa_tree_add_190_195_groupi_g36372(csa_tree_add_190_195_groupi_n_12531 ,csa_tree_add_190_195_groupi_n_12461 ,csa_tree_add_190_195_groupi_n_12482);
  xnor csa_tree_add_190_195_groupi_g36373(csa_tree_add_190_195_groupi_n_12529 ,csa_tree_add_190_195_groupi_n_12479 ,csa_tree_add_190_195_groupi_n_12483);
  not csa_tree_add_190_195_groupi_g36375(csa_tree_add_190_195_groupi_n_12524 ,csa_tree_add_190_195_groupi_n_12523);
  not csa_tree_add_190_195_groupi_g36376(csa_tree_add_190_195_groupi_n_12521 ,csa_tree_add_190_195_groupi_n_12520);
  not csa_tree_add_190_195_groupi_g36377(csa_tree_add_190_195_groupi_n_12518 ,csa_tree_add_190_195_groupi_n_12519);
  or csa_tree_add_190_195_groupi_g36378(csa_tree_add_190_195_groupi_n_12517 ,csa_tree_add_190_195_groupi_n_12420 ,csa_tree_add_190_195_groupi_n_12490);
  or csa_tree_add_190_195_groupi_g36379(csa_tree_add_190_195_groupi_n_12516 ,csa_tree_add_190_195_groupi_n_12498 ,csa_tree_add_190_195_groupi_n_12444);
  nor csa_tree_add_190_195_groupi_g36380(csa_tree_add_190_195_groupi_n_12515 ,csa_tree_add_190_195_groupi_n_12487 ,csa_tree_add_190_195_groupi_n_12478);
  or csa_tree_add_190_195_groupi_g36381(csa_tree_add_190_195_groupi_n_12514 ,csa_tree_add_190_195_groupi_n_12486 ,csa_tree_add_190_195_groupi_n_12500);
  and csa_tree_add_190_195_groupi_g36382(csa_tree_add_190_195_groupi_n_12525 ,csa_tree_add_190_195_groupi_n_12496 ,csa_tree_add_190_195_groupi_n_12430);
  and csa_tree_add_190_195_groupi_g36383(csa_tree_add_190_195_groupi_n_12523 ,csa_tree_add_190_195_groupi_n_12463 ,csa_tree_add_190_195_groupi_n_12493);
  and csa_tree_add_190_195_groupi_g36384(csa_tree_add_190_195_groupi_n_12522 ,csa_tree_add_190_195_groupi_n_12465 ,csa_tree_add_190_195_groupi_n_12494);
  and csa_tree_add_190_195_groupi_g36385(csa_tree_add_190_195_groupi_n_12520 ,csa_tree_add_190_195_groupi_n_12499 ,csa_tree_add_190_195_groupi_n_12472);
  or csa_tree_add_190_195_groupi_g36386(csa_tree_add_190_195_groupi_n_12519 ,csa_tree_add_190_195_groupi_n_12497 ,csa_tree_add_190_195_groupi_n_12474);
  not csa_tree_add_190_195_groupi_g36387(csa_tree_add_190_195_groupi_n_12513 ,csa_tree_add_190_195_groupi_n_12512);
  not csa_tree_add_190_195_groupi_g36388(csa_tree_add_190_195_groupi_n_12511 ,csa_tree_add_190_195_groupi_n_12510);
  not csa_tree_add_190_195_groupi_g36389(csa_tree_add_190_195_groupi_n_12509 ,csa_tree_add_190_195_groupi_n_12508);
  not csa_tree_add_190_195_groupi_g36390(csa_tree_add_190_195_groupi_n_12507 ,csa_tree_add_190_195_groupi_n_12506);
  and csa_tree_add_190_195_groupi_g36391(csa_tree_add_190_195_groupi_n_12505 ,csa_tree_add_190_195_groupi_n_12487 ,csa_tree_add_190_195_groupi_n_12478);
  and csa_tree_add_190_195_groupi_g36392(csa_tree_add_190_195_groupi_n_12504 ,csa_tree_add_190_195_groupi_n_12486 ,csa_tree_add_190_195_groupi_n_12500);
  xnor csa_tree_add_190_195_groupi_g36393(csa_tree_add_190_195_groupi_n_12503 ,csa_tree_add_190_195_groupi_n_12459 ,csa_tree_add_190_195_groupi_n_12440);
  xnor csa_tree_add_190_195_groupi_g36395(csa_tree_add_190_195_groupi_n_12502 ,csa_tree_add_190_195_groupi_n_12344 ,csa_tree_add_190_195_groupi_n_12456);
  xnor csa_tree_add_190_195_groupi_g36396(csa_tree_add_190_195_groupi_n_12501 ,csa_tree_add_190_195_groupi_n_12462 ,csa_tree_add_190_195_groupi_n_12388);
  xnor csa_tree_add_190_195_groupi_g36397(csa_tree_add_190_195_groupi_n_12512 ,csa_tree_add_190_195_groupi_n_12445 ,csa_tree_add_190_195_groupi_n_12447);
  xnor csa_tree_add_190_195_groupi_g36398(csa_tree_add_190_195_groupi_n_12510 ,csa_tree_add_190_195_groupi_n_12427 ,csa_tree_add_190_195_groupi_n_12450);
  xnor csa_tree_add_190_195_groupi_g36399(csa_tree_add_190_195_groupi_n_12508 ,csa_tree_add_190_195_groupi_n_12423 ,csa_tree_add_190_195_groupi_n_12446);
  xnor csa_tree_add_190_195_groupi_g36400(csa_tree_add_190_195_groupi_n_12506 ,csa_tree_add_190_195_groupi_n_12460 ,csa_tree_add_190_195_groupi_n_12448);
  or csa_tree_add_190_195_groupi_g36402(csa_tree_add_190_195_groupi_n_12499 ,csa_tree_add_190_195_groupi_n_12462 ,csa_tree_add_190_195_groupi_n_12473);
  nor csa_tree_add_190_195_groupi_g36403(csa_tree_add_190_195_groupi_n_12498 ,csa_tree_add_190_195_groupi_n_12344 ,csa_tree_add_190_195_groupi_n_12456);
  nor csa_tree_add_190_195_groupi_g36404(csa_tree_add_190_195_groupi_n_12497 ,csa_tree_add_190_195_groupi_n_12469 ,csa_tree_add_190_195_groupi_n_12461);
  or csa_tree_add_190_195_groupi_g36405(csa_tree_add_190_195_groupi_n_12496 ,csa_tree_add_190_195_groupi_n_12434 ,csa_tree_add_190_195_groupi_n_12460);
  nor csa_tree_add_190_195_groupi_g36406(csa_tree_add_190_195_groupi_n_12495 ,csa_tree_add_190_195_groupi_n_12459 ,csa_tree_add_190_195_groupi_n_12440);
  or csa_tree_add_190_195_groupi_g36407(csa_tree_add_190_195_groupi_n_12494 ,csa_tree_add_190_195_groupi_n_12464 ,csa_tree_add_190_195_groupi_n_12412);
  or csa_tree_add_190_195_groupi_g36408(csa_tree_add_190_195_groupi_n_12493 ,csa_tree_add_190_195_groupi_n_12479 ,csa_tree_add_190_195_groupi_n_12451);
  or csa_tree_add_190_195_groupi_g36409(csa_tree_add_190_195_groupi_n_12492 ,csa_tree_add_190_195_groupi_n_12454 ,csa_tree_add_190_195_groupi_n_12457);
  or csa_tree_add_190_195_groupi_g36410(csa_tree_add_190_195_groupi_n_12491 ,csa_tree_add_190_195_groupi_n_12458 ,csa_tree_add_190_195_groupi_n_12439);
  and csa_tree_add_190_195_groupi_g36411(csa_tree_add_190_195_groupi_n_12500 ,csa_tree_add_190_195_groupi_n_12433 ,csa_tree_add_190_195_groupi_n_12466);
  not csa_tree_add_190_195_groupi_g36413(csa_tree_add_190_195_groupi_n_12489 ,csa_tree_add_190_195_groupi_n_12488);
  or csa_tree_add_190_195_groupi_g36414(csa_tree_add_190_195_groupi_n_12485 ,csa_tree_add_190_195_groupi_n_12343 ,csa_tree_add_190_195_groupi_n_12455);
  and csa_tree_add_190_195_groupi_g36416(csa_tree_add_190_195_groupi_n_12484 ,csa_tree_add_190_195_groupi_n_12454 ,csa_tree_add_190_195_groupi_n_12457);
  xnor csa_tree_add_190_195_groupi_g36417(csa_tree_add_190_195_groupi_n_12483 ,csa_tree_add_190_195_groupi_n_12426 ,csa_tree_add_190_195_groupi_n_12345);
  xnor csa_tree_add_190_195_groupi_g36418(csa_tree_add_190_195_groupi_n_12482 ,csa_tree_add_190_195_groupi_n_12342 ,csa_tree_add_190_195_groupi_n_12443);
  xnor csa_tree_add_190_195_groupi_g36419(csa_tree_add_190_195_groupi_n_12481 ,csa_tree_add_190_195_groupi_n_12442 ,csa_tree_add_190_195_groupi_n_12295);
  xnor csa_tree_add_190_195_groupi_g36420(csa_tree_add_190_195_groupi_n_12480 ,csa_tree_add_190_195_groupi_n_12425 ,csa_tree_add_190_195_groupi_n_12407);
  and csa_tree_add_190_195_groupi_g36421(csa_tree_add_190_195_groupi_n_12490 ,csa_tree_add_190_195_groupi_n_12453 ,csa_tree_add_190_195_groupi_n_12384);
  and csa_tree_add_190_195_groupi_g36422(csa_tree_add_190_195_groupi_n_12488 ,csa_tree_add_190_195_groupi_n_12418 ,csa_tree_add_190_195_groupi_n_12452);
  xnor csa_tree_add_190_195_groupi_g36423(csa_tree_add_190_195_groupi_n_12487 ,csa_tree_add_190_195_groupi_n_12391 ,csa_tree_add_190_195_groupi_n_12415);
  xnor csa_tree_add_190_195_groupi_g36424(csa_tree_add_190_195_groupi_n_12486 ,csa_tree_add_190_195_groupi_n_12413 ,csa_tree_add_190_195_groupi_n_12414);
  not csa_tree_add_190_195_groupi_g36425(csa_tree_add_190_195_groupi_n_12478 ,csa_tree_add_190_195_groupi_n_12477);
  not csa_tree_add_190_195_groupi_g36426(csa_tree_add_190_195_groupi_n_12476 ,csa_tree_add_190_195_groupi_n_12475);
  and csa_tree_add_190_195_groupi_g36427(csa_tree_add_190_195_groupi_n_12474 ,csa_tree_add_190_195_groupi_n_12342 ,csa_tree_add_190_195_groupi_n_12443);
  nor csa_tree_add_190_195_groupi_g36428(csa_tree_add_190_195_groupi_n_12473 ,csa_tree_add_190_195_groupi_n_12388 ,csa_tree_add_190_195_groupi_n_12438);
  or csa_tree_add_190_195_groupi_g36429(csa_tree_add_190_195_groupi_n_12472 ,csa_tree_add_190_195_groupi_n_12387 ,csa_tree_add_190_195_groupi_n_12437);
  or csa_tree_add_190_195_groupi_g36430(csa_tree_add_190_195_groupi_n_12471 ,csa_tree_add_190_195_groupi_n_12424 ,csa_tree_add_190_195_groupi_n_12407);
  nor csa_tree_add_190_195_groupi_g36431(csa_tree_add_190_195_groupi_n_12470 ,csa_tree_add_190_195_groupi_n_12425 ,csa_tree_add_190_195_groupi_n_12406);
  nor csa_tree_add_190_195_groupi_g36432(csa_tree_add_190_195_groupi_n_12469 ,csa_tree_add_190_195_groupi_n_12342 ,csa_tree_add_190_195_groupi_n_12443);
  or csa_tree_add_190_195_groupi_g36433(csa_tree_add_190_195_groupi_n_12468 ,csa_tree_add_190_195_groupi_n_12442 ,csa_tree_add_190_195_groupi_n_176);
  nor csa_tree_add_190_195_groupi_g36434(csa_tree_add_190_195_groupi_n_12467 ,csa_tree_add_190_195_groupi_n_12441 ,csa_tree_add_190_195_groupi_n_12295);
  or csa_tree_add_190_195_groupi_g36435(csa_tree_add_190_195_groupi_n_12466 ,csa_tree_add_190_195_groupi_n_12432 ,csa_tree_add_190_195_groupi_n_12445);
  or csa_tree_add_190_195_groupi_g36436(csa_tree_add_190_195_groupi_n_12465 ,csa_tree_add_190_195_groupi_n_12296 ,csa_tree_add_190_195_groupi_n_12422);
  nor csa_tree_add_190_195_groupi_g36437(csa_tree_add_190_195_groupi_n_12464 ,csa_tree_add_190_195_groupi_n_12297 ,csa_tree_add_190_195_groupi_n_12423);
  or csa_tree_add_190_195_groupi_g36438(csa_tree_add_190_195_groupi_n_12463 ,csa_tree_add_190_195_groupi_n_12426 ,csa_tree_add_190_195_groupi_n_12346);
  and csa_tree_add_190_195_groupi_g36439(csa_tree_add_190_195_groupi_n_12479 ,csa_tree_add_190_195_groupi_n_12366 ,csa_tree_add_190_195_groupi_n_12421);
  or csa_tree_add_190_195_groupi_g36440(csa_tree_add_190_195_groupi_n_12477 ,csa_tree_add_190_195_groupi_n_12305 ,csa_tree_add_190_195_groupi_n_12431);
  and csa_tree_add_190_195_groupi_g36441(csa_tree_add_190_195_groupi_n_12475 ,csa_tree_add_190_195_groupi_n_12435 ,csa_tree_add_190_195_groupi_n_12402);
  not csa_tree_add_190_195_groupi_g36442(csa_tree_add_190_195_groupi_n_12459 ,csa_tree_add_190_195_groupi_n_12458);
  not csa_tree_add_190_195_groupi_g36444(csa_tree_add_190_195_groupi_n_12456 ,csa_tree_add_190_195_groupi_n_12455);
  or csa_tree_add_190_195_groupi_g36445(csa_tree_add_190_195_groupi_n_12453 ,csa_tree_add_190_195_groupi_n_12382 ,csa_tree_add_190_195_groupi_n_12429);
  or csa_tree_add_190_195_groupi_g36446(csa_tree_add_190_195_groupi_n_12452 ,csa_tree_add_190_195_groupi_n_12417 ,csa_tree_add_190_195_groupi_n_12428);
  and csa_tree_add_190_195_groupi_g36447(csa_tree_add_190_195_groupi_n_12451 ,csa_tree_add_190_195_groupi_n_12426 ,csa_tree_add_190_195_groupi_n_12346);
  xnor csa_tree_add_190_195_groupi_g36448(csa_tree_add_190_195_groupi_n_12450 ,csa_tree_add_190_195_groupi_n_12352 ,csa_tree_add_190_195_groupi_n_12409);
  xnor csa_tree_add_190_195_groupi_g36449(csa_tree_add_190_195_groupi_n_12449 ,csa_tree_add_190_195_groupi_n_12369 ,csa_tree_add_190_195_groupi_n_12386);
  xnor csa_tree_add_190_195_groupi_g36450(csa_tree_add_190_195_groupi_n_12448 ,csa_tree_add_190_195_groupi_n_12341 ,csa_tree_add_190_195_groupi_n_12411);
  xnor csa_tree_add_190_195_groupi_g36451(csa_tree_add_190_195_groupi_n_12447 ,csa_tree_add_190_195_groupi_n_12325 ,csa_tree_add_190_195_groupi_n_12390);
  xnor csa_tree_add_190_195_groupi_g36452(csa_tree_add_190_195_groupi_n_12446 ,csa_tree_add_190_195_groupi_n_12297 ,csa_tree_add_190_195_groupi_n_12412);
  xnor csa_tree_add_190_195_groupi_g36453(csa_tree_add_190_195_groupi_n_12462 ,csa_tree_add_190_195_groupi_n_12393 ,csa_tree_add_190_195_groupi_n_177);
  xnor csa_tree_add_190_195_groupi_g36454(csa_tree_add_190_195_groupi_n_12461 ,csa_tree_add_190_195_groupi_n_12326 ,csa_tree_add_190_195_groupi_n_12379);
  xnor csa_tree_add_190_195_groupi_g36455(csa_tree_add_190_195_groupi_n_12460 ,csa_tree_add_190_195_groupi_n_12373 ,csa_tree_add_190_195_groupi_n_12377);
  xnor csa_tree_add_190_195_groupi_g36456(csa_tree_add_190_195_groupi_n_12458 ,csa_tree_add_190_195_groupi_n_12395 ,csa_tree_add_190_195_groupi_n_12330);
  and csa_tree_add_190_195_groupi_g36457(csa_tree_add_190_195_groupi_n_12457 ,csa_tree_add_190_195_groupi_n_12436 ,csa_tree_add_190_195_groupi_n_12400);
  xnor csa_tree_add_190_195_groupi_g36458(csa_tree_add_190_195_groupi_n_12455 ,csa_tree_add_190_195_groupi_n_12372 ,csa_tree_add_190_195_groupi_n_12380);
  xnor csa_tree_add_190_195_groupi_g36459(csa_tree_add_190_195_groupi_n_12454 ,csa_tree_add_190_195_groupi_n_12374 ,csa_tree_add_190_195_groupi_n_12376);
  not csa_tree_add_190_195_groupi_g36460(csa_tree_add_190_195_groupi_n_12442 ,csa_tree_add_190_195_groupi_n_12441);
  not csa_tree_add_190_195_groupi_g36461(csa_tree_add_190_195_groupi_n_12439 ,csa_tree_add_190_195_groupi_n_12440);
  not csa_tree_add_190_195_groupi_g36462(csa_tree_add_190_195_groupi_n_12437 ,csa_tree_add_190_195_groupi_n_12438);
  or csa_tree_add_190_195_groupi_g36463(csa_tree_add_190_195_groupi_n_12436 ,csa_tree_add_190_195_groupi_n_12413 ,csa_tree_add_190_195_groupi_n_12396);
  or csa_tree_add_190_195_groupi_g36464(csa_tree_add_190_195_groupi_n_12435 ,csa_tree_add_190_195_groupi_n_12392 ,csa_tree_add_190_195_groupi_n_12403);
  nor csa_tree_add_190_195_groupi_g36465(csa_tree_add_190_195_groupi_n_12434 ,csa_tree_add_190_195_groupi_n_12341 ,csa_tree_add_190_195_groupi_n_12411);
  or csa_tree_add_190_195_groupi_g36466(csa_tree_add_190_195_groupi_n_12433 ,csa_tree_add_190_195_groupi_n_12324 ,csa_tree_add_190_195_groupi_n_12389);
  nor csa_tree_add_190_195_groupi_g36467(csa_tree_add_190_195_groupi_n_12432 ,csa_tree_add_190_195_groupi_n_12325 ,csa_tree_add_190_195_groupi_n_12390);
  nor csa_tree_add_190_195_groupi_g36468(csa_tree_add_190_195_groupi_n_12431 ,csa_tree_add_190_195_groupi_n_12304 ,csa_tree_add_190_195_groupi_n_12395);
  or csa_tree_add_190_195_groupi_g36469(csa_tree_add_190_195_groupi_n_12430 ,csa_tree_add_190_195_groupi_n_12340 ,csa_tree_add_190_195_groupi_n_12410);
  and csa_tree_add_190_195_groupi_g36470(csa_tree_add_190_195_groupi_n_12445 ,csa_tree_add_190_195_groupi_n_12401 ,csa_tree_add_190_195_groupi_n_12306);
  and csa_tree_add_190_195_groupi_g36471(csa_tree_add_190_195_groupi_n_12444 ,csa_tree_add_190_195_groupi_n_12361 ,csa_tree_add_190_195_groupi_n_12399);
  or csa_tree_add_190_195_groupi_g36472(csa_tree_add_190_195_groupi_n_12443 ,csa_tree_add_190_195_groupi_n_12357 ,csa_tree_add_190_195_groupi_n_12405);
  or csa_tree_add_190_195_groupi_g36473(csa_tree_add_190_195_groupi_n_12441 ,csa_tree_add_190_195_groupi_n_12397 ,csa_tree_add_190_195_groupi_n_12337);
  or csa_tree_add_190_195_groupi_g36474(csa_tree_add_190_195_groupi_n_12440 ,csa_tree_add_190_195_groupi_n_12334 ,csa_tree_add_190_195_groupi_n_12404);
  or csa_tree_add_190_195_groupi_g36475(csa_tree_add_190_195_groupi_n_12438 ,csa_tree_add_190_195_groupi_n_12398 ,csa_tree_add_190_195_groupi_n_12358);
  not csa_tree_add_190_195_groupi_g36477(csa_tree_add_190_195_groupi_n_12428 ,csa_tree_add_190_195_groupi_n_12427);
  not csa_tree_add_190_195_groupi_g36478(csa_tree_add_190_195_groupi_n_12425 ,csa_tree_add_190_195_groupi_n_12424);
  not csa_tree_add_190_195_groupi_g36479(csa_tree_add_190_195_groupi_n_12423 ,csa_tree_add_190_195_groupi_n_12422);
  or csa_tree_add_190_195_groupi_g36481(csa_tree_add_190_195_groupi_n_12421 ,csa_tree_add_190_195_groupi_n_12336 ,csa_tree_add_190_195_groupi_n_12394);
  nor csa_tree_add_190_195_groupi_g36482(csa_tree_add_190_195_groupi_n_12420 ,csa_tree_add_190_195_groupi_n_12369 ,csa_tree_add_190_195_groupi_n_12386);
  or csa_tree_add_190_195_groupi_g36483(csa_tree_add_190_195_groupi_n_12419 ,csa_tree_add_190_195_groupi_n_12368 ,csa_tree_add_190_195_groupi_n_12385);
  or csa_tree_add_190_195_groupi_g36484(csa_tree_add_190_195_groupi_n_12418 ,csa_tree_add_190_195_groupi_n_12351 ,csa_tree_add_190_195_groupi_n_12408);
  nor csa_tree_add_190_195_groupi_g36485(csa_tree_add_190_195_groupi_n_12417 ,csa_tree_add_190_195_groupi_n_12352 ,csa_tree_add_190_195_groupi_n_12409);
  xnor csa_tree_add_190_195_groupi_g36486(csa_tree_add_190_195_groupi_n_12416 ,csa_tree_add_190_195_groupi_n_12348 ,csa_tree_add_190_195_groupi_n_12291);
  xnor csa_tree_add_190_195_groupi_g36487(csa_tree_add_190_195_groupi_n_12415 ,csa_tree_add_190_195_groupi_n_12371 ,csa_tree_add_190_195_groupi_n_12275);
  xnor csa_tree_add_190_195_groupi_g36488(csa_tree_add_190_195_groupi_n_12414 ,csa_tree_add_190_195_groupi_n_12269 ,csa_tree_add_190_195_groupi_n_12350);
  and csa_tree_add_190_195_groupi_g36489(csa_tree_add_190_195_groupi_n_12429 ,csa_tree_add_190_195_groupi_n_12285 ,csa_tree_add_190_195_groupi_n_12383);
  xnor csa_tree_add_190_195_groupi_g36490(csa_tree_add_190_195_groupi_n_12427 ,csa_tree_add_190_195_groupi_n_12276 ,csa_tree_add_190_195_groupi_n_12327);
  xnor csa_tree_add_190_195_groupi_g36491(csa_tree_add_190_195_groupi_n_12426 ,csa_tree_add_190_195_groupi_n_12375 ,csa_tree_add_190_195_groupi_n_12328);
  xnor csa_tree_add_190_195_groupi_g36492(csa_tree_add_190_195_groupi_n_12424 ,csa_tree_add_190_195_groupi_n_12298 ,csa_tree_add_190_195_groupi_n_12331);
  xnor csa_tree_add_190_195_groupi_g36493(csa_tree_add_190_195_groupi_n_12422 ,csa_tree_add_190_195_groupi_n_12243 ,csa_tree_add_190_195_groupi_n_12329);
  not csa_tree_add_190_195_groupi_g36494(csa_tree_add_190_195_groupi_n_12411 ,csa_tree_add_190_195_groupi_n_12410);
  not csa_tree_add_190_195_groupi_g36495(csa_tree_add_190_195_groupi_n_12409 ,csa_tree_add_190_195_groupi_n_12408);
  not csa_tree_add_190_195_groupi_g36496(csa_tree_add_190_195_groupi_n_12406 ,csa_tree_add_190_195_groupi_n_12407);
  nor csa_tree_add_190_195_groupi_g36497(csa_tree_add_190_195_groupi_n_12405 ,csa_tree_add_190_195_groupi_n_12356 ,csa_tree_add_190_195_groupi_n_12373);
  nor csa_tree_add_190_195_groupi_g36498(csa_tree_add_190_195_groupi_n_12404 ,csa_tree_add_190_195_groupi_n_12339 ,csa_tree_add_190_195_groupi_n_12190);
  nor csa_tree_add_190_195_groupi_g36499(csa_tree_add_190_195_groupi_n_12403 ,csa_tree_add_190_195_groupi_n_12370 ,csa_tree_add_190_195_groupi_n_12275);
  or csa_tree_add_190_195_groupi_g36500(csa_tree_add_190_195_groupi_n_12402 ,csa_tree_add_190_195_groupi_n_12371 ,csa_tree_add_190_195_groupi_n_12274);
  or csa_tree_add_190_195_groupi_g36501(csa_tree_add_190_195_groupi_n_12401 ,csa_tree_add_190_195_groupi_n_12375 ,csa_tree_add_190_195_groupi_n_12312);
  or csa_tree_add_190_195_groupi_g36502(csa_tree_add_190_195_groupi_n_12400 ,csa_tree_add_190_195_groupi_n_12268 ,csa_tree_add_190_195_groupi_n_12349);
  or csa_tree_add_190_195_groupi_g36503(csa_tree_add_190_195_groupi_n_12399 ,csa_tree_add_190_195_groupi_n_12360 ,csa_tree_add_190_195_groupi_n_12326);
  and csa_tree_add_190_195_groupi_g36504(csa_tree_add_190_195_groupi_n_12398 ,csa_tree_add_190_195_groupi_n_12372 ,csa_tree_add_190_195_groupi_n_12359);
  nor csa_tree_add_190_195_groupi_g36505(csa_tree_add_190_195_groupi_n_12397 ,csa_tree_add_190_195_groupi_n_12374 ,csa_tree_add_190_195_groupi_n_12338);
  nor csa_tree_add_190_195_groupi_g36506(csa_tree_add_190_195_groupi_n_12396 ,csa_tree_add_190_195_groupi_n_12269 ,csa_tree_add_190_195_groupi_n_12350);
  and csa_tree_add_190_195_groupi_g36507(csa_tree_add_190_195_groupi_n_12413 ,csa_tree_add_190_195_groupi_n_12365 ,csa_tree_add_190_195_groupi_n_12264);
  and csa_tree_add_190_195_groupi_g36508(csa_tree_add_190_195_groupi_n_12412 ,csa_tree_add_190_195_groupi_n_12367 ,csa_tree_add_190_195_groupi_n_12206);
  and csa_tree_add_190_195_groupi_g36509(csa_tree_add_190_195_groupi_n_12410 ,csa_tree_add_190_195_groupi_n_12315 ,csa_tree_add_190_195_groupi_n_12355);
  and csa_tree_add_190_195_groupi_g36510(csa_tree_add_190_195_groupi_n_12408 ,csa_tree_add_190_195_groupi_n_12308 ,csa_tree_add_190_195_groupi_n_12364);
  and csa_tree_add_190_195_groupi_g36511(csa_tree_add_190_195_groupi_n_12407 ,csa_tree_add_190_195_groupi_n_12362 ,csa_tree_add_190_195_groupi_n_12314);
  not csa_tree_add_190_195_groupi_g36512(csa_tree_add_190_195_groupi_n_12394 ,csa_tree_add_190_195_groupi_n_12393);
  not csa_tree_add_190_195_groupi_g36513(csa_tree_add_190_195_groupi_n_12392 ,csa_tree_add_190_195_groupi_n_12391);
  not csa_tree_add_190_195_groupi_g36514(csa_tree_add_190_195_groupi_n_12390 ,csa_tree_add_190_195_groupi_n_12389);
  not csa_tree_add_190_195_groupi_g36515(csa_tree_add_190_195_groupi_n_12388 ,csa_tree_add_190_195_groupi_n_12387);
  not csa_tree_add_190_195_groupi_g36516(csa_tree_add_190_195_groupi_n_12386 ,csa_tree_add_190_195_groupi_n_12385);
  or csa_tree_add_190_195_groupi_g36517(csa_tree_add_190_195_groupi_n_12384 ,csa_tree_add_190_195_groupi_n_12347 ,csa_tree_add_190_195_groupi_n_12290);
  or csa_tree_add_190_195_groupi_g36518(csa_tree_add_190_195_groupi_n_12383 ,csa_tree_add_190_195_groupi_n_12286 ,csa_tree_add_190_195_groupi_n_12353);
  nor csa_tree_add_190_195_groupi_g36519(csa_tree_add_190_195_groupi_n_12382 ,csa_tree_add_190_195_groupi_n_12348 ,csa_tree_add_190_195_groupi_n_12291);
  xnor csa_tree_add_190_195_groupi_g36520(out1[7] ,csa_tree_add_190_195_groupi_n_12247 ,csa_tree_add_190_195_groupi_n_12282);
  xnor csa_tree_add_190_195_groupi_g36522(csa_tree_add_190_195_groupi_n_12380 ,csa_tree_add_190_195_groupi_n_12233 ,csa_tree_add_190_195_groupi_n_12289);
  xnor csa_tree_add_190_195_groupi_g36523(csa_tree_add_190_195_groupi_n_12379 ,csa_tree_add_190_195_groupi_n_12293 ,csa_tree_add_190_195_groupi_n_12271);
  xnor csa_tree_add_190_195_groupi_g36524(csa_tree_add_190_195_groupi_n_12378 ,csa_tree_add_190_195_groupi_n_12237 ,csa_tree_add_190_195_groupi_n_12323);
  xnor csa_tree_add_190_195_groupi_g36525(csa_tree_add_190_195_groupi_n_12377 ,csa_tree_add_190_195_groupi_n_12189 ,csa_tree_add_190_195_groupi_n_12299);
  xnor csa_tree_add_190_195_groupi_g36526(csa_tree_add_190_195_groupi_n_12376 ,csa_tree_add_190_195_groupi_n_12188 ,csa_tree_add_190_195_groupi_n_12294);
  xnor csa_tree_add_190_195_groupi_g36527(csa_tree_add_190_195_groupi_n_12395 ,csa_tree_add_190_195_groupi_n_12218 ,csa_tree_add_190_195_groupi_n_12280);
  or csa_tree_add_190_195_groupi_g36528(csa_tree_add_190_195_groupi_n_12393 ,csa_tree_add_190_195_groupi_n_12321 ,csa_tree_add_190_195_groupi_n_12335);
  xnor csa_tree_add_190_195_groupi_g36529(csa_tree_add_190_195_groupi_n_12391 ,csa_tree_add_190_195_groupi_n_12303 ,csa_tree_add_190_195_groupi_n_12220);
  xnor csa_tree_add_190_195_groupi_g36530(csa_tree_add_190_195_groupi_n_12389 ,csa_tree_add_190_195_groupi_n_12301 ,csa_tree_add_190_195_groupi_n_12278);
  xnor csa_tree_add_190_195_groupi_g36531(csa_tree_add_190_195_groupi_n_12387 ,csa_tree_add_190_195_groupi_n_12191 ,csa_tree_add_190_195_groupi_n_12279);
  xnor csa_tree_add_190_195_groupi_g36532(csa_tree_add_190_195_groupi_n_12385 ,csa_tree_add_190_195_groupi_n_12244 ,csa_tree_add_190_195_groupi_n_12281);
  not csa_tree_add_190_195_groupi_g36533(csa_tree_add_190_195_groupi_n_12370 ,csa_tree_add_190_195_groupi_n_12371);
  not csa_tree_add_190_195_groupi_g36534(csa_tree_add_190_195_groupi_n_12368 ,csa_tree_add_190_195_groupi_n_12369);
  or csa_tree_add_190_195_groupi_g36535(csa_tree_add_190_195_groupi_n_12367 ,csa_tree_add_190_195_groupi_n_12303 ,csa_tree_add_190_195_groupi_n_12207);
  or csa_tree_add_190_195_groupi_g36536(csa_tree_add_190_195_groupi_n_12366 ,csa_tree_add_190_195_groupi_n_12300 ,csa_tree_add_190_195_groupi_n_12273);
  or csa_tree_add_190_195_groupi_g36537(csa_tree_add_190_195_groupi_n_12365 ,csa_tree_add_190_195_groupi_n_12302 ,csa_tree_add_190_195_groupi_n_12263);
  or csa_tree_add_190_195_groupi_g36538(csa_tree_add_190_195_groupi_n_12364 ,csa_tree_add_190_195_groupi_n_12277 ,csa_tree_add_190_195_groupi_n_12307);
  or csa_tree_add_190_195_groupi_g36539(csa_tree_add_190_195_groupi_n_12363 ,csa_tree_add_190_195_groupi_n_12237 ,csa_tree_add_190_195_groupi_n_12322);
  or csa_tree_add_190_195_groupi_g36540(csa_tree_add_190_195_groupi_n_12362 ,csa_tree_add_190_195_groupi_n_12217 ,csa_tree_add_190_195_groupi_n_12311);
  or csa_tree_add_190_195_groupi_g36541(csa_tree_add_190_195_groupi_n_12361 ,csa_tree_add_190_195_groupi_n_12292 ,csa_tree_add_190_195_groupi_n_12270);
  nor csa_tree_add_190_195_groupi_g36542(csa_tree_add_190_195_groupi_n_12360 ,csa_tree_add_190_195_groupi_n_12293 ,csa_tree_add_190_195_groupi_n_12271);
  or csa_tree_add_190_195_groupi_g36543(csa_tree_add_190_195_groupi_n_12359 ,csa_tree_add_190_195_groupi_n_12232 ,csa_tree_add_190_195_groupi_n_12289);
  nor csa_tree_add_190_195_groupi_g36544(csa_tree_add_190_195_groupi_n_12358 ,csa_tree_add_190_195_groupi_n_12233 ,csa_tree_add_190_195_groupi_n_12288);
  and csa_tree_add_190_195_groupi_g36545(csa_tree_add_190_195_groupi_n_12357 ,csa_tree_add_190_195_groupi_n_12189 ,csa_tree_add_190_195_groupi_n_12299);
  nor csa_tree_add_190_195_groupi_g36546(csa_tree_add_190_195_groupi_n_12356 ,csa_tree_add_190_195_groupi_n_12189 ,csa_tree_add_190_195_groupi_n_12299);
  or csa_tree_add_190_195_groupi_g36547(csa_tree_add_190_195_groupi_n_12355 ,csa_tree_add_190_195_groupi_n_12313 ,csa_tree_add_190_195_groupi_n_12276);
  nor csa_tree_add_190_195_groupi_g36548(csa_tree_add_190_195_groupi_n_12354 ,csa_tree_add_190_195_groupi_n_12236 ,csa_tree_add_190_195_groupi_n_12323);
  and csa_tree_add_190_195_groupi_g36549(csa_tree_add_190_195_groupi_n_12375 ,csa_tree_add_190_195_groupi_n_12254 ,csa_tree_add_190_195_groupi_n_12309);
  and csa_tree_add_190_195_groupi_g36550(csa_tree_add_190_195_groupi_n_12374 ,csa_tree_add_190_195_groupi_n_12258 ,csa_tree_add_190_195_groupi_n_12310);
  and csa_tree_add_190_195_groupi_g36551(csa_tree_add_190_195_groupi_n_12373 ,csa_tree_add_190_195_groupi_n_12259 ,csa_tree_add_190_195_groupi_n_12316);
  or csa_tree_add_190_195_groupi_g36552(csa_tree_add_190_195_groupi_n_12372 ,csa_tree_add_190_195_groupi_n_12320 ,csa_tree_add_190_195_groupi_n_12230);
  and csa_tree_add_190_195_groupi_g36553(csa_tree_add_190_195_groupi_n_12371 ,csa_tree_add_190_195_groupi_n_12317 ,csa_tree_add_190_195_groupi_n_12253);
  or csa_tree_add_190_195_groupi_g36554(csa_tree_add_190_195_groupi_n_12369 ,csa_tree_add_190_195_groupi_n_12319 ,csa_tree_add_190_195_groupi_n_12202);
  not csa_tree_add_190_195_groupi_g36556(csa_tree_add_190_195_groupi_n_12352 ,csa_tree_add_190_195_groupi_n_12351);
  not csa_tree_add_190_195_groupi_g36557(csa_tree_add_190_195_groupi_n_12350 ,csa_tree_add_190_195_groupi_n_12349);
  not csa_tree_add_190_195_groupi_g36558(csa_tree_add_190_195_groupi_n_12348 ,csa_tree_add_190_195_groupi_n_12347);
  not csa_tree_add_190_195_groupi_g36559(csa_tree_add_190_195_groupi_n_12346 ,csa_tree_add_190_195_groupi_n_12345);
  not csa_tree_add_190_195_groupi_g36560(csa_tree_add_190_195_groupi_n_12344 ,csa_tree_add_190_195_groupi_n_12343);
  not csa_tree_add_190_195_groupi_g36561(csa_tree_add_190_195_groupi_n_12341 ,csa_tree_add_190_195_groupi_n_12340);
  and csa_tree_add_190_195_groupi_g36562(csa_tree_add_190_195_groupi_n_12339 ,csa_tree_add_190_195_groupi_n_12245 ,csa_tree_add_190_195_groupi_n_12298);
  nor csa_tree_add_190_195_groupi_g36563(csa_tree_add_190_195_groupi_n_12338 ,csa_tree_add_190_195_groupi_n_12188 ,csa_tree_add_190_195_groupi_n_12294);
  and csa_tree_add_190_195_groupi_g36564(csa_tree_add_190_195_groupi_n_12337 ,csa_tree_add_190_195_groupi_n_12188 ,csa_tree_add_190_195_groupi_n_12294);
  and csa_tree_add_190_195_groupi_g36565(csa_tree_add_190_195_groupi_n_12336 ,csa_tree_add_190_195_groupi_n_12300 ,csa_tree_add_190_195_groupi_n_12273);
  nor csa_tree_add_190_195_groupi_g36566(csa_tree_add_190_195_groupi_n_12335 ,csa_tree_add_190_195_groupi_n_12127 ,csa_tree_add_190_195_groupi_n_12284);
  nor csa_tree_add_190_195_groupi_g36567(csa_tree_add_190_195_groupi_n_12334 ,csa_tree_add_190_195_groupi_n_12245 ,csa_tree_add_190_195_groupi_n_12298);
  xnor csa_tree_add_190_195_groupi_g36568(csa_tree_add_190_195_groupi_n_12333 ,csa_tree_add_190_195_groupi_n_12239 ,csa_tree_add_190_195_groupi_n_12156);
  xnor csa_tree_add_190_195_groupi_g36569(csa_tree_add_190_195_groupi_n_12332 ,csa_tree_add_190_195_groupi_n_12267 ,csa_tree_add_190_195_groupi_n_11630);
  xnor csa_tree_add_190_195_groupi_g36570(csa_tree_add_190_195_groupi_n_12331 ,csa_tree_add_190_195_groupi_n_12190 ,csa_tree_add_190_195_groupi_n_12245);
  xnor csa_tree_add_190_195_groupi_g36571(csa_tree_add_190_195_groupi_n_12330 ,csa_tree_add_190_195_groupi_n_12272 ,csa_tree_add_190_195_groupi_n_12246);
  xnor csa_tree_add_190_195_groupi_g36572(csa_tree_add_190_195_groupi_n_12329 ,csa_tree_add_190_195_groupi_n_12078 ,csa_tree_add_190_195_groupi_n_12277);
  xnor csa_tree_add_190_195_groupi_g36573(csa_tree_add_190_195_groupi_n_12328 ,csa_tree_add_190_195_groupi_n_12241 ,csa_tree_add_190_195_groupi_n_12266);
  xnor csa_tree_add_190_195_groupi_g36574(csa_tree_add_190_195_groupi_n_12327 ,csa_tree_add_190_195_groupi_n_12211 ,csa_tree_add_190_195_groupi_n_12235);
  and csa_tree_add_190_195_groupi_g36575(csa_tree_add_190_195_groupi_n_12353 ,csa_tree_add_190_195_groupi_n_12287 ,csa_tree_add_190_195_groupi_n_12228);
  xnor csa_tree_add_190_195_groupi_g36576(csa_tree_add_190_195_groupi_n_12351 ,csa_tree_add_190_195_groupi_n_12187 ,csa_tree_add_190_195_groupi_n_12221);
  xnor csa_tree_add_190_195_groupi_g36577(csa_tree_add_190_195_groupi_n_12349 ,csa_tree_add_190_195_groupi_n_12179 ,csa_tree_add_190_195_groupi_n_12225);
  xnor csa_tree_add_190_195_groupi_g36578(csa_tree_add_190_195_groupi_n_12347 ,csa_tree_add_190_195_groupi_n_12249 ,csa_tree_add_190_195_groupi_n_12223);
  xnor csa_tree_add_190_195_groupi_g36579(csa_tree_add_190_195_groupi_n_12345 ,csa_tree_add_190_195_groupi_n_12214 ,csa_tree_add_190_195_groupi_n_12222);
  xnor csa_tree_add_190_195_groupi_g36580(csa_tree_add_190_195_groupi_n_12343 ,csa_tree_add_190_195_groupi_n_12242 ,csa_tree_add_190_195_groupi_n_12224);
  xnor csa_tree_add_190_195_groupi_g36581(csa_tree_add_190_195_groupi_n_12342 ,csa_tree_add_190_195_groupi_n_12181 ,csa_tree_add_190_195_groupi_n_12227);
  xnor csa_tree_add_190_195_groupi_g36582(csa_tree_add_190_195_groupi_n_12340 ,csa_tree_add_190_195_groupi_n_12216 ,csa_tree_add_190_195_groupi_n_12226);
  not csa_tree_add_190_195_groupi_g36583(csa_tree_add_190_195_groupi_n_12325 ,csa_tree_add_190_195_groupi_n_12324);
  not csa_tree_add_190_195_groupi_g36584(csa_tree_add_190_195_groupi_n_12323 ,csa_tree_add_190_195_groupi_n_12322);
  nor csa_tree_add_190_195_groupi_g36585(csa_tree_add_190_195_groupi_n_12321 ,csa_tree_add_190_195_groupi_n_12119 ,csa_tree_add_190_195_groupi_n_12242);
  and csa_tree_add_190_195_groupi_g36586(csa_tree_add_190_195_groupi_n_12320 ,csa_tree_add_190_195_groupi_n_12229 ,csa_tree_add_190_195_groupi_n_12161);
  and csa_tree_add_190_195_groupi_g36587(csa_tree_add_190_195_groupi_n_12319 ,csa_tree_add_190_195_groupi_n_12249 ,csa_tree_add_190_195_groupi_n_12203);
  or csa_tree_add_190_195_groupi_g36588(csa_tree_add_190_195_groupi_n_12318 ,csa_tree_add_190_195_groupi_n_12267 ,csa_tree_add_190_195_groupi_n_11631);
  or csa_tree_add_190_195_groupi_g36589(csa_tree_add_190_195_groupi_n_12317 ,csa_tree_add_190_195_groupi_n_12218 ,csa_tree_add_190_195_groupi_n_12252);
  or csa_tree_add_190_195_groupi_g36590(csa_tree_add_190_195_groupi_n_12316 ,csa_tree_add_190_195_groupi_n_12088 ,csa_tree_add_190_195_groupi_n_12257);
  or csa_tree_add_190_195_groupi_g36591(csa_tree_add_190_195_groupi_n_12315 ,csa_tree_add_190_195_groupi_n_12211 ,csa_tree_add_190_195_groupi_n_12234);
  or csa_tree_add_190_195_groupi_g36592(csa_tree_add_190_195_groupi_n_12314 ,csa_tree_add_190_195_groupi_n_174 ,csa_tree_add_190_195_groupi_n_12122);
  nor csa_tree_add_190_195_groupi_g36593(csa_tree_add_190_195_groupi_n_12313 ,csa_tree_add_190_195_groupi_n_12210 ,csa_tree_add_190_195_groupi_n_12235);
  nor csa_tree_add_190_195_groupi_g36594(csa_tree_add_190_195_groupi_n_12312 ,csa_tree_add_190_195_groupi_n_12241 ,csa_tree_add_190_195_groupi_n_12266);
  nor csa_tree_add_190_195_groupi_g36595(csa_tree_add_190_195_groupi_n_12311 ,csa_tree_add_190_195_groupi_n_12244 ,csa_tree_add_190_195_groupi_n_12123);
  or csa_tree_add_190_195_groupi_g36596(csa_tree_add_190_195_groupi_n_12310 ,csa_tree_add_190_195_groupi_n_12162 ,csa_tree_add_190_195_groupi_n_12256);
  or csa_tree_add_190_195_groupi_g36597(csa_tree_add_190_195_groupi_n_12309 ,csa_tree_add_190_195_groupi_n_12250 ,csa_tree_add_190_195_groupi_n_12191);
  or csa_tree_add_190_195_groupi_g36598(csa_tree_add_190_195_groupi_n_12308 ,csa_tree_add_190_195_groupi_n_12243 ,csa_tree_add_190_195_groupi_n_12078);
  and csa_tree_add_190_195_groupi_g36599(csa_tree_add_190_195_groupi_n_12307 ,csa_tree_add_190_195_groupi_n_12243 ,csa_tree_add_190_195_groupi_n_12078);
  or csa_tree_add_190_195_groupi_g36600(csa_tree_add_190_195_groupi_n_12306 ,csa_tree_add_190_195_groupi_n_12240 ,csa_tree_add_190_195_groupi_n_12265);
  and csa_tree_add_190_195_groupi_g36601(csa_tree_add_190_195_groupi_n_12305 ,csa_tree_add_190_195_groupi_n_12272 ,csa_tree_add_190_195_groupi_n_12246);
  nor csa_tree_add_190_195_groupi_g36602(csa_tree_add_190_195_groupi_n_12304 ,csa_tree_add_190_195_groupi_n_12272 ,csa_tree_add_190_195_groupi_n_12246);
  and csa_tree_add_190_195_groupi_g36603(csa_tree_add_190_195_groupi_n_12326 ,csa_tree_add_190_195_groupi_n_12198 ,csa_tree_add_190_195_groupi_n_12260);
  and csa_tree_add_190_195_groupi_g36604(csa_tree_add_190_195_groupi_n_12324 ,csa_tree_add_190_195_groupi_n_12255 ,csa_tree_add_190_195_groupi_n_12194);
  and csa_tree_add_190_195_groupi_g36605(csa_tree_add_190_195_groupi_n_12322 ,csa_tree_add_190_195_groupi_n_12251 ,csa_tree_add_190_195_groupi_n_12135);
  not csa_tree_add_190_195_groupi_g36606(csa_tree_add_190_195_groupi_n_12302 ,csa_tree_add_190_195_groupi_n_12301);
  not csa_tree_add_190_195_groupi_g36607(csa_tree_add_190_195_groupi_n_12297 ,csa_tree_add_190_195_groupi_n_12296);
  not csa_tree_add_190_195_groupi_g36608(csa_tree_add_190_195_groupi_n_12295 ,csa_tree_add_190_195_groupi_n_176);
  not csa_tree_add_190_195_groupi_g36609(csa_tree_add_190_195_groupi_n_12293 ,csa_tree_add_190_195_groupi_n_12292);
  not csa_tree_add_190_195_groupi_g36610(csa_tree_add_190_195_groupi_n_12291 ,csa_tree_add_190_195_groupi_n_12290);
  not csa_tree_add_190_195_groupi_g36611(csa_tree_add_190_195_groupi_n_12289 ,csa_tree_add_190_195_groupi_n_12288);
  or csa_tree_add_190_195_groupi_g36612(csa_tree_add_190_195_groupi_n_12287 ,csa_tree_add_190_195_groupi_n_12262 ,csa_tree_add_190_195_groupi_n_12248);
  nor csa_tree_add_190_195_groupi_g36613(csa_tree_add_190_195_groupi_n_12286 ,csa_tree_add_190_195_groupi_n_12239 ,csa_tree_add_190_195_groupi_n_12156);
  or csa_tree_add_190_195_groupi_g36614(csa_tree_add_190_195_groupi_n_12285 ,csa_tree_add_190_195_groupi_n_12238 ,csa_tree_add_190_195_groupi_n_12155);
  and csa_tree_add_190_195_groupi_g36615(csa_tree_add_190_195_groupi_n_12284 ,csa_tree_add_190_195_groupi_n_12119 ,csa_tree_add_190_195_groupi_n_12242);
  and csa_tree_add_190_195_groupi_g36616(csa_tree_add_190_195_groupi_n_12283 ,csa_tree_add_190_195_groupi_n_12267 ,csa_tree_add_190_195_groupi_n_11631);
  xnor csa_tree_add_190_195_groupi_g36617(csa_tree_add_190_195_groupi_n_12282 ,csa_tree_add_190_195_groupi_n_12183 ,csa_tree_add_190_195_groupi_n_11936);
  xnor csa_tree_add_190_195_groupi_g36618(csa_tree_add_190_195_groupi_n_12281 ,csa_tree_add_190_195_groupi_n_12217 ,csa_tree_add_190_195_groupi_n_12123);
  xnor csa_tree_add_190_195_groupi_g36619(csa_tree_add_190_195_groupi_n_12280 ,csa_tree_add_190_195_groupi_n_12116 ,csa_tree_add_190_195_groupi_n_12185);
  xnor csa_tree_add_190_195_groupi_g36620(csa_tree_add_190_195_groupi_n_12279 ,csa_tree_add_190_195_groupi_n_12031 ,csa_tree_add_190_195_groupi_n_12209);
  xnor csa_tree_add_190_195_groupi_g36621(csa_tree_add_190_195_groupi_n_12278 ,csa_tree_add_190_195_groupi_n_12213 ,csa_tree_add_190_195_groupi_n_12114);
  xnor csa_tree_add_190_195_groupi_g36622(csa_tree_add_190_195_groupi_n_12303 ,csa_tree_add_190_195_groupi_n_12043 ,csa_tree_add_190_195_groupi_n_12168);
  xnor csa_tree_add_190_195_groupi_g36623(csa_tree_add_190_195_groupi_n_12301 ,csa_tree_add_190_195_groupi_n_12125 ,csa_tree_add_190_195_groupi_n_12169);
  xnor csa_tree_add_190_195_groupi_g36624(csa_tree_add_190_195_groupi_n_12300 ,csa_tree_add_190_195_groupi_n_12042 ,csa_tree_add_190_195_groupi_n_12167);
  xnor csa_tree_add_190_195_groupi_g36625(csa_tree_add_190_195_groupi_n_12299 ,csa_tree_add_190_195_groupi_n_12033 ,csa_tree_add_190_195_groupi_n_12171);
  xnor csa_tree_add_190_195_groupi_g36626(csa_tree_add_190_195_groupi_n_12298 ,csa_tree_add_190_195_groupi_n_12079 ,csa_tree_add_190_195_groupi_n_12166);
  xnor csa_tree_add_190_195_groupi_g36627(csa_tree_add_190_195_groupi_n_12296 ,csa_tree_add_190_195_groupi_n_12128 ,csa_tree_add_190_195_groupi_n_12170);
  xnor csa_tree_add_190_195_groupi_g36629(csa_tree_add_190_195_groupi_n_12294 ,csa_tree_add_190_195_groupi_n_11938 ,csa_tree_add_190_195_groupi_n_12165);
  xnor csa_tree_add_190_195_groupi_g36630(csa_tree_add_190_195_groupi_n_12292 ,csa_tree_add_190_195_groupi_n_12025 ,csa_tree_add_190_195_groupi_n_12172);
  and csa_tree_add_190_195_groupi_g36631(csa_tree_add_190_195_groupi_n_12290 ,csa_tree_add_190_195_groupi_n_12261 ,csa_tree_add_190_195_groupi_n_12176);
  xnor csa_tree_add_190_195_groupi_g36632(csa_tree_add_190_195_groupi_n_12288 ,csa_tree_add_190_195_groupi_n_12037 ,csa_tree_add_190_195_groupi_n_175);
  not csa_tree_add_190_195_groupi_g36633(csa_tree_add_190_195_groupi_n_12275 ,csa_tree_add_190_195_groupi_n_12274);
  not csa_tree_add_190_195_groupi_g36635(csa_tree_add_190_195_groupi_n_12271 ,csa_tree_add_190_195_groupi_n_12270);
  not csa_tree_add_190_195_groupi_g36636(csa_tree_add_190_195_groupi_n_12269 ,csa_tree_add_190_195_groupi_n_12268);
  not csa_tree_add_190_195_groupi_g36637(csa_tree_add_190_195_groupi_n_12266 ,csa_tree_add_190_195_groupi_n_12265);
  or csa_tree_add_190_195_groupi_g36638(csa_tree_add_190_195_groupi_n_12264 ,csa_tree_add_190_195_groupi_n_12212 ,csa_tree_add_190_195_groupi_n_12114);
  nor csa_tree_add_190_195_groupi_g36639(csa_tree_add_190_195_groupi_n_12263 ,csa_tree_add_190_195_groupi_n_12213 ,csa_tree_add_190_195_groupi_n_12113);
  nor csa_tree_add_190_195_groupi_g36640(csa_tree_add_190_195_groupi_n_12262 ,csa_tree_add_190_195_groupi_n_12183 ,csa_tree_add_190_195_groupi_n_11936);
  or csa_tree_add_190_195_groupi_g36641(csa_tree_add_190_195_groupi_n_12261 ,csa_tree_add_190_195_groupi_n_11871 ,csa_tree_add_190_195_groupi_n_12177);
  or csa_tree_add_190_195_groupi_g36642(csa_tree_add_190_195_groupi_n_12260 ,csa_tree_add_190_195_groupi_n_12216 ,csa_tree_add_190_195_groupi_n_12195);
  or csa_tree_add_190_195_groupi_g36643(csa_tree_add_190_195_groupi_n_12259 ,csa_tree_add_190_195_groupi_n_12186 ,csa_tree_add_190_195_groupi_n_12108);
  or csa_tree_add_190_195_groupi_g36644(csa_tree_add_190_195_groupi_n_12258 ,csa_tree_add_190_195_groupi_n_12110 ,csa_tree_add_190_195_groupi_n_12179);
  nor csa_tree_add_190_195_groupi_g36645(csa_tree_add_190_195_groupi_n_12257 ,csa_tree_add_190_195_groupi_n_12187 ,csa_tree_add_190_195_groupi_n_12109);
  and csa_tree_add_190_195_groupi_g36646(csa_tree_add_190_195_groupi_n_12256 ,csa_tree_add_190_195_groupi_n_12110 ,csa_tree_add_190_195_groupi_n_12179);
  or csa_tree_add_190_195_groupi_g36647(csa_tree_add_190_195_groupi_n_12255 ,csa_tree_add_190_195_groupi_n_12192 ,csa_tree_add_190_195_groupi_n_12215);
  or csa_tree_add_190_195_groupi_g36648(csa_tree_add_190_195_groupi_n_12254 ,csa_tree_add_190_195_groupi_n_12030 ,csa_tree_add_190_195_groupi_n_12208);
  or csa_tree_add_190_195_groupi_g36649(csa_tree_add_190_195_groupi_n_12253 ,csa_tree_add_190_195_groupi_n_12115 ,csa_tree_add_190_195_groupi_n_12184);
  nor csa_tree_add_190_195_groupi_g36650(csa_tree_add_190_195_groupi_n_12252 ,csa_tree_add_190_195_groupi_n_12116 ,csa_tree_add_190_195_groupi_n_12185);
  or csa_tree_add_190_195_groupi_g36651(csa_tree_add_190_195_groupi_n_12251 ,csa_tree_add_190_195_groupi_n_12219 ,csa_tree_add_190_195_groupi_n_12137);
  nor csa_tree_add_190_195_groupi_g36652(csa_tree_add_190_195_groupi_n_12250 ,csa_tree_add_190_195_groupi_n_12031 ,csa_tree_add_190_195_groupi_n_12209);
  and csa_tree_add_190_195_groupi_g36653(csa_tree_add_190_195_groupi_n_12277 ,csa_tree_add_190_195_groupi_n_12144 ,csa_tree_add_190_195_groupi_n_12201);
  and csa_tree_add_190_195_groupi_g36654(csa_tree_add_190_195_groupi_n_12276 ,csa_tree_add_190_195_groupi_n_12139 ,csa_tree_add_190_195_groupi_n_12196);
  and csa_tree_add_190_195_groupi_g36655(csa_tree_add_190_195_groupi_n_12274 ,csa_tree_add_190_195_groupi_n_12054 ,csa_tree_add_190_195_groupi_n_12205);
  and csa_tree_add_190_195_groupi_g36656(csa_tree_add_190_195_groupi_n_12273 ,csa_tree_add_190_195_groupi_n_12105 ,csa_tree_add_190_195_groupi_n_12173);
  or csa_tree_add_190_195_groupi_g36657(csa_tree_add_190_195_groupi_n_12272 ,csa_tree_add_190_195_groupi_n_12104 ,csa_tree_add_190_195_groupi_n_12174);
  and csa_tree_add_190_195_groupi_g36658(csa_tree_add_190_195_groupi_n_12270 ,csa_tree_add_190_195_groupi_n_12141 ,csa_tree_add_190_195_groupi_n_12199);
  and csa_tree_add_190_195_groupi_g36659(csa_tree_add_190_195_groupi_n_12268 ,csa_tree_add_190_195_groupi_n_12193 ,csa_tree_add_190_195_groupi_n_12134);
  and csa_tree_add_190_195_groupi_g36660(csa_tree_add_190_195_groupi_n_12267 ,csa_tree_add_190_195_groupi_n_12197 ,csa_tree_add_190_195_groupi_n_11793);
  and csa_tree_add_190_195_groupi_g36661(csa_tree_add_190_195_groupi_n_12265 ,csa_tree_add_190_195_groupi_n_12204 ,csa_tree_add_190_195_groupi_n_12150);
  not csa_tree_add_190_195_groupi_g36662(csa_tree_add_190_195_groupi_n_12248 ,csa_tree_add_190_195_groupi_n_12247);
  not csa_tree_add_190_195_groupi_g36663(csa_tree_add_190_195_groupi_n_12244 ,csa_tree_add_190_195_groupi_n_174);
  not csa_tree_add_190_195_groupi_g36664(csa_tree_add_190_195_groupi_n_12241 ,csa_tree_add_190_195_groupi_n_12240);
  not csa_tree_add_190_195_groupi_g36665(csa_tree_add_190_195_groupi_n_12239 ,csa_tree_add_190_195_groupi_n_12238);
  not csa_tree_add_190_195_groupi_g36666(csa_tree_add_190_195_groupi_n_12237 ,csa_tree_add_190_195_groupi_n_12236);
  not csa_tree_add_190_195_groupi_g36667(csa_tree_add_190_195_groupi_n_12235 ,csa_tree_add_190_195_groupi_n_12234);
  not csa_tree_add_190_195_groupi_g36668(csa_tree_add_190_195_groupi_n_12232 ,csa_tree_add_190_195_groupi_n_12233);
  xnor csa_tree_add_190_195_groupi_g36669(out1[6] ,csa_tree_add_190_195_groupi_n_12160 ,csa_tree_add_190_195_groupi_n_12098);
  nor csa_tree_add_190_195_groupi_g36670(csa_tree_add_190_195_groupi_n_12230 ,csa_tree_add_190_195_groupi_n_12181 ,csa_tree_add_190_195_groupi_n_12112);
  or csa_tree_add_190_195_groupi_g36671(csa_tree_add_190_195_groupi_n_12229 ,csa_tree_add_190_195_groupi_n_12180 ,csa_tree_add_190_195_groupi_n_12111);
  or csa_tree_add_190_195_groupi_g36672(csa_tree_add_190_195_groupi_n_12228 ,csa_tree_add_190_195_groupi_n_12182 ,csa_tree_add_190_195_groupi_n_11935);
  xnor csa_tree_add_190_195_groupi_g36673(csa_tree_add_190_195_groupi_n_12227 ,csa_tree_add_190_195_groupi_n_12112 ,csa_tree_add_190_195_groupi_n_12161);
  xnor csa_tree_add_190_195_groupi_g36674(csa_tree_add_190_195_groupi_n_12226 ,csa_tree_add_190_195_groupi_n_12107 ,csa_tree_add_190_195_groupi_n_12158);
  xnor csa_tree_add_190_195_groupi_g36675(csa_tree_add_190_195_groupi_n_12225 ,csa_tree_add_190_195_groupi_n_12110 ,csa_tree_add_190_195_groupi_n_12162);
  xnor csa_tree_add_190_195_groupi_g36676(csa_tree_add_190_195_groupi_n_12224 ,csa_tree_add_190_195_groupi_n_12119 ,csa_tree_add_190_195_groupi_n_12127);
  xnor csa_tree_add_190_195_groupi_g36677(csa_tree_add_190_195_groupi_n_12223 ,csa_tree_add_190_195_groupi_n_12035 ,csa_tree_add_190_195_groupi_n_12154);
  xnor csa_tree_add_190_195_groupi_g36678(csa_tree_add_190_195_groupi_n_12222 ,csa_tree_add_190_195_groupi_n_12041 ,csa_tree_add_190_195_groupi_n_12118);
  xnor csa_tree_add_190_195_groupi_g36679(csa_tree_add_190_195_groupi_n_12221 ,csa_tree_add_190_195_groupi_n_12109 ,csa_tree_add_190_195_groupi_n_12088);
  xnor csa_tree_add_190_195_groupi_g36680(csa_tree_add_190_195_groupi_n_12220 ,csa_tree_add_190_195_groupi_n_12152 ,csa_tree_add_190_195_groupi_n_12121);
  xnor csa_tree_add_190_195_groupi_g36681(csa_tree_add_190_195_groupi_n_12249 ,csa_tree_add_190_195_groupi_n_12003 ,csa_tree_add_190_195_groupi_n_12095);
  or csa_tree_add_190_195_groupi_g36682(csa_tree_add_190_195_groupi_n_12247 ,csa_tree_add_190_195_groupi_n_12019 ,csa_tree_add_190_195_groupi_n_12175);
  xnor csa_tree_add_190_195_groupi_g36683(csa_tree_add_190_195_groupi_n_12246 ,csa_tree_add_190_195_groupi_n_12163 ,csa_tree_add_190_195_groupi_n_12089);
  xnor csa_tree_add_190_195_groupi_g36684(csa_tree_add_190_195_groupi_n_12245 ,csa_tree_add_190_195_groupi_n_12087 ,csa_tree_add_190_195_groupi_n_12090);
  xnor csa_tree_add_190_195_groupi_g36686(csa_tree_add_190_195_groupi_n_12243 ,csa_tree_add_190_195_groupi_n_12050 ,csa_tree_add_190_195_groupi_n_12092);
  xnor csa_tree_add_190_195_groupi_g36687(csa_tree_add_190_195_groupi_n_12242 ,csa_tree_add_190_195_groupi_n_11950 ,csa_tree_add_190_195_groupi_n_12096);
  xnor csa_tree_add_190_195_groupi_g36688(csa_tree_add_190_195_groupi_n_12240 ,csa_tree_add_190_195_groupi_n_12084 ,csa_tree_add_190_195_groupi_n_12093);
  xnor csa_tree_add_190_195_groupi_g36689(csa_tree_add_190_195_groupi_n_12238 ,csa_tree_add_190_195_groupi_n_12124 ,csa_tree_add_190_195_groupi_n_12097);
  xnor csa_tree_add_190_195_groupi_g36690(csa_tree_add_190_195_groupi_n_12236 ,csa_tree_add_190_195_groupi_n_12159 ,csa_tree_add_190_195_groupi_n_11828);
  xnor csa_tree_add_190_195_groupi_g36691(csa_tree_add_190_195_groupi_n_12234 ,csa_tree_add_190_195_groupi_n_11914 ,csa_tree_add_190_195_groupi_n_12094);
  and csa_tree_add_190_195_groupi_g36692(csa_tree_add_190_195_groupi_n_12233 ,csa_tree_add_190_195_groupi_n_12099 ,csa_tree_add_190_195_groupi_n_12200);
  not csa_tree_add_190_195_groupi_g36694(csa_tree_add_190_195_groupi_n_12215 ,csa_tree_add_190_195_groupi_n_12214);
  not csa_tree_add_190_195_groupi_g36695(csa_tree_add_190_195_groupi_n_12212 ,csa_tree_add_190_195_groupi_n_12213);
  not csa_tree_add_190_195_groupi_g36696(csa_tree_add_190_195_groupi_n_12211 ,csa_tree_add_190_195_groupi_n_12210);
  not csa_tree_add_190_195_groupi_g36697(csa_tree_add_190_195_groupi_n_12209 ,csa_tree_add_190_195_groupi_n_12208);
  nor csa_tree_add_190_195_groupi_g36698(csa_tree_add_190_195_groupi_n_12207 ,csa_tree_add_190_195_groupi_n_12152 ,csa_tree_add_190_195_groupi_n_12120);
  or csa_tree_add_190_195_groupi_g36699(csa_tree_add_190_195_groupi_n_12206 ,csa_tree_add_190_195_groupi_n_12151 ,csa_tree_add_190_195_groupi_n_12121);
  or csa_tree_add_190_195_groupi_g36700(csa_tree_add_190_195_groupi_n_12205 ,csa_tree_add_190_195_groupi_n_12163 ,csa_tree_add_190_195_groupi_n_12052);
  or csa_tree_add_190_195_groupi_g36701(csa_tree_add_190_195_groupi_n_12204 ,csa_tree_add_190_195_groupi_n_12147 ,csa_tree_add_190_195_groupi_n_12083);
  or csa_tree_add_190_195_groupi_g36702(csa_tree_add_190_195_groupi_n_12203 ,csa_tree_add_190_195_groupi_n_12034 ,csa_tree_add_190_195_groupi_n_12154);
  nor csa_tree_add_190_195_groupi_g36703(csa_tree_add_190_195_groupi_n_12202 ,csa_tree_add_190_195_groupi_n_12035 ,csa_tree_add_190_195_groupi_n_12153);
  or csa_tree_add_190_195_groupi_g36704(csa_tree_add_190_195_groupi_n_12201 ,csa_tree_add_190_195_groupi_n_12145 ,csa_tree_add_190_195_groupi_n_12004);
  or csa_tree_add_190_195_groupi_g36705(csa_tree_add_190_195_groupi_n_12200 ,csa_tree_add_190_195_groupi_n_12051 ,csa_tree_add_190_195_groupi_n_12142);
  or csa_tree_add_190_195_groupi_g36706(csa_tree_add_190_195_groupi_n_12199 ,csa_tree_add_190_195_groupi_n_12082 ,csa_tree_add_190_195_groupi_n_12140);
  or csa_tree_add_190_195_groupi_g36707(csa_tree_add_190_195_groupi_n_12198 ,csa_tree_add_190_195_groupi_n_12106 ,csa_tree_add_190_195_groupi_n_12157);
  or csa_tree_add_190_195_groupi_g36708(csa_tree_add_190_195_groupi_n_12197 ,csa_tree_add_190_195_groupi_n_12159 ,csa_tree_add_190_195_groupi_n_11789);
  or csa_tree_add_190_195_groupi_g36709(csa_tree_add_190_195_groupi_n_12196 ,csa_tree_add_190_195_groupi_n_12138 ,csa_tree_add_190_195_groupi_n_12129);
  nor csa_tree_add_190_195_groupi_g36710(csa_tree_add_190_195_groupi_n_12195 ,csa_tree_add_190_195_groupi_n_12107 ,csa_tree_add_190_195_groupi_n_12158);
  or csa_tree_add_190_195_groupi_g36711(csa_tree_add_190_195_groupi_n_12194 ,csa_tree_add_190_195_groupi_n_12040 ,csa_tree_add_190_195_groupi_n_12117);
  or csa_tree_add_190_195_groupi_g36712(csa_tree_add_190_195_groupi_n_12193 ,csa_tree_add_190_195_groupi_n_12133 ,csa_tree_add_190_195_groupi_n_12126);
  nor csa_tree_add_190_195_groupi_g36713(csa_tree_add_190_195_groupi_n_12192 ,csa_tree_add_190_195_groupi_n_12041 ,csa_tree_add_190_195_groupi_n_12118);
  and csa_tree_add_190_195_groupi_g36714(csa_tree_add_190_195_groupi_n_12219 ,csa_tree_add_190_195_groupi_n_12146 ,csa_tree_add_190_195_groupi_n_12063);
  and csa_tree_add_190_195_groupi_g36715(csa_tree_add_190_195_groupi_n_12218 ,csa_tree_add_190_195_groupi_n_12056 ,csa_tree_add_190_195_groupi_n_12148);
  and csa_tree_add_190_195_groupi_g36716(csa_tree_add_190_195_groupi_n_12217 ,csa_tree_add_190_195_groupi_n_12143 ,csa_tree_add_190_195_groupi_n_12021);
  and csa_tree_add_190_195_groupi_g36717(csa_tree_add_190_195_groupi_n_12216 ,csa_tree_add_190_195_groupi_n_12136 ,csa_tree_add_190_195_groupi_n_12064);
  or csa_tree_add_190_195_groupi_g36718(csa_tree_add_190_195_groupi_n_12214 ,csa_tree_add_190_195_groupi_n_11978 ,csa_tree_add_190_195_groupi_n_12132);
  or csa_tree_add_190_195_groupi_g36719(csa_tree_add_190_195_groupi_n_12213 ,csa_tree_add_190_195_groupi_n_12015 ,csa_tree_add_190_195_groupi_n_12149);
  or csa_tree_add_190_195_groupi_g36720(csa_tree_add_190_195_groupi_n_12210 ,csa_tree_add_190_195_groupi_n_12061 ,csa_tree_add_190_195_groupi_n_12130);
  and csa_tree_add_190_195_groupi_g36721(csa_tree_add_190_195_groupi_n_12208 ,csa_tree_add_190_195_groupi_n_12131 ,csa_tree_add_190_195_groupi_n_12058);
  not csa_tree_add_190_195_groupi_g36722(csa_tree_add_190_195_groupi_n_12187 ,csa_tree_add_190_195_groupi_n_12186);
  not csa_tree_add_190_195_groupi_g36723(csa_tree_add_190_195_groupi_n_12185 ,csa_tree_add_190_195_groupi_n_12184);
  not csa_tree_add_190_195_groupi_g36724(csa_tree_add_190_195_groupi_n_12183 ,csa_tree_add_190_195_groupi_n_12182);
  not csa_tree_add_190_195_groupi_g36725(csa_tree_add_190_195_groupi_n_12181 ,csa_tree_add_190_195_groupi_n_12180);
  xnor csa_tree_add_190_195_groupi_g36726(out1[5] ,csa_tree_add_190_195_groupi_n_11869 ,csa_tree_add_190_195_groupi_n_12007);
  and csa_tree_add_190_195_groupi_g36727(csa_tree_add_190_195_groupi_n_12177 ,csa_tree_add_190_195_groupi_n_11945 ,csa_tree_add_190_195_groupi_n_12124);
  or csa_tree_add_190_195_groupi_g36728(csa_tree_add_190_195_groupi_n_12176 ,csa_tree_add_190_195_groupi_n_11945 ,csa_tree_add_190_195_groupi_n_12124);
  nor csa_tree_add_190_195_groupi_g36729(csa_tree_add_190_195_groupi_n_12175 ,csa_tree_add_190_195_groupi_n_12160 ,csa_tree_add_190_195_groupi_n_12018);
  and csa_tree_add_190_195_groupi_g36730(csa_tree_add_190_195_groupi_n_12174 ,csa_tree_add_190_195_groupi_n_12079 ,csa_tree_add_190_195_groupi_n_12102);
  or csa_tree_add_190_195_groupi_g36731(csa_tree_add_190_195_groupi_n_12173 ,csa_tree_add_190_195_groupi_n_12103 ,csa_tree_add_190_195_groupi_n_12081);
  xnor csa_tree_add_190_195_groupi_g36732(csa_tree_add_190_195_groupi_n_12172 ,csa_tree_add_190_195_groupi_n_12051 ,csa_tree_add_190_195_groupi_n_12046);
  xnor csa_tree_add_190_195_groupi_g36733(csa_tree_add_190_195_groupi_n_12171 ,csa_tree_add_190_195_groupi_n_11908 ,csa_tree_add_190_195_groupi_n_12082);
  xnor csa_tree_add_190_195_groupi_g36734(csa_tree_add_190_195_groupi_n_12170 ,csa_tree_add_190_195_groupi_n_12048 ,csa_tree_add_190_195_groupi_n_12077);
  xnor csa_tree_add_190_195_groupi_g36736(csa_tree_add_190_195_groupi_n_12169 ,csa_tree_add_190_195_groupi_n_12000 ,csa_tree_add_190_195_groupi_n_12027);
  xnor csa_tree_add_190_195_groupi_g36737(csa_tree_add_190_195_groupi_n_12168 ,csa_tree_add_190_195_groupi_n_12044 ,csa_tree_add_190_195_groupi_n_12004);
  xnor csa_tree_add_190_195_groupi_g36738(csa_tree_add_190_195_groupi_n_12167 ,csa_tree_add_190_195_groupi_n_12083 ,csa_tree_add_190_195_groupi_n_11909);
  xnor csa_tree_add_190_195_groupi_g36739(csa_tree_add_190_195_groupi_n_12166 ,csa_tree_add_190_195_groupi_n_11957 ,csa_tree_add_190_195_groupi_n_12039);
  xnor csa_tree_add_190_195_groupi_g36740(csa_tree_add_190_195_groupi_n_12165 ,csa_tree_add_190_195_groupi_n_12085 ,csa_tree_add_190_195_groupi_n_11758);
  xnor csa_tree_add_190_195_groupi_g36741(csa_tree_add_190_195_groupi_n_12164 ,csa_tree_add_190_195_groupi_n_12029 ,csa_tree_add_190_195_groupi_n_12075);
  xnor csa_tree_add_190_195_groupi_g36742(csa_tree_add_190_195_groupi_n_12191 ,csa_tree_add_190_195_groupi_n_12049 ,csa_tree_add_190_195_groupi_n_12011);
  and csa_tree_add_190_195_groupi_g36743(csa_tree_add_190_195_groupi_n_12190 ,csa_tree_add_190_195_groupi_n_12101 ,csa_tree_add_190_195_groupi_n_12023);
  xnor csa_tree_add_190_195_groupi_g36744(csa_tree_add_190_195_groupi_n_12189 ,csa_tree_add_190_195_groupi_n_11853 ,csa_tree_add_190_195_groupi_n_12010);
  or csa_tree_add_190_195_groupi_g36745(csa_tree_add_190_195_groupi_n_12188 ,csa_tree_add_190_195_groupi_n_12100 ,csa_tree_add_190_195_groupi_n_11976);
  xnor csa_tree_add_190_195_groupi_g36746(csa_tree_add_190_195_groupi_n_12186 ,csa_tree_add_190_195_groupi_n_11915 ,csa_tree_add_190_195_groupi_n_12013);
  xnor csa_tree_add_190_195_groupi_g36747(csa_tree_add_190_195_groupi_n_12184 ,csa_tree_add_190_195_groupi_n_11905 ,csa_tree_add_190_195_groupi_n_12014);
  xnor csa_tree_add_190_195_groupi_g36748(csa_tree_add_190_195_groupi_n_12182 ,csa_tree_add_190_195_groupi_n_11962 ,csa_tree_add_190_195_groupi_n_12009);
  xnor csa_tree_add_190_195_groupi_g36749(csa_tree_add_190_195_groupi_n_12180 ,csa_tree_add_190_195_groupi_n_11964 ,csa_tree_add_190_195_groupi_n_12008);
  xnor csa_tree_add_190_195_groupi_g36750(csa_tree_add_190_195_groupi_n_12179 ,csa_tree_add_190_195_groupi_n_12080 ,csa_tree_add_190_195_groupi_n_12012);
  not csa_tree_add_190_195_groupi_g36751(csa_tree_add_190_195_groupi_n_12157 ,csa_tree_add_190_195_groupi_n_12158);
  not csa_tree_add_190_195_groupi_g36752(csa_tree_add_190_195_groupi_n_12156 ,csa_tree_add_190_195_groupi_n_12155);
  not csa_tree_add_190_195_groupi_g36753(csa_tree_add_190_195_groupi_n_12153 ,csa_tree_add_190_195_groupi_n_12154);
  not csa_tree_add_190_195_groupi_g36754(csa_tree_add_190_195_groupi_n_12151 ,csa_tree_add_190_195_groupi_n_12152);
  or csa_tree_add_190_195_groupi_g36755(csa_tree_add_190_195_groupi_n_12150 ,csa_tree_add_190_195_groupi_n_11909 ,csa_tree_add_190_195_groupi_n_12042);
  and csa_tree_add_190_195_groupi_g36756(csa_tree_add_190_195_groupi_n_12149 ,csa_tree_add_190_195_groupi_n_12066 ,csa_tree_add_190_195_groupi_n_12084);
  or csa_tree_add_190_195_groupi_g36757(csa_tree_add_190_195_groupi_n_12148 ,csa_tree_add_190_195_groupi_n_12055 ,csa_tree_add_190_195_groupi_n_12087);
  and csa_tree_add_190_195_groupi_g36758(csa_tree_add_190_195_groupi_n_12147 ,csa_tree_add_190_195_groupi_n_11909 ,csa_tree_add_190_195_groupi_n_12042);
  or csa_tree_add_190_195_groupi_g36759(csa_tree_add_190_195_groupi_n_12146 ,csa_tree_add_190_195_groupi_n_12086 ,csa_tree_add_190_195_groupi_n_12068);
  and csa_tree_add_190_195_groupi_g36760(csa_tree_add_190_195_groupi_n_12145 ,csa_tree_add_190_195_groupi_n_12043 ,csa_tree_add_190_195_groupi_n_12044);
  or csa_tree_add_190_195_groupi_g36761(csa_tree_add_190_195_groupi_n_12144 ,csa_tree_add_190_195_groupi_n_12043 ,csa_tree_add_190_195_groupi_n_12044);
  or csa_tree_add_190_195_groupi_g36762(csa_tree_add_190_195_groupi_n_12143 ,csa_tree_add_190_195_groupi_n_12022 ,csa_tree_add_190_195_groupi_n_12003);
  nor csa_tree_add_190_195_groupi_g36763(csa_tree_add_190_195_groupi_n_12142 ,csa_tree_add_190_195_groupi_n_12025 ,csa_tree_add_190_195_groupi_n_12046);
  or csa_tree_add_190_195_groupi_g36764(csa_tree_add_190_195_groupi_n_12141 ,csa_tree_add_190_195_groupi_n_11908 ,csa_tree_add_190_195_groupi_n_12032);
  nor csa_tree_add_190_195_groupi_g36765(csa_tree_add_190_195_groupi_n_12140 ,csa_tree_add_190_195_groupi_n_11907 ,csa_tree_add_190_195_groupi_n_12033);
  or csa_tree_add_190_195_groupi_g36766(csa_tree_add_190_195_groupi_n_12139 ,csa_tree_add_190_195_groupi_n_12048 ,csa_tree_add_190_195_groupi_n_12076);
  nor csa_tree_add_190_195_groupi_g36767(csa_tree_add_190_195_groupi_n_12138 ,csa_tree_add_190_195_groupi_n_12047 ,csa_tree_add_190_195_groupi_n_12077);
  nor csa_tree_add_190_195_groupi_g36768(csa_tree_add_190_195_groupi_n_12137 ,csa_tree_add_190_195_groupi_n_12028 ,csa_tree_add_190_195_groupi_n_12075);
  or csa_tree_add_190_195_groupi_g36769(csa_tree_add_190_195_groupi_n_12136 ,csa_tree_add_190_195_groupi_n_12065 ,csa_tree_add_190_195_groupi_n_11914);
  or csa_tree_add_190_195_groupi_g36770(csa_tree_add_190_195_groupi_n_12135 ,csa_tree_add_190_195_groupi_n_12029 ,csa_tree_add_190_195_groupi_n_12074);
  or csa_tree_add_190_195_groupi_g36771(csa_tree_add_190_195_groupi_n_12134 ,csa_tree_add_190_195_groupi_n_11999 ,csa_tree_add_190_195_groupi_n_12026);
  nor csa_tree_add_190_195_groupi_g36772(csa_tree_add_190_195_groupi_n_12133 ,csa_tree_add_190_195_groupi_n_12000 ,csa_tree_add_190_195_groupi_n_12027);
  nor csa_tree_add_190_195_groupi_g36773(csa_tree_add_190_195_groupi_n_12132 ,csa_tree_add_190_195_groupi_n_11977 ,csa_tree_add_190_195_groupi_n_12049);
  or csa_tree_add_190_195_groupi_g36774(csa_tree_add_190_195_groupi_n_12131 ,csa_tree_add_190_195_groupi_n_12005 ,csa_tree_add_190_195_groupi_n_12059);
  and csa_tree_add_190_195_groupi_g36775(csa_tree_add_190_195_groupi_n_12130 ,csa_tree_add_190_195_groupi_n_12050 ,csa_tree_add_190_195_groupi_n_12060);
  and csa_tree_add_190_195_groupi_g36776(csa_tree_add_190_195_groupi_n_12163 ,csa_tree_add_190_195_groupi_n_12053 ,csa_tree_add_190_195_groupi_n_11966);
  and csa_tree_add_190_195_groupi_g36777(csa_tree_add_190_195_groupi_n_12162 ,csa_tree_add_190_195_groupi_n_12057 ,csa_tree_add_190_195_groupi_n_11979);
  or csa_tree_add_190_195_groupi_g36778(csa_tree_add_190_195_groupi_n_12161 ,csa_tree_add_190_195_groupi_n_12071 ,csa_tree_add_190_195_groupi_n_11929);
  and csa_tree_add_190_195_groupi_g36779(csa_tree_add_190_195_groupi_n_12160 ,csa_tree_add_190_195_groupi_n_11991 ,csa_tree_add_190_195_groupi_n_12072);
  and csa_tree_add_190_195_groupi_g36780(csa_tree_add_190_195_groupi_n_12159 ,csa_tree_add_190_195_groupi_n_11984 ,csa_tree_add_190_195_groupi_n_12017);
  or csa_tree_add_190_195_groupi_g36781(csa_tree_add_190_195_groupi_n_12158 ,csa_tree_add_190_195_groupi_n_12067 ,csa_tree_add_190_195_groupi_n_11982);
  and csa_tree_add_190_195_groupi_g36782(csa_tree_add_190_195_groupi_n_12155 ,csa_tree_add_190_195_groupi_n_11988 ,csa_tree_add_190_195_groupi_n_12069);
  or csa_tree_add_190_195_groupi_g36783(csa_tree_add_190_195_groupi_n_12154 ,csa_tree_add_190_195_groupi_n_12070 ,csa_tree_add_190_195_groupi_n_11934);
  or csa_tree_add_190_195_groupi_g36784(csa_tree_add_190_195_groupi_n_12152 ,csa_tree_add_190_195_groupi_n_12062 ,csa_tree_add_190_195_groupi_n_11969);
  not csa_tree_add_190_195_groupi_g36785(csa_tree_add_190_195_groupi_n_12129 ,csa_tree_add_190_195_groupi_n_12128);
  not csa_tree_add_190_195_groupi_g36786(csa_tree_add_190_195_groupi_n_12126 ,csa_tree_add_190_195_groupi_n_12125);
  not csa_tree_add_190_195_groupi_g36787(csa_tree_add_190_195_groupi_n_12123 ,csa_tree_add_190_195_groupi_n_12122);
  not csa_tree_add_190_195_groupi_g36788(csa_tree_add_190_195_groupi_n_12121 ,csa_tree_add_190_195_groupi_n_12120);
  not csa_tree_add_190_195_groupi_g36789(csa_tree_add_190_195_groupi_n_12118 ,csa_tree_add_190_195_groupi_n_12117);
  not csa_tree_add_190_195_groupi_g36790(csa_tree_add_190_195_groupi_n_12116 ,csa_tree_add_190_195_groupi_n_12115);
  not csa_tree_add_190_195_groupi_g36791(csa_tree_add_190_195_groupi_n_12114 ,csa_tree_add_190_195_groupi_n_12113);
  not csa_tree_add_190_195_groupi_g36792(csa_tree_add_190_195_groupi_n_12112 ,csa_tree_add_190_195_groupi_n_12111);
  not csa_tree_add_190_195_groupi_g36793(csa_tree_add_190_195_groupi_n_12109 ,csa_tree_add_190_195_groupi_n_12108);
  not csa_tree_add_190_195_groupi_g36794(csa_tree_add_190_195_groupi_n_12107 ,csa_tree_add_190_195_groupi_n_12106);
  or csa_tree_add_190_195_groupi_g36795(csa_tree_add_190_195_groupi_n_12105 ,csa_tree_add_190_195_groupi_n_11997 ,csa_tree_add_190_195_groupi_n_12037);
  nor csa_tree_add_190_195_groupi_g36796(csa_tree_add_190_195_groupi_n_12104 ,csa_tree_add_190_195_groupi_n_11957 ,csa_tree_add_190_195_groupi_n_12038);
  nor csa_tree_add_190_195_groupi_g36797(csa_tree_add_190_195_groupi_n_12103 ,csa_tree_add_190_195_groupi_n_11998 ,csa_tree_add_190_195_groupi_n_12036);
  or csa_tree_add_190_195_groupi_g36798(csa_tree_add_190_195_groupi_n_12102 ,csa_tree_add_190_195_groupi_n_11956 ,csa_tree_add_190_195_groupi_n_12039);
  or csa_tree_add_190_195_groupi_g36799(csa_tree_add_190_195_groupi_n_12101 ,csa_tree_add_190_195_groupi_n_12006 ,csa_tree_add_190_195_groupi_n_12073);
  nor csa_tree_add_190_195_groupi_g36800(csa_tree_add_190_195_groupi_n_12100 ,csa_tree_add_190_195_groupi_n_12080 ,csa_tree_add_190_195_groupi_n_11986);
  or csa_tree_add_190_195_groupi_g36801(csa_tree_add_190_195_groupi_n_12099 ,csa_tree_add_190_195_groupi_n_12024 ,csa_tree_add_190_195_groupi_n_12045);
  xnor csa_tree_add_190_195_groupi_g36802(csa_tree_add_190_195_groupi_n_12098 ,csa_tree_add_190_195_groupi_n_11761 ,csa_tree_add_190_195_groupi_n_11941);
  xnor csa_tree_add_190_195_groupi_g36803(csa_tree_add_190_195_groupi_n_12097 ,csa_tree_add_190_195_groupi_n_11871 ,csa_tree_add_190_195_groupi_n_11945);
  xnor csa_tree_add_190_195_groupi_g36804(csa_tree_add_190_195_groupi_n_12096 ,csa_tree_add_190_195_groupi_n_11960 ,csa_tree_add_190_195_groupi_n_12005);
  xnor csa_tree_add_190_195_groupi_g36805(csa_tree_add_190_195_groupi_n_12095 ,csa_tree_add_190_195_groupi_n_11952 ,csa_tree_add_190_195_groupi_n_11864);
  xnor csa_tree_add_190_195_groupi_g36806(csa_tree_add_190_195_groupi_n_12094 ,csa_tree_add_190_195_groupi_n_11940 ,csa_tree_add_190_195_groupi_n_11944);
  xnor csa_tree_add_190_195_groupi_g36807(csa_tree_add_190_195_groupi_n_12093 ,csa_tree_add_190_195_groupi_n_11995 ,csa_tree_add_190_195_groupi_n_11855);
  xnor csa_tree_add_190_195_groupi_g36808(csa_tree_add_190_195_groupi_n_12092 ,csa_tree_add_190_195_groupi_n_11947 ,csa_tree_add_190_195_groupi_n_12002);
  xnor csa_tree_add_190_195_groupi_g36809(csa_tree_add_190_195_groupi_n_12091 ,csa_tree_add_190_195_groupi_n_11954 ,csa_tree_add_190_195_groupi_n_11955);
  xnor csa_tree_add_190_195_groupi_g36810(csa_tree_add_190_195_groupi_n_12090 ,csa_tree_add_190_195_groupi_n_11903 ,csa_tree_add_190_195_groupi_n_11949);
  xnor csa_tree_add_190_195_groupi_g36811(csa_tree_add_190_195_groupi_n_12089 ,csa_tree_add_190_195_groupi_n_11959 ,csa_tree_add_190_195_groupi_n_11852);
  xnor csa_tree_add_190_195_groupi_g36812(csa_tree_add_190_195_groupi_n_12128 ,csa_tree_add_190_195_groupi_n_11812 ,csa_tree_add_190_195_groupi_n_11920);
  and csa_tree_add_190_195_groupi_g36813(csa_tree_add_190_195_groupi_n_12127 ,csa_tree_add_190_195_groupi_n_12020 ,csa_tree_add_190_195_groupi_n_11931);
  or csa_tree_add_190_195_groupi_g36814(csa_tree_add_190_195_groupi_n_12125 ,csa_tree_add_190_195_groupi_n_11848 ,csa_tree_add_190_195_groupi_n_12016);
  xnor csa_tree_add_190_195_groupi_g36815(csa_tree_add_190_195_groupi_n_12124 ,csa_tree_add_190_195_groupi_n_11861 ,csa_tree_add_190_195_groupi_n_11925);
  xnor csa_tree_add_190_195_groupi_g36816(csa_tree_add_190_195_groupi_n_12122 ,csa_tree_add_190_195_groupi_n_11910 ,csa_tree_add_190_195_groupi_n_11919);
  xnor csa_tree_add_190_195_groupi_g36817(csa_tree_add_190_195_groupi_n_12120 ,csa_tree_add_190_195_groupi_n_11821 ,csa_tree_add_190_195_groupi_n_11918);
  xnor csa_tree_add_190_195_groupi_g36818(csa_tree_add_190_195_groupi_n_12119 ,csa_tree_add_190_195_groupi_n_11815 ,csa_tree_add_190_195_groupi_n_11922);
  xnor csa_tree_add_190_195_groupi_g36819(csa_tree_add_190_195_groupi_n_12117 ,csa_tree_add_190_195_groupi_n_11961 ,csa_tree_add_190_195_groupi_n_11926);
  xnor csa_tree_add_190_195_groupi_g36820(csa_tree_add_190_195_groupi_n_12115 ,csa_tree_add_190_195_groupi_n_11644 ,csa_tree_add_190_195_groupi_n_173);
  xnor csa_tree_add_190_195_groupi_g36821(csa_tree_add_190_195_groupi_n_12113 ,csa_tree_add_190_195_groupi_n_11867 ,csa_tree_add_190_195_groupi_n_11921);
  xnor csa_tree_add_190_195_groupi_g36822(csa_tree_add_190_195_groupi_n_12111 ,csa_tree_add_190_195_groupi_n_11721 ,csa_tree_add_190_195_groupi_n_11917);
  xnor csa_tree_add_190_195_groupi_g36823(csa_tree_add_190_195_groupi_n_12110 ,csa_tree_add_190_195_groupi_n_11822 ,csa_tree_add_190_195_groupi_n_11923);
  xnor csa_tree_add_190_195_groupi_g36824(csa_tree_add_190_195_groupi_n_12108 ,csa_tree_add_190_195_groupi_n_11913 ,csa_tree_add_190_195_groupi_n_11924);
  xnor csa_tree_add_190_195_groupi_g36825(csa_tree_add_190_195_groupi_n_12106 ,csa_tree_add_190_195_groupi_n_11754 ,csa_tree_add_190_195_groupi_n_172);
  not csa_tree_add_190_195_groupi_g36826(csa_tree_add_190_195_groupi_n_12086 ,csa_tree_add_190_195_groupi_n_12085);
  not csa_tree_add_190_195_groupi_g36828(csa_tree_add_190_195_groupi_n_12076 ,csa_tree_add_190_195_groupi_n_12077);
  not csa_tree_add_190_195_groupi_g36829(csa_tree_add_190_195_groupi_n_12075 ,csa_tree_add_190_195_groupi_n_12074);
  nor csa_tree_add_190_195_groupi_g36830(csa_tree_add_190_195_groupi_n_12073 ,csa_tree_add_190_195_groupi_n_11953 ,csa_tree_add_190_195_groupi_n_11955);
  or csa_tree_add_190_195_groupi_g36831(csa_tree_add_190_195_groupi_n_12072 ,csa_tree_add_190_195_groupi_n_11990 ,csa_tree_add_190_195_groupi_n_11870);
  and csa_tree_add_190_195_groupi_g36832(csa_tree_add_190_195_groupi_n_12071 ,csa_tree_add_190_195_groupi_n_11912 ,csa_tree_add_190_195_groupi_n_11928);
  nor csa_tree_add_190_195_groupi_g36833(csa_tree_add_190_195_groupi_n_12070 ,csa_tree_add_190_195_groupi_n_11989 ,csa_tree_add_190_195_groupi_n_11825);
  or csa_tree_add_190_195_groupi_g36834(csa_tree_add_190_195_groupi_n_12069 ,csa_tree_add_190_195_groupi_n_11963 ,csa_tree_add_190_195_groupi_n_11987);
  nor csa_tree_add_190_195_groupi_g36835(csa_tree_add_190_195_groupi_n_12068 ,csa_tree_add_190_195_groupi_n_11758 ,csa_tree_add_190_195_groupi_n_11938);
  and csa_tree_add_190_195_groupi_g36836(csa_tree_add_190_195_groupi_n_12067 ,csa_tree_add_190_195_groupi_n_11915 ,csa_tree_add_190_195_groupi_n_11983);
  or csa_tree_add_190_195_groupi_g36837(csa_tree_add_190_195_groupi_n_12066 ,csa_tree_add_190_195_groupi_n_11996 ,csa_tree_add_190_195_groupi_n_11855);
  nor csa_tree_add_190_195_groupi_g36838(csa_tree_add_190_195_groupi_n_12065 ,csa_tree_add_190_195_groupi_n_11940 ,csa_tree_add_190_195_groupi_n_11944);
  or csa_tree_add_190_195_groupi_g36839(csa_tree_add_190_195_groupi_n_12064 ,csa_tree_add_190_195_groupi_n_11939 ,csa_tree_add_190_195_groupi_n_11943);
  or csa_tree_add_190_195_groupi_g36840(csa_tree_add_190_195_groupi_n_12063 ,csa_tree_add_190_195_groupi_n_168 ,csa_tree_add_190_195_groupi_n_11937);
  and csa_tree_add_190_195_groupi_g36841(csa_tree_add_190_195_groupi_n_12062 ,csa_tree_add_190_195_groupi_n_11916 ,csa_tree_add_190_195_groupi_n_11970);
  nor csa_tree_add_190_195_groupi_g36842(csa_tree_add_190_195_groupi_n_12061 ,csa_tree_add_190_195_groupi_n_11947 ,csa_tree_add_190_195_groupi_n_12001);
  or csa_tree_add_190_195_groupi_g36843(csa_tree_add_190_195_groupi_n_12060 ,csa_tree_add_190_195_groupi_n_11946 ,csa_tree_add_190_195_groupi_n_12002);
  and csa_tree_add_190_195_groupi_g36844(csa_tree_add_190_195_groupi_n_12059 ,csa_tree_add_190_195_groupi_n_11960 ,csa_tree_add_190_195_groupi_n_11950);
  or csa_tree_add_190_195_groupi_g36845(csa_tree_add_190_195_groupi_n_12058 ,csa_tree_add_190_195_groupi_n_11960 ,csa_tree_add_190_195_groupi_n_11950);
  or csa_tree_add_190_195_groupi_g36846(csa_tree_add_190_195_groupi_n_12057 ,csa_tree_add_190_195_groupi_n_11971 ,csa_tree_add_190_195_groupi_n_11823);
  or csa_tree_add_190_195_groupi_g36847(csa_tree_add_190_195_groupi_n_12056 ,csa_tree_add_190_195_groupi_n_11902 ,csa_tree_add_190_195_groupi_n_11948);
  nor csa_tree_add_190_195_groupi_g36848(csa_tree_add_190_195_groupi_n_12055 ,csa_tree_add_190_195_groupi_n_11903 ,csa_tree_add_190_195_groupi_n_11949);
  or csa_tree_add_190_195_groupi_g36849(csa_tree_add_190_195_groupi_n_12054 ,csa_tree_add_190_195_groupi_n_11959 ,csa_tree_add_190_195_groupi_n_11851);
  or csa_tree_add_190_195_groupi_g36850(csa_tree_add_190_195_groupi_n_12053 ,csa_tree_add_190_195_groupi_n_11968 ,csa_tree_add_190_195_groupi_n_11719);
  nor csa_tree_add_190_195_groupi_g36851(csa_tree_add_190_195_groupi_n_12052 ,csa_tree_add_190_195_groupi_n_11958 ,csa_tree_add_190_195_groupi_n_11852);
  and csa_tree_add_190_195_groupi_g36852(csa_tree_add_190_195_groupi_n_12088 ,csa_tree_add_190_195_groupi_n_11981 ,csa_tree_add_190_195_groupi_n_11884);
  and csa_tree_add_190_195_groupi_g36853(csa_tree_add_190_195_groupi_n_12087 ,csa_tree_add_190_195_groupi_n_11992 ,csa_tree_add_190_195_groupi_n_11875);
  or csa_tree_add_190_195_groupi_g36854(csa_tree_add_190_195_groupi_n_12085 ,csa_tree_add_190_195_groupi_n_11879 ,csa_tree_add_190_195_groupi_n_11974);
  or csa_tree_add_190_195_groupi_g36855(csa_tree_add_190_195_groupi_n_12084 ,csa_tree_add_190_195_groupi_n_11994 ,csa_tree_add_190_195_groupi_n_11785);
  and csa_tree_add_190_195_groupi_g36856(csa_tree_add_190_195_groupi_n_12083 ,csa_tree_add_190_195_groupi_n_11993 ,csa_tree_add_190_195_groupi_n_11898);
  and csa_tree_add_190_195_groupi_g36857(csa_tree_add_190_195_groupi_n_12082 ,csa_tree_add_190_195_groupi_n_11985 ,csa_tree_add_190_195_groupi_n_11889);
  and csa_tree_add_190_195_groupi_g36858(csa_tree_add_190_195_groupi_n_12081 ,csa_tree_add_190_195_groupi_n_11888 ,csa_tree_add_190_195_groupi_n_11967);
  and csa_tree_add_190_195_groupi_g36859(csa_tree_add_190_195_groupi_n_12080 ,csa_tree_add_190_195_groupi_n_11787 ,csa_tree_add_190_195_groupi_n_11972);
  or csa_tree_add_190_195_groupi_g36860(csa_tree_add_190_195_groupi_n_12079 ,csa_tree_add_190_195_groupi_n_11965 ,csa_tree_add_190_195_groupi_n_11890);
  and csa_tree_add_190_195_groupi_g36861(csa_tree_add_190_195_groupi_n_12078 ,csa_tree_add_190_195_groupi_n_11973 ,csa_tree_add_190_195_groupi_n_11877);
  or csa_tree_add_190_195_groupi_g36862(csa_tree_add_190_195_groupi_n_12077 ,csa_tree_add_190_195_groupi_n_11975 ,csa_tree_add_190_195_groupi_n_11778);
  and csa_tree_add_190_195_groupi_g36863(csa_tree_add_190_195_groupi_n_12074 ,csa_tree_add_190_195_groupi_n_11980 ,csa_tree_add_190_195_groupi_n_11886);
  not csa_tree_add_190_195_groupi_g36864(csa_tree_add_190_195_groupi_n_12048 ,csa_tree_add_190_195_groupi_n_12047);
  not csa_tree_add_190_195_groupi_g36865(csa_tree_add_190_195_groupi_n_12046 ,csa_tree_add_190_195_groupi_n_12045);
  not csa_tree_add_190_195_groupi_g36866(csa_tree_add_190_195_groupi_n_12041 ,csa_tree_add_190_195_groupi_n_12040);
  not csa_tree_add_190_195_groupi_g36867(csa_tree_add_190_195_groupi_n_12039 ,csa_tree_add_190_195_groupi_n_12038);
  not csa_tree_add_190_195_groupi_g36868(csa_tree_add_190_195_groupi_n_12037 ,csa_tree_add_190_195_groupi_n_12036);
  not csa_tree_add_190_195_groupi_g36869(csa_tree_add_190_195_groupi_n_12035 ,csa_tree_add_190_195_groupi_n_12034);
  not csa_tree_add_190_195_groupi_g36870(csa_tree_add_190_195_groupi_n_12033 ,csa_tree_add_190_195_groupi_n_12032);
  not csa_tree_add_190_195_groupi_g36871(csa_tree_add_190_195_groupi_n_12031 ,csa_tree_add_190_195_groupi_n_12030);
  not csa_tree_add_190_195_groupi_g36872(csa_tree_add_190_195_groupi_n_12029 ,csa_tree_add_190_195_groupi_n_12028);
  not csa_tree_add_190_195_groupi_g36873(csa_tree_add_190_195_groupi_n_12027 ,csa_tree_add_190_195_groupi_n_12026);
  not csa_tree_add_190_195_groupi_g36874(csa_tree_add_190_195_groupi_n_12025 ,csa_tree_add_190_195_groupi_n_12024);
  or csa_tree_add_190_195_groupi_g36875(csa_tree_add_190_195_groupi_n_12023 ,csa_tree_add_190_195_groupi_n_11954 ,csa_tree_add_190_195_groupi_n_170);
  nor csa_tree_add_190_195_groupi_g36876(csa_tree_add_190_195_groupi_n_12022 ,csa_tree_add_190_195_groupi_n_11951 ,csa_tree_add_190_195_groupi_n_11864);
  or csa_tree_add_190_195_groupi_g36877(csa_tree_add_190_195_groupi_n_12021 ,csa_tree_add_190_195_groupi_n_11952 ,csa_tree_add_190_195_groupi_n_11863);
  or csa_tree_add_190_195_groupi_g36878(csa_tree_add_190_195_groupi_n_12020 ,csa_tree_add_190_195_groupi_n_11964 ,csa_tree_add_190_195_groupi_n_11932);
  nor csa_tree_add_190_195_groupi_g36879(csa_tree_add_190_195_groupi_n_12019 ,csa_tree_add_190_195_groupi_n_11761 ,csa_tree_add_190_195_groupi_n_11942);
  and csa_tree_add_190_195_groupi_g36880(csa_tree_add_190_195_groupi_n_12018 ,csa_tree_add_190_195_groupi_n_11761 ,csa_tree_add_190_195_groupi_n_11942);
  or csa_tree_add_190_195_groupi_g36881(csa_tree_add_190_195_groupi_n_12017 ,csa_tree_add_190_195_groupi_n_11930 ,csa_tree_add_190_195_groupi_n_11720);
  and csa_tree_add_190_195_groupi_g36882(csa_tree_add_190_195_groupi_n_12016 ,csa_tree_add_190_195_groupi_n_11961 ,csa_tree_add_190_195_groupi_n_11846);
  and csa_tree_add_190_195_groupi_g36883(csa_tree_add_190_195_groupi_n_12015 ,csa_tree_add_190_195_groupi_n_11996 ,csa_tree_add_190_195_groupi_n_11855);
  xnor csa_tree_add_190_195_groupi_g36884(csa_tree_add_190_195_groupi_n_12014 ,csa_tree_add_190_195_groupi_n_11916 ,csa_tree_add_190_195_groupi_n_11662);
  xnor csa_tree_add_190_195_groupi_g36885(csa_tree_add_190_195_groupi_n_12013 ,csa_tree_add_190_195_groupi_n_11866 ,csa_tree_add_190_195_groupi_n_11760);
  xnor csa_tree_add_190_195_groupi_g36886(csa_tree_add_190_195_groupi_n_12012 ,csa_tree_add_190_195_groupi_n_11814 ,csa_tree_add_190_195_groupi_n_11850);
  xnor csa_tree_add_190_195_groupi_g36887(csa_tree_add_190_195_groupi_n_12011 ,csa_tree_add_190_195_groupi_n_11763 ,csa_tree_add_190_195_groupi_n_11906);
  xnor csa_tree_add_190_195_groupi_g36888(csa_tree_add_190_195_groupi_n_12010 ,csa_tree_add_190_195_groupi_n_11755 ,csa_tree_add_190_195_groupi_n_11912);
  xnor csa_tree_add_190_195_groupi_g36889(csa_tree_add_190_195_groupi_n_12009 ,csa_tree_add_190_195_groupi_n_11860 ,csa_tree_add_190_195_groupi_n_11817);
  xnor csa_tree_add_190_195_groupi_g36890(csa_tree_add_190_195_groupi_n_12008 ,csa_tree_add_190_195_groupi_n_11857 ,csa_tree_add_190_195_groupi_n_11752);
  xnor csa_tree_add_190_195_groupi_g36891(csa_tree_add_190_195_groupi_n_12007 ,csa_tree_add_190_195_groupi_n_11858 ,csa_tree_add_190_195_groupi_n_11460);
  xnor csa_tree_add_190_195_groupi_g36892(csa_tree_add_190_195_groupi_n_12051 ,csa_tree_add_190_195_groupi_n_11660 ,csa_tree_add_190_195_groupi_n_11841);
  xnor csa_tree_add_190_195_groupi_g36893(csa_tree_add_190_195_groupi_n_12050 ,csa_tree_add_190_195_groupi_n_11584 ,csa_tree_add_190_195_groupi_n_11833);
  xnor csa_tree_add_190_195_groupi_g36894(csa_tree_add_190_195_groupi_n_12049 ,csa_tree_add_190_195_groupi_n_11632 ,csa_tree_add_190_195_groupi_n_11835);
  xnor csa_tree_add_190_195_groupi_g36895(csa_tree_add_190_195_groupi_n_12047 ,csa_tree_add_190_195_groupi_n_11590 ,csa_tree_add_190_195_groupi_n_11832);
  xnor csa_tree_add_190_195_groupi_g36896(csa_tree_add_190_195_groupi_n_12045 ,csa_tree_add_190_195_groupi_n_11713 ,csa_tree_add_190_195_groupi_n_11842);
  xnor csa_tree_add_190_195_groupi_g36897(csa_tree_add_190_195_groupi_n_12044 ,csa_tree_add_190_195_groupi_n_11716 ,csa_tree_add_190_195_groupi_n_11829);
  xnor csa_tree_add_190_195_groupi_g36898(csa_tree_add_190_195_groupi_n_12043 ,csa_tree_add_190_195_groupi_n_11868 ,csa_tree_add_190_195_groupi_n_11844);
  xnor csa_tree_add_190_195_groupi_g36899(csa_tree_add_190_195_groupi_n_12042 ,csa_tree_add_190_195_groupi_n_11472 ,csa_tree_add_190_195_groupi_n_11831);
  xnor csa_tree_add_190_195_groupi_g36900(csa_tree_add_190_195_groupi_n_12040 ,csa_tree_add_190_195_groupi_n_11665 ,csa_tree_add_190_195_groupi_n_11836);
  xnor csa_tree_add_190_195_groupi_g36901(csa_tree_add_190_195_groupi_n_12038 ,csa_tree_add_190_195_groupi_n_11854 ,csa_tree_add_190_195_groupi_n_11838);
  xnor csa_tree_add_190_195_groupi_g36902(csa_tree_add_190_195_groupi_n_12036 ,csa_tree_add_190_195_groupi_n_159 ,csa_tree_add_190_195_groupi_n_171);
  xnor csa_tree_add_190_195_groupi_g36903(csa_tree_add_190_195_groupi_n_12034 ,csa_tree_add_190_195_groupi_n_11773 ,csa_tree_add_190_195_groupi_n_11839);
  xnor csa_tree_add_190_195_groupi_g36904(csa_tree_add_190_195_groupi_n_12032 ,csa_tree_add_190_195_groupi_n_11775 ,csa_tree_add_190_195_groupi_n_11840);
  xnor csa_tree_add_190_195_groupi_g36905(csa_tree_add_190_195_groupi_n_12030 ,csa_tree_add_190_195_groupi_n_11911 ,csa_tree_add_190_195_groupi_n_11834);
  xnor csa_tree_add_190_195_groupi_g36906(csa_tree_add_190_195_groupi_n_12028 ,csa_tree_add_190_195_groupi_n_11862 ,csa_tree_add_190_195_groupi_n_11837);
  xnor csa_tree_add_190_195_groupi_g36907(csa_tree_add_190_195_groupi_n_12026 ,csa_tree_add_190_195_groupi_n_11872 ,csa_tree_add_190_195_groupi_n_11830);
  and csa_tree_add_190_195_groupi_g36908(csa_tree_add_190_195_groupi_n_12024 ,csa_tree_add_190_195_groupi_n_11927 ,csa_tree_add_190_195_groupi_n_11892);
  not csa_tree_add_190_195_groupi_g36910(csa_tree_add_190_195_groupi_n_12002 ,csa_tree_add_190_195_groupi_n_12001);
  not csa_tree_add_190_195_groupi_g36911(csa_tree_add_190_195_groupi_n_12000 ,csa_tree_add_190_195_groupi_n_11999);
  not csa_tree_add_190_195_groupi_g36912(csa_tree_add_190_195_groupi_n_11998 ,csa_tree_add_190_195_groupi_n_11997);
  not csa_tree_add_190_195_groupi_g36913(csa_tree_add_190_195_groupi_n_11996 ,csa_tree_add_190_195_groupi_n_11995);
  and csa_tree_add_190_195_groupi_g36914(csa_tree_add_190_195_groupi_n_11994 ,csa_tree_add_190_195_groupi_n_11911 ,csa_tree_add_190_195_groupi_n_11786);
  or csa_tree_add_190_195_groupi_g36915(csa_tree_add_190_195_groupi_n_11993 ,csa_tree_add_190_195_groupi_n_11776 ,csa_tree_add_190_195_groupi_n_11899);
  or csa_tree_add_190_195_groupi_g36916(csa_tree_add_190_195_groupi_n_11992 ,csa_tree_add_190_195_groupi_n_11594 ,csa_tree_add_190_195_groupi_n_11876);
  or csa_tree_add_190_195_groupi_g36917(csa_tree_add_190_195_groupi_n_11991 ,csa_tree_add_190_195_groupi_n_11460 ,csa_tree_add_190_195_groupi_n_11858);
  and csa_tree_add_190_195_groupi_g36918(csa_tree_add_190_195_groupi_n_11990 ,csa_tree_add_190_195_groupi_n_11460 ,csa_tree_add_190_195_groupi_n_11858);
  and csa_tree_add_190_195_groupi_g36919(csa_tree_add_190_195_groupi_n_11989 ,csa_tree_add_190_195_groupi_n_11861 ,csa_tree_add_190_195_groupi_n_161);
  or csa_tree_add_190_195_groupi_g36920(csa_tree_add_190_195_groupi_n_11988 ,csa_tree_add_190_195_groupi_n_11859 ,csa_tree_add_190_195_groupi_n_11817);
  nor csa_tree_add_190_195_groupi_g36921(csa_tree_add_190_195_groupi_n_11987 ,csa_tree_add_190_195_groupi_n_11860 ,csa_tree_add_190_195_groupi_n_11816);
  nor csa_tree_add_190_195_groupi_g36922(csa_tree_add_190_195_groupi_n_11986 ,csa_tree_add_190_195_groupi_n_11814 ,csa_tree_add_190_195_groupi_n_11850);
  or csa_tree_add_190_195_groupi_g36923(csa_tree_add_190_195_groupi_n_11985 ,csa_tree_add_190_195_groupi_n_11891 ,csa_tree_add_190_195_groupi_n_11913);
  or csa_tree_add_190_195_groupi_g36924(csa_tree_add_190_195_groupi_n_11984 ,csa_tree_add_190_195_groupi_n_11862 ,csa_tree_add_190_195_groupi_n_11255);
  or csa_tree_add_190_195_groupi_g36925(csa_tree_add_190_195_groupi_n_11983 ,csa_tree_add_190_195_groupi_n_11865 ,csa_tree_add_190_195_groupi_n_11760);
  nor csa_tree_add_190_195_groupi_g36926(csa_tree_add_190_195_groupi_n_11982 ,csa_tree_add_190_195_groupi_n_11866 ,csa_tree_add_190_195_groupi_n_11759);
  or csa_tree_add_190_195_groupi_g36927(csa_tree_add_190_195_groupi_n_11981 ,csa_tree_add_190_195_groupi_n_11887 ,csa_tree_add_190_195_groupi_n_11826);
  or csa_tree_add_190_195_groupi_g36928(csa_tree_add_190_195_groupi_n_11980 ,csa_tree_add_190_195_groupi_n_11601 ,csa_tree_add_190_195_groupi_n_11885);
  or csa_tree_add_190_195_groupi_g36929(csa_tree_add_190_195_groupi_n_11979 ,csa_tree_add_190_195_groupi_n_11820 ,csa_tree_add_190_195_groupi_n_11867);
  and csa_tree_add_190_195_groupi_g36930(csa_tree_add_190_195_groupi_n_11978 ,csa_tree_add_190_195_groupi_n_11763 ,csa_tree_add_190_195_groupi_n_11906);
  nor csa_tree_add_190_195_groupi_g36931(csa_tree_add_190_195_groupi_n_11977 ,csa_tree_add_190_195_groupi_n_11763 ,csa_tree_add_190_195_groupi_n_11906);
  and csa_tree_add_190_195_groupi_g36932(csa_tree_add_190_195_groupi_n_11976 ,csa_tree_add_190_195_groupi_n_11814 ,csa_tree_add_190_195_groupi_n_11850);
  and csa_tree_add_190_195_groupi_g36933(csa_tree_add_190_195_groupi_n_11975 ,csa_tree_add_190_195_groupi_n_11779 ,csa_tree_add_190_195_groupi_n_11868);
  and csa_tree_add_190_195_groupi_g36934(csa_tree_add_190_195_groupi_n_11974 ,csa_tree_add_190_195_groupi_n_11822 ,csa_tree_add_190_195_groupi_n_11894);
  or csa_tree_add_190_195_groupi_g36935(csa_tree_add_190_195_groupi_n_11973 ,csa_tree_add_190_195_groupi_n_11821 ,csa_tree_add_190_195_groupi_n_11878);
  or csa_tree_add_190_195_groupi_g36936(csa_tree_add_190_195_groupi_n_11972 ,csa_tree_add_190_195_groupi_n_11873 ,csa_tree_add_190_195_groupi_n_11794);
  and csa_tree_add_190_195_groupi_g36937(csa_tree_add_190_195_groupi_n_11971 ,csa_tree_add_190_195_groupi_n_11820 ,csa_tree_add_190_195_groupi_n_11867);
  or csa_tree_add_190_195_groupi_g36938(csa_tree_add_190_195_groupi_n_11970 ,csa_tree_add_190_195_groupi_n_11662 ,csa_tree_add_190_195_groupi_n_11904);
  nor csa_tree_add_190_195_groupi_g36939(csa_tree_add_190_195_groupi_n_11969 ,csa_tree_add_190_195_groupi_n_11661 ,csa_tree_add_190_195_groupi_n_11905);
  nor csa_tree_add_190_195_groupi_g36940(csa_tree_add_190_195_groupi_n_11968 ,csa_tree_add_190_195_groupi_n_11659 ,csa_tree_add_190_195_groupi_n_11854);
  or csa_tree_add_190_195_groupi_g36941(csa_tree_add_190_195_groupi_n_11967 ,csa_tree_add_190_195_groupi_n_11721 ,csa_tree_add_190_195_groupi_n_11900);
  or csa_tree_add_190_195_groupi_g36942(csa_tree_add_190_195_groupi_n_11966 ,csa_tree_add_190_195_groupi_n_11658 ,csa_tree_add_190_195_groupi_n_169);
  nor csa_tree_add_190_195_groupi_g36943(csa_tree_add_190_195_groupi_n_11965 ,csa_tree_add_190_195_groupi_n_11910 ,csa_tree_add_190_195_groupi_n_11883);
  and csa_tree_add_190_195_groupi_g36944(csa_tree_add_190_195_groupi_n_12006 ,csa_tree_add_190_195_groupi_n_11750 ,csa_tree_add_190_195_groupi_n_11897);
  and csa_tree_add_190_195_groupi_g36945(csa_tree_add_190_195_groupi_n_12005 ,csa_tree_add_190_195_groupi_n_11781 ,csa_tree_add_190_195_groupi_n_11881);
  and csa_tree_add_190_195_groupi_g36946(csa_tree_add_190_195_groupi_n_12004 ,csa_tree_add_190_195_groupi_n_11777 ,csa_tree_add_190_195_groupi_n_11880);
  and csa_tree_add_190_195_groupi_g36947(csa_tree_add_190_195_groupi_n_12003 ,csa_tree_add_190_195_groupi_n_11747 ,csa_tree_add_190_195_groupi_n_11895);
  and csa_tree_add_190_195_groupi_g36948(csa_tree_add_190_195_groupi_n_12001 ,csa_tree_add_190_195_groupi_n_11807 ,csa_tree_add_190_195_groupi_n_11882);
  and csa_tree_add_190_195_groupi_g36949(csa_tree_add_190_195_groupi_n_11999 ,csa_tree_add_190_195_groupi_n_11745 ,csa_tree_add_190_195_groupi_n_11845);
  and csa_tree_add_190_195_groupi_g36950(csa_tree_add_190_195_groupi_n_11997 ,csa_tree_add_190_195_groupi_n_11874 ,csa_tree_add_190_195_groupi_n_11804);
  and csa_tree_add_190_195_groupi_g36951(csa_tree_add_190_195_groupi_n_11995 ,csa_tree_add_190_195_groupi_n_11798 ,csa_tree_add_190_195_groupi_n_11896);
  not csa_tree_add_190_195_groupi_g36952(csa_tree_add_190_195_groupi_n_11963 ,csa_tree_add_190_195_groupi_n_11962);
  not csa_tree_add_190_195_groupi_g36953(csa_tree_add_190_195_groupi_n_11959 ,csa_tree_add_190_195_groupi_n_11958);
  not csa_tree_add_190_195_groupi_g36954(csa_tree_add_190_195_groupi_n_11957 ,csa_tree_add_190_195_groupi_n_11956);
  not csa_tree_add_190_195_groupi_g36955(csa_tree_add_190_195_groupi_n_11955 ,csa_tree_add_190_195_groupi_n_170);
  not csa_tree_add_190_195_groupi_g36956(csa_tree_add_190_195_groupi_n_11954 ,csa_tree_add_190_195_groupi_n_11953);
  not csa_tree_add_190_195_groupi_g36957(csa_tree_add_190_195_groupi_n_11952 ,csa_tree_add_190_195_groupi_n_11951);
  not csa_tree_add_190_195_groupi_g36958(csa_tree_add_190_195_groupi_n_11949 ,csa_tree_add_190_195_groupi_n_11948);
  not csa_tree_add_190_195_groupi_g36959(csa_tree_add_190_195_groupi_n_11947 ,csa_tree_add_190_195_groupi_n_11946);
  not csa_tree_add_190_195_groupi_g36960(csa_tree_add_190_195_groupi_n_11944 ,csa_tree_add_190_195_groupi_n_11943);
  not csa_tree_add_190_195_groupi_g36961(csa_tree_add_190_195_groupi_n_11942 ,csa_tree_add_190_195_groupi_n_11941);
  not csa_tree_add_190_195_groupi_g36962(csa_tree_add_190_195_groupi_n_11940 ,csa_tree_add_190_195_groupi_n_11939);
  not csa_tree_add_190_195_groupi_g36963(csa_tree_add_190_195_groupi_n_11938 ,csa_tree_add_190_195_groupi_n_11937);
  not csa_tree_add_190_195_groupi_g36964(csa_tree_add_190_195_groupi_n_11936 ,csa_tree_add_190_195_groupi_n_11935);
  nor csa_tree_add_190_195_groupi_g36965(csa_tree_add_190_195_groupi_n_11934 ,csa_tree_add_190_195_groupi_n_11861 ,csa_tree_add_190_195_groupi_n_161);
  xnor csa_tree_add_190_195_groupi_g36966(out1[4] ,csa_tree_add_190_195_groupi_n_11541 ,csa_tree_add_190_195_groupi_n_11722);
  nor csa_tree_add_190_195_groupi_g36967(csa_tree_add_190_195_groupi_n_11932 ,csa_tree_add_190_195_groupi_n_11856 ,csa_tree_add_190_195_groupi_n_11752);
  or csa_tree_add_190_195_groupi_g36968(csa_tree_add_190_195_groupi_n_11931 ,csa_tree_add_190_195_groupi_n_11857 ,csa_tree_add_190_195_groupi_n_11751);
  and csa_tree_add_190_195_groupi_g36969(csa_tree_add_190_195_groupi_n_11930 ,csa_tree_add_190_195_groupi_n_11862 ,csa_tree_add_190_195_groupi_n_11255);
  and csa_tree_add_190_195_groupi_g36970(csa_tree_add_190_195_groupi_n_11929 ,csa_tree_add_190_195_groupi_n_11755 ,csa_tree_add_190_195_groupi_n_11853);
  or csa_tree_add_190_195_groupi_g36971(csa_tree_add_190_195_groupi_n_11928 ,csa_tree_add_190_195_groupi_n_11755 ,csa_tree_add_190_195_groupi_n_11853);
  or csa_tree_add_190_195_groupi_g36972(csa_tree_add_190_195_groupi_n_11927 ,csa_tree_add_190_195_groupi_n_11824 ,csa_tree_add_190_195_groupi_n_11893);
  xnor csa_tree_add_190_195_groupi_g36973(csa_tree_add_190_195_groupi_n_11926 ,csa_tree_add_190_195_groupi_n_11636 ,csa_tree_add_190_195_groupi_n_11757);
  xnor csa_tree_add_190_195_groupi_g36974(csa_tree_add_190_195_groupi_n_11925 ,csa_tree_add_190_195_groupi_n_161 ,csa_tree_add_190_195_groupi_n_11825);
  xnor csa_tree_add_190_195_groupi_g36975(csa_tree_add_190_195_groupi_n_11924 ,csa_tree_add_190_195_groupi_n_11640 ,csa_tree_add_190_195_groupi_n_11819);
  xnor csa_tree_add_190_195_groupi_g36976(csa_tree_add_190_195_groupi_n_11923 ,csa_tree_add_190_195_groupi_n_11765 ,csa_tree_add_190_195_groupi_n_11527);
  xnor csa_tree_add_190_195_groupi_g36977(csa_tree_add_190_195_groupi_n_11922 ,csa_tree_add_190_195_groupi_n_11776 ,csa_tree_add_190_195_groupi_n_11762);
  xor csa_tree_add_190_195_groupi_g36978(csa_tree_add_190_195_groupi_n_11921 ,csa_tree_add_190_195_groupi_n_11823 ,csa_tree_add_190_195_groupi_n_11820);
  xnor csa_tree_add_190_195_groupi_g36980(csa_tree_add_190_195_groupi_n_11920 ,csa_tree_add_190_195_groupi_n_11772 ,csa_tree_add_190_195_groupi_n_11826);
  xnor csa_tree_add_190_195_groupi_g36981(csa_tree_add_190_195_groupi_n_11919 ,csa_tree_add_190_195_groupi_n_11813 ,csa_tree_add_190_195_groupi_n_11769);
  xnor csa_tree_add_190_195_groupi_g36983(csa_tree_add_190_195_groupi_n_11918 ,csa_tree_add_190_195_groupi_n_11767 ,csa_tree_add_190_195_groupi_n_11810);
  xnor csa_tree_add_190_195_groupi_g36984(csa_tree_add_190_195_groupi_n_11917 ,csa_tree_add_190_195_groupi_n_11523 ,csa_tree_add_190_195_groupi_n_11770);
  and csa_tree_add_190_195_groupi_g36985(csa_tree_add_190_195_groupi_n_11964 ,csa_tree_add_190_195_groupi_n_11901 ,csa_tree_add_190_195_groupi_n_11738);
  xnor csa_tree_add_190_195_groupi_g36986(csa_tree_add_190_195_groupi_n_11962 ,csa_tree_add_190_195_groupi_n_11538 ,csa_tree_add_190_195_groupi_n_11734);
  or csa_tree_add_190_195_groupi_g36987(csa_tree_add_190_195_groupi_n_11961 ,csa_tree_add_190_195_groupi_n_11849 ,csa_tree_add_190_195_groupi_n_11749);
  xnor csa_tree_add_190_195_groupi_g36988(csa_tree_add_190_195_groupi_n_11960 ,csa_tree_add_190_195_groupi_n_11241 ,csa_tree_add_190_195_groupi_n_11728);
  xnor csa_tree_add_190_195_groupi_g36989(csa_tree_add_190_195_groupi_n_11958 ,csa_tree_add_190_195_groupi_n_11447 ,csa_tree_add_190_195_groupi_n_11737);
  xnor csa_tree_add_190_195_groupi_g36990(csa_tree_add_190_195_groupi_n_11956 ,csa_tree_add_190_195_groupi_n_11509 ,csa_tree_add_190_195_groupi_n_11723);
  xnor csa_tree_add_190_195_groupi_g36992(csa_tree_add_190_195_groupi_n_11953 ,csa_tree_add_190_195_groupi_n_11768 ,csa_tree_add_190_195_groupi_n_11725);
  xnor csa_tree_add_190_195_groupi_g36993(csa_tree_add_190_195_groupi_n_11951 ,csa_tree_add_190_195_groupi_n_11597 ,csa_tree_add_190_195_groupi_n_11729);
  xnor csa_tree_add_190_195_groupi_g36994(csa_tree_add_190_195_groupi_n_11950 ,csa_tree_add_190_195_groupi_n_11478 ,csa_tree_add_190_195_groupi_n_11727);
  xnor csa_tree_add_190_195_groupi_g36995(csa_tree_add_190_195_groupi_n_11948 ,csa_tree_add_190_195_groupi_n_11339 ,csa_tree_add_190_195_groupi_n_11724);
  xnor csa_tree_add_190_195_groupi_g36996(csa_tree_add_190_195_groupi_n_11946 ,csa_tree_add_190_195_groupi_n_11506 ,csa_tree_add_190_195_groupi_n_11730);
  xnor csa_tree_add_190_195_groupi_g36997(csa_tree_add_190_195_groupi_n_11945 ,csa_tree_add_190_195_groupi_n_11647 ,csa_tree_add_190_195_groupi_n_11731);
  xnor csa_tree_add_190_195_groupi_g36998(csa_tree_add_190_195_groupi_n_11943 ,csa_tree_add_190_195_groupi_n_11595 ,csa_tree_add_190_195_groupi_n_11732);
  xnor csa_tree_add_190_195_groupi_g36999(csa_tree_add_190_195_groupi_n_11941 ,csa_tree_add_190_195_groupi_n_11774 ,csa_tree_add_190_195_groupi_n_11736);
  xnor csa_tree_add_190_195_groupi_g37000(csa_tree_add_190_195_groupi_n_11939 ,csa_tree_add_190_195_groupi_n_11521 ,csa_tree_add_190_195_groupi_n_11733);
  xnor csa_tree_add_190_195_groupi_g37001(csa_tree_add_190_195_groupi_n_11937 ,csa_tree_add_190_195_groupi_n_11808 ,csa_tree_add_190_195_groupi_n_11735);
  and csa_tree_add_190_195_groupi_g37002(csa_tree_add_190_195_groupi_n_11935 ,csa_tree_add_190_195_groupi_n_11628 ,csa_tree_add_190_195_groupi_n_11847);
  not csa_tree_add_190_195_groupi_g37003(csa_tree_add_190_195_groupi_n_11908 ,csa_tree_add_190_195_groupi_n_11907);
  not csa_tree_add_190_195_groupi_g37004(csa_tree_add_190_195_groupi_n_11905 ,csa_tree_add_190_195_groupi_n_11904);
  not csa_tree_add_190_195_groupi_g37005(csa_tree_add_190_195_groupi_n_11903 ,csa_tree_add_190_195_groupi_n_11902);
  or csa_tree_add_190_195_groupi_g37006(csa_tree_add_190_195_groupi_n_11901 ,csa_tree_add_190_195_groupi_n_11744 ,csa_tree_add_190_195_groupi_n_11775);
  nor csa_tree_add_190_195_groupi_g37007(csa_tree_add_190_195_groupi_n_11900 ,csa_tree_add_190_195_groupi_n_11522 ,csa_tree_add_190_195_groupi_n_11770);
  and csa_tree_add_190_195_groupi_g37008(csa_tree_add_190_195_groupi_n_11899 ,csa_tree_add_190_195_groupi_n_11815 ,csa_tree_add_190_195_groupi_n_11762);
  or csa_tree_add_190_195_groupi_g37009(csa_tree_add_190_195_groupi_n_11898 ,csa_tree_add_190_195_groupi_n_11815 ,csa_tree_add_190_195_groupi_n_11762);
  or csa_tree_add_190_195_groupi_g37010(csa_tree_add_190_195_groupi_n_11897 ,csa_tree_add_190_195_groupi_n_11773 ,csa_tree_add_190_195_groupi_n_11748);
  or csa_tree_add_190_195_groupi_g37011(csa_tree_add_190_195_groupi_n_11896 ,csa_tree_add_190_195_groupi_n_11799 ,csa_tree_add_190_195_groupi_n_11472);
  or csa_tree_add_190_195_groupi_g37012(csa_tree_add_190_195_groupi_n_11895 ,csa_tree_add_190_195_groupi_n_11746 ,csa_tree_add_190_195_groupi_n_11600);
  or csa_tree_add_190_195_groupi_g37013(csa_tree_add_190_195_groupi_n_11894 ,csa_tree_add_190_195_groupi_n_11764 ,csa_tree_add_190_195_groupi_n_11527);
  nor csa_tree_add_190_195_groupi_g37014(csa_tree_add_190_195_groupi_n_11893 ,csa_tree_add_190_195_groupi_n_11753 ,csa_tree_add_190_195_groupi_n_11638);
  or csa_tree_add_190_195_groupi_g37015(csa_tree_add_190_195_groupi_n_11892 ,csa_tree_add_190_195_groupi_n_11754 ,csa_tree_add_190_195_groupi_n_163);
  nor csa_tree_add_190_195_groupi_g37016(csa_tree_add_190_195_groupi_n_11891 ,csa_tree_add_190_195_groupi_n_11640 ,csa_tree_add_190_195_groupi_n_11819);
  and csa_tree_add_190_195_groupi_g37017(csa_tree_add_190_195_groupi_n_11890 ,csa_tree_add_190_195_groupi_n_11813 ,csa_tree_add_190_195_groupi_n_11769);
  or csa_tree_add_190_195_groupi_g37018(csa_tree_add_190_195_groupi_n_11889 ,csa_tree_add_190_195_groupi_n_11639 ,csa_tree_add_190_195_groupi_n_11818);
  or csa_tree_add_190_195_groupi_g37019(csa_tree_add_190_195_groupi_n_11888 ,csa_tree_add_190_195_groupi_n_11523 ,csa_tree_add_190_195_groupi_n_162);
  nor csa_tree_add_190_195_groupi_g37020(csa_tree_add_190_195_groupi_n_11887 ,csa_tree_add_190_195_groupi_n_11812 ,csa_tree_add_190_195_groupi_n_11771);
  or csa_tree_add_190_195_groupi_g37021(csa_tree_add_190_195_groupi_n_11886 ,csa_tree_add_190_195_groupi_n_11808 ,csa_tree_add_190_195_groupi_n_11515);
  and csa_tree_add_190_195_groupi_g37022(csa_tree_add_190_195_groupi_n_11885 ,csa_tree_add_190_195_groupi_n_11808 ,csa_tree_add_190_195_groupi_n_11515);
  or csa_tree_add_190_195_groupi_g37023(csa_tree_add_190_195_groupi_n_11884 ,csa_tree_add_190_195_groupi_n_11811 ,csa_tree_add_190_195_groupi_n_11772);
  nor csa_tree_add_190_195_groupi_g37024(csa_tree_add_190_195_groupi_n_11883 ,csa_tree_add_190_195_groupi_n_11813 ,csa_tree_add_190_195_groupi_n_11769);
  or csa_tree_add_190_195_groupi_g37025(csa_tree_add_190_195_groupi_n_11882 ,csa_tree_add_190_195_groupi_n_11782 ,csa_tree_add_190_195_groupi_n_11716);
  or csa_tree_add_190_195_groupi_g37026(csa_tree_add_190_195_groupi_n_11881 ,csa_tree_add_190_195_groupi_n_11780 ,csa_tree_add_190_195_groupi_n_11593);
  or csa_tree_add_190_195_groupi_g37027(csa_tree_add_190_195_groupi_n_11880 ,csa_tree_add_190_195_groupi_n_11827 ,csa_tree_add_190_195_groupi_n_11788);
  nor csa_tree_add_190_195_groupi_g37028(csa_tree_add_190_195_groupi_n_11879 ,csa_tree_add_190_195_groupi_n_11765 ,csa_tree_add_190_195_groupi_n_11526);
  nor csa_tree_add_190_195_groupi_g37029(csa_tree_add_190_195_groupi_n_11878 ,csa_tree_add_190_195_groupi_n_11766 ,csa_tree_add_190_195_groupi_n_11810);
  or csa_tree_add_190_195_groupi_g37030(csa_tree_add_190_195_groupi_n_11877 ,csa_tree_add_190_195_groupi_n_11767 ,csa_tree_add_190_195_groupi_n_11809);
  and csa_tree_add_190_195_groupi_g37031(csa_tree_add_190_195_groupi_n_11876 ,csa_tree_add_190_195_groupi_n_11378 ,csa_tree_add_190_195_groupi_n_11768);
  or csa_tree_add_190_195_groupi_g37032(csa_tree_add_190_195_groupi_n_11875 ,csa_tree_add_190_195_groupi_n_11378 ,csa_tree_add_190_195_groupi_n_11768);
  or csa_tree_add_190_195_groupi_g37033(csa_tree_add_190_195_groupi_n_11874 ,csa_tree_add_190_195_groupi_n_11717 ,csa_tree_add_190_195_groupi_n_11803);
  or csa_tree_add_190_195_groupi_g37034(csa_tree_add_190_195_groupi_n_11916 ,csa_tree_add_190_195_groupi_n_11680 ,csa_tree_add_190_195_groupi_n_11805);
  or csa_tree_add_190_195_groupi_g37035(csa_tree_add_190_195_groupi_n_11915 ,csa_tree_add_190_195_groupi_n_11687 ,csa_tree_add_190_195_groupi_n_11806);
  and csa_tree_add_190_195_groupi_g37036(csa_tree_add_190_195_groupi_n_11914 ,csa_tree_add_190_195_groupi_n_11790 ,csa_tree_add_190_195_groupi_n_11692);
  and csa_tree_add_190_195_groupi_g37037(csa_tree_add_190_195_groupi_n_11913 ,csa_tree_add_190_195_groupi_n_11697 ,csa_tree_add_190_195_groupi_n_11792);
  or csa_tree_add_190_195_groupi_g37038(csa_tree_add_190_195_groupi_n_11912 ,csa_tree_add_190_195_groupi_n_11801 ,csa_tree_add_190_195_groupi_n_11701);
  or csa_tree_add_190_195_groupi_g37039(csa_tree_add_190_195_groupi_n_11911 ,csa_tree_add_190_195_groupi_n_11784 ,csa_tree_add_190_195_groupi_n_11688);
  and csa_tree_add_190_195_groupi_g37040(csa_tree_add_190_195_groupi_n_11910 ,csa_tree_add_190_195_groupi_n_11802 ,csa_tree_add_190_195_groupi_n_11678);
  and csa_tree_add_190_195_groupi_g37041(csa_tree_add_190_195_groupi_n_11909 ,csa_tree_add_190_195_groupi_n_11682 ,csa_tree_add_190_195_groupi_n_11796);
  or csa_tree_add_190_195_groupi_g37042(csa_tree_add_190_195_groupi_n_11907 ,csa_tree_add_190_195_groupi_n_11700 ,csa_tree_add_190_195_groupi_n_11795);
  or csa_tree_add_190_195_groupi_g37043(csa_tree_add_190_195_groupi_n_11906 ,csa_tree_add_190_195_groupi_n_11783 ,csa_tree_add_190_195_groupi_n_11686);
  or csa_tree_add_190_195_groupi_g37044(csa_tree_add_190_195_groupi_n_11904 ,csa_tree_add_190_195_groupi_n_11797 ,csa_tree_add_190_195_groupi_n_11675);
  and csa_tree_add_190_195_groupi_g37045(csa_tree_add_190_195_groupi_n_11902 ,csa_tree_add_190_195_groupi_n_11674 ,csa_tree_add_190_195_groupi_n_11800);
  not csa_tree_add_190_195_groupi_g37046(csa_tree_add_190_195_groupi_n_11873 ,csa_tree_add_190_195_groupi_n_11872);
  not csa_tree_add_190_195_groupi_g37047(csa_tree_add_190_195_groupi_n_11870 ,csa_tree_add_190_195_groupi_n_11869);
  not csa_tree_add_190_195_groupi_g37048(csa_tree_add_190_195_groupi_n_11866 ,csa_tree_add_190_195_groupi_n_11865);
  not csa_tree_add_190_195_groupi_g37049(csa_tree_add_190_195_groupi_n_11864 ,csa_tree_add_190_195_groupi_n_11863);
  not csa_tree_add_190_195_groupi_g37050(csa_tree_add_190_195_groupi_n_11860 ,csa_tree_add_190_195_groupi_n_11859);
  not csa_tree_add_190_195_groupi_g37051(csa_tree_add_190_195_groupi_n_11857 ,csa_tree_add_190_195_groupi_n_11856);
  not csa_tree_add_190_195_groupi_g37052(csa_tree_add_190_195_groupi_n_11854 ,csa_tree_add_190_195_groupi_n_169);
  not csa_tree_add_190_195_groupi_g37053(csa_tree_add_190_195_groupi_n_11852 ,csa_tree_add_190_195_groupi_n_11851);
  nor csa_tree_add_190_195_groupi_g37054(csa_tree_add_190_195_groupi_n_11849 ,csa_tree_add_190_195_groupi_n_11670 ,csa_tree_add_190_195_groupi_n_11741);
  nor csa_tree_add_190_195_groupi_g37055(csa_tree_add_190_195_groupi_n_11848 ,csa_tree_add_190_195_groupi_n_11636 ,csa_tree_add_190_195_groupi_n_11756);
  or csa_tree_add_190_195_groupi_g37056(csa_tree_add_190_195_groupi_n_11847 ,csa_tree_add_190_195_groupi_n_11627 ,csa_tree_add_190_195_groupi_n_11774);
  or csa_tree_add_190_195_groupi_g37057(csa_tree_add_190_195_groupi_n_11846 ,csa_tree_add_190_195_groupi_n_11635 ,csa_tree_add_190_195_groupi_n_11757);
  or csa_tree_add_190_195_groupi_g37058(csa_tree_add_190_195_groupi_n_11845 ,csa_tree_add_190_195_groupi_n_11742 ,csa_tree_add_190_195_groupi_n_11665);
  xnor csa_tree_add_190_195_groupi_g37059(csa_tree_add_190_195_groupi_n_11844 ,csa_tree_add_190_195_groupi_n_11634 ,csa_tree_add_190_195_groupi_n_11519);
  xnor csa_tree_add_190_195_groupi_g37060(csa_tree_add_190_195_groupi_n_11843 ,csa_tree_add_190_195_groupi_n_11637 ,csa_tree_add_190_195_groupi_n_8314);
  xnor csa_tree_add_190_195_groupi_g37061(csa_tree_add_190_195_groupi_n_11842 ,csa_tree_add_190_195_groupi_n_11653 ,csa_tree_add_190_195_groupi_n_11717);
  xnor csa_tree_add_190_195_groupi_g37062(csa_tree_add_190_195_groupi_n_11841 ,csa_tree_add_190_195_groupi_n_11663 ,csa_tree_add_190_195_groupi_n_11593);
  xnor csa_tree_add_190_195_groupi_g37063(csa_tree_add_190_195_groupi_n_11840 ,csa_tree_add_190_195_groupi_n_11642 ,csa_tree_add_190_195_groupi_n_11531);
  xnor csa_tree_add_190_195_groupi_g37064(csa_tree_add_190_195_groupi_n_11839 ,csa_tree_add_190_195_groupi_n_11652 ,csa_tree_add_190_195_groupi_n_11650);
  xnor csa_tree_add_190_195_groupi_g37066(csa_tree_add_190_195_groupi_n_11838 ,csa_tree_add_190_195_groupi_n_11659 ,csa_tree_add_190_195_groupi_n_11719);
  xor csa_tree_add_190_195_groupi_g37067(csa_tree_add_190_195_groupi_n_11837 ,csa_tree_add_190_195_groupi_n_11720 ,csa_tree_add_190_195_groupi_n_11255);
  xnor csa_tree_add_190_195_groupi_g37068(csa_tree_add_190_195_groupi_n_11836 ,csa_tree_add_190_195_groupi_n_11646 ,csa_tree_add_190_195_groupi_n_11537);
  xnor csa_tree_add_190_195_groupi_g37069(csa_tree_add_190_195_groupi_n_11835 ,csa_tree_add_190_195_groupi_n_11669 ,csa_tree_add_190_195_groupi_n_11025);
  xnor csa_tree_add_190_195_groupi_g37070(csa_tree_add_190_195_groupi_n_11834 ,csa_tree_add_190_195_groupi_n_11655 ,csa_tree_add_190_195_groupi_n_11581);
  xnor csa_tree_add_190_195_groupi_g37071(csa_tree_add_190_195_groupi_n_11833 ,csa_tree_add_190_195_groupi_n_11668 ,csa_tree_add_190_195_groupi_n_11393);
  xnor csa_tree_add_190_195_groupi_g37072(csa_tree_add_190_195_groupi_n_11832 ,csa_tree_add_190_195_groupi_n_11666 ,csa_tree_add_190_195_groupi_n_11533);
  xnor csa_tree_add_190_195_groupi_g37073(csa_tree_add_190_195_groupi_n_11831 ,csa_tree_add_190_195_groupi_n_11641 ,csa_tree_add_190_195_groupi_n_11459);
  xnor csa_tree_add_190_195_groupi_g37074(csa_tree_add_190_195_groupi_n_11830 ,csa_tree_add_190_195_groupi_n_11588 ,csa_tree_add_190_195_groupi_n_11664);
  xnor csa_tree_add_190_195_groupi_g37075(csa_tree_add_190_195_groupi_n_11829 ,csa_tree_add_190_195_groupi_n_11657 ,csa_tree_add_190_195_groupi_n_11579);
  xnor csa_tree_add_190_195_groupi_g37076(csa_tree_add_190_195_groupi_n_11828 ,csa_tree_add_190_195_groupi_n_11406 ,csa_tree_add_190_195_groupi_n_11715);
  xnor csa_tree_add_190_195_groupi_g37077(csa_tree_add_190_195_groupi_n_11872 ,csa_tree_add_190_195_groupi_n_11327 ,csa_tree_add_190_195_groupi_n_11609);
  and csa_tree_add_190_195_groupi_g37078(csa_tree_add_190_195_groupi_n_11871 ,csa_tree_add_190_195_groupi_n_11743 ,csa_tree_add_190_195_groupi_n_11621);
  or csa_tree_add_190_195_groupi_g37079(csa_tree_add_190_195_groupi_n_11869 ,csa_tree_add_190_195_groupi_n_11625 ,csa_tree_add_190_195_groupi_n_11740);
  xnor csa_tree_add_190_195_groupi_g37080(csa_tree_add_190_195_groupi_n_11868 ,csa_tree_add_190_195_groupi_n_11540 ,csa_tree_add_190_195_groupi_n_11607);
  xnor csa_tree_add_190_195_groupi_g37081(csa_tree_add_190_195_groupi_n_11867 ,csa_tree_add_190_195_groupi_n_11474 ,csa_tree_add_190_195_groupi_n_11613);
  xnor csa_tree_add_190_195_groupi_g37082(csa_tree_add_190_195_groupi_n_11865 ,csa_tree_add_190_195_groupi_n_11382 ,csa_tree_add_190_195_groupi_n_11619);
  xnor csa_tree_add_190_195_groupi_g37083(csa_tree_add_190_195_groupi_n_11863 ,csa_tree_add_190_195_groupi_n_11385 ,csa_tree_add_190_195_groupi_n_11614);
  xnor csa_tree_add_190_195_groupi_g37084(csa_tree_add_190_195_groupi_n_11862 ,csa_tree_add_190_195_groupi_n_11260 ,csa_tree_add_190_195_groupi_n_11612);
  xnor csa_tree_add_190_195_groupi_g37085(csa_tree_add_190_195_groupi_n_11861 ,csa_tree_add_190_195_groupi_n_11464 ,csa_tree_add_190_195_groupi_n_11616);
  xnor csa_tree_add_190_195_groupi_g37086(csa_tree_add_190_195_groupi_n_11859 ,csa_tree_add_190_195_groupi_n_11398 ,csa_tree_add_190_195_groupi_n_11617);
  xnor csa_tree_add_190_195_groupi_g37087(csa_tree_add_190_195_groupi_n_11858 ,csa_tree_add_190_195_groupi_n_11544 ,csa_tree_add_190_195_groupi_n_11618);
  xnor csa_tree_add_190_195_groupi_g37088(csa_tree_add_190_195_groupi_n_11856 ,csa_tree_add_190_195_groupi_n_11232 ,csa_tree_add_190_195_groupi_n_11620);
  xnor csa_tree_add_190_195_groupi_g37089(csa_tree_add_190_195_groupi_n_11855 ,csa_tree_add_190_195_groupi_n_11384 ,csa_tree_add_190_195_groupi_n_11615);
  xnor csa_tree_add_190_195_groupi_g37091(csa_tree_add_190_195_groupi_n_11853 ,csa_tree_add_190_195_groupi_n_11036 ,csa_tree_add_190_195_groupi_n_166);
  xnor csa_tree_add_190_195_groupi_g37092(csa_tree_add_190_195_groupi_n_11851 ,csa_tree_add_190_195_groupi_n_11468 ,csa_tree_add_190_195_groupi_n_11610);
  xnor csa_tree_add_190_195_groupi_g37093(csa_tree_add_190_195_groupi_n_11850 ,csa_tree_add_190_195_groupi_n_11603 ,csa_tree_add_190_195_groupi_n_11608);
  not csa_tree_add_190_195_groupi_g37096(csa_tree_add_190_195_groupi_n_11819 ,csa_tree_add_190_195_groupi_n_11818);
  not csa_tree_add_190_195_groupi_g37097(csa_tree_add_190_195_groupi_n_11816 ,csa_tree_add_190_195_groupi_n_11817);
  not csa_tree_add_190_195_groupi_g37098(csa_tree_add_190_195_groupi_n_11812 ,csa_tree_add_190_195_groupi_n_11811);
  not csa_tree_add_190_195_groupi_g37099(csa_tree_add_190_195_groupi_n_11809 ,csa_tree_add_190_195_groupi_n_11810);
  or csa_tree_add_190_195_groupi_g37100(csa_tree_add_190_195_groupi_n_11807 ,csa_tree_add_190_195_groupi_n_11656 ,csa_tree_add_190_195_groupi_n_11578);
  nor csa_tree_add_190_195_groupi_g37101(csa_tree_add_190_195_groupi_n_11806 ,csa_tree_add_190_195_groupi_n_11668 ,csa_tree_add_190_195_groupi_n_11711);
  and csa_tree_add_190_195_groupi_g37102(csa_tree_add_190_195_groupi_n_11805 ,csa_tree_add_190_195_groupi_n_11339 ,csa_tree_add_190_195_groupi_n_11677);
  or csa_tree_add_190_195_groupi_g37103(csa_tree_add_190_195_groupi_n_11804 ,csa_tree_add_190_195_groupi_n_11713 ,csa_tree_add_190_195_groupi_n_11653);
  and csa_tree_add_190_195_groupi_g37104(csa_tree_add_190_195_groupi_n_11803 ,csa_tree_add_190_195_groupi_n_11713 ,csa_tree_add_190_195_groupi_n_11653);
  or csa_tree_add_190_195_groupi_g37105(csa_tree_add_190_195_groupi_n_11802 ,csa_tree_add_190_195_groupi_n_11672 ,csa_tree_add_190_195_groupi_n_11598);
  and csa_tree_add_190_195_groupi_g37106(csa_tree_add_190_195_groupi_n_11801 ,csa_tree_add_190_195_groupi_n_11595 ,csa_tree_add_190_195_groupi_n_11702);
  or csa_tree_add_190_195_groupi_g37107(csa_tree_add_190_195_groupi_n_11800 ,csa_tree_add_190_195_groupi_n_11596 ,csa_tree_add_190_195_groupi_n_11673);
  and csa_tree_add_190_195_groupi_g37108(csa_tree_add_190_195_groupi_n_11799 ,csa_tree_add_190_195_groupi_n_11459 ,csa_tree_add_190_195_groupi_n_11641);
  or csa_tree_add_190_195_groupi_g37109(csa_tree_add_190_195_groupi_n_11798 ,csa_tree_add_190_195_groupi_n_11459 ,csa_tree_add_190_195_groupi_n_11641);
  nor csa_tree_add_190_195_groupi_g37110(csa_tree_add_190_195_groupi_n_11797 ,csa_tree_add_190_195_groupi_n_11676 ,csa_tree_add_190_195_groupi_n_11604);
  or csa_tree_add_190_195_groupi_g37111(csa_tree_add_190_195_groupi_n_11796 ,csa_tree_add_190_195_groupi_n_11679 ,csa_tree_add_190_195_groupi_n_11718);
  nor csa_tree_add_190_195_groupi_g37112(csa_tree_add_190_195_groupi_n_11795 ,csa_tree_add_190_195_groupi_n_11699 ,csa_tree_add_190_195_groupi_n_11599);
  nor csa_tree_add_190_195_groupi_g37113(csa_tree_add_190_195_groupi_n_11794 ,csa_tree_add_190_195_groupi_n_11587 ,csa_tree_add_190_195_groupi_n_11664);
  or csa_tree_add_190_195_groupi_g37114(csa_tree_add_190_195_groupi_n_11793 ,csa_tree_add_190_195_groupi_n_11406 ,csa_tree_add_190_195_groupi_n_11714);
  or csa_tree_add_190_195_groupi_g37115(csa_tree_add_190_195_groupi_n_11792 ,csa_tree_add_190_195_groupi_n_11696 ,csa_tree_add_190_195_groupi_n_11602);
  nor csa_tree_add_190_195_groupi_g37116(csa_tree_add_190_195_groupi_n_11791 ,csa_tree_add_190_195_groupi_n_8313 ,csa_tree_add_190_195_groupi_n_11637);
  or csa_tree_add_190_195_groupi_g37117(csa_tree_add_190_195_groupi_n_11790 ,csa_tree_add_190_195_groupi_n_11667 ,csa_tree_add_190_195_groupi_n_11693);
  nor csa_tree_add_190_195_groupi_g37118(csa_tree_add_190_195_groupi_n_11789 ,csa_tree_add_190_195_groupi_n_11405 ,csa_tree_add_190_195_groupi_n_11715);
  nor csa_tree_add_190_195_groupi_g37119(csa_tree_add_190_195_groupi_n_11788 ,csa_tree_add_190_195_groupi_n_11648 ,csa_tree_add_190_195_groupi_n_11643);
  or csa_tree_add_190_195_groupi_g37120(csa_tree_add_190_195_groupi_n_11787 ,csa_tree_add_190_195_groupi_n_11588 ,csa_tree_add_190_195_groupi_n_158);
  or csa_tree_add_190_195_groupi_g37121(csa_tree_add_190_195_groupi_n_11786 ,csa_tree_add_190_195_groupi_n_11654 ,csa_tree_add_190_195_groupi_n_11581);
  nor csa_tree_add_190_195_groupi_g37122(csa_tree_add_190_195_groupi_n_11785 ,csa_tree_add_190_195_groupi_n_11655 ,csa_tree_add_190_195_groupi_n_11580);
  and csa_tree_add_190_195_groupi_g37123(csa_tree_add_190_195_groupi_n_11784 ,csa_tree_add_190_195_groupi_n_11606 ,csa_tree_add_190_195_groupi_n_11694);
  nor csa_tree_add_190_195_groupi_g37124(csa_tree_add_190_195_groupi_n_11783 ,csa_tree_add_190_195_groupi_n_11478 ,csa_tree_add_190_195_groupi_n_11712);
  nor csa_tree_add_190_195_groupi_g37125(csa_tree_add_190_195_groupi_n_11782 ,csa_tree_add_190_195_groupi_n_11657 ,csa_tree_add_190_195_groupi_n_11579);
  or csa_tree_add_190_195_groupi_g37126(csa_tree_add_190_195_groupi_n_11781 ,csa_tree_add_190_195_groupi_n_11660 ,csa_tree_add_190_195_groupi_n_11663);
  and csa_tree_add_190_195_groupi_g37127(csa_tree_add_190_195_groupi_n_11780 ,csa_tree_add_190_195_groupi_n_11660 ,csa_tree_add_190_195_groupi_n_11663);
  or csa_tree_add_190_195_groupi_g37128(csa_tree_add_190_195_groupi_n_11779 ,csa_tree_add_190_195_groupi_n_11633 ,csa_tree_add_190_195_groupi_n_11519);
  nor csa_tree_add_190_195_groupi_g37129(csa_tree_add_190_195_groupi_n_11778 ,csa_tree_add_190_195_groupi_n_11634 ,csa_tree_add_190_195_groupi_n_11518);
  or csa_tree_add_190_195_groupi_g37130(csa_tree_add_190_195_groupi_n_11777 ,csa_tree_add_190_195_groupi_n_157 ,csa_tree_add_190_195_groupi_n_11644);
  and csa_tree_add_190_195_groupi_g37131(csa_tree_add_190_195_groupi_n_11827 ,csa_tree_add_190_195_groupi_n_11685 ,csa_tree_add_190_195_groupi_n_11549);
  and csa_tree_add_190_195_groupi_g37132(csa_tree_add_190_195_groupi_n_11826 ,csa_tree_add_190_195_groupi_n_11690 ,csa_tree_add_190_195_groupi_n_11411);
  and csa_tree_add_190_195_groupi_g37133(csa_tree_add_190_195_groupi_n_11825 ,csa_tree_add_190_195_groupi_n_11705 ,csa_tree_add_190_195_groupi_n_11502);
  and csa_tree_add_190_195_groupi_g37134(csa_tree_add_190_195_groupi_n_11824 ,csa_tree_add_190_195_groupi_n_11568 ,csa_tree_add_190_195_groupi_n_11706);
  and csa_tree_add_190_195_groupi_g37135(csa_tree_add_190_195_groupi_n_11823 ,csa_tree_add_190_195_groupi_n_11709 ,csa_tree_add_190_195_groupi_n_11570);
  or csa_tree_add_190_195_groupi_g37136(csa_tree_add_190_195_groupi_n_11822 ,csa_tree_add_190_195_groupi_n_11572 ,csa_tree_add_190_195_groupi_n_11707);
  and csa_tree_add_190_195_groupi_g37137(csa_tree_add_190_195_groupi_n_11821 ,csa_tree_add_190_195_groupi_n_11548 ,csa_tree_add_190_195_groupi_n_11684);
  and csa_tree_add_190_195_groupi_g37138(csa_tree_add_190_195_groupi_n_11820 ,csa_tree_add_190_195_groupi_n_11427 ,csa_tree_add_190_195_groupi_n_11671);
  and csa_tree_add_190_195_groupi_g37139(csa_tree_add_190_195_groupi_n_11818 ,csa_tree_add_190_195_groupi_n_11563 ,csa_tree_add_190_195_groupi_n_11698);
  and csa_tree_add_190_195_groupi_g37140(csa_tree_add_190_195_groupi_n_11817 ,csa_tree_add_190_195_groupi_n_11703 ,csa_tree_add_190_195_groupi_n_11500);
  and csa_tree_add_190_195_groupi_g37141(csa_tree_add_190_195_groupi_n_11815 ,csa_tree_add_190_195_groupi_n_11562 ,csa_tree_add_190_195_groupi_n_11710);
  or csa_tree_add_190_195_groupi_g37142(csa_tree_add_190_195_groupi_n_11814 ,csa_tree_add_190_195_groupi_n_11552 ,csa_tree_add_190_195_groupi_n_11689);
  or csa_tree_add_190_195_groupi_g37143(csa_tree_add_190_195_groupi_n_11813 ,csa_tree_add_190_195_groupi_n_11683 ,csa_tree_add_190_195_groupi_n_11576);
  and csa_tree_add_190_195_groupi_g37144(csa_tree_add_190_195_groupi_n_11811 ,csa_tree_add_190_195_groupi_n_11555 ,csa_tree_add_190_195_groupi_n_11691);
  or csa_tree_add_190_195_groupi_g37145(csa_tree_add_190_195_groupi_n_11810 ,csa_tree_add_190_195_groupi_n_11553 ,csa_tree_add_190_195_groupi_n_11681);
  and csa_tree_add_190_195_groupi_g37146(csa_tree_add_190_195_groupi_n_11808 ,csa_tree_add_190_195_groupi_n_11561 ,csa_tree_add_190_195_groupi_n_11695);
  not csa_tree_add_190_195_groupi_g37147(csa_tree_add_190_195_groupi_n_11772 ,csa_tree_add_190_195_groupi_n_11771);
  not csa_tree_add_190_195_groupi_g37148(csa_tree_add_190_195_groupi_n_11770 ,csa_tree_add_190_195_groupi_n_162);
  not csa_tree_add_190_195_groupi_g37149(csa_tree_add_190_195_groupi_n_11767 ,csa_tree_add_190_195_groupi_n_11766);
  not csa_tree_add_190_195_groupi_g37150(csa_tree_add_190_195_groupi_n_11765 ,csa_tree_add_190_195_groupi_n_11764);
  not csa_tree_add_190_195_groupi_g37151(csa_tree_add_190_195_groupi_n_11760 ,csa_tree_add_190_195_groupi_n_11759);
  not csa_tree_add_190_195_groupi_g37152(csa_tree_add_190_195_groupi_n_11758 ,csa_tree_add_190_195_groupi_n_168);
  not csa_tree_add_190_195_groupi_g37153(csa_tree_add_190_195_groupi_n_11757 ,csa_tree_add_190_195_groupi_n_11756);
  not csa_tree_add_190_195_groupi_g37154(csa_tree_add_190_195_groupi_n_11754 ,csa_tree_add_190_195_groupi_n_11753);
  not csa_tree_add_190_195_groupi_g37155(csa_tree_add_190_195_groupi_n_11752 ,csa_tree_add_190_195_groupi_n_11751);
  or csa_tree_add_190_195_groupi_g37156(csa_tree_add_190_195_groupi_n_11750 ,csa_tree_add_190_195_groupi_n_11652 ,csa_tree_add_190_195_groupi_n_11649);
  nor csa_tree_add_190_195_groupi_g37157(csa_tree_add_190_195_groupi_n_11749 ,csa_tree_add_190_195_groupi_n_11026 ,csa_tree_add_190_195_groupi_n_11632);
  nor csa_tree_add_190_195_groupi_g37158(csa_tree_add_190_195_groupi_n_11748 ,csa_tree_add_190_195_groupi_n_11651 ,csa_tree_add_190_195_groupi_n_11650);
  or csa_tree_add_190_195_groupi_g37159(csa_tree_add_190_195_groupi_n_11747 ,csa_tree_add_190_195_groupi_n_11647 ,csa_tree_add_190_195_groupi_n_11399);
  and csa_tree_add_190_195_groupi_g37160(csa_tree_add_190_195_groupi_n_11746 ,csa_tree_add_190_195_groupi_n_11647 ,csa_tree_add_190_195_groupi_n_11399);
  or csa_tree_add_190_195_groupi_g37161(csa_tree_add_190_195_groupi_n_11745 ,csa_tree_add_190_195_groupi_n_11645 ,csa_tree_add_190_195_groupi_n_11536);
  nor csa_tree_add_190_195_groupi_g37162(csa_tree_add_190_195_groupi_n_11744 ,csa_tree_add_190_195_groupi_n_11642 ,csa_tree_add_190_195_groupi_n_11531);
  or csa_tree_add_190_195_groupi_g37163(csa_tree_add_190_195_groupi_n_11743 ,csa_tree_add_190_195_groupi_n_11708 ,csa_tree_add_190_195_groupi_n_11539);
  nor csa_tree_add_190_195_groupi_g37164(csa_tree_add_190_195_groupi_n_11742 ,csa_tree_add_190_195_groupi_n_11646 ,csa_tree_add_190_195_groupi_n_11537);
  and csa_tree_add_190_195_groupi_g37165(csa_tree_add_190_195_groupi_n_11741 ,csa_tree_add_190_195_groupi_n_11026 ,csa_tree_add_190_195_groupi_n_11632);
  nor csa_tree_add_190_195_groupi_g37166(csa_tree_add_190_195_groupi_n_11740 ,csa_tree_add_190_195_groupi_n_11541 ,csa_tree_add_190_195_groupi_n_11622);
  and csa_tree_add_190_195_groupi_g37167(csa_tree_add_190_195_groupi_n_11739 ,csa_tree_add_190_195_groupi_n_1332 ,csa_tree_add_190_195_groupi_n_11637);
  or csa_tree_add_190_195_groupi_g37168(csa_tree_add_190_195_groupi_n_11738 ,csa_tree_add_190_195_groupi_n_167 ,csa_tree_add_190_195_groupi_n_11530);
  xnor csa_tree_add_190_195_groupi_g37169(csa_tree_add_190_195_groupi_n_11737 ,csa_tree_add_190_195_groupi_n_11591 ,csa_tree_add_190_195_groupi_n_11251);
  xnor csa_tree_add_190_195_groupi_g37170(csa_tree_add_190_195_groupi_n_11736 ,csa_tree_add_190_195_groupi_n_11529 ,csa_tree_add_190_195_groupi_n_11380);
  xnor csa_tree_add_190_195_groupi_g37171(csa_tree_add_190_195_groupi_n_11735 ,csa_tree_add_190_195_groupi_n_11601 ,csa_tree_add_190_195_groupi_n_11515);
  xnor csa_tree_add_190_195_groupi_g37172(csa_tree_add_190_195_groupi_n_11734 ,csa_tree_add_190_195_groupi_n_11583 ,csa_tree_add_190_195_groupi_n_11517);
  xnor csa_tree_add_190_195_groupi_g37173(csa_tree_add_190_195_groupi_n_11733 ,csa_tree_add_190_195_groupi_n_11261 ,csa_tree_add_190_195_groupi_n_11599);
  xnor csa_tree_add_190_195_groupi_g37174(csa_tree_add_190_195_groupi_n_11732 ,csa_tree_add_190_195_groupi_n_11331 ,csa_tree_add_190_195_groupi_n_11508);
  xnor csa_tree_add_190_195_groupi_g37175(csa_tree_add_190_195_groupi_n_11731 ,csa_tree_add_190_195_groupi_n_11600 ,csa_tree_add_190_195_groupi_n_11399);
  xnor csa_tree_add_190_195_groupi_g37176(csa_tree_add_190_195_groupi_n_11730 ,csa_tree_add_190_195_groupi_n_11449 ,csa_tree_add_190_195_groupi_n_11602);
  xnor csa_tree_add_190_195_groupi_g37177(csa_tree_add_190_195_groupi_n_11729 ,csa_tree_add_190_195_groupi_n_11525 ,csa_tree_add_190_195_groupi_n_11452);
  xnor csa_tree_add_190_195_groupi_g37178(csa_tree_add_190_195_groupi_n_11728 ,csa_tree_add_190_195_groupi_n_11586 ,csa_tree_add_190_195_groupi_n_11606);
  xnor csa_tree_add_190_195_groupi_g37179(csa_tree_add_190_195_groupi_n_11727 ,csa_tree_add_190_195_groupi_n_11256 ,csa_tree_add_190_195_groupi_n_11520);
  xnor csa_tree_add_190_195_groupi_g37180(csa_tree_add_190_195_groupi_n_11726 ,csa_tree_add_190_195_groupi_n_11535 ,csa_tree_add_190_195_groupi_n_11377);
  xor csa_tree_add_190_195_groupi_g37181(csa_tree_add_190_195_groupi_n_11725 ,csa_tree_add_190_195_groupi_n_11594 ,csa_tree_add_190_195_groupi_n_11378);
  xnor csa_tree_add_190_195_groupi_g37182(csa_tree_add_190_195_groupi_n_11724 ,csa_tree_add_190_195_groupi_n_11512 ,csa_tree_add_190_195_groupi_n_11458);
  xnor csa_tree_add_190_195_groupi_g37183(csa_tree_add_190_195_groupi_n_11723 ,csa_tree_add_190_195_groupi_n_11240 ,csa_tree_add_190_195_groupi_n_11604);
  xnor csa_tree_add_190_195_groupi_g37184(csa_tree_add_190_195_groupi_n_11722 ,csa_tree_add_190_195_groupi_n_11239 ,csa_tree_add_190_195_groupi_n_11513);
  xnor csa_tree_add_190_195_groupi_g37185(csa_tree_add_190_195_groupi_n_11776 ,csa_tree_add_190_195_groupi_n_11151 ,csa_tree_add_190_195_groupi_n_164);
  and csa_tree_add_190_195_groupi_g37186(csa_tree_add_190_195_groupi_n_11775 ,csa_tree_add_190_195_groupi_n_11494 ,csa_tree_add_190_195_groupi_n_11624);
  and csa_tree_add_190_195_groupi_g37187(csa_tree_add_190_195_groupi_n_11774 ,csa_tree_add_190_195_groupi_n_11626 ,csa_tree_add_190_195_groupi_n_11498);
  and csa_tree_add_190_195_groupi_g37188(csa_tree_add_190_195_groupi_n_11773 ,csa_tree_add_190_195_groupi_n_11497 ,csa_tree_add_190_195_groupi_n_11704);
  xnor csa_tree_add_190_195_groupi_g37189(csa_tree_add_190_195_groupi_n_11771 ,csa_tree_add_190_195_groupi_n_11387 ,csa_tree_add_190_195_groupi_n_11491);
  xnor csa_tree_add_190_195_groupi_g37191(csa_tree_add_190_195_groupi_n_11769 ,csa_tree_add_190_195_groupi_n_11469 ,csa_tree_add_190_195_groupi_n_11483);
  xnor csa_tree_add_190_195_groupi_g37192(csa_tree_add_190_195_groupi_n_11768 ,csa_tree_add_190_195_groupi_n_11071 ,csa_tree_add_190_195_groupi_n_165);
  xnor csa_tree_add_190_195_groupi_g37193(csa_tree_add_190_195_groupi_n_11766 ,csa_tree_add_190_195_groupi_n_11605 ,csa_tree_add_190_195_groupi_n_11488);
  xnor csa_tree_add_190_195_groupi_g37194(csa_tree_add_190_195_groupi_n_11764 ,csa_tree_add_190_195_groupi_n_10969 ,csa_tree_add_190_195_groupi_n_11487);
  xnor csa_tree_add_190_195_groupi_g37195(csa_tree_add_190_195_groupi_n_11763 ,csa_tree_add_190_195_groupi_n_11038 ,csa_tree_add_190_195_groupi_n_11490);
  xnor csa_tree_add_190_195_groupi_g37196(csa_tree_add_190_195_groupi_n_11762 ,csa_tree_add_190_195_groupi_n_10845 ,csa_tree_add_190_195_groupi_n_11485);
  xnor csa_tree_add_190_195_groupi_g37197(csa_tree_add_190_195_groupi_n_11761 ,csa_tree_add_190_195_groupi_n_11392 ,csa_tree_add_190_195_groupi_n_11482);
  xnor csa_tree_add_190_195_groupi_g37198(csa_tree_add_190_195_groupi_n_11759 ,csa_tree_add_190_195_groupi_n_11389 ,csa_tree_add_190_195_groupi_n_11486);
  xnor csa_tree_add_190_195_groupi_g37200(csa_tree_add_190_195_groupi_n_11756 ,csa_tree_add_190_195_groupi_n_11542 ,csa_tree_add_190_195_groupi_n_11481);
  xnor csa_tree_add_190_195_groupi_g37201(csa_tree_add_190_195_groupi_n_11755 ,csa_tree_add_190_195_groupi_n_153 ,csa_tree_add_190_195_groupi_n_11480);
  xnor csa_tree_add_190_195_groupi_g37202(csa_tree_add_190_195_groupi_n_11753 ,csa_tree_add_190_195_groupi_n_11262 ,csa_tree_add_190_195_groupi_n_11489);
  and csa_tree_add_190_195_groupi_g37203(csa_tree_add_190_195_groupi_n_11751 ,csa_tree_add_190_195_groupi_n_11623 ,csa_tree_add_190_195_groupi_n_11367);
  not csa_tree_add_190_195_groupi_g37205(csa_tree_add_190_195_groupi_n_11715 ,csa_tree_add_190_195_groupi_n_11714);
  nor csa_tree_add_190_195_groupi_g37206(csa_tree_add_190_195_groupi_n_11712 ,csa_tree_add_190_195_groupi_n_11256 ,csa_tree_add_190_195_groupi_n_11520);
  and csa_tree_add_190_195_groupi_g37207(csa_tree_add_190_195_groupi_n_11711 ,csa_tree_add_190_195_groupi_n_11394 ,csa_tree_add_190_195_groupi_n_11584);
  or csa_tree_add_190_195_groupi_g37208(csa_tree_add_190_195_groupi_n_11710 ,csa_tree_add_190_195_groupi_n_11178 ,csa_tree_add_190_195_groupi_n_11564);
  or csa_tree_add_190_195_groupi_g37209(csa_tree_add_190_195_groupi_n_11709 ,csa_tree_add_190_195_groupi_n_11467 ,csa_tree_add_190_195_groupi_n_11571);
  nor csa_tree_add_190_195_groupi_g37210(csa_tree_add_190_195_groupi_n_11708 ,csa_tree_add_190_195_groupi_n_11583 ,csa_tree_add_190_195_groupi_n_11517);
  nor csa_tree_add_190_195_groupi_g37211(csa_tree_add_190_195_groupi_n_11707 ,csa_tree_add_190_195_groupi_n_11408 ,csa_tree_add_190_195_groupi_n_11554);
  or csa_tree_add_190_195_groupi_g37212(csa_tree_add_190_195_groupi_n_11706 ,csa_tree_add_190_195_groupi_n_11336 ,csa_tree_add_190_195_groupi_n_11556);
  or csa_tree_add_190_195_groupi_g37213(csa_tree_add_190_195_groupi_n_11705 ,csa_tree_add_190_195_groupi_n_11503 ,csa_tree_add_190_195_groupi_n_11465);
  or csa_tree_add_190_195_groupi_g37214(csa_tree_add_190_195_groupi_n_11704 ,csa_tree_add_190_195_groupi_n_11464 ,csa_tree_add_190_195_groupi_n_11504);
  or csa_tree_add_190_195_groupi_g37215(csa_tree_add_190_195_groupi_n_11703 ,csa_tree_add_190_195_groupi_n_11501 ,csa_tree_add_190_195_groupi_n_11337);
  or csa_tree_add_190_195_groupi_g37216(csa_tree_add_190_195_groupi_n_11702 ,csa_tree_add_190_195_groupi_n_11331 ,csa_tree_add_190_195_groupi_n_11507);
  nor csa_tree_add_190_195_groupi_g37217(csa_tree_add_190_195_groupi_n_11701 ,csa_tree_add_190_195_groupi_n_11330 ,csa_tree_add_190_195_groupi_n_11508);
  and csa_tree_add_190_195_groupi_g37218(csa_tree_add_190_195_groupi_n_11700 ,csa_tree_add_190_195_groupi_n_11261 ,csa_tree_add_190_195_groupi_n_11521);
  nor csa_tree_add_190_195_groupi_g37219(csa_tree_add_190_195_groupi_n_11699 ,csa_tree_add_190_195_groupi_n_11261 ,csa_tree_add_190_195_groupi_n_11521);
  or csa_tree_add_190_195_groupi_g37220(csa_tree_add_190_195_groupi_n_11698 ,csa_tree_add_190_195_groupi_n_11172 ,csa_tree_add_190_195_groupi_n_11560);
  or csa_tree_add_190_195_groupi_g37221(csa_tree_add_190_195_groupi_n_11697 ,csa_tree_add_190_195_groupi_n_11449 ,csa_tree_add_190_195_groupi_n_11505);
  nor csa_tree_add_190_195_groupi_g37222(csa_tree_add_190_195_groupi_n_11696 ,csa_tree_add_190_195_groupi_n_11448 ,csa_tree_add_190_195_groupi_n_11506);
  or csa_tree_add_190_195_groupi_g37223(csa_tree_add_190_195_groupi_n_11695 ,csa_tree_add_190_195_groupi_n_11558 ,csa_tree_add_190_195_groupi_n_11603);
  or csa_tree_add_190_195_groupi_g37224(csa_tree_add_190_195_groupi_n_11694 ,csa_tree_add_190_195_groupi_n_11241 ,csa_tree_add_190_195_groupi_n_11585);
  nor csa_tree_add_190_195_groupi_g37225(csa_tree_add_190_195_groupi_n_11693 ,csa_tree_add_190_195_groupi_n_11533 ,csa_tree_add_190_195_groupi_n_11590);
  or csa_tree_add_190_195_groupi_g37226(csa_tree_add_190_195_groupi_n_11692 ,csa_tree_add_190_195_groupi_n_11532 ,csa_tree_add_190_195_groupi_n_11589);
  or csa_tree_add_190_195_groupi_g37227(csa_tree_add_190_195_groupi_n_11691 ,csa_tree_add_190_195_groupi_n_11540 ,csa_tree_add_190_195_groupi_n_11577);
  or csa_tree_add_190_195_groupi_g37228(csa_tree_add_190_195_groupi_n_11690 ,csa_tree_add_190_195_groupi_n_11605 ,csa_tree_add_190_195_groupi_n_11413);
  nor csa_tree_add_190_195_groupi_g37229(csa_tree_add_190_195_groupi_n_11689 ,csa_tree_add_190_195_groupi_n_11474 ,csa_tree_add_190_195_groupi_n_11551);
  nor csa_tree_add_190_195_groupi_g37230(csa_tree_add_190_195_groupi_n_11688 ,csa_tree_add_190_195_groupi_n_151 ,csa_tree_add_190_195_groupi_n_11586);
  nor csa_tree_add_190_195_groupi_g37231(csa_tree_add_190_195_groupi_n_11687 ,csa_tree_add_190_195_groupi_n_11394 ,csa_tree_add_190_195_groupi_n_11584);
  and csa_tree_add_190_195_groupi_g37232(csa_tree_add_190_195_groupi_n_11686 ,csa_tree_add_190_195_groupi_n_11256 ,csa_tree_add_190_195_groupi_n_11520);
  or csa_tree_add_190_195_groupi_g37233(csa_tree_add_190_195_groupi_n_11685 ,csa_tree_add_190_195_groupi_n_11477 ,csa_tree_add_190_195_groupi_n_11550);
  or csa_tree_add_190_195_groupi_g37234(csa_tree_add_190_195_groupi_n_11684 ,csa_tree_add_190_195_groupi_n_11592 ,csa_tree_add_190_195_groupi_n_11547);
  nor csa_tree_add_190_195_groupi_g37235(csa_tree_add_190_195_groupi_n_11683 ,csa_tree_add_190_195_groupi_n_11573 ,csa_tree_add_190_195_groupi_n_11410);
  or csa_tree_add_190_195_groupi_g37236(csa_tree_add_190_195_groupi_n_11682 ,csa_tree_add_190_195_groupi_n_159 ,csa_tree_add_190_195_groupi_n_11450);
  nor csa_tree_add_190_195_groupi_g37237(csa_tree_add_190_195_groupi_n_11681 ,csa_tree_add_190_195_groupi_n_11557 ,csa_tree_add_190_195_groupi_n_11468);
  nor csa_tree_add_190_195_groupi_g37238(csa_tree_add_190_195_groupi_n_11680 ,csa_tree_add_190_195_groupi_n_11512 ,csa_tree_add_190_195_groupi_n_11457);
  and csa_tree_add_190_195_groupi_g37239(csa_tree_add_190_195_groupi_n_11679 ,csa_tree_add_190_195_groupi_n_159 ,csa_tree_add_190_195_groupi_n_11450);
  or csa_tree_add_190_195_groupi_g37240(csa_tree_add_190_195_groupi_n_11678 ,csa_tree_add_190_195_groupi_n_11524 ,csa_tree_add_190_195_groupi_n_11451);
  or csa_tree_add_190_195_groupi_g37241(csa_tree_add_190_195_groupi_n_11677 ,csa_tree_add_190_195_groupi_n_11511 ,csa_tree_add_190_195_groupi_n_11458);
  and csa_tree_add_190_195_groupi_g37242(csa_tree_add_190_195_groupi_n_11676 ,csa_tree_add_190_195_groupi_n_11240 ,csa_tree_add_190_195_groupi_n_11510);
  nor csa_tree_add_190_195_groupi_g37243(csa_tree_add_190_195_groupi_n_11675 ,csa_tree_add_190_195_groupi_n_11240 ,csa_tree_add_190_195_groupi_n_11510);
  or csa_tree_add_190_195_groupi_g37244(csa_tree_add_190_195_groupi_n_11674 ,csa_tree_add_190_195_groupi_n_11535 ,csa_tree_add_190_195_groupi_n_11376);
  nor csa_tree_add_190_195_groupi_g37245(csa_tree_add_190_195_groupi_n_11673 ,csa_tree_add_190_195_groupi_n_11534 ,csa_tree_add_190_195_groupi_n_11377);
  nor csa_tree_add_190_195_groupi_g37246(csa_tree_add_190_195_groupi_n_11672 ,csa_tree_add_190_195_groupi_n_11525 ,csa_tree_add_190_195_groupi_n_11452);
  or csa_tree_add_190_195_groupi_g37247(csa_tree_add_190_195_groupi_n_11671 ,csa_tree_add_190_195_groupi_n_11437 ,csa_tree_add_190_195_groupi_n_11543);
  and csa_tree_add_190_195_groupi_g37248(csa_tree_add_190_195_groupi_n_11721 ,csa_tree_add_190_195_groupi_n_11373 ,csa_tree_add_190_195_groupi_n_11574);
  and csa_tree_add_190_195_groupi_g37249(csa_tree_add_190_195_groupi_n_11720 ,csa_tree_add_190_195_groupi_n_11433 ,csa_tree_add_190_195_groupi_n_11575);
  and csa_tree_add_190_195_groupi_g37250(csa_tree_add_190_195_groupi_n_11719 ,csa_tree_add_190_195_groupi_n_11436 ,csa_tree_add_190_195_groupi_n_11566);
  and csa_tree_add_190_195_groupi_g37251(csa_tree_add_190_195_groupi_n_11718 ,csa_tree_add_190_195_groupi_n_11430 ,csa_tree_add_190_195_groupi_n_11559);
  and csa_tree_add_190_195_groupi_g37252(csa_tree_add_190_195_groupi_n_11717 ,csa_tree_add_190_195_groupi_n_11207 ,csa_tree_add_190_195_groupi_n_11567);
  and csa_tree_add_190_195_groupi_g37253(csa_tree_add_190_195_groupi_n_11716 ,csa_tree_add_190_195_groupi_n_11425 ,csa_tree_add_190_195_groupi_n_11565);
  and csa_tree_add_190_195_groupi_g37254(csa_tree_add_190_195_groupi_n_11714 ,csa_tree_add_190_195_groupi_n_11415 ,csa_tree_add_190_195_groupi_n_11546);
  and csa_tree_add_190_195_groupi_g37255(csa_tree_add_190_195_groupi_n_11713 ,csa_tree_add_190_195_groupi_n_11375 ,csa_tree_add_190_195_groupi_n_11569);
  not csa_tree_add_190_195_groupi_g37256(csa_tree_add_190_195_groupi_n_11670 ,csa_tree_add_190_195_groupi_n_11669);
  not csa_tree_add_190_195_groupi_g37257(csa_tree_add_190_195_groupi_n_11667 ,csa_tree_add_190_195_groupi_n_11666);
  not csa_tree_add_190_195_groupi_g37258(csa_tree_add_190_195_groupi_n_11664 ,csa_tree_add_190_195_groupi_n_158);
  not csa_tree_add_190_195_groupi_g37259(csa_tree_add_190_195_groupi_n_11662 ,csa_tree_add_190_195_groupi_n_11661);
  not csa_tree_add_190_195_groupi_g37260(csa_tree_add_190_195_groupi_n_11659 ,csa_tree_add_190_195_groupi_n_11658);
  not csa_tree_add_190_195_groupi_g37261(csa_tree_add_190_195_groupi_n_11657 ,csa_tree_add_190_195_groupi_n_11656);
  not csa_tree_add_190_195_groupi_g37262(csa_tree_add_190_195_groupi_n_11655 ,csa_tree_add_190_195_groupi_n_11654);
  not csa_tree_add_190_195_groupi_g37263(csa_tree_add_190_195_groupi_n_11652 ,csa_tree_add_190_195_groupi_n_11651);
  not csa_tree_add_190_195_groupi_g37264(csa_tree_add_190_195_groupi_n_11650 ,csa_tree_add_190_195_groupi_n_11649);
  not csa_tree_add_190_195_groupi_g37265(csa_tree_add_190_195_groupi_n_11648 ,csa_tree_add_190_195_groupi_n_157);
  not csa_tree_add_190_195_groupi_g37266(csa_tree_add_190_195_groupi_n_11646 ,csa_tree_add_190_195_groupi_n_11645);
  not csa_tree_add_190_195_groupi_g37267(csa_tree_add_190_195_groupi_n_11644 ,csa_tree_add_190_195_groupi_n_11643);
  not csa_tree_add_190_195_groupi_g37268(csa_tree_add_190_195_groupi_n_11642 ,csa_tree_add_190_195_groupi_n_167);
  not csa_tree_add_190_195_groupi_g37269(csa_tree_add_190_195_groupi_n_11640 ,csa_tree_add_190_195_groupi_n_11639);
  not csa_tree_add_190_195_groupi_g37270(csa_tree_add_190_195_groupi_n_11638 ,csa_tree_add_190_195_groupi_n_163);
  not csa_tree_add_190_195_groupi_g37271(csa_tree_add_190_195_groupi_n_11636 ,csa_tree_add_190_195_groupi_n_11635);
  not csa_tree_add_190_195_groupi_g37272(csa_tree_add_190_195_groupi_n_11634 ,csa_tree_add_190_195_groupi_n_11633);
  not csa_tree_add_190_195_groupi_g37273(csa_tree_add_190_195_groupi_n_11631 ,csa_tree_add_190_195_groupi_n_11630);
  xnor csa_tree_add_190_195_groupi_g37274(out1[3] ,csa_tree_add_190_195_groupi_n_10785 ,csa_tree_add_190_195_groupi_n_11359);
  or csa_tree_add_190_195_groupi_g37275(csa_tree_add_190_195_groupi_n_11628 ,csa_tree_add_190_195_groupi_n_11529 ,csa_tree_add_190_195_groupi_n_11379);
  nor csa_tree_add_190_195_groupi_g37276(csa_tree_add_190_195_groupi_n_11627 ,csa_tree_add_190_195_groupi_n_11528 ,csa_tree_add_190_195_groupi_n_11380);
  or csa_tree_add_190_195_groupi_g37277(csa_tree_add_190_195_groupi_n_11626 ,csa_tree_add_190_195_groupi_n_11545 ,csa_tree_add_190_195_groupi_n_11499);
  nor csa_tree_add_190_195_groupi_g37278(csa_tree_add_190_195_groupi_n_11625 ,csa_tree_add_190_195_groupi_n_11239 ,csa_tree_add_190_195_groupi_n_11514);
  or csa_tree_add_190_195_groupi_g37279(csa_tree_add_190_195_groupi_n_11624 ,csa_tree_add_190_195_groupi_n_11263 ,csa_tree_add_190_195_groupi_n_11496);
  or csa_tree_add_190_195_groupi_g37280(csa_tree_add_190_195_groupi_n_11623 ,csa_tree_add_190_195_groupi_n_11368 ,csa_tree_add_190_195_groupi_n_153);
  and csa_tree_add_190_195_groupi_g37281(csa_tree_add_190_195_groupi_n_11622 ,csa_tree_add_190_195_groupi_n_11239 ,csa_tree_add_190_195_groupi_n_11514);
  or csa_tree_add_190_195_groupi_g37282(csa_tree_add_190_195_groupi_n_11621 ,csa_tree_add_190_195_groupi_n_11582 ,csa_tree_add_190_195_groupi_n_11516);
  xnor csa_tree_add_190_195_groupi_g37284(csa_tree_add_190_195_groupi_n_11620 ,csa_tree_add_190_195_groupi_n_11178 ,csa_tree_add_190_195_groupi_n_11456);
  xor csa_tree_add_190_195_groupi_g37285(csa_tree_add_190_195_groupi_n_11619 ,csa_tree_add_190_195_groupi_n_11461 ,csa_tree_add_190_195_groupi_n_11336);
  xnor csa_tree_add_190_195_groupi_g37286(csa_tree_add_190_195_groupi_n_11618 ,csa_tree_add_190_195_groupi_n_11391 ,csa_tree_add_190_195_groupi_n_11055);
  xnor csa_tree_add_190_195_groupi_g37287(csa_tree_add_190_195_groupi_n_11617 ,csa_tree_add_190_195_groupi_n_11048 ,csa_tree_add_190_195_groupi_n_11465);
  xnor csa_tree_add_190_195_groupi_g37288(csa_tree_add_190_195_groupi_n_11616 ,csa_tree_add_190_195_groupi_n_11402 ,csa_tree_add_190_195_groupi_n_11249);
  xnor csa_tree_add_190_195_groupi_g37289(csa_tree_add_190_195_groupi_n_11615 ,csa_tree_add_190_195_groupi_n_11463 ,csa_tree_add_190_195_groupi_n_11467);
  xnor csa_tree_add_190_195_groupi_g37290(csa_tree_add_190_195_groupi_n_11614 ,csa_tree_add_190_195_groupi_n_11410 ,csa_tree_add_190_195_groupi_n_11252);
  xnor csa_tree_add_190_195_groupi_g37291(csa_tree_add_190_195_groupi_n_11613 ,csa_tree_add_190_195_groupi_n_11051 ,csa_tree_add_190_195_groupi_n_11400);
  xnor csa_tree_add_190_195_groupi_g37292(csa_tree_add_190_195_groupi_n_11612 ,csa_tree_add_190_195_groupi_n_9930 ,csa_tree_add_190_195_groupi_n_11475);
  xnor csa_tree_add_190_195_groupi_g37293(csa_tree_add_190_195_groupi_n_11611 ,csa_tree_add_190_195_groupi_n_11022 ,csa_tree_add_190_195_groupi_n_11404);
  xnor csa_tree_add_190_195_groupi_g37294(csa_tree_add_190_195_groupi_n_11610 ,csa_tree_add_190_195_groupi_n_11407 ,csa_tree_add_190_195_groupi_n_11243);
  xnor csa_tree_add_190_195_groupi_g37295(csa_tree_add_190_195_groupi_n_11609 ,csa_tree_add_190_195_groupi_n_11408 ,csa_tree_add_190_195_groupi_n_11381);
  xnor csa_tree_add_190_195_groupi_g37296(csa_tree_add_190_195_groupi_n_11608 ,csa_tree_add_190_195_groupi_n_11050 ,csa_tree_add_190_195_groupi_n_11454);
  xnor csa_tree_add_190_195_groupi_g37297(csa_tree_add_190_195_groupi_n_11607 ,csa_tree_add_190_195_groupi_n_11396 ,csa_tree_add_190_195_groupi_n_11169);
  xnor csa_tree_add_190_195_groupi_g37298(csa_tree_add_190_195_groupi_n_11669 ,csa_tree_add_190_195_groupi_n_10656 ,csa_tree_add_190_195_groupi_n_160);
  xnor csa_tree_add_190_195_groupi_g37299(csa_tree_add_190_195_groupi_n_11668 ,csa_tree_add_190_195_groupi_n_11159 ,csa_tree_add_190_195_groupi_n_11353);
  xnor csa_tree_add_190_195_groupi_g37300(csa_tree_add_190_195_groupi_n_11666 ,csa_tree_add_190_195_groupi_n_10786 ,csa_tree_add_190_195_groupi_n_11352);
  and csa_tree_add_190_195_groupi_g37301(csa_tree_add_190_195_groupi_n_11665 ,csa_tree_add_190_195_groupi_n_11370 ,csa_tree_add_190_195_groupi_n_11495);
  xnor csa_tree_add_190_195_groupi_g37303(csa_tree_add_190_195_groupi_n_11663 ,csa_tree_add_190_195_groupi_n_10795 ,csa_tree_add_190_195_groupi_n_11347);
  xnor csa_tree_add_190_195_groupi_g37304(csa_tree_add_190_195_groupi_n_11661 ,csa_tree_add_190_195_groupi_n_11329 ,csa_tree_add_190_195_groupi_n_11340);
  xnor csa_tree_add_190_195_groupi_g37305(csa_tree_add_190_195_groupi_n_11660 ,csa_tree_add_190_195_groupi_n_10771 ,csa_tree_add_190_195_groupi_n_11361);
  xnor csa_tree_add_190_195_groupi_g37306(csa_tree_add_190_195_groupi_n_11658 ,csa_tree_add_190_195_groupi_n_11183 ,csa_tree_add_190_195_groupi_n_11341);
  xnor csa_tree_add_190_195_groupi_g37307(csa_tree_add_190_195_groupi_n_11656 ,csa_tree_add_190_195_groupi_n_10959 ,csa_tree_add_190_195_groupi_n_11348);
  xnor csa_tree_add_190_195_groupi_g37308(csa_tree_add_190_195_groupi_n_11654 ,csa_tree_add_190_195_groupi_n_10891 ,csa_tree_add_190_195_groupi_n_11349);
  xnor csa_tree_add_190_195_groupi_g37309(csa_tree_add_190_195_groupi_n_11653 ,csa_tree_add_190_195_groupi_n_10886 ,csa_tree_add_190_195_groupi_n_11343);
  xnor csa_tree_add_190_195_groupi_g37310(csa_tree_add_190_195_groupi_n_11651 ,csa_tree_add_190_195_groupi_n_11067 ,csa_tree_add_190_195_groupi_n_11344);
  xnor csa_tree_add_190_195_groupi_g37311(csa_tree_add_190_195_groupi_n_11649 ,csa_tree_add_190_195_groupi_n_11333 ,csa_tree_add_190_195_groupi_n_11350);
  xnor csa_tree_add_190_195_groupi_g37313(csa_tree_add_190_195_groupi_n_11647 ,csa_tree_add_190_195_groupi_n_11265 ,csa_tree_add_190_195_groupi_n_11351);
  xnor csa_tree_add_190_195_groupi_g37314(csa_tree_add_190_195_groupi_n_11645 ,csa_tree_add_190_195_groupi_n_10574 ,csa_tree_add_190_195_groupi_n_11354);
  xnor csa_tree_add_190_195_groupi_g37315(csa_tree_add_190_195_groupi_n_11643 ,csa_tree_add_190_195_groupi_n_10972 ,csa_tree_add_190_195_groupi_n_11345);
  xnor csa_tree_add_190_195_groupi_g37317(csa_tree_add_190_195_groupi_n_11641 ,csa_tree_add_190_195_groupi_n_10666 ,csa_tree_add_190_195_groupi_n_11355);
  xnor csa_tree_add_190_195_groupi_g37318(csa_tree_add_190_195_groupi_n_11639 ,csa_tree_add_190_195_groupi_n_11084 ,csa_tree_add_190_195_groupi_n_11357);
  or csa_tree_add_190_195_groupi_g37320(csa_tree_add_190_195_groupi_n_11637 ,csa_tree_add_190_195_groupi_n_10397 ,csa_tree_add_190_195_groupi_n_11493);
  xnor csa_tree_add_190_195_groupi_g37321(csa_tree_add_190_195_groupi_n_11635 ,csa_tree_add_190_195_groupi_n_10970 ,csa_tree_add_190_195_groupi_n_11362);
  xnor csa_tree_add_190_195_groupi_g37322(csa_tree_add_190_195_groupi_n_11633 ,csa_tree_add_190_195_groupi_n_11078 ,csa_tree_add_190_195_groupi_n_11346);
  and csa_tree_add_190_195_groupi_g37323(csa_tree_add_190_195_groupi_n_11632 ,csa_tree_add_190_195_groupi_n_11365 ,csa_tree_add_190_195_groupi_n_11492);
  xnor csa_tree_add_190_195_groupi_g37324(csa_tree_add_190_195_groupi_n_11630 ,csa_tree_add_190_195_groupi_n_11409 ,csa_tree_add_190_195_groupi_n_10600);
  not csa_tree_add_190_195_groupi_g37325(csa_tree_add_190_195_groupi_n_11598 ,csa_tree_add_190_195_groupi_n_11597);
  not csa_tree_add_190_195_groupi_g37327(csa_tree_add_190_195_groupi_n_11592 ,csa_tree_add_190_195_groupi_n_11591);
  not csa_tree_add_190_195_groupi_g37328(csa_tree_add_190_195_groupi_n_11590 ,csa_tree_add_190_195_groupi_n_11589);
  not csa_tree_add_190_195_groupi_g37329(csa_tree_add_190_195_groupi_n_11588 ,csa_tree_add_190_195_groupi_n_11587);
  not csa_tree_add_190_195_groupi_g37330(csa_tree_add_190_195_groupi_n_11585 ,csa_tree_add_190_195_groupi_n_11586);
  not csa_tree_add_190_195_groupi_g37331(csa_tree_add_190_195_groupi_n_11583 ,csa_tree_add_190_195_groupi_n_11582);
  not csa_tree_add_190_195_groupi_g37332(csa_tree_add_190_195_groupi_n_11581 ,csa_tree_add_190_195_groupi_n_11580);
  not csa_tree_add_190_195_groupi_g37333(csa_tree_add_190_195_groupi_n_11579 ,csa_tree_add_190_195_groupi_n_11578);
  nor csa_tree_add_190_195_groupi_g37334(csa_tree_add_190_195_groupi_n_11577 ,csa_tree_add_190_195_groupi_n_11395 ,csa_tree_add_190_195_groupi_n_11169);
  nor csa_tree_add_190_195_groupi_g37335(csa_tree_add_190_195_groupi_n_11576 ,csa_tree_add_190_195_groupi_n_11252 ,csa_tree_add_190_195_groupi_n_11385);
  or csa_tree_add_190_195_groupi_g37336(csa_tree_add_190_195_groupi_n_11575 ,csa_tree_add_190_195_groupi_n_11473 ,csa_tree_add_190_195_groupi_n_11439);
  or csa_tree_add_190_195_groupi_g37337(csa_tree_add_190_195_groupi_n_11574 ,csa_tree_add_190_195_groupi_n_11466 ,csa_tree_add_190_195_groupi_n_11372);
  and csa_tree_add_190_195_groupi_g37338(csa_tree_add_190_195_groupi_n_11573 ,csa_tree_add_190_195_groupi_n_11252 ,csa_tree_add_190_195_groupi_n_11385);
  nor csa_tree_add_190_195_groupi_g37339(csa_tree_add_190_195_groupi_n_11572 ,csa_tree_add_190_195_groupi_n_11328 ,csa_tree_add_190_195_groupi_n_11381);
  nor csa_tree_add_190_195_groupi_g37340(csa_tree_add_190_195_groupi_n_11571 ,csa_tree_add_190_195_groupi_n_11383 ,csa_tree_add_190_195_groupi_n_11463);
  or csa_tree_add_190_195_groupi_g37341(csa_tree_add_190_195_groupi_n_11570 ,csa_tree_add_190_195_groupi_n_11384 ,csa_tree_add_190_195_groupi_n_11462);
  or csa_tree_add_190_195_groupi_g37342(csa_tree_add_190_195_groupi_n_11569 ,csa_tree_add_190_195_groupi_n_11262 ,csa_tree_add_190_195_groupi_n_11374);
  or csa_tree_add_190_195_groupi_g37343(csa_tree_add_190_195_groupi_n_11568 ,csa_tree_add_190_195_groupi_n_11461 ,csa_tree_add_190_195_groupi_n_11382);
  or csa_tree_add_190_195_groupi_g37344(csa_tree_add_190_195_groupi_n_11567 ,csa_tree_add_190_195_groupi_n_11471 ,csa_tree_add_190_195_groupi_n_11220);
  or csa_tree_add_190_195_groupi_g37345(csa_tree_add_190_195_groupi_n_11566 ,csa_tree_add_190_195_groupi_n_11443 ,csa_tree_add_190_195_groupi_n_11470);
  or csa_tree_add_190_195_groupi_g37346(csa_tree_add_190_195_groupi_n_11565 ,csa_tree_add_190_195_groupi_n_11179 ,csa_tree_add_190_195_groupi_n_11424);
  nor csa_tree_add_190_195_groupi_g37347(csa_tree_add_190_195_groupi_n_11564 ,csa_tree_add_190_195_groupi_n_11231 ,csa_tree_add_190_195_groupi_n_11456);
  or csa_tree_add_190_195_groupi_g37348(csa_tree_add_190_195_groupi_n_11563 ,csa_tree_add_190_195_groupi_n_11238 ,csa_tree_add_190_195_groupi_n_11386);
  or csa_tree_add_190_195_groupi_g37349(csa_tree_add_190_195_groupi_n_11562 ,csa_tree_add_190_195_groupi_n_11232 ,csa_tree_add_190_195_groupi_n_11455);
  or csa_tree_add_190_195_groupi_g37350(csa_tree_add_190_195_groupi_n_11561 ,csa_tree_add_190_195_groupi_n_11050 ,csa_tree_add_190_195_groupi_n_11453);
  nor csa_tree_add_190_195_groupi_g37351(csa_tree_add_190_195_groupi_n_11560 ,csa_tree_add_190_195_groupi_n_11237 ,csa_tree_add_190_195_groupi_n_11387);
  or csa_tree_add_190_195_groupi_g37352(csa_tree_add_190_195_groupi_n_11559 ,csa_tree_add_190_195_groupi_n_11175 ,csa_tree_add_190_195_groupi_n_11432);
  nor csa_tree_add_190_195_groupi_g37353(csa_tree_add_190_195_groupi_n_11558 ,csa_tree_add_190_195_groupi_n_11049 ,csa_tree_add_190_195_groupi_n_11454);
  nor csa_tree_add_190_195_groupi_g37354(csa_tree_add_190_195_groupi_n_11557 ,csa_tree_add_190_195_groupi_n_11407 ,csa_tree_add_190_195_groupi_n_11243);
  and csa_tree_add_190_195_groupi_g37355(csa_tree_add_190_195_groupi_n_11556 ,csa_tree_add_190_195_groupi_n_11461 ,csa_tree_add_190_195_groupi_n_11382);
  or csa_tree_add_190_195_groupi_g37356(csa_tree_add_190_195_groupi_n_11555 ,csa_tree_add_190_195_groupi_n_11396 ,csa_tree_add_190_195_groupi_n_11168);
  and csa_tree_add_190_195_groupi_g37357(csa_tree_add_190_195_groupi_n_11554 ,csa_tree_add_190_195_groupi_n_11328 ,csa_tree_add_190_195_groupi_n_11381);
  and csa_tree_add_190_195_groupi_g37358(csa_tree_add_190_195_groupi_n_11553 ,csa_tree_add_190_195_groupi_n_11407 ,csa_tree_add_190_195_groupi_n_11243);
  and csa_tree_add_190_195_groupi_g37359(csa_tree_add_190_195_groupi_n_11552 ,csa_tree_add_190_195_groupi_n_11051 ,csa_tree_add_190_195_groupi_n_11400);
  nor csa_tree_add_190_195_groupi_g37360(csa_tree_add_190_195_groupi_n_11551 ,csa_tree_add_190_195_groupi_n_11051 ,csa_tree_add_190_195_groupi_n_11400);
  nor csa_tree_add_190_195_groupi_g37361(csa_tree_add_190_195_groupi_n_11550 ,csa_tree_add_190_195_groupi_n_11021 ,csa_tree_add_190_195_groupi_n_11404);
  or csa_tree_add_190_195_groupi_g37362(csa_tree_add_190_195_groupi_n_11549 ,csa_tree_add_190_195_groupi_n_11022 ,csa_tree_add_190_195_groupi_n_11403);
  or csa_tree_add_190_195_groupi_g37363(csa_tree_add_190_195_groupi_n_11548 ,csa_tree_add_190_195_groupi_n_11250 ,csa_tree_add_190_195_groupi_n_11446);
  nor csa_tree_add_190_195_groupi_g37364(csa_tree_add_190_195_groupi_n_11547 ,csa_tree_add_190_195_groupi_n_11251 ,csa_tree_add_190_195_groupi_n_11447);
  or csa_tree_add_190_195_groupi_g37365(csa_tree_add_190_195_groupi_n_11546 ,csa_tree_add_190_195_groupi_n_11476 ,csa_tree_add_190_195_groupi_n_11419);
  or csa_tree_add_190_195_groupi_g37366(csa_tree_add_190_195_groupi_n_11606 ,csa_tree_add_190_195_groupi_n_11285 ,csa_tree_add_190_195_groupi_n_11444);
  and csa_tree_add_190_195_groupi_g37367(csa_tree_add_190_195_groupi_n_11605 ,csa_tree_add_190_195_groupi_n_11279 ,csa_tree_add_190_195_groupi_n_11414);
  and csa_tree_add_190_195_groupi_g37368(csa_tree_add_190_195_groupi_n_11604 ,csa_tree_add_190_195_groupi_n_11431 ,csa_tree_add_190_195_groupi_n_11313);
  and csa_tree_add_190_195_groupi_g37369(csa_tree_add_190_195_groupi_n_11603 ,csa_tree_add_190_195_groupi_n_11284 ,csa_tree_add_190_195_groupi_n_11416);
  and csa_tree_add_190_195_groupi_g37370(csa_tree_add_190_195_groupi_n_11602 ,csa_tree_add_190_195_groupi_n_11289 ,csa_tree_add_190_195_groupi_n_11418);
  and csa_tree_add_190_195_groupi_g37371(csa_tree_add_190_195_groupi_n_11601 ,csa_tree_add_190_195_groupi_n_11293 ,csa_tree_add_190_195_groupi_n_11422);
  and csa_tree_add_190_195_groupi_g37372(csa_tree_add_190_195_groupi_n_11600 ,csa_tree_add_190_195_groupi_n_11423 ,csa_tree_add_190_195_groupi_n_11013);
  and csa_tree_add_190_195_groupi_g37373(csa_tree_add_190_195_groupi_n_11599 ,csa_tree_add_190_195_groupi_n_11300 ,csa_tree_add_190_195_groupi_n_11426);
  or csa_tree_add_190_195_groupi_g37374(csa_tree_add_190_195_groupi_n_11597 ,csa_tree_add_190_195_groupi_n_11363 ,csa_tree_add_190_195_groupi_n_11219);
  and csa_tree_add_190_195_groupi_g37375(csa_tree_add_190_195_groupi_n_11596 ,csa_tree_add_190_195_groupi_n_11303 ,csa_tree_add_190_195_groupi_n_11428);
  or csa_tree_add_190_195_groupi_g37376(csa_tree_add_190_195_groupi_n_11595 ,csa_tree_add_190_195_groupi_n_11210 ,csa_tree_add_190_195_groupi_n_11434);
  and csa_tree_add_190_195_groupi_g37377(csa_tree_add_190_195_groupi_n_11594 ,csa_tree_add_190_195_groupi_n_11438 ,csa_tree_add_190_195_groupi_n_11315);
  and csa_tree_add_190_195_groupi_g37378(csa_tree_add_190_195_groupi_n_11593 ,csa_tree_add_190_195_groupi_n_11317 ,csa_tree_add_190_195_groupi_n_11440);
  or csa_tree_add_190_195_groupi_g37379(csa_tree_add_190_195_groupi_n_11591 ,csa_tree_add_190_195_groupi_n_11266 ,csa_tree_add_190_195_groupi_n_11420);
  and csa_tree_add_190_195_groupi_g37380(csa_tree_add_190_195_groupi_n_11589 ,csa_tree_add_190_195_groupi_n_11282 ,csa_tree_add_190_195_groupi_n_11417);
  or csa_tree_add_190_195_groupi_g37381(csa_tree_add_190_195_groupi_n_11587 ,csa_tree_add_190_195_groupi_n_11270 ,csa_tree_add_190_195_groupi_n_11421);
  and csa_tree_add_190_195_groupi_g37382(csa_tree_add_190_195_groupi_n_11586 ,csa_tree_add_190_195_groupi_n_11322 ,csa_tree_add_190_195_groupi_n_11442);
  and csa_tree_add_190_195_groupi_g37383(csa_tree_add_190_195_groupi_n_11584 ,csa_tree_add_190_195_groupi_n_11286 ,csa_tree_add_190_195_groupi_n_11445);
  and csa_tree_add_190_195_groupi_g37384(csa_tree_add_190_195_groupi_n_11582 ,csa_tree_add_190_195_groupi_n_11429 ,csa_tree_add_190_195_groupi_n_11305);
  and csa_tree_add_190_195_groupi_g37385(csa_tree_add_190_195_groupi_n_11580 ,csa_tree_add_190_195_groupi_n_11319 ,csa_tree_add_190_195_groupi_n_11441);
  and csa_tree_add_190_195_groupi_g37386(csa_tree_add_190_195_groupi_n_11578 ,csa_tree_add_190_195_groupi_n_11274 ,csa_tree_add_190_195_groupi_n_11412);
  not csa_tree_add_190_195_groupi_g37387(csa_tree_add_190_195_groupi_n_11545 ,csa_tree_add_190_195_groupi_n_11544);
  not csa_tree_add_190_195_groupi_g37388(csa_tree_add_190_195_groupi_n_11543 ,csa_tree_add_190_195_groupi_n_11542);
  not csa_tree_add_190_195_groupi_g37389(csa_tree_add_190_195_groupi_n_11539 ,csa_tree_add_190_195_groupi_n_11538);
  not csa_tree_add_190_195_groupi_g37390(csa_tree_add_190_195_groupi_n_11537 ,csa_tree_add_190_195_groupi_n_11536);
  not csa_tree_add_190_195_groupi_g37391(csa_tree_add_190_195_groupi_n_11535 ,csa_tree_add_190_195_groupi_n_11534);
  not csa_tree_add_190_195_groupi_g37392(csa_tree_add_190_195_groupi_n_11533 ,csa_tree_add_190_195_groupi_n_11532);
  not csa_tree_add_190_195_groupi_g37393(csa_tree_add_190_195_groupi_n_11531 ,csa_tree_add_190_195_groupi_n_11530);
  not csa_tree_add_190_195_groupi_g37394(csa_tree_add_190_195_groupi_n_11529 ,csa_tree_add_190_195_groupi_n_11528);
  not csa_tree_add_190_195_groupi_g37395(csa_tree_add_190_195_groupi_n_11527 ,csa_tree_add_190_195_groupi_n_11526);
  not csa_tree_add_190_195_groupi_g37396(csa_tree_add_190_195_groupi_n_11525 ,csa_tree_add_190_195_groupi_n_11524);
  not csa_tree_add_190_195_groupi_g37397(csa_tree_add_190_195_groupi_n_11523 ,csa_tree_add_190_195_groupi_n_11522);
  not csa_tree_add_190_195_groupi_g37398(csa_tree_add_190_195_groupi_n_11519 ,csa_tree_add_190_195_groupi_n_11518);
  not csa_tree_add_190_195_groupi_g37399(csa_tree_add_190_195_groupi_n_11517 ,csa_tree_add_190_195_groupi_n_11516);
  not csa_tree_add_190_195_groupi_g37400(csa_tree_add_190_195_groupi_n_11514 ,csa_tree_add_190_195_groupi_n_11513);
  not csa_tree_add_190_195_groupi_g37401(csa_tree_add_190_195_groupi_n_11512 ,csa_tree_add_190_195_groupi_n_11511);
  not csa_tree_add_190_195_groupi_g37402(csa_tree_add_190_195_groupi_n_11510 ,csa_tree_add_190_195_groupi_n_11509);
  not csa_tree_add_190_195_groupi_g37403(csa_tree_add_190_195_groupi_n_11508 ,csa_tree_add_190_195_groupi_n_11507);
  not csa_tree_add_190_195_groupi_g37404(csa_tree_add_190_195_groupi_n_11506 ,csa_tree_add_190_195_groupi_n_11505);
  nor csa_tree_add_190_195_groupi_g37405(csa_tree_add_190_195_groupi_n_11504 ,csa_tree_add_190_195_groupi_n_11402 ,csa_tree_add_190_195_groupi_n_11249);
  nor csa_tree_add_190_195_groupi_g37406(csa_tree_add_190_195_groupi_n_11503 ,csa_tree_add_190_195_groupi_n_11398 ,csa_tree_add_190_195_groupi_n_11048);
  or csa_tree_add_190_195_groupi_g37407(csa_tree_add_190_195_groupi_n_11502 ,csa_tree_add_190_195_groupi_n_11397 ,csa_tree_add_190_195_groupi_n_11047);
  and csa_tree_add_190_195_groupi_g37408(csa_tree_add_190_195_groupi_n_11501 ,csa_tree_add_190_195_groupi_n_11392 ,csa_tree_add_190_195_groupi_n_11242);
  or csa_tree_add_190_195_groupi_g37409(csa_tree_add_190_195_groupi_n_11500 ,csa_tree_add_190_195_groupi_n_11392 ,csa_tree_add_190_195_groupi_n_11242);
  nor csa_tree_add_190_195_groupi_g37410(csa_tree_add_190_195_groupi_n_11499 ,csa_tree_add_190_195_groupi_n_11390 ,csa_tree_add_190_195_groupi_n_11055);
  or csa_tree_add_190_195_groupi_g37411(csa_tree_add_190_195_groupi_n_11498 ,csa_tree_add_190_195_groupi_n_11391 ,csa_tree_add_190_195_groupi_n_11054);
  or csa_tree_add_190_195_groupi_g37412(csa_tree_add_190_195_groupi_n_11497 ,csa_tree_add_190_195_groupi_n_11401 ,csa_tree_add_190_195_groupi_n_11248);
  nor csa_tree_add_190_195_groupi_g37413(csa_tree_add_190_195_groupi_n_11496 ,csa_tree_add_190_195_groupi_n_10852 ,csa_tree_add_190_195_groupi_n_11389);
  or csa_tree_add_190_195_groupi_g37414(csa_tree_add_190_195_groupi_n_11495 ,csa_tree_add_190_195_groupi_n_11086 ,csa_tree_add_190_195_groupi_n_11366);
  or csa_tree_add_190_195_groupi_g37415(csa_tree_add_190_195_groupi_n_11494 ,csa_tree_add_190_195_groupi_n_139 ,csa_tree_add_190_195_groupi_n_11388);
  and csa_tree_add_190_195_groupi_g37416(csa_tree_add_190_195_groupi_n_11493 ,csa_tree_add_190_195_groupi_n_10415 ,csa_tree_add_190_195_groupi_n_11409);
  or csa_tree_add_190_195_groupi_g37417(csa_tree_add_190_195_groupi_n_11492 ,csa_tree_add_190_195_groupi_n_10697 ,csa_tree_add_190_195_groupi_n_11364);
  xnor csa_tree_add_190_195_groupi_g37419(csa_tree_add_190_195_groupi_n_11491 ,csa_tree_add_190_195_groupi_n_11172 ,csa_tree_add_190_195_groupi_n_11238);
  xnor csa_tree_add_190_195_groupi_g37420(csa_tree_add_190_195_groupi_n_11490 ,csa_tree_add_190_195_groupi_n_11086 ,csa_tree_add_190_195_groupi_n_11326);
  xnor csa_tree_add_190_195_groupi_g37421(csa_tree_add_190_195_groupi_n_11489 ,csa_tree_add_190_195_groupi_n_10880 ,csa_tree_add_190_195_groupi_n_11254);
  xnor csa_tree_add_190_195_groupi_g37422(csa_tree_add_190_195_groupi_n_11488 ,csa_tree_add_190_195_groupi_n_11324 ,csa_tree_add_190_195_groupi_n_11228);
  xnor csa_tree_add_190_195_groupi_g37423(csa_tree_add_190_195_groupi_n_11487 ,csa_tree_add_190_195_groupi_n_11074 ,csa_tree_add_190_195_groupi_n_11334);
  xnor csa_tree_add_190_195_groupi_g37425(csa_tree_add_190_195_groupi_n_11486 ,csa_tree_add_190_195_groupi_n_10852 ,csa_tree_add_190_195_groupi_n_11263);
  xnor csa_tree_add_190_195_groupi_g37426(csa_tree_add_190_195_groupi_n_11485 ,csa_tree_add_190_195_groupi_n_10697 ,csa_tree_add_190_195_groupi_n_11230);
  xnor csa_tree_add_190_195_groupi_g37427(csa_tree_add_190_195_groupi_n_11484 ,csa_tree_add_190_195_groupi_n_11155 ,csa_tree_add_190_195_groupi_n_11236);
  xnor csa_tree_add_190_195_groupi_g37428(csa_tree_add_190_195_groupi_n_11483 ,csa_tree_add_190_195_groupi_n_11161 ,csa_tree_add_190_195_groupi_n_11258);
  xnor csa_tree_add_190_195_groupi_g37429(csa_tree_add_190_195_groupi_n_11482 ,csa_tree_add_190_195_groupi_n_11242 ,csa_tree_add_190_195_groupi_n_11337);
  xnor csa_tree_add_190_195_groupi_g37430(csa_tree_add_190_195_groupi_n_11481 ,csa_tree_add_190_195_groupi_n_11148 ,csa_tree_add_190_195_groupi_n_11227);
  xnor csa_tree_add_190_195_groupi_g37431(csa_tree_add_190_195_groupi_n_11480 ,csa_tree_add_190_195_groupi_n_11234 ,csa_tree_add_190_195_groupi_n_11030);
  xnor csa_tree_add_190_195_groupi_g37432(csa_tree_add_190_195_groupi_n_11479 ,csa_tree_add_190_195_groupi_n_11163 ,csa_tree_add_190_195_groupi_n_11245);
  xnor csa_tree_add_190_195_groupi_g37433(csa_tree_add_190_195_groupi_n_11544 ,csa_tree_add_190_195_groupi_n_11091 ,csa_tree_add_190_195_groupi_n_11186);
  xnor csa_tree_add_190_195_groupi_g37434(csa_tree_add_190_195_groupi_n_11542 ,csa_tree_add_190_195_groupi_n_10842 ,csa_tree_add_190_195_groupi_n_11194);
  and csa_tree_add_190_195_groupi_g37436(csa_tree_add_190_195_groupi_n_11541 ,csa_tree_add_190_195_groupi_n_11435 ,csa_tree_add_190_195_groupi_n_11211);
  xnor csa_tree_add_190_195_groupi_g37437(csa_tree_add_190_195_groupi_n_11540 ,csa_tree_add_190_195_groupi_n_11020 ,csa_tree_add_190_195_groupi_n_11202);
  xnor csa_tree_add_190_195_groupi_g37438(csa_tree_add_190_195_groupi_n_11538 ,csa_tree_add_190_195_groupi_n_11332 ,csa_tree_add_190_195_groupi_n_11192);
  and csa_tree_add_190_195_groupi_g37439(csa_tree_add_190_195_groupi_n_11536 ,csa_tree_add_190_195_groupi_n_11217 ,csa_tree_add_190_195_groupi_n_11371);
  xnor csa_tree_add_190_195_groupi_g37440(csa_tree_add_190_195_groupi_n_11534 ,csa_tree_add_190_195_groupi_n_10165 ,csa_tree_add_190_195_groupi_n_11195);
  xnor csa_tree_add_190_195_groupi_g37441(csa_tree_add_190_195_groupi_n_11532 ,csa_tree_add_190_195_groupi_n_10653 ,csa_tree_add_190_195_groupi_n_11203);
  and csa_tree_add_190_195_groupi_g37442(csa_tree_add_190_195_groupi_n_11530 ,csa_tree_add_190_195_groupi_n_11225 ,csa_tree_add_190_195_groupi_n_11369);
  xnor csa_tree_add_190_195_groupi_g37443(csa_tree_add_190_195_groupi_n_11528 ,csa_tree_add_190_195_groupi_n_11044 ,csa_tree_add_190_195_groupi_n_11187);
  xnor csa_tree_add_190_195_groupi_g37444(csa_tree_add_190_195_groupi_n_11526 ,csa_tree_add_190_195_groupi_n_10875 ,csa_tree_add_190_195_groupi_n_11193);
  xnor csa_tree_add_190_195_groupi_g37445(csa_tree_add_190_195_groupi_n_11524 ,csa_tree_add_190_195_groupi_n_10703 ,csa_tree_add_190_195_groupi_n_11191);
  xnor csa_tree_add_190_195_groupi_g37446(csa_tree_add_190_195_groupi_n_11522 ,csa_tree_add_190_195_groupi_n_11090 ,csa_tree_add_190_195_groupi_n_11190);
  xnor csa_tree_add_190_195_groupi_g37447(csa_tree_add_190_195_groupi_n_11521 ,csa_tree_add_190_195_groupi_n_10677 ,csa_tree_add_190_195_groupi_n_11204);
  xnor csa_tree_add_190_195_groupi_g37448(csa_tree_add_190_195_groupi_n_11520 ,csa_tree_add_190_195_groupi_n_10794 ,csa_tree_add_190_195_groupi_n_11200);
  xnor csa_tree_add_190_195_groupi_g37450(csa_tree_add_190_195_groupi_n_11518 ,csa_tree_add_190_195_groupi_n_11061 ,csa_tree_add_190_195_groupi_n_11199);
  xnor csa_tree_add_190_195_groupi_g37451(csa_tree_add_190_195_groupi_n_11516 ,csa_tree_add_190_195_groupi_n_10980 ,csa_tree_add_190_195_groupi_n_11188);
  xnor csa_tree_add_190_195_groupi_g37453(csa_tree_add_190_195_groupi_n_11515 ,csa_tree_add_190_195_groupi_n_10670 ,csa_tree_add_190_195_groupi_n_156);
  xnor csa_tree_add_190_195_groupi_g37454(csa_tree_add_190_195_groupi_n_11513 ,csa_tree_add_190_195_groupi_n_10977 ,csa_tree_add_190_195_groupi_n_11185);
  xnor csa_tree_add_190_195_groupi_g37455(csa_tree_add_190_195_groupi_n_11511 ,csa_tree_add_190_195_groupi_n_10693 ,csa_tree_add_190_195_groupi_n_11197);
  xnor csa_tree_add_190_195_groupi_g37456(csa_tree_add_190_195_groupi_n_11509 ,csa_tree_add_190_195_groupi_n_11089 ,csa_tree_add_190_195_groupi_n_11196);
  xnor csa_tree_add_190_195_groupi_g37457(csa_tree_add_190_195_groupi_n_11507 ,csa_tree_add_190_195_groupi_n_10691 ,csa_tree_add_190_195_groupi_n_11205);
  xnor csa_tree_add_190_195_groupi_g37458(csa_tree_add_190_195_groupi_n_11505 ,csa_tree_add_190_195_groupi_n_10153 ,csa_tree_add_190_195_groupi_n_11206);
  not csa_tree_add_190_195_groupi_g37460(csa_tree_add_190_195_groupi_n_11476 ,csa_tree_add_190_195_groupi_n_11475);
  not csa_tree_add_190_195_groupi_g37463(csa_tree_add_190_195_groupi_n_11470 ,csa_tree_add_190_195_groupi_n_11469);
  not csa_tree_add_190_195_groupi_g37465(csa_tree_add_190_195_groupi_n_11462 ,csa_tree_add_190_195_groupi_n_11463);
  not csa_tree_add_190_195_groupi_g37466(csa_tree_add_190_195_groupi_n_11458 ,csa_tree_add_190_195_groupi_n_11457);
  not csa_tree_add_190_195_groupi_g37467(csa_tree_add_190_195_groupi_n_11456 ,csa_tree_add_190_195_groupi_n_11455);
  not csa_tree_add_190_195_groupi_g37468(csa_tree_add_190_195_groupi_n_11454 ,csa_tree_add_190_195_groupi_n_11453);
  not csa_tree_add_190_195_groupi_g37469(csa_tree_add_190_195_groupi_n_11452 ,csa_tree_add_190_195_groupi_n_11451);
  not csa_tree_add_190_195_groupi_g37470(csa_tree_add_190_195_groupi_n_11449 ,csa_tree_add_190_195_groupi_n_11448);
  not csa_tree_add_190_195_groupi_g37471(csa_tree_add_190_195_groupi_n_11447 ,csa_tree_add_190_195_groupi_n_11446);
  or csa_tree_add_190_195_groupi_g37472(csa_tree_add_190_195_groupi_n_11445 ,csa_tree_add_190_195_groupi_n_11174 ,csa_tree_add_190_195_groupi_n_11283);
  and csa_tree_add_190_195_groupi_g37473(csa_tree_add_190_195_groupi_n_11444 ,csa_tree_add_190_195_groupi_n_10795 ,csa_tree_add_190_195_groupi_n_11281);
  nor csa_tree_add_190_195_groupi_g37474(csa_tree_add_190_195_groupi_n_11443 ,csa_tree_add_190_195_groupi_n_11161 ,csa_tree_add_190_195_groupi_n_11258);
  or csa_tree_add_190_195_groupi_g37475(csa_tree_add_190_195_groupi_n_11442 ,csa_tree_add_190_195_groupi_n_10771 ,csa_tree_add_190_195_groupi_n_11320);
  or csa_tree_add_190_195_groupi_g37476(csa_tree_add_190_195_groupi_n_11441 ,csa_tree_add_190_195_groupi_n_11264 ,csa_tree_add_190_195_groupi_n_11318);
  or csa_tree_add_190_195_groupi_g37477(csa_tree_add_190_195_groupi_n_11440 ,csa_tree_add_190_195_groupi_n_11182 ,csa_tree_add_190_195_groupi_n_11316);
  nor csa_tree_add_190_195_groupi_g37478(csa_tree_add_190_195_groupi_n_11439 ,csa_tree_add_190_195_groupi_n_11162 ,csa_tree_add_190_195_groupi_n_11245);
  or csa_tree_add_190_195_groupi_g37479(csa_tree_add_190_195_groupi_n_11438 ,csa_tree_add_190_195_groupi_n_11333 ,csa_tree_add_190_195_groupi_n_11314);
  nor csa_tree_add_190_195_groupi_g37480(csa_tree_add_190_195_groupi_n_11437 ,csa_tree_add_190_195_groupi_n_11147 ,csa_tree_add_190_195_groupi_n_11227);
  or csa_tree_add_190_195_groupi_g37481(csa_tree_add_190_195_groupi_n_11436 ,csa_tree_add_190_195_groupi_n_11160 ,csa_tree_add_190_195_groupi_n_11257);
  or csa_tree_add_190_195_groupi_g37482(csa_tree_add_190_195_groupi_n_11435 ,csa_tree_add_190_195_groupi_n_10785 ,csa_tree_add_190_195_groupi_n_11212);
  and csa_tree_add_190_195_groupi_g37483(csa_tree_add_190_195_groupi_n_11434 ,csa_tree_add_190_195_groupi_n_10786 ,csa_tree_add_190_195_groupi_n_11209);
  or csa_tree_add_190_195_groupi_g37484(csa_tree_add_190_195_groupi_n_11433 ,csa_tree_add_190_195_groupi_n_11163 ,csa_tree_add_190_195_groupi_n_11244);
  nor csa_tree_add_190_195_groupi_g37485(csa_tree_add_190_195_groupi_n_11432 ,csa_tree_add_190_195_groupi_n_11154 ,csa_tree_add_190_195_groupi_n_11236);
  or csa_tree_add_190_195_groupi_g37486(csa_tree_add_190_195_groupi_n_11431 ,csa_tree_add_190_195_groupi_n_11338 ,csa_tree_add_190_195_groupi_n_11308);
  or csa_tree_add_190_195_groupi_g37487(csa_tree_add_190_195_groupi_n_11430 ,csa_tree_add_190_195_groupi_n_11155 ,csa_tree_add_190_195_groupi_n_11235);
  or csa_tree_add_190_195_groupi_g37488(csa_tree_add_190_195_groupi_n_11429 ,csa_tree_add_190_195_groupi_n_10986 ,csa_tree_add_190_195_groupi_n_11304);
  or csa_tree_add_190_195_groupi_g37489(csa_tree_add_190_195_groupi_n_11428 ,csa_tree_add_190_195_groupi_n_11184 ,csa_tree_add_190_195_groupi_n_11302);
  or csa_tree_add_190_195_groupi_g37490(csa_tree_add_190_195_groupi_n_11427 ,csa_tree_add_190_195_groupi_n_11148 ,csa_tree_add_190_195_groupi_n_11226);
  or csa_tree_add_190_195_groupi_g37491(csa_tree_add_190_195_groupi_n_11426 ,csa_tree_add_190_195_groupi_n_11087 ,csa_tree_add_190_195_groupi_n_11299);
  or csa_tree_add_190_195_groupi_g37492(csa_tree_add_190_195_groupi_n_11425 ,csa_tree_add_190_195_groupi_n_11027 ,csa_tree_add_190_195_groupi_n_11329);
  and csa_tree_add_190_195_groupi_g37493(csa_tree_add_190_195_groupi_n_11424 ,csa_tree_add_190_195_groupi_n_11027 ,csa_tree_add_190_195_groupi_n_11329);
  or csa_tree_add_190_195_groupi_g37494(csa_tree_add_190_195_groupi_n_11423 ,csa_tree_add_190_195_groupi_n_11332 ,csa_tree_add_190_195_groupi_n_11014);
  or csa_tree_add_190_195_groupi_g37495(csa_tree_add_190_195_groupi_n_11422 ,csa_tree_add_190_195_groupi_n_11335 ,csa_tree_add_190_195_groupi_n_11292);
  nor csa_tree_add_190_195_groupi_g37496(csa_tree_add_190_195_groupi_n_11421 ,csa_tree_add_190_195_groupi_n_10903 ,csa_tree_add_190_195_groupi_n_11275);
  and csa_tree_add_190_195_groupi_g37497(csa_tree_add_190_195_groupi_n_11420 ,csa_tree_add_190_195_groupi_n_11183 ,csa_tree_add_190_195_groupi_n_11294);
  nor csa_tree_add_190_195_groupi_g37498(csa_tree_add_190_195_groupi_n_11419 ,csa_tree_add_190_195_groupi_n_9929 ,csa_tree_add_190_195_groupi_n_11260);
  or csa_tree_add_190_195_groupi_g37499(csa_tree_add_190_195_groupi_n_11418 ,csa_tree_add_190_195_groupi_n_10984 ,csa_tree_add_190_195_groupi_n_11287);
  or csa_tree_add_190_195_groupi_g37500(csa_tree_add_190_195_groupi_n_11417 ,csa_tree_add_190_195_groupi_n_10979 ,csa_tree_add_190_195_groupi_n_11280);
  or csa_tree_add_190_195_groupi_g37501(csa_tree_add_190_195_groupi_n_11416 ,csa_tree_add_190_195_groupi_n_10978 ,csa_tree_add_190_195_groupi_n_11277);
  or csa_tree_add_190_195_groupi_g37502(csa_tree_add_190_195_groupi_n_11415 ,csa_tree_add_190_195_groupi_n_9930 ,csa_tree_add_190_195_groupi_n_11259);
  or csa_tree_add_190_195_groupi_g37503(csa_tree_add_190_195_groupi_n_11414 ,csa_tree_add_190_195_groupi_n_10975 ,csa_tree_add_190_195_groupi_n_11276);
  nor csa_tree_add_190_195_groupi_g37504(csa_tree_add_190_195_groupi_n_11413 ,csa_tree_add_190_195_groupi_n_11323 ,csa_tree_add_190_195_groupi_n_11228);
  or csa_tree_add_190_195_groupi_g37505(csa_tree_add_190_195_groupi_n_11412 ,csa_tree_add_190_195_groupi_n_10972 ,csa_tree_add_190_195_groupi_n_11272);
  or csa_tree_add_190_195_groupi_g37506(csa_tree_add_190_195_groupi_n_11411 ,csa_tree_add_190_195_groupi_n_11324 ,csa_tree_add_190_195_groupi_n_150);
  and csa_tree_add_190_195_groupi_g37507(csa_tree_add_190_195_groupi_n_11478 ,csa_tree_add_190_195_groupi_n_11105 ,csa_tree_add_190_195_groupi_n_11273);
  and csa_tree_add_190_195_groupi_g37508(csa_tree_add_190_195_groupi_n_11477 ,csa_tree_add_190_195_groupi_n_11100 ,csa_tree_add_190_195_groupi_n_11269);
  or csa_tree_add_190_195_groupi_g37509(csa_tree_add_190_195_groupi_n_11475 ,csa_tree_add_190_195_groupi_n_11144 ,csa_tree_add_190_195_groupi_n_11321);
  and csa_tree_add_190_195_groupi_g37510(csa_tree_add_190_195_groupi_n_11474 ,csa_tree_add_190_195_groupi_n_10717 ,csa_tree_add_190_195_groupi_n_11271);
  and csa_tree_add_190_195_groupi_g37511(csa_tree_add_190_195_groupi_n_11473 ,csa_tree_add_190_195_groupi_n_11146 ,csa_tree_add_190_195_groupi_n_11278);
  and csa_tree_add_190_195_groupi_g37512(csa_tree_add_190_195_groupi_n_11472 ,csa_tree_add_190_195_groupi_n_11112 ,csa_tree_add_190_195_groupi_n_11288);
  and csa_tree_add_190_195_groupi_g37513(csa_tree_add_190_195_groupi_n_11471 ,csa_tree_add_190_195_groupi_n_11138 ,csa_tree_add_190_195_groupi_n_11222);
  or csa_tree_add_190_195_groupi_g37514(csa_tree_add_190_195_groupi_n_11469 ,csa_tree_add_190_195_groupi_n_11126 ,csa_tree_add_190_195_groupi_n_11216);
  and csa_tree_add_190_195_groupi_g37515(csa_tree_add_190_195_groupi_n_11468 ,csa_tree_add_190_195_groupi_n_11097 ,csa_tree_add_190_195_groupi_n_11295);
  and csa_tree_add_190_195_groupi_g37516(csa_tree_add_190_195_groupi_n_11467 ,csa_tree_add_190_195_groupi_n_11125 ,csa_tree_add_190_195_groupi_n_11223);
  and csa_tree_add_190_195_groupi_g37517(csa_tree_add_190_195_groupi_n_11466 ,csa_tree_add_190_195_groupi_n_11135 ,csa_tree_add_190_195_groupi_n_11311);
  and csa_tree_add_190_195_groupi_g37518(csa_tree_add_190_195_groupi_n_11465 ,csa_tree_add_190_195_groupi_n_11012 ,csa_tree_add_190_195_groupi_n_11301);
  and csa_tree_add_190_195_groupi_g37519(csa_tree_add_190_195_groupi_n_11464 ,csa_tree_add_190_195_groupi_n_11128 ,csa_tree_add_190_195_groupi_n_11306);
  or csa_tree_add_190_195_groupi_g37520(csa_tree_add_190_195_groupi_n_11463 ,csa_tree_add_190_195_groupi_n_11145 ,csa_tree_add_190_195_groupi_n_11312);
  and csa_tree_add_190_195_groupi_g37521(csa_tree_add_190_195_groupi_n_11461 ,csa_tree_add_190_195_groupi_n_11130 ,csa_tree_add_190_195_groupi_n_11309);
  and csa_tree_add_190_195_groupi_g37522(csa_tree_add_190_195_groupi_n_11460 ,csa_tree_add_190_195_groupi_n_11007 ,csa_tree_add_190_195_groupi_n_11310);
  and csa_tree_add_190_195_groupi_g37523(csa_tree_add_190_195_groupi_n_11459 ,csa_tree_add_190_195_groupi_n_11004 ,csa_tree_add_190_195_groupi_n_11307);
  and csa_tree_add_190_195_groupi_g37524(csa_tree_add_190_195_groupi_n_11457 ,csa_tree_add_190_195_groupi_n_11103 ,csa_tree_add_190_195_groupi_n_11296);
  and csa_tree_add_190_195_groupi_g37525(csa_tree_add_190_195_groupi_n_11455 ,csa_tree_add_190_195_groupi_n_11117 ,csa_tree_add_190_195_groupi_n_11298);
  and csa_tree_add_190_195_groupi_g37526(csa_tree_add_190_195_groupi_n_11453 ,csa_tree_add_190_195_groupi_n_11115 ,csa_tree_add_190_195_groupi_n_11291);
  and csa_tree_add_190_195_groupi_g37527(csa_tree_add_190_195_groupi_n_11451 ,csa_tree_add_190_195_groupi_n_11134 ,csa_tree_add_190_195_groupi_n_11224);
  and csa_tree_add_190_195_groupi_g37528(csa_tree_add_190_195_groupi_n_11450 ,csa_tree_add_190_195_groupi_n_11094 ,csa_tree_add_190_195_groupi_n_11297);
  or csa_tree_add_190_195_groupi_g37529(csa_tree_add_190_195_groupi_n_11448 ,csa_tree_add_190_195_groupi_n_11114 ,csa_tree_add_190_195_groupi_n_11290);
  and csa_tree_add_190_195_groupi_g37530(csa_tree_add_190_195_groupi_n_11446 ,csa_tree_add_190_195_groupi_n_11098 ,csa_tree_add_190_195_groupi_n_11267);
  not csa_tree_add_190_195_groupi_g37531(csa_tree_add_190_195_groupi_n_11406 ,csa_tree_add_190_195_groupi_n_11405);
  not csa_tree_add_190_195_groupi_g37532(csa_tree_add_190_195_groupi_n_11404 ,csa_tree_add_190_195_groupi_n_11403);
  not csa_tree_add_190_195_groupi_g37533(csa_tree_add_190_195_groupi_n_11402 ,csa_tree_add_190_195_groupi_n_11401);
  not csa_tree_add_190_195_groupi_g37534(csa_tree_add_190_195_groupi_n_11398 ,csa_tree_add_190_195_groupi_n_11397);
  not csa_tree_add_190_195_groupi_g37535(csa_tree_add_190_195_groupi_n_11396 ,csa_tree_add_190_195_groupi_n_11395);
  not csa_tree_add_190_195_groupi_g37536(csa_tree_add_190_195_groupi_n_11394 ,csa_tree_add_190_195_groupi_n_11393);
  not csa_tree_add_190_195_groupi_g37537(csa_tree_add_190_195_groupi_n_11391 ,csa_tree_add_190_195_groupi_n_11390);
  not csa_tree_add_190_195_groupi_g37538(csa_tree_add_190_195_groupi_n_11389 ,csa_tree_add_190_195_groupi_n_11388);
  not csa_tree_add_190_195_groupi_g37539(csa_tree_add_190_195_groupi_n_11387 ,csa_tree_add_190_195_groupi_n_11386);
  not csa_tree_add_190_195_groupi_g37540(csa_tree_add_190_195_groupi_n_11384 ,csa_tree_add_190_195_groupi_n_11383);
  not csa_tree_add_190_195_groupi_g37541(csa_tree_add_190_195_groupi_n_11380 ,csa_tree_add_190_195_groupi_n_11379);
  not csa_tree_add_190_195_groupi_g37542(csa_tree_add_190_195_groupi_n_11377 ,csa_tree_add_190_195_groupi_n_11376);
  or csa_tree_add_190_195_groupi_g37543(csa_tree_add_190_195_groupi_n_11375 ,csa_tree_add_190_195_groupi_n_10880 ,csa_tree_add_190_195_groupi_n_11253);
  nor csa_tree_add_190_195_groupi_g37544(csa_tree_add_190_195_groupi_n_11374 ,csa_tree_add_190_195_groupi_n_10879 ,csa_tree_add_190_195_groupi_n_11254);
  or csa_tree_add_190_195_groupi_g37545(csa_tree_add_190_195_groupi_n_11373 ,csa_tree_add_190_195_groupi_n_11035 ,csa_tree_add_190_195_groupi_n_11246);
  nor csa_tree_add_190_195_groupi_g37546(csa_tree_add_190_195_groupi_n_11372 ,csa_tree_add_190_195_groupi_n_11036 ,csa_tree_add_190_195_groupi_n_11247);
  or csa_tree_add_190_195_groupi_g37547(csa_tree_add_190_195_groupi_n_11371 ,csa_tree_add_190_195_groupi_n_11093 ,csa_tree_add_190_195_groupi_n_11215);
  or csa_tree_add_190_195_groupi_g37548(csa_tree_add_190_195_groupi_n_11370 ,csa_tree_add_190_195_groupi_n_11038 ,csa_tree_add_190_195_groupi_n_11325);
  or csa_tree_add_190_195_groupi_g37549(csa_tree_add_190_195_groupi_n_11369 ,csa_tree_add_190_195_groupi_n_11085 ,csa_tree_add_190_195_groupi_n_11213);
  nor csa_tree_add_190_195_groupi_g37550(csa_tree_add_190_195_groupi_n_11368 ,csa_tree_add_190_195_groupi_n_11233 ,csa_tree_add_190_195_groupi_n_11030);
  or csa_tree_add_190_195_groupi_g37551(csa_tree_add_190_195_groupi_n_11367 ,csa_tree_add_190_195_groupi_n_11234 ,csa_tree_add_190_195_groupi_n_11029);
  nor csa_tree_add_190_195_groupi_g37552(csa_tree_add_190_195_groupi_n_11366 ,csa_tree_add_190_195_groupi_n_11037 ,csa_tree_add_190_195_groupi_n_11326);
  or csa_tree_add_190_195_groupi_g37553(csa_tree_add_190_195_groupi_n_11365 ,csa_tree_add_190_195_groupi_n_140 ,csa_tree_add_190_195_groupi_n_11229);
  nor csa_tree_add_190_195_groupi_g37554(csa_tree_add_190_195_groupi_n_11364 ,csa_tree_add_190_195_groupi_n_10845 ,csa_tree_add_190_195_groupi_n_11230);
  and csa_tree_add_190_195_groupi_g37555(csa_tree_add_190_195_groupi_n_11363 ,csa_tree_add_190_195_groupi_n_11221 ,csa_tree_add_190_195_groupi_n_11265);
  xnor csa_tree_add_190_195_groupi_g37556(csa_tree_add_190_195_groupi_n_11362 ,csa_tree_add_190_195_groupi_n_11023 ,csa_tree_add_190_195_groupi_n_10903);
  xnor csa_tree_add_190_195_groupi_g37557(csa_tree_add_190_195_groupi_n_11361 ,csa_tree_add_190_195_groupi_n_10841 ,csa_tree_add_190_195_groupi_n_11149);
  xnor csa_tree_add_190_195_groupi_g37558(csa_tree_add_190_195_groupi_n_11360 ,csa_tree_add_190_195_groupi_n_10669 ,csa_tree_add_190_195_groupi_n_11053);
  xnor csa_tree_add_190_195_groupi_g37559(csa_tree_add_190_195_groupi_n_11359 ,csa_tree_add_190_195_groupi_n_10675 ,csa_tree_add_190_195_groupi_n_11032);
  xnor csa_tree_add_190_195_groupi_g37560(csa_tree_add_190_195_groupi_n_11358 ,csa_tree_add_190_195_groupi_n_11153 ,csa_tree_add_190_195_groupi_n_10893);
  xnor csa_tree_add_190_195_groupi_g37561(csa_tree_add_190_195_groupi_n_11357 ,csa_tree_add_190_195_groupi_n_11057 ,csa_tree_add_190_195_groupi_n_11034);
  xnor csa_tree_add_190_195_groupi_g37562(csa_tree_add_190_195_groupi_n_11356 ,csa_tree_add_190_195_groupi_n_11167 ,csa_tree_add_190_195_groupi_n_11059);
  xnor csa_tree_add_190_195_groupi_g37563(csa_tree_add_190_195_groupi_n_11355 ,csa_tree_add_190_195_groupi_n_10866 ,csa_tree_add_190_195_groupi_n_11173);
  xnor csa_tree_add_190_195_groupi_g37564(csa_tree_add_190_195_groupi_n_11354 ,csa_tree_add_190_195_groupi_n_10572 ,csa_tree_add_190_195_groupi_n_11180);
  xnor csa_tree_add_190_195_groupi_g37565(csa_tree_add_190_195_groupi_n_11353 ,csa_tree_add_190_195_groupi_n_11087 ,csa_tree_add_190_195_groupi_n_10840);
  xnor csa_tree_add_190_195_groupi_g37566(csa_tree_add_190_195_groupi_n_11352 ,csa_tree_add_190_195_groupi_n_10847 ,csa_tree_add_190_195_groupi_n_11028);
  xnor csa_tree_add_190_195_groupi_g37567(csa_tree_add_190_195_groupi_n_11351 ,csa_tree_add_190_195_groupi_n_11157 ,csa_tree_add_190_195_groupi_n_10877);
  xnor csa_tree_add_190_195_groupi_g37568(csa_tree_add_190_195_groupi_n_11350 ,csa_tree_add_190_195_groupi_n_11065 ,csa_tree_add_190_195_groupi_n_11063);
  xnor csa_tree_add_190_195_groupi_g37569(csa_tree_add_190_195_groupi_n_11349 ,csa_tree_add_190_195_groupi_n_11093 ,csa_tree_add_190_195_groupi_n_11046);
  xnor csa_tree_add_190_195_groupi_g37570(csa_tree_add_190_195_groupi_n_11348 ,csa_tree_add_190_195_groupi_n_10849 ,csa_tree_add_190_195_groupi_n_11088);
  xnor csa_tree_add_190_195_groupi_g37571(csa_tree_add_190_195_groupi_n_11347 ,csa_tree_add_190_195_groupi_n_10869 ,csa_tree_add_190_195_groupi_n_11076);
  xnor csa_tree_add_190_195_groupi_g37572(csa_tree_add_190_195_groupi_n_11346 ,csa_tree_add_190_195_groupi_n_10770 ,csa_tree_add_190_195_groupi_n_11174);
  xnor csa_tree_add_190_195_groupi_g37574(csa_tree_add_190_195_groupi_n_11345 ,csa_tree_add_190_195_groupi_n_11040 ,csa_tree_add_190_195_groupi_n_11082);
  xnor csa_tree_add_190_195_groupi_g37575(csa_tree_add_190_195_groupi_n_11344 ,csa_tree_add_190_195_groupi_n_11165 ,csa_tree_add_190_195_groupi_n_11184);
  xnor csa_tree_add_190_195_groupi_g37576(csa_tree_add_190_195_groupi_n_11343 ,csa_tree_add_190_195_groupi_n_10889 ,csa_tree_add_190_195_groupi_n_11176);
  xnor csa_tree_add_190_195_groupi_g37577(csa_tree_add_190_195_groupi_n_11342 ,csa_tree_add_190_195_groupi_n_11069 ,csa_tree_add_190_195_groupi_n_10961);
  xnor csa_tree_add_190_195_groupi_g37578(csa_tree_add_190_195_groupi_n_11341 ,csa_tree_add_190_195_groupi_n_10968 ,csa_tree_add_190_195_groupi_n_11080);
  xnor csa_tree_add_190_195_groupi_g37579(csa_tree_add_190_195_groupi_n_11340 ,csa_tree_add_190_195_groupi_n_11027 ,csa_tree_add_190_195_groupi_n_11179);
  and csa_tree_add_190_195_groupi_g37580(csa_tree_add_190_195_groupi_n_11410 ,csa_tree_add_190_195_groupi_n_11011 ,csa_tree_add_190_195_groupi_n_11218);
  or csa_tree_add_190_195_groupi_g37581(csa_tree_add_190_195_groupi_n_11409 ,csa_tree_add_190_195_groupi_n_10408 ,csa_tree_add_190_195_groupi_n_11268);
  and csa_tree_add_190_195_groupi_g37582(csa_tree_add_190_195_groupi_n_11408 ,csa_tree_add_190_195_groupi_n_11005 ,csa_tree_add_190_195_groupi_n_11208);
  xnor csa_tree_add_190_195_groupi_g37583(csa_tree_add_190_195_groupi_n_11407 ,csa_tree_add_190_195_groupi_n_10462 ,csa_tree_add_190_195_groupi_n_10993);
  xnor csa_tree_add_190_195_groupi_g37584(csa_tree_add_190_195_groupi_n_11405 ,csa_tree_add_190_195_groupi_n_11170 ,csa_tree_add_190_195_groupi_n_10620);
  xnor csa_tree_add_190_195_groupi_g37585(csa_tree_add_190_195_groupi_n_11403 ,csa_tree_add_190_195_groupi_n_10328 ,csa_tree_add_190_195_groupi_n_155);
  xnor csa_tree_add_190_195_groupi_g37586(csa_tree_add_190_195_groupi_n_11401 ,csa_tree_add_190_195_groupi_n_10433 ,csa_tree_add_190_195_groupi_n_10989);
  xnor csa_tree_add_190_195_groupi_g37587(csa_tree_add_190_195_groupi_n_11400 ,csa_tree_add_190_195_groupi_n_10844 ,csa_tree_add_190_195_groupi_n_10996);
  xnor csa_tree_add_190_195_groupi_g37588(csa_tree_add_190_195_groupi_n_11399 ,csa_tree_add_190_195_groupi_n_10873 ,csa_tree_add_190_195_groupi_n_10992);
  xnor csa_tree_add_190_195_groupi_g37589(csa_tree_add_190_195_groupi_n_11397 ,csa_tree_add_190_195_groupi_n_10686 ,csa_tree_add_190_195_groupi_n_154);
  xnor csa_tree_add_190_195_groupi_g37590(csa_tree_add_190_195_groupi_n_11395 ,csa_tree_add_190_195_groupi_n_9860 ,csa_tree_add_190_195_groupi_n_152);
  xnor csa_tree_add_190_195_groupi_g37591(csa_tree_add_190_195_groupi_n_11393 ,csa_tree_add_190_195_groupi_n_10789 ,csa_tree_add_190_195_groupi_n_10998);
  xnor csa_tree_add_190_195_groupi_g37592(csa_tree_add_190_195_groupi_n_11392 ,csa_tree_add_190_195_groupi_n_10860 ,csa_tree_add_190_195_groupi_n_10994);
  xnor csa_tree_add_190_195_groupi_g37593(csa_tree_add_190_195_groupi_n_11390 ,csa_tree_add_190_195_groupi_n_10586 ,csa_tree_add_190_195_groupi_n_10999);
  xnor csa_tree_add_190_195_groupi_g37594(csa_tree_add_190_195_groupi_n_11388 ,csa_tree_add_190_195_groupi_n_9768 ,csa_tree_add_190_195_groupi_n_10997);
  xnor csa_tree_add_190_195_groupi_g37595(csa_tree_add_190_195_groupi_n_11386 ,csa_tree_add_190_195_groupi_n_10435 ,csa_tree_add_190_195_groupi_n_11000);
  xnor csa_tree_add_190_195_groupi_g37596(csa_tree_add_190_195_groupi_n_11385 ,csa_tree_add_190_195_groupi_n_10775 ,csa_tree_add_190_195_groupi_n_10987);
  xnor csa_tree_add_190_195_groupi_g37597(csa_tree_add_190_195_groupi_n_11383 ,csa_tree_add_190_195_groupi_n_10681 ,csa_tree_add_190_195_groupi_n_10988);
  xnor csa_tree_add_190_195_groupi_g37598(csa_tree_add_190_195_groupi_n_11382 ,csa_tree_add_190_195_groupi_n_10157 ,csa_tree_add_190_195_groupi_n_10995);
  xnor csa_tree_add_190_195_groupi_g37599(csa_tree_add_190_195_groupi_n_11381 ,csa_tree_add_190_195_groupi_n_10346 ,csa_tree_add_190_195_groupi_n_11001);
  and csa_tree_add_190_195_groupi_g37600(csa_tree_add_190_195_groupi_n_11379 ,csa_tree_add_190_195_groupi_n_11214 ,csa_tree_add_190_195_groupi_n_11008);
  xnor csa_tree_add_190_195_groupi_g37601(csa_tree_add_190_195_groupi_n_11378 ,csa_tree_add_190_195_groupi_n_10662 ,csa_tree_add_190_195_groupi_n_10990);
  xnor csa_tree_add_190_195_groupi_g37602(csa_tree_add_190_195_groupi_n_11376 ,csa_tree_add_190_195_groupi_n_10964 ,csa_tree_add_190_195_groupi_n_10991);
  not csa_tree_add_190_195_groupi_g37604(csa_tree_add_190_195_groupi_n_11335 ,csa_tree_add_190_195_groupi_n_11334);
  not csa_tree_add_190_195_groupi_g37605(csa_tree_add_190_195_groupi_n_11330 ,csa_tree_add_190_195_groupi_n_11331);
  not csa_tree_add_190_195_groupi_g37606(csa_tree_add_190_195_groupi_n_11328 ,csa_tree_add_190_195_groupi_n_11327);
  not csa_tree_add_190_195_groupi_g37607(csa_tree_add_190_195_groupi_n_11326 ,csa_tree_add_190_195_groupi_n_11325);
  not csa_tree_add_190_195_groupi_g37608(csa_tree_add_190_195_groupi_n_11324 ,csa_tree_add_190_195_groupi_n_11323);
  or csa_tree_add_190_195_groupi_g37609(csa_tree_add_190_195_groupi_n_11322 ,csa_tree_add_190_195_groupi_n_11149 ,csa_tree_add_190_195_groupi_n_10841);
  nor csa_tree_add_190_195_groupi_g37610(csa_tree_add_190_195_groupi_n_11321 ,csa_tree_add_190_195_groupi_n_10581 ,csa_tree_add_190_195_groupi_n_11137);
  and csa_tree_add_190_195_groupi_g37611(csa_tree_add_190_195_groupi_n_11320 ,csa_tree_add_190_195_groupi_n_11149 ,csa_tree_add_190_195_groupi_n_10841);
  or csa_tree_add_190_195_groupi_g37612(csa_tree_add_190_195_groupi_n_11319 ,csa_tree_add_190_195_groupi_n_11151 ,csa_tree_add_190_195_groupi_n_11041);
  nor csa_tree_add_190_195_groupi_g37613(csa_tree_add_190_195_groupi_n_11318 ,csa_tree_add_190_195_groupi_n_11150 ,csa_tree_add_190_195_groupi_n_11042);
  or csa_tree_add_190_195_groupi_g37614(csa_tree_add_190_195_groupi_n_11317 ,csa_tree_add_190_195_groupi_n_11152 ,csa_tree_add_190_195_groupi_n_10893);
  nor csa_tree_add_190_195_groupi_g37615(csa_tree_add_190_195_groupi_n_11316 ,csa_tree_add_190_195_groupi_n_11153 ,csa_tree_add_190_195_groupi_n_10892);
  or csa_tree_add_190_195_groupi_g37616(csa_tree_add_190_195_groupi_n_11315 ,csa_tree_add_190_195_groupi_n_11064 ,csa_tree_add_190_195_groupi_n_11062);
  nor csa_tree_add_190_195_groupi_g37617(csa_tree_add_190_195_groupi_n_11314 ,csa_tree_add_190_195_groupi_n_11065 ,csa_tree_add_190_195_groupi_n_11063);
  or csa_tree_add_190_195_groupi_g37618(csa_tree_add_190_195_groupi_n_11313 ,csa_tree_add_190_195_groupi_n_11070 ,csa_tree_add_190_195_groupi_n_11073);
  and csa_tree_add_190_195_groupi_g37619(csa_tree_add_190_195_groupi_n_11312 ,csa_tree_add_190_195_groupi_n_11173 ,csa_tree_add_190_195_groupi_n_11015);
  or csa_tree_add_190_195_groupi_g37620(csa_tree_add_190_195_groupi_n_11311 ,csa_tree_add_190_195_groupi_n_10985 ,csa_tree_add_190_195_groupi_n_11133);
  or csa_tree_add_190_195_groupi_g37621(csa_tree_add_190_195_groupi_n_11310 ,csa_tree_add_190_195_groupi_n_10977 ,csa_tree_add_190_195_groupi_n_11006);
  or csa_tree_add_190_195_groupi_g37622(csa_tree_add_190_195_groupi_n_11309 ,csa_tree_add_190_195_groupi_n_10788 ,csa_tree_add_190_195_groupi_n_11129);
  nor csa_tree_add_190_195_groupi_g37623(csa_tree_add_190_195_groupi_n_11308 ,csa_tree_add_190_195_groupi_n_11071 ,csa_tree_add_190_195_groupi_n_11072);
  or csa_tree_add_190_195_groupi_g37624(csa_tree_add_190_195_groupi_n_11307 ,csa_tree_add_190_195_groupi_n_10794 ,csa_tree_add_190_195_groupi_n_11113);
  or csa_tree_add_190_195_groupi_g37625(csa_tree_add_190_195_groupi_n_11306 ,csa_tree_add_190_195_groupi_n_10981 ,csa_tree_add_190_195_groupi_n_11127);
  or csa_tree_add_190_195_groupi_g37626(csa_tree_add_190_195_groupi_n_11305 ,csa_tree_add_190_195_groupi_n_10837 ,csa_tree_add_190_195_groupi_n_11043);
  nor csa_tree_add_190_195_groupi_g37627(csa_tree_add_190_195_groupi_n_11304 ,csa_tree_add_190_195_groupi_n_10836 ,csa_tree_add_190_195_groupi_n_11044);
  or csa_tree_add_190_195_groupi_g37628(csa_tree_add_190_195_groupi_n_11303 ,csa_tree_add_190_195_groupi_n_11164 ,csa_tree_add_190_195_groupi_n_11067);
  nor csa_tree_add_190_195_groupi_g37629(csa_tree_add_190_195_groupi_n_11302 ,csa_tree_add_190_195_groupi_n_11165 ,csa_tree_add_190_195_groupi_n_11066);
  or csa_tree_add_190_195_groupi_g37630(csa_tree_add_190_195_groupi_n_11301 ,csa_tree_add_190_195_groupi_n_10798 ,csa_tree_add_190_195_groupi_n_11010);
  or csa_tree_add_190_195_groupi_g37631(csa_tree_add_190_195_groupi_n_11300 ,csa_tree_add_190_195_groupi_n_11158 ,csa_tree_add_190_195_groupi_n_10839);
  nor csa_tree_add_190_195_groupi_g37632(csa_tree_add_190_195_groupi_n_11299 ,csa_tree_add_190_195_groupi_n_11159 ,csa_tree_add_190_195_groupi_n_10840);
  or csa_tree_add_190_195_groupi_g37633(csa_tree_add_190_195_groupi_n_11298 ,csa_tree_add_190_195_groupi_n_10778 ,csa_tree_add_190_195_groupi_n_11120);
  or csa_tree_add_190_195_groupi_g37634(csa_tree_add_190_195_groupi_n_11297 ,csa_tree_add_190_195_groupi_n_11090 ,csa_tree_add_190_195_groupi_n_11104);
  or csa_tree_add_190_195_groupi_g37635(csa_tree_add_190_195_groupi_n_11296 ,csa_tree_add_190_195_groupi_n_10973 ,csa_tree_add_190_195_groupi_n_11107);
  or csa_tree_add_190_195_groupi_g37636(csa_tree_add_190_195_groupi_n_11295 ,csa_tree_add_190_195_groupi_n_10781 ,csa_tree_add_190_195_groupi_n_11102);
  or csa_tree_add_190_195_groupi_g37637(csa_tree_add_190_195_groupi_n_11294 ,csa_tree_add_190_195_groupi_n_10967 ,csa_tree_add_190_195_groupi_n_11080);
  or csa_tree_add_190_195_groupi_g37638(csa_tree_add_190_195_groupi_n_11293 ,csa_tree_add_190_195_groupi_n_10969 ,csa_tree_add_190_195_groupi_n_11074);
  and csa_tree_add_190_195_groupi_g37639(csa_tree_add_190_195_groupi_n_11292 ,csa_tree_add_190_195_groupi_n_10969 ,csa_tree_add_190_195_groupi_n_11074);
  or csa_tree_add_190_195_groupi_g37640(csa_tree_add_190_195_groupi_n_11291 ,csa_tree_add_190_195_groupi_n_10801 ,csa_tree_add_190_195_groupi_n_11109);
  and csa_tree_add_190_195_groupi_g37641(csa_tree_add_190_195_groupi_n_11290 ,csa_tree_add_190_195_groupi_n_11088 ,csa_tree_add_190_195_groupi_n_11111);
  or csa_tree_add_190_195_groupi_g37642(csa_tree_add_190_195_groupi_n_11289 ,csa_tree_add_190_195_groupi_n_11019 ,csa_tree_add_190_195_groupi_n_10850);
  or csa_tree_add_190_195_groupi_g37643(csa_tree_add_190_195_groupi_n_11288 ,csa_tree_add_190_195_groupi_n_11110 ,csa_tree_add_190_195_groupi_n_10983);
  nor csa_tree_add_190_195_groupi_g37644(csa_tree_add_190_195_groupi_n_11287 ,csa_tree_add_190_195_groupi_n_11020 ,csa_tree_add_190_195_groupi_n_10851);
  or csa_tree_add_190_195_groupi_g37645(csa_tree_add_190_195_groupi_n_11286 ,csa_tree_add_190_195_groupi_n_10769 ,csa_tree_add_190_195_groupi_n_11078);
  nor csa_tree_add_190_195_groupi_g37646(csa_tree_add_190_195_groupi_n_11285 ,csa_tree_add_190_195_groupi_n_10869 ,csa_tree_add_190_195_groupi_n_11075);
  or csa_tree_add_190_195_groupi_g37647(csa_tree_add_190_195_groupi_n_11284 ,csa_tree_add_190_195_groupi_n_11069 ,csa_tree_add_190_195_groupi_n_10960);
  nor csa_tree_add_190_195_groupi_g37648(csa_tree_add_190_195_groupi_n_11283 ,csa_tree_add_190_195_groupi_n_10770 ,csa_tree_add_190_195_groupi_n_11077);
  or csa_tree_add_190_195_groupi_g37649(csa_tree_add_190_195_groupi_n_11282 ,csa_tree_add_190_195_groupi_n_10870 ,csa_tree_add_190_195_groupi_n_11060);
  or csa_tree_add_190_195_groupi_g37650(csa_tree_add_190_195_groupi_n_11281 ,csa_tree_add_190_195_groupi_n_10868 ,csa_tree_add_190_195_groupi_n_11076);
  nor csa_tree_add_190_195_groupi_g37651(csa_tree_add_190_195_groupi_n_11280 ,csa_tree_add_190_195_groupi_n_10871 ,csa_tree_add_190_195_groupi_n_11061);
  or csa_tree_add_190_195_groupi_g37652(csa_tree_add_190_195_groupi_n_11279 ,csa_tree_add_190_195_groupi_n_10669 ,csa_tree_add_190_195_groupi_n_11052);
  or csa_tree_add_190_195_groupi_g37653(csa_tree_add_190_195_groupi_n_11278 ,csa_tree_add_190_195_groupi_n_10976 ,csa_tree_add_190_195_groupi_n_11096);
  nor csa_tree_add_190_195_groupi_g37654(csa_tree_add_190_195_groupi_n_11277 ,csa_tree_add_190_195_groupi_n_11068 ,csa_tree_add_190_195_groupi_n_10961);
  nor csa_tree_add_190_195_groupi_g37655(csa_tree_add_190_195_groupi_n_11276 ,csa_tree_add_190_195_groupi_n_10668 ,csa_tree_add_190_195_groupi_n_11053);
  and csa_tree_add_190_195_groupi_g37656(csa_tree_add_190_195_groupi_n_11275 ,csa_tree_add_190_195_groupi_n_11024 ,csa_tree_add_190_195_groupi_n_10970);
  or csa_tree_add_190_195_groupi_g37657(csa_tree_add_190_195_groupi_n_11274 ,csa_tree_add_190_195_groupi_n_11040 ,csa_tree_add_190_195_groupi_n_11081);
  or csa_tree_add_190_195_groupi_g37658(csa_tree_add_190_195_groupi_n_11273 ,csa_tree_add_190_195_groupi_n_11177 ,csa_tree_add_190_195_groupi_n_11101);
  nor csa_tree_add_190_195_groupi_g37659(csa_tree_add_190_195_groupi_n_11272 ,csa_tree_add_190_195_groupi_n_11039 ,csa_tree_add_190_195_groupi_n_11082);
  or csa_tree_add_190_195_groupi_g37660(csa_tree_add_190_195_groupi_n_11271 ,csa_tree_add_190_195_groupi_n_10730 ,csa_tree_add_190_195_groupi_n_11181);
  nor csa_tree_add_190_195_groupi_g37661(csa_tree_add_190_195_groupi_n_11270 ,csa_tree_add_190_195_groupi_n_11024 ,csa_tree_add_190_195_groupi_n_10970);
  or csa_tree_add_190_195_groupi_g37662(csa_tree_add_190_195_groupi_n_11269 ,csa_tree_add_190_195_groupi_n_10793 ,csa_tree_add_190_195_groupi_n_11099);
  and csa_tree_add_190_195_groupi_g37663(csa_tree_add_190_195_groupi_n_11268 ,csa_tree_add_190_195_groupi_n_10521 ,csa_tree_add_190_195_groupi_n_11170);
  or csa_tree_add_190_195_groupi_g37664(csa_tree_add_190_195_groupi_n_11267 ,csa_tree_add_190_195_groupi_n_11089 ,csa_tree_add_190_195_groupi_n_11095);
  nor csa_tree_add_190_195_groupi_g37665(csa_tree_add_190_195_groupi_n_11266 ,csa_tree_add_190_195_groupi_n_10968 ,csa_tree_add_190_195_groupi_n_11079);
  or csa_tree_add_190_195_groupi_g37666(csa_tree_add_190_195_groupi_n_11339 ,csa_tree_add_190_195_groupi_n_10920 ,csa_tree_add_190_195_groupi_n_11139);
  and csa_tree_add_190_195_groupi_g37667(csa_tree_add_190_195_groupi_n_11338 ,csa_tree_add_190_195_groupi_n_10917 ,csa_tree_add_190_195_groupi_n_11108);
  and csa_tree_add_190_195_groupi_g37668(csa_tree_add_190_195_groupi_n_11337 ,csa_tree_add_190_195_groupi_n_10940 ,csa_tree_add_190_195_groupi_n_11123);
  and csa_tree_add_190_195_groupi_g37669(csa_tree_add_190_195_groupi_n_11336 ,csa_tree_add_190_195_groupi_n_10828 ,csa_tree_add_190_195_groupi_n_11131);
  or csa_tree_add_190_195_groupi_g37670(csa_tree_add_190_195_groupi_n_11334 ,csa_tree_add_190_195_groupi_n_10914 ,csa_tree_add_190_195_groupi_n_11118);
  and csa_tree_add_190_195_groupi_g37671(csa_tree_add_190_195_groupi_n_11333 ,csa_tree_add_190_195_groupi_n_10912 ,csa_tree_add_190_195_groupi_n_11136);
  and csa_tree_add_190_195_groupi_g37672(csa_tree_add_190_195_groupi_n_11332 ,csa_tree_add_190_195_groupi_n_10934 ,csa_tree_add_190_195_groupi_n_11119);
  or csa_tree_add_190_195_groupi_g37673(csa_tree_add_190_195_groupi_n_11331 ,csa_tree_add_190_195_groupi_n_10831 ,csa_tree_add_190_195_groupi_n_11122);
  and csa_tree_add_190_195_groupi_g37674(csa_tree_add_190_195_groupi_n_11329 ,csa_tree_add_190_195_groupi_n_10931 ,csa_tree_add_190_195_groupi_n_11124);
  or csa_tree_add_190_195_groupi_g37675(csa_tree_add_190_195_groupi_n_11327 ,csa_tree_add_190_195_groupi_n_10906 ,csa_tree_add_190_195_groupi_n_11141);
  and csa_tree_add_190_195_groupi_g37676(csa_tree_add_190_195_groupi_n_11325 ,csa_tree_add_190_195_groupi_n_10745 ,csa_tree_add_190_195_groupi_n_11121);
  or csa_tree_add_190_195_groupi_g37677(csa_tree_add_190_195_groupi_n_11323 ,csa_tree_add_190_195_groupi_n_10705 ,csa_tree_add_190_195_groupi_n_11106);
  not csa_tree_add_190_195_groupi_g37679(csa_tree_add_190_195_groupi_n_11260 ,csa_tree_add_190_195_groupi_n_11259);
  not csa_tree_add_190_195_groupi_g37680(csa_tree_add_190_195_groupi_n_11258 ,csa_tree_add_190_195_groupi_n_11257);
  not csa_tree_add_190_195_groupi_g37681(csa_tree_add_190_195_groupi_n_11254 ,csa_tree_add_190_195_groupi_n_11253);
  not csa_tree_add_190_195_groupi_g37682(csa_tree_add_190_195_groupi_n_11251 ,csa_tree_add_190_195_groupi_n_11250);
  not csa_tree_add_190_195_groupi_g37683(csa_tree_add_190_195_groupi_n_11249 ,csa_tree_add_190_195_groupi_n_11248);
  not csa_tree_add_190_195_groupi_g37684(csa_tree_add_190_195_groupi_n_11247 ,csa_tree_add_190_195_groupi_n_11246);
  not csa_tree_add_190_195_groupi_g37685(csa_tree_add_190_195_groupi_n_11245 ,csa_tree_add_190_195_groupi_n_11244);
  not csa_tree_add_190_195_groupi_g37686(csa_tree_add_190_195_groupi_n_11241 ,csa_tree_add_190_195_groupi_n_151);
  not csa_tree_add_190_195_groupi_g37687(csa_tree_add_190_195_groupi_n_11238 ,csa_tree_add_190_195_groupi_n_11237);
  not csa_tree_add_190_195_groupi_g37688(csa_tree_add_190_195_groupi_n_11236 ,csa_tree_add_190_195_groupi_n_11235);
  not csa_tree_add_190_195_groupi_g37689(csa_tree_add_190_195_groupi_n_11234 ,csa_tree_add_190_195_groupi_n_11233);
  not csa_tree_add_190_195_groupi_g37690(csa_tree_add_190_195_groupi_n_11232 ,csa_tree_add_190_195_groupi_n_11231);
  not csa_tree_add_190_195_groupi_g37691(csa_tree_add_190_195_groupi_n_11230 ,csa_tree_add_190_195_groupi_n_11229);
  not csa_tree_add_190_195_groupi_g37692(csa_tree_add_190_195_groupi_n_11228 ,csa_tree_add_190_195_groupi_n_150);
  not csa_tree_add_190_195_groupi_g37693(csa_tree_add_190_195_groupi_n_11227 ,csa_tree_add_190_195_groupi_n_11226);
  or csa_tree_add_190_195_groupi_g37694(csa_tree_add_190_195_groupi_n_11225 ,csa_tree_add_190_195_groupi_n_11057 ,csa_tree_add_190_195_groupi_n_11033);
  or csa_tree_add_190_195_groupi_g37695(csa_tree_add_190_195_groupi_n_11224 ,csa_tree_add_190_195_groupi_n_11171 ,csa_tree_add_190_195_groupi_n_11142);
  or csa_tree_add_190_195_groupi_g37696(csa_tree_add_190_195_groupi_n_11223 ,csa_tree_add_190_195_groupi_n_11143 ,csa_tree_add_190_195_groupi_n_11083);
  or csa_tree_add_190_195_groupi_g37697(csa_tree_add_190_195_groupi_n_11222 ,csa_tree_add_190_195_groupi_n_10780 ,csa_tree_add_190_195_groupi_n_11140);
  or csa_tree_add_190_195_groupi_g37698(csa_tree_add_190_195_groupi_n_11221 ,csa_tree_add_190_195_groupi_n_11156 ,csa_tree_add_190_195_groupi_n_10877);
  nor csa_tree_add_190_195_groupi_g37699(csa_tree_add_190_195_groupi_n_11220 ,csa_tree_add_190_195_groupi_n_11166 ,csa_tree_add_190_195_groupi_n_11059);
  nor csa_tree_add_190_195_groupi_g37700(csa_tree_add_190_195_groupi_n_11219 ,csa_tree_add_190_195_groupi_n_11157 ,csa_tree_add_190_195_groupi_n_10876);
  or csa_tree_add_190_195_groupi_g37701(csa_tree_add_190_195_groupi_n_11218 ,csa_tree_add_190_195_groupi_n_10797 ,csa_tree_add_190_195_groupi_n_11017);
  or csa_tree_add_190_195_groupi_g37702(csa_tree_add_190_195_groupi_n_11217 ,csa_tree_add_190_195_groupi_n_10891 ,csa_tree_add_190_195_groupi_n_11045);
  and csa_tree_add_190_195_groupi_g37703(csa_tree_add_190_195_groupi_n_11216 ,csa_tree_add_190_195_groupi_n_10703 ,csa_tree_add_190_195_groupi_n_11132);
  nor csa_tree_add_190_195_groupi_g37704(csa_tree_add_190_195_groupi_n_11215 ,csa_tree_add_190_195_groupi_n_10890 ,csa_tree_add_190_195_groupi_n_11046);
  or csa_tree_add_190_195_groupi_g37705(csa_tree_add_190_195_groupi_n_11214 ,csa_tree_add_190_195_groupi_n_11092 ,csa_tree_add_190_195_groupi_n_11009);
  nor csa_tree_add_190_195_groupi_g37706(csa_tree_add_190_195_groupi_n_11213 ,csa_tree_add_190_195_groupi_n_11056 ,csa_tree_add_190_195_groupi_n_11034);
  nor csa_tree_add_190_195_groupi_g37707(csa_tree_add_190_195_groupi_n_11212 ,csa_tree_add_190_195_groupi_n_10674 ,csa_tree_add_190_195_groupi_n_11032);
  or csa_tree_add_190_195_groupi_g37708(csa_tree_add_190_195_groupi_n_11211 ,csa_tree_add_190_195_groupi_n_10675 ,csa_tree_add_190_195_groupi_n_11031);
  and csa_tree_add_190_195_groupi_g37709(csa_tree_add_190_195_groupi_n_11210 ,csa_tree_add_190_195_groupi_n_10847 ,csa_tree_add_190_195_groupi_n_11028);
  or csa_tree_add_190_195_groupi_g37710(csa_tree_add_190_195_groupi_n_11209 ,csa_tree_add_190_195_groupi_n_10847 ,csa_tree_add_190_195_groupi_n_11028);
  or csa_tree_add_190_195_groupi_g37711(csa_tree_add_190_195_groupi_n_11208 ,csa_tree_add_190_195_groupi_n_10792 ,csa_tree_add_190_195_groupi_n_11116);
  or csa_tree_add_190_195_groupi_g37712(csa_tree_add_190_195_groupi_n_11207 ,csa_tree_add_190_195_groupi_n_11167 ,csa_tree_add_190_195_groupi_n_11058);
  xnor csa_tree_add_190_195_groupi_g37713(csa_tree_add_190_195_groupi_n_11206 ,csa_tree_add_190_195_groupi_n_10838 ,csa_tree_add_190_195_groupi_n_10788);
  xnor csa_tree_add_190_195_groupi_g37714(csa_tree_add_190_195_groupi_n_11205 ,csa_tree_add_190_195_groupi_n_10780 ,csa_tree_add_190_195_groupi_n_10882);
  xnor csa_tree_add_190_195_groupi_g37715(csa_tree_add_190_195_groupi_n_11204 ,csa_tree_add_190_195_groupi_n_10955 ,csa_tree_add_190_195_groupi_n_10985);
  xnor csa_tree_add_190_195_groupi_g37717(csa_tree_add_190_195_groupi_n_11203 ,csa_tree_add_190_195_groupi_n_10658 ,csa_tree_add_190_195_groupi_n_10982);
  xnor csa_tree_add_190_195_groupi_g37718(csa_tree_add_190_195_groupi_n_11202 ,csa_tree_add_190_195_groupi_n_10984 ,csa_tree_add_190_195_groupi_n_10851);
  xnor csa_tree_add_190_195_groupi_g37719(csa_tree_add_190_195_groupi_n_11201 ,csa_tree_add_190_195_groupi_n_10645 ,csa_tree_add_190_195_groupi_n_10895);
  xnor csa_tree_add_190_195_groupi_g37720(csa_tree_add_190_195_groupi_n_11200 ,csa_tree_add_190_195_groupi_n_9871 ,csa_tree_add_190_195_groupi_n_10957);
  xnor csa_tree_add_190_195_groupi_g37721(csa_tree_add_190_195_groupi_n_11199 ,csa_tree_add_190_195_groupi_n_10979 ,csa_tree_add_190_195_groupi_n_10871);
  xnor csa_tree_add_190_195_groupi_g37722(csa_tree_add_190_195_groupi_n_11198 ,csa_tree_add_190_195_groupi_n_10553 ,csa_tree_add_190_195_groupi_n_10858);
  xnor csa_tree_add_190_195_groupi_g37723(csa_tree_add_190_195_groupi_n_11197 ,csa_tree_add_190_195_groupi_n_10781 ,csa_tree_add_190_195_groupi_n_10901);
  xnor csa_tree_add_190_195_groupi_g37724(csa_tree_add_190_195_groupi_n_11196 ,csa_tree_add_190_195_groupi_n_10966 ,csa_tree_add_190_195_groupi_n_10897);
  xnor csa_tree_add_190_195_groupi_g37725(csa_tree_add_190_195_groupi_n_11195 ,csa_tree_add_190_195_groupi_n_10973 ,csa_tree_add_190_195_groupi_n_10899);
  xnor csa_tree_add_190_195_groupi_g37726(csa_tree_add_190_195_groupi_n_11194 ,csa_tree_add_190_195_groupi_n_10843 ,csa_tree_add_190_195_groupi_n_10791);
  xnor csa_tree_add_190_195_groupi_g37727(csa_tree_add_190_195_groupi_n_11193 ,csa_tree_add_190_195_groupi_n_10448 ,csa_tree_add_190_195_groupi_n_10976);
  xnor csa_tree_add_190_195_groupi_g37728(csa_tree_add_190_195_groupi_n_11192 ,csa_tree_add_190_195_groupi_n_10864 ,csa_tree_add_190_195_groupi_n_10862);
  xnor csa_tree_add_190_195_groupi_g37729(csa_tree_add_190_195_groupi_n_11191 ,csa_tree_add_190_195_groupi_n_10425 ,csa_tree_add_190_195_groupi_n_10887);
  xnor csa_tree_add_190_195_groupi_g37730(csa_tree_add_190_195_groupi_n_11190 ,csa_tree_add_190_195_groupi_n_10768 ,csa_tree_add_190_195_groupi_n_10846);
  xnor csa_tree_add_190_195_groupi_g37731(csa_tree_add_190_195_groupi_n_11189 ,csa_tree_add_190_195_groupi_n_10884 ,csa_tree_add_190_195_groupi_n_10655);
  xnor csa_tree_add_190_195_groupi_g37732(csa_tree_add_190_195_groupi_n_11188 ,csa_tree_add_190_195_groupi_n_10953 ,csa_tree_add_190_195_groupi_n_10867);
  xnor csa_tree_add_190_195_groupi_g37733(csa_tree_add_190_195_groupi_n_11187 ,csa_tree_add_190_195_groupi_n_10837 ,csa_tree_add_190_195_groupi_n_10986);
  xnor csa_tree_add_190_195_groupi_g37734(csa_tree_add_190_195_groupi_n_11186 ,csa_tree_add_190_195_groupi_n_10765 ,csa_tree_add_190_195_groupi_n_10856);
  xnor csa_tree_add_190_195_groupi_g37735(csa_tree_add_190_195_groupi_n_11185 ,csa_tree_add_190_195_groupi_n_10551 ,csa_tree_add_190_195_groupi_n_10854);
  or csa_tree_add_190_195_groupi_g37736(csa_tree_add_190_195_groupi_n_11265 ,csa_tree_add_190_195_groupi_n_10921 ,csa_tree_add_190_195_groupi_n_11002);
  xnor csa_tree_add_190_195_groupi_g37737(csa_tree_add_190_195_groupi_n_11264 ,csa_tree_add_190_195_groupi_n_10469 ,csa_tree_add_190_195_groupi_n_10811);
  xnor csa_tree_add_190_195_groupi_g37738(csa_tree_add_190_195_groupi_n_11263 ,csa_tree_add_190_195_groupi_n_9869 ,csa_tree_add_190_195_groupi_n_10821);
  and csa_tree_add_190_195_groupi_g37739(csa_tree_add_190_195_groupi_n_11262 ,csa_tree_add_190_195_groupi_n_10905 ,csa_tree_add_190_195_groupi_n_11018);
  xnor csa_tree_add_190_195_groupi_g37740(csa_tree_add_190_195_groupi_n_11261 ,csa_tree_add_190_195_groupi_n_10704 ,csa_tree_add_190_195_groupi_n_10824);
  xnor csa_tree_add_190_195_groupi_g37741(csa_tree_add_190_195_groupi_n_11259 ,csa_tree_add_190_195_groupi_n_10350 ,csa_tree_add_190_195_groupi_n_10817);
  xnor csa_tree_add_190_195_groupi_g37742(csa_tree_add_190_195_groupi_n_11257 ,csa_tree_add_190_195_groupi_n_10463 ,csa_tree_add_190_195_groupi_n_10809);
  xnor csa_tree_add_190_195_groupi_g37743(csa_tree_add_190_195_groupi_n_11256 ,csa_tree_add_190_195_groupi_n_10902 ,csa_tree_add_190_195_groupi_n_10826);
  and csa_tree_add_190_195_groupi_g37744(csa_tree_add_190_195_groupi_n_11255 ,csa_tree_add_190_195_groupi_n_10909 ,csa_tree_add_190_195_groupi_n_11016);
  xnor csa_tree_add_190_195_groupi_g37745(csa_tree_add_190_195_groupi_n_11253 ,csa_tree_add_190_195_groupi_n_10583 ,csa_tree_add_190_195_groupi_n_10813);
  xnor csa_tree_add_190_195_groupi_g37746(csa_tree_add_190_195_groupi_n_11252 ,csa_tree_add_190_195_groupi_n_10782 ,csa_tree_add_190_195_groupi_n_10816);
  xnor csa_tree_add_190_195_groupi_g37747(csa_tree_add_190_195_groupi_n_11250 ,csa_tree_add_190_195_groupi_n_10700 ,csa_tree_add_190_195_groupi_n_10807);
  xnor csa_tree_add_190_195_groupi_g37748(csa_tree_add_190_195_groupi_n_11248 ,csa_tree_add_190_195_groupi_n_10441 ,csa_tree_add_190_195_groupi_n_10818);
  xnor csa_tree_add_190_195_groupi_g37749(csa_tree_add_190_195_groupi_n_11246 ,csa_tree_add_190_195_groupi_n_9625 ,csa_tree_add_190_195_groupi_n_10819);
  xnor csa_tree_add_190_195_groupi_g37750(csa_tree_add_190_195_groupi_n_11244 ,csa_tree_add_190_195_groupi_n_10878 ,csa_tree_add_190_195_groupi_n_10814);
  xnor csa_tree_add_190_195_groupi_g37751(csa_tree_add_190_195_groupi_n_11243 ,csa_tree_add_190_195_groupi_n_10974 ,csa_tree_add_190_195_groupi_n_10803);
  xnor csa_tree_add_190_195_groupi_g37752(csa_tree_add_190_195_groupi_n_11242 ,csa_tree_add_190_195_groupi_n_10679 ,csa_tree_add_190_195_groupi_n_10820);
  xnor csa_tree_add_190_195_groupi_g37754(csa_tree_add_190_195_groupi_n_11240 ,csa_tree_add_190_195_groupi_n_10673 ,csa_tree_add_190_195_groupi_n_10804);
  xnor csa_tree_add_190_195_groupi_g37755(csa_tree_add_190_195_groupi_n_11239 ,csa_tree_add_190_195_groupi_n_10699 ,csa_tree_add_190_195_groupi_n_10810);
  xnor csa_tree_add_190_195_groupi_g37756(csa_tree_add_190_195_groupi_n_11237 ,csa_tree_add_190_195_groupi_n_10047 ,csa_tree_add_190_195_groupi_n_10823);
  xnor csa_tree_add_190_195_groupi_g37757(csa_tree_add_190_195_groupi_n_11235 ,csa_tree_add_190_195_groupi_n_10468 ,csa_tree_add_190_195_groupi_n_10805);
  xnor csa_tree_add_190_195_groupi_g37758(csa_tree_add_190_195_groupi_n_11233 ,csa_tree_add_190_195_groupi_n_10777 ,csa_tree_add_190_195_groupi_n_10822);
  xnor csa_tree_add_190_195_groupi_g37759(csa_tree_add_190_195_groupi_n_11231 ,csa_tree_add_190_195_groupi_n_10215 ,csa_tree_add_190_195_groupi_n_10806);
  xnor csa_tree_add_190_195_groupi_g37760(csa_tree_add_190_195_groupi_n_11229 ,csa_tree_add_190_195_groupi_n_9609 ,csa_tree_add_190_195_groupi_n_10825);
  xnor csa_tree_add_190_195_groupi_g37762(csa_tree_add_190_195_groupi_n_11226 ,csa_tree_add_190_195_groupi_n_10326 ,csa_tree_add_190_195_groupi_n_10808);
  not csa_tree_add_190_195_groupi_g37764(csa_tree_add_190_195_groupi_n_11181 ,csa_tree_add_190_195_groupi_n_11180);
  not csa_tree_add_190_195_groupi_g37765(csa_tree_add_190_195_groupi_n_11177 ,csa_tree_add_190_195_groupi_n_11176);
  not csa_tree_add_190_195_groupi_g37768(csa_tree_add_190_195_groupi_n_11169 ,csa_tree_add_190_195_groupi_n_11168);
  not csa_tree_add_190_195_groupi_g37769(csa_tree_add_190_195_groupi_n_11166 ,csa_tree_add_190_195_groupi_n_11167);
  not csa_tree_add_190_195_groupi_g37770(csa_tree_add_190_195_groupi_n_11164 ,csa_tree_add_190_195_groupi_n_11165);
  not csa_tree_add_190_195_groupi_g37771(csa_tree_add_190_195_groupi_n_11162 ,csa_tree_add_190_195_groupi_n_11163);
  not csa_tree_add_190_195_groupi_g37772(csa_tree_add_190_195_groupi_n_11160 ,csa_tree_add_190_195_groupi_n_11161);
  not csa_tree_add_190_195_groupi_g37773(csa_tree_add_190_195_groupi_n_11159 ,csa_tree_add_190_195_groupi_n_11158);
  not csa_tree_add_190_195_groupi_g37774(csa_tree_add_190_195_groupi_n_11157 ,csa_tree_add_190_195_groupi_n_11156);
  not csa_tree_add_190_195_groupi_g37775(csa_tree_add_190_195_groupi_n_11155 ,csa_tree_add_190_195_groupi_n_11154);
  not csa_tree_add_190_195_groupi_g37776(csa_tree_add_190_195_groupi_n_11152 ,csa_tree_add_190_195_groupi_n_11153);
  not csa_tree_add_190_195_groupi_g37777(csa_tree_add_190_195_groupi_n_11150 ,csa_tree_add_190_195_groupi_n_11151);
  not csa_tree_add_190_195_groupi_g37778(csa_tree_add_190_195_groupi_n_11148 ,csa_tree_add_190_195_groupi_n_11147);
  or csa_tree_add_190_195_groupi_g37779(csa_tree_add_190_195_groupi_n_11146 ,csa_tree_add_190_195_groupi_n_138 ,csa_tree_add_190_195_groupi_n_10874);
  nor csa_tree_add_190_195_groupi_g37780(csa_tree_add_190_195_groupi_n_11145 ,csa_tree_add_190_195_groupi_n_10665 ,csa_tree_add_190_195_groupi_n_10866);
  nor csa_tree_add_190_195_groupi_g37781(csa_tree_add_190_195_groupi_n_11144 ,csa_tree_add_190_195_groupi_n_8505 ,csa_tree_add_190_195_groupi_n_10878);
  and csa_tree_add_190_195_groupi_g37782(csa_tree_add_190_195_groupi_n_11143 ,csa_tree_add_190_195_groupi_n_10656 ,csa_tree_add_190_195_groupi_n_10962);
  nor csa_tree_add_190_195_groupi_g37783(csa_tree_add_190_195_groupi_n_11142 ,csa_tree_add_190_195_groupi_n_10883 ,csa_tree_add_190_195_groupi_n_10655);
  and csa_tree_add_190_195_groupi_g37784(csa_tree_add_190_195_groupi_n_11141 ,csa_tree_add_190_195_groupi_n_10827 ,csa_tree_add_190_195_groupi_n_10787);
  nor csa_tree_add_190_195_groupi_g37785(csa_tree_add_190_195_groupi_n_11140 ,csa_tree_add_190_195_groupi_n_10690 ,csa_tree_add_190_195_groupi_n_10882);
  and csa_tree_add_190_195_groupi_g37786(csa_tree_add_190_195_groupi_n_11139 ,csa_tree_add_190_195_groupi_n_10773 ,csa_tree_add_190_195_groupi_n_10919);
  or csa_tree_add_190_195_groupi_g37787(csa_tree_add_190_195_groupi_n_11138 ,csa_tree_add_190_195_groupi_n_10691 ,csa_tree_add_190_195_groupi_n_10881);
  and csa_tree_add_190_195_groupi_g37788(csa_tree_add_190_195_groupi_n_11137 ,csa_tree_add_190_195_groupi_n_8505 ,csa_tree_add_190_195_groupi_n_10878);
  or csa_tree_add_190_195_groupi_g37789(csa_tree_add_190_195_groupi_n_11136 ,csa_tree_add_190_195_groupi_n_10584 ,csa_tree_add_190_195_groupi_n_10911);
  or csa_tree_add_190_195_groupi_g37790(csa_tree_add_190_195_groupi_n_11135 ,csa_tree_add_190_195_groupi_n_10954 ,csa_tree_add_190_195_groupi_n_10677);
  or csa_tree_add_190_195_groupi_g37791(csa_tree_add_190_195_groupi_n_11134 ,csa_tree_add_190_195_groupi_n_10884 ,csa_tree_add_190_195_groupi_n_10654);
  nor csa_tree_add_190_195_groupi_g37792(csa_tree_add_190_195_groupi_n_11133 ,csa_tree_add_190_195_groupi_n_10955 ,csa_tree_add_190_195_groupi_n_10676);
  or csa_tree_add_190_195_groupi_g37793(csa_tree_add_190_195_groupi_n_11132 ,csa_tree_add_190_195_groupi_n_10424 ,csa_tree_add_190_195_groupi_n_10887);
  or csa_tree_add_190_195_groupi_g37794(csa_tree_add_190_195_groupi_n_11131 ,csa_tree_add_190_195_groupi_n_10790 ,csa_tree_add_190_195_groupi_n_10937);
  or csa_tree_add_190_195_groupi_g37795(csa_tree_add_190_195_groupi_n_11130 ,csa_tree_add_190_195_groupi_n_10153 ,csa_tree_add_190_195_groupi_n_10838);
  and csa_tree_add_190_195_groupi_g37796(csa_tree_add_190_195_groupi_n_11129 ,csa_tree_add_190_195_groupi_n_10153 ,csa_tree_add_190_195_groupi_n_10838);
  or csa_tree_add_190_195_groupi_g37797(csa_tree_add_190_195_groupi_n_11128 ,csa_tree_add_190_195_groupi_n_10953 ,csa_tree_add_190_195_groupi_n_144);
  nor csa_tree_add_190_195_groupi_g37798(csa_tree_add_190_195_groupi_n_11127 ,csa_tree_add_190_195_groupi_n_10952 ,csa_tree_add_190_195_groupi_n_10867);
  nor csa_tree_add_190_195_groupi_g37799(csa_tree_add_190_195_groupi_n_11126 ,csa_tree_add_190_195_groupi_n_10425 ,csa_tree_add_190_195_groupi_n_137);
  or csa_tree_add_190_195_groupi_g37800(csa_tree_add_190_195_groupi_n_11125 ,csa_tree_add_190_195_groupi_n_10656 ,csa_tree_add_190_195_groupi_n_10962);
  or csa_tree_add_190_195_groupi_g37801(csa_tree_add_190_195_groupi_n_11124 ,csa_tree_add_190_195_groupi_n_10589 ,csa_tree_add_190_195_groupi_n_10930);
  or csa_tree_add_190_195_groupi_g37802(csa_tree_add_190_195_groupi_n_11123 ,csa_tree_add_190_195_groupi_n_10586 ,csa_tree_add_190_195_groupi_n_10939);
  and csa_tree_add_190_195_groupi_g37803(csa_tree_add_190_195_groupi_n_11122 ,csa_tree_add_190_195_groupi_n_10982 ,csa_tree_add_190_195_groupi_n_10829);
  or csa_tree_add_190_195_groupi_g37804(csa_tree_add_190_195_groupi_n_11121 ,csa_tree_add_190_195_groupi_n_10740 ,csa_tree_add_190_195_groupi_n_10902);
  nor csa_tree_add_190_195_groupi_g37805(csa_tree_add_190_195_groupi_n_11120 ,csa_tree_add_190_195_groupi_n_10644 ,csa_tree_add_190_195_groupi_n_10895);
  or csa_tree_add_190_195_groupi_g37806(csa_tree_add_190_195_groupi_n_11119 ,csa_tree_add_190_195_groupi_n_10587 ,csa_tree_add_190_195_groupi_n_10938);
  and csa_tree_add_190_195_groupi_g37807(csa_tree_add_190_195_groupi_n_11118 ,csa_tree_add_190_195_groupi_n_10346 ,csa_tree_add_190_195_groupi_n_10908);
  or csa_tree_add_190_195_groupi_g37808(csa_tree_add_190_195_groupi_n_11117 ,csa_tree_add_190_195_groupi_n_10645 ,csa_tree_add_190_195_groupi_n_10894);
  and csa_tree_add_190_195_groupi_g37809(csa_tree_add_190_195_groupi_n_11116 ,csa_tree_add_190_195_groupi_n_10843 ,csa_tree_add_190_195_groupi_n_10842);
  or csa_tree_add_190_195_groupi_g37810(csa_tree_add_190_195_groupi_n_11115 ,csa_tree_add_190_195_groupi_n_10315 ,csa_tree_add_190_195_groupi_n_10844);
  nor csa_tree_add_190_195_groupi_g37811(csa_tree_add_190_195_groupi_n_11114 ,csa_tree_add_190_195_groupi_n_10958 ,csa_tree_add_190_195_groupi_n_10849);
  nor csa_tree_add_190_195_groupi_g37812(csa_tree_add_190_195_groupi_n_11113 ,csa_tree_add_190_195_groupi_n_9870 ,csa_tree_add_190_195_groupi_n_10957);
  or csa_tree_add_190_195_groupi_g37813(csa_tree_add_190_195_groupi_n_11112 ,csa_tree_add_190_195_groupi_n_10553 ,csa_tree_add_190_195_groupi_n_10857);
  or csa_tree_add_190_195_groupi_g37814(csa_tree_add_190_195_groupi_n_11111 ,csa_tree_add_190_195_groupi_n_10959 ,csa_tree_add_190_195_groupi_n_10848);
  nor csa_tree_add_190_195_groupi_g37815(csa_tree_add_190_195_groupi_n_11110 ,csa_tree_add_190_195_groupi_n_10552 ,csa_tree_add_190_195_groupi_n_10858);
  and csa_tree_add_190_195_groupi_g37816(csa_tree_add_190_195_groupi_n_11109 ,csa_tree_add_190_195_groupi_n_10315 ,csa_tree_add_190_195_groupi_n_10844);
  or csa_tree_add_190_195_groupi_g37817(csa_tree_add_190_195_groupi_n_11108 ,csa_tree_add_190_195_groupi_n_10776 ,csa_tree_add_190_195_groupi_n_10915);
  nor csa_tree_add_190_195_groupi_g37818(csa_tree_add_190_195_groupi_n_11107 ,csa_tree_add_190_195_groupi_n_10164 ,csa_tree_add_190_195_groupi_n_10899);
  nor csa_tree_add_190_195_groupi_g37819(csa_tree_add_190_195_groupi_n_11106 ,csa_tree_add_190_195_groupi_n_10718 ,csa_tree_add_190_195_groupi_n_10974);
  or csa_tree_add_190_195_groupi_g37820(csa_tree_add_190_195_groupi_n_11105 ,csa_tree_add_190_195_groupi_n_10885 ,csa_tree_add_190_195_groupi_n_10889);
  nor csa_tree_add_190_195_groupi_g37821(csa_tree_add_190_195_groupi_n_11104 ,csa_tree_add_190_195_groupi_n_10767 ,csa_tree_add_190_195_groupi_n_10846);
  or csa_tree_add_190_195_groupi_g37822(csa_tree_add_190_195_groupi_n_11103 ,csa_tree_add_190_195_groupi_n_10165 ,csa_tree_add_190_195_groupi_n_10898);
  nor csa_tree_add_190_195_groupi_g37823(csa_tree_add_190_195_groupi_n_11102 ,csa_tree_add_190_195_groupi_n_10901 ,csa_tree_add_190_195_groupi_n_10692);
  nor csa_tree_add_190_195_groupi_g37824(csa_tree_add_190_195_groupi_n_11101 ,csa_tree_add_190_195_groupi_n_10886 ,csa_tree_add_190_195_groupi_n_10888);
  or csa_tree_add_190_195_groupi_g37825(csa_tree_add_190_195_groupi_n_11100 ,csa_tree_add_190_195_groupi_n_10560 ,csa_tree_add_190_195_groupi_n_10963);
  nor csa_tree_add_190_195_groupi_g37826(csa_tree_add_190_195_groupi_n_11099 ,csa_tree_add_190_195_groupi_n_10561 ,csa_tree_add_190_195_groupi_n_10964);
  or csa_tree_add_190_195_groupi_g37827(csa_tree_add_190_195_groupi_n_11098 ,csa_tree_add_190_195_groupi_n_10966 ,csa_tree_add_190_195_groupi_n_10896);
  or csa_tree_add_190_195_groupi_g37828(csa_tree_add_190_195_groupi_n_11097 ,csa_tree_add_190_195_groupi_n_10900 ,csa_tree_add_190_195_groupi_n_10693);
  nor csa_tree_add_190_195_groupi_g37829(csa_tree_add_190_195_groupi_n_11096 ,csa_tree_add_190_195_groupi_n_10448 ,csa_tree_add_190_195_groupi_n_10875);
  nor csa_tree_add_190_195_groupi_g37830(csa_tree_add_190_195_groupi_n_11095 ,csa_tree_add_190_195_groupi_n_10965 ,csa_tree_add_190_195_groupi_n_10897);
  or csa_tree_add_190_195_groupi_g37831(csa_tree_add_190_195_groupi_n_11094 ,csa_tree_add_190_195_groupi_n_10768 ,csa_tree_add_190_195_groupi_n_148);
  and csa_tree_add_190_195_groupi_g37832(csa_tree_add_190_195_groupi_n_11184 ,csa_tree_add_190_195_groupi_n_10758 ,csa_tree_add_190_195_groupi_n_10913);
  or csa_tree_add_190_195_groupi_g37833(csa_tree_add_190_195_groupi_n_11183 ,csa_tree_add_190_195_groupi_n_10743 ,csa_tree_add_190_195_groupi_n_10922);
  and csa_tree_add_190_195_groupi_g37834(csa_tree_add_190_195_groupi_n_11182 ,csa_tree_add_190_195_groupi_n_10741 ,csa_tree_add_190_195_groupi_n_10924);
  or csa_tree_add_190_195_groupi_g37835(csa_tree_add_190_195_groupi_n_11180 ,csa_tree_add_190_195_groupi_n_10477 ,csa_tree_add_190_195_groupi_n_10928);
  and csa_tree_add_190_195_groupi_g37836(csa_tree_add_190_195_groupi_n_11179 ,csa_tree_add_190_195_groupi_n_10476 ,csa_tree_add_190_195_groupi_n_10929);
  and csa_tree_add_190_195_groupi_g37837(csa_tree_add_190_195_groupi_n_11178 ,csa_tree_add_190_195_groupi_n_10754 ,csa_tree_add_190_195_groupi_n_10946);
  or csa_tree_add_190_195_groupi_g37838(csa_tree_add_190_195_groupi_n_11176 ,csa_tree_add_190_195_groupi_n_10728 ,csa_tree_add_190_195_groupi_n_10932);
  and csa_tree_add_190_195_groupi_g37839(csa_tree_add_190_195_groupi_n_11175 ,csa_tree_add_190_195_groupi_n_10538 ,csa_tree_add_190_195_groupi_n_10916);
  and csa_tree_add_190_195_groupi_g37840(csa_tree_add_190_195_groupi_n_11174 ,csa_tree_add_190_195_groupi_n_10714 ,csa_tree_add_190_195_groupi_n_10951);
  or csa_tree_add_190_195_groupi_g37841(csa_tree_add_190_195_groupi_n_11173 ,csa_tree_add_190_195_groupi_n_10638 ,csa_tree_add_190_195_groupi_n_10944);
  and csa_tree_add_190_195_groupi_g37842(csa_tree_add_190_195_groupi_n_11172 ,csa_tree_add_190_195_groupi_n_10720 ,csa_tree_add_190_195_groupi_n_10935);
  and csa_tree_add_190_195_groupi_g37843(csa_tree_add_190_195_groupi_n_11171 ,csa_tree_add_190_195_groupi_n_10642 ,csa_tree_add_190_195_groupi_n_10904);
  or csa_tree_add_190_195_groupi_g37844(csa_tree_add_190_195_groupi_n_11170 ,csa_tree_add_190_195_groupi_n_10749 ,csa_tree_add_190_195_groupi_n_10830);
  and csa_tree_add_190_195_groupi_g37845(csa_tree_add_190_195_groupi_n_11168 ,csa_tree_add_190_195_groupi_n_10709 ,csa_tree_add_190_195_groupi_n_10933);
  and csa_tree_add_190_195_groupi_g37846(csa_tree_add_190_195_groupi_n_11167 ,csa_tree_add_190_195_groupi_n_10732 ,csa_tree_add_190_195_groupi_n_10942);
  or csa_tree_add_190_195_groupi_g37847(csa_tree_add_190_195_groupi_n_11165 ,csa_tree_add_190_195_groupi_n_10753 ,csa_tree_add_190_195_groupi_n_10943);
  and csa_tree_add_190_195_groupi_g37848(csa_tree_add_190_195_groupi_n_11163 ,csa_tree_add_190_195_groupi_n_10403 ,csa_tree_add_190_195_groupi_n_10927);
  or csa_tree_add_190_195_groupi_g37849(csa_tree_add_190_195_groupi_n_11161 ,csa_tree_add_190_195_groupi_n_10760 ,csa_tree_add_190_195_groupi_n_10910);
  and csa_tree_add_190_195_groupi_g37850(csa_tree_add_190_195_groupi_n_11158 ,csa_tree_add_190_195_groupi_n_10236 ,csa_tree_add_190_195_groupi_n_10936);
  or csa_tree_add_190_195_groupi_g37851(csa_tree_add_190_195_groupi_n_11156 ,csa_tree_add_190_195_groupi_n_10724 ,csa_tree_add_190_195_groupi_n_10941);
  or csa_tree_add_190_195_groupi_g37852(csa_tree_add_190_195_groupi_n_11154 ,csa_tree_add_190_195_groupi_n_10757 ,csa_tree_add_190_195_groupi_n_10947);
  or csa_tree_add_190_195_groupi_g37853(csa_tree_add_190_195_groupi_n_11153 ,csa_tree_add_190_195_groupi_n_10297 ,csa_tree_add_190_195_groupi_n_10948);
  and csa_tree_add_190_195_groupi_g37854(csa_tree_add_190_195_groupi_n_11151 ,csa_tree_add_190_195_groupi_n_10727 ,csa_tree_add_190_195_groupi_n_10949);
  and csa_tree_add_190_195_groupi_g37855(csa_tree_add_190_195_groupi_n_11149 ,csa_tree_add_190_195_groupi_n_10735 ,csa_tree_add_190_195_groupi_n_10950);
  or csa_tree_add_190_195_groupi_g37856(csa_tree_add_190_195_groupi_n_11147 ,csa_tree_add_190_195_groupi_n_10308 ,csa_tree_add_190_195_groupi_n_10918);
  not csa_tree_add_190_195_groupi_g37857(csa_tree_add_190_195_groupi_n_11092 ,csa_tree_add_190_195_groupi_n_11091);
  not csa_tree_add_190_195_groupi_g37858(csa_tree_add_190_195_groupi_n_11085 ,csa_tree_add_190_195_groupi_n_11084);
  not csa_tree_add_190_195_groupi_g37860(csa_tree_add_190_195_groupi_n_11082 ,csa_tree_add_190_195_groupi_n_11081);
  not csa_tree_add_190_195_groupi_g37861(csa_tree_add_190_195_groupi_n_11080 ,csa_tree_add_190_195_groupi_n_11079);
  not csa_tree_add_190_195_groupi_g37862(csa_tree_add_190_195_groupi_n_11078 ,csa_tree_add_190_195_groupi_n_11077);
  not csa_tree_add_190_195_groupi_g37863(csa_tree_add_190_195_groupi_n_11076 ,csa_tree_add_190_195_groupi_n_11075);
  not csa_tree_add_190_195_groupi_g37864(csa_tree_add_190_195_groupi_n_11073 ,csa_tree_add_190_195_groupi_n_11072);
  not csa_tree_add_190_195_groupi_g37865(csa_tree_add_190_195_groupi_n_11071 ,csa_tree_add_190_195_groupi_n_11070);
  not csa_tree_add_190_195_groupi_g37866(csa_tree_add_190_195_groupi_n_11069 ,csa_tree_add_190_195_groupi_n_11068);
  not csa_tree_add_190_195_groupi_g37867(csa_tree_add_190_195_groupi_n_11067 ,csa_tree_add_190_195_groupi_n_11066);
  not csa_tree_add_190_195_groupi_g37868(csa_tree_add_190_195_groupi_n_11065 ,csa_tree_add_190_195_groupi_n_11064);
  not csa_tree_add_190_195_groupi_g37869(csa_tree_add_190_195_groupi_n_11063 ,csa_tree_add_190_195_groupi_n_11062);
  not csa_tree_add_190_195_groupi_g37870(csa_tree_add_190_195_groupi_n_11061 ,csa_tree_add_190_195_groupi_n_11060);
  not csa_tree_add_190_195_groupi_g37871(csa_tree_add_190_195_groupi_n_11059 ,csa_tree_add_190_195_groupi_n_11058);
  not csa_tree_add_190_195_groupi_g37872(csa_tree_add_190_195_groupi_n_11056 ,csa_tree_add_190_195_groupi_n_11057);
  not csa_tree_add_190_195_groupi_g37873(csa_tree_add_190_195_groupi_n_11054 ,csa_tree_add_190_195_groupi_n_11055);
  not csa_tree_add_190_195_groupi_g37874(csa_tree_add_190_195_groupi_n_11053 ,csa_tree_add_190_195_groupi_n_11052);
  not csa_tree_add_190_195_groupi_g37875(csa_tree_add_190_195_groupi_n_11050 ,csa_tree_add_190_195_groupi_n_11049);
  not csa_tree_add_190_195_groupi_g37876(csa_tree_add_190_195_groupi_n_11048 ,csa_tree_add_190_195_groupi_n_11047);
  not csa_tree_add_190_195_groupi_g37877(csa_tree_add_190_195_groupi_n_11046 ,csa_tree_add_190_195_groupi_n_11045);
  not csa_tree_add_190_195_groupi_g37878(csa_tree_add_190_195_groupi_n_11044 ,csa_tree_add_190_195_groupi_n_11043);
  not csa_tree_add_190_195_groupi_g37879(csa_tree_add_190_195_groupi_n_11042 ,csa_tree_add_190_195_groupi_n_11041);
  not csa_tree_add_190_195_groupi_g37880(csa_tree_add_190_195_groupi_n_11040 ,csa_tree_add_190_195_groupi_n_11039);
  not csa_tree_add_190_195_groupi_g37881(csa_tree_add_190_195_groupi_n_11038 ,csa_tree_add_190_195_groupi_n_11037);
  not csa_tree_add_190_195_groupi_g37882(csa_tree_add_190_195_groupi_n_11036 ,csa_tree_add_190_195_groupi_n_11035);
  not csa_tree_add_190_195_groupi_g37883(csa_tree_add_190_195_groupi_n_11034 ,csa_tree_add_190_195_groupi_n_11033);
  not csa_tree_add_190_195_groupi_g37884(csa_tree_add_190_195_groupi_n_11032 ,csa_tree_add_190_195_groupi_n_11031);
  not csa_tree_add_190_195_groupi_g37885(csa_tree_add_190_195_groupi_n_11030 ,csa_tree_add_190_195_groupi_n_11029);
  not csa_tree_add_190_195_groupi_g37886(csa_tree_add_190_195_groupi_n_11026 ,csa_tree_add_190_195_groupi_n_11025);
  not csa_tree_add_190_195_groupi_g37887(csa_tree_add_190_195_groupi_n_11024 ,csa_tree_add_190_195_groupi_n_11023);
  not csa_tree_add_190_195_groupi_g37888(csa_tree_add_190_195_groupi_n_11022 ,csa_tree_add_190_195_groupi_n_11021);
  not csa_tree_add_190_195_groupi_g37889(csa_tree_add_190_195_groupi_n_11020 ,csa_tree_add_190_195_groupi_n_11019);
  or csa_tree_add_190_195_groupi_g37890(csa_tree_add_190_195_groupi_n_11018 ,csa_tree_add_190_195_groupi_n_10702 ,csa_tree_add_190_195_groupi_n_10925);
  nor csa_tree_add_190_195_groupi_g37891(csa_tree_add_190_195_groupi_n_11017 ,csa_tree_add_190_195_groupi_n_10651 ,csa_tree_add_190_195_groupi_n_10873);
  or csa_tree_add_190_195_groupi_g37892(csa_tree_add_190_195_groupi_n_11016 ,csa_tree_add_190_195_groupi_n_10971 ,csa_tree_add_190_195_groupi_n_10832);
  or csa_tree_add_190_195_groupi_g37893(csa_tree_add_190_195_groupi_n_11015 ,csa_tree_add_190_195_groupi_n_10666 ,csa_tree_add_190_195_groupi_n_10865);
  nor csa_tree_add_190_195_groupi_g37894(csa_tree_add_190_195_groupi_n_11014 ,csa_tree_add_190_195_groupi_n_10863 ,csa_tree_add_190_195_groupi_n_10862);
  or csa_tree_add_190_195_groupi_g37895(csa_tree_add_190_195_groupi_n_11013 ,csa_tree_add_190_195_groupi_n_10864 ,csa_tree_add_190_195_groupi_n_10861);
  or csa_tree_add_190_195_groupi_g37896(csa_tree_add_190_195_groupi_n_11012 ,csa_tree_add_190_195_groupi_n_10456 ,csa_tree_add_190_195_groupi_n_10859);
  or csa_tree_add_190_195_groupi_g37897(csa_tree_add_190_195_groupi_n_11011 ,csa_tree_add_190_195_groupi_n_10650 ,csa_tree_add_190_195_groupi_n_10872);
  nor csa_tree_add_190_195_groupi_g37898(csa_tree_add_190_195_groupi_n_11010 ,csa_tree_add_190_195_groupi_n_10457 ,csa_tree_add_190_195_groupi_n_10860);
  nor csa_tree_add_190_195_groupi_g37899(csa_tree_add_190_195_groupi_n_11009 ,csa_tree_add_190_195_groupi_n_10765 ,csa_tree_add_190_195_groupi_n_10856);
  or csa_tree_add_190_195_groupi_g37900(csa_tree_add_190_195_groupi_n_11008 ,csa_tree_add_190_195_groupi_n_10764 ,csa_tree_add_190_195_groupi_n_10855);
  or csa_tree_add_190_195_groupi_g37901(csa_tree_add_190_195_groupi_n_11007 ,csa_tree_add_190_195_groupi_n_10551 ,csa_tree_add_190_195_groupi_n_10853);
  nor csa_tree_add_190_195_groupi_g37902(csa_tree_add_190_195_groupi_n_11006 ,csa_tree_add_190_195_groupi_n_10550 ,csa_tree_add_190_195_groupi_n_10854);
  or csa_tree_add_190_195_groupi_g37903(csa_tree_add_190_195_groupi_n_11005 ,csa_tree_add_190_195_groupi_n_10843 ,csa_tree_add_190_195_groupi_n_10842);
  or csa_tree_add_190_195_groupi_g37904(csa_tree_add_190_195_groupi_n_11004 ,csa_tree_add_190_195_groupi_n_9871 ,csa_tree_add_190_195_groupi_n_10956);
  xnor csa_tree_add_190_195_groupi_g37905(out1[2] ,csa_tree_add_190_195_groupi_n_9775 ,csa_tree_add_190_195_groupi_n_146);
  nor csa_tree_add_190_195_groupi_g37906(csa_tree_add_190_195_groupi_n_11002 ,csa_tree_add_190_195_groupi_n_10783 ,csa_tree_add_190_195_groupi_n_10923);
  xnor csa_tree_add_190_195_groupi_g37907(csa_tree_add_190_195_groupi_n_11001 ,csa_tree_add_190_195_groupi_n_10445 ,csa_tree_add_190_195_groupi_n_10685);
  xnor csa_tree_add_190_195_groupi_g37909(csa_tree_add_190_195_groupi_n_11000 ,csa_tree_add_190_195_groupi_n_10437 ,csa_tree_add_190_195_groupi_n_10800);
  xnor csa_tree_add_190_195_groupi_g37910(csa_tree_add_190_195_groupi_n_10999 ,csa_tree_add_190_195_groupi_n_10647 ,csa_tree_add_190_195_groupi_n_10667);
  xnor csa_tree_add_190_195_groupi_g37911(csa_tree_add_190_195_groupi_n_10998 ,csa_tree_add_190_195_groupi_n_10460 ,csa_tree_add_190_195_groupi_n_10649);
  xnor csa_tree_add_190_195_groupi_g37912(csa_tree_add_190_195_groupi_n_10997 ,csa_tree_add_190_195_groupi_n_10037 ,csa_tree_add_190_195_groupi_n_10772);
  xor csa_tree_add_190_195_groupi_g37914(csa_tree_add_190_195_groupi_n_10996 ,csa_tree_add_190_195_groupi_n_10801 ,csa_tree_add_190_195_groupi_n_10315);
  xnor csa_tree_add_190_195_groupi_g37915(csa_tree_add_190_195_groupi_n_10995 ,csa_tree_add_190_195_groupi_n_10702 ,csa_tree_add_190_195_groupi_n_10683);
  xnor csa_tree_add_190_195_groupi_g37917(csa_tree_add_190_195_groupi_n_10994 ,csa_tree_add_190_195_groupi_n_10457 ,csa_tree_add_190_195_groupi_n_10798);
  xnor csa_tree_add_190_195_groupi_g37918(csa_tree_add_190_195_groupi_n_10993 ,csa_tree_add_190_195_groupi_n_10321 ,csa_tree_add_190_195_groupi_n_10779);
  xnor csa_tree_add_190_195_groupi_g37919(csa_tree_add_190_195_groupi_n_10992 ,csa_tree_add_190_195_groupi_n_10651 ,csa_tree_add_190_195_groupi_n_10797);
  xnor csa_tree_add_190_195_groupi_g37920(csa_tree_add_190_195_groupi_n_10991 ,csa_tree_add_190_195_groupi_n_10561 ,csa_tree_add_190_195_groupi_n_10793);
  xnor csa_tree_add_190_195_groupi_g37921(csa_tree_add_190_195_groupi_n_10990 ,csa_tree_add_190_195_groupi_n_10660 ,csa_tree_add_190_195_groupi_n_10773);
  xnor csa_tree_add_190_195_groupi_g37922(csa_tree_add_190_195_groupi_n_10989 ,csa_tree_add_190_195_groupi_n_10584 ,csa_tree_add_190_195_groupi_n_10664);
  xnor csa_tree_add_190_195_groupi_g37923(csa_tree_add_190_195_groupi_n_10988 ,csa_tree_add_190_195_groupi_n_9782 ,csa_tree_add_190_195_groupi_n_10787);
  xnor csa_tree_add_190_195_groupi_g37924(csa_tree_add_190_195_groupi_n_10987 ,csa_tree_add_190_195_groupi_n_10564 ,csa_tree_add_190_195_groupi_n_10689);
  and csa_tree_add_190_195_groupi_g37925(csa_tree_add_190_195_groupi_n_11093 ,csa_tree_add_190_195_groupi_n_9852 ,csa_tree_add_190_195_groupi_n_10945);
  xnor csa_tree_add_190_195_groupi_g37926(csa_tree_add_190_195_groupi_n_11091 ,csa_tree_add_190_195_groupi_n_10231 ,csa_tree_add_190_195_groupi_n_10618);
  xnor csa_tree_add_190_195_groupi_g37927(csa_tree_add_190_195_groupi_n_11090 ,csa_tree_add_190_195_groupi_n_9949 ,csa_tree_add_190_195_groupi_n_10597);
  xnor csa_tree_add_190_195_groupi_g37928(csa_tree_add_190_195_groupi_n_11089 ,csa_tree_add_190_195_groupi_n_9915 ,csa_tree_add_190_195_groupi_n_10601);
  xnor csa_tree_add_190_195_groupi_g37929(csa_tree_add_190_195_groupi_n_11088 ,csa_tree_add_190_195_groupi_n_9611 ,csa_tree_add_190_195_groupi_n_10615);
  xnor csa_tree_add_190_195_groupi_g37930(csa_tree_add_190_195_groupi_n_11087 ,csa_tree_add_190_195_groupi_n_8683 ,csa_tree_add_190_195_groupi_n_10617);
  and csa_tree_add_190_195_groupi_g37931(csa_tree_add_190_195_groupi_n_11086 ,csa_tree_add_190_195_groupi_n_10628 ,csa_tree_add_190_195_groupi_n_10833);
  or csa_tree_add_190_195_groupi_g37932(csa_tree_add_190_195_groupi_n_11084 ,csa_tree_add_190_195_groupi_n_10630 ,csa_tree_add_190_195_groupi_n_10834);
  xnor csa_tree_add_190_195_groupi_g37933(csa_tree_add_190_195_groupi_n_11083 ,csa_tree_add_190_195_groupi_n_7640 ,csa_tree_add_190_195_groupi_n_10603);
  xnor csa_tree_add_190_195_groupi_g37934(csa_tree_add_190_195_groupi_n_11081 ,csa_tree_add_190_195_groupi_n_10167 ,csa_tree_add_190_195_groupi_n_10606);
  xnor csa_tree_add_190_195_groupi_g37935(csa_tree_add_190_195_groupi_n_11079 ,csa_tree_add_190_195_groupi_n_10228 ,csa_tree_add_190_195_groupi_n_10599);
  xnor csa_tree_add_190_195_groupi_g37936(csa_tree_add_190_195_groupi_n_11077 ,csa_tree_add_190_195_groupi_n_9874 ,csa_tree_add_190_195_groupi_n_10614);
  xnor csa_tree_add_190_195_groupi_g37937(csa_tree_add_190_195_groupi_n_11075 ,csa_tree_add_190_195_groupi_n_9503 ,csa_tree_add_190_195_groupi_n_145);
  xnor csa_tree_add_190_195_groupi_g37938(csa_tree_add_190_195_groupi_n_11074 ,csa_tree_add_190_195_groupi_n_9660 ,csa_tree_add_190_195_groupi_n_10592);
  xnor csa_tree_add_190_195_groupi_g37939(csa_tree_add_190_195_groupi_n_11072 ,csa_tree_add_190_195_groupi_n_10473 ,csa_tree_add_190_195_groupi_n_10594);
  xnor csa_tree_add_190_195_groupi_g37940(csa_tree_add_190_195_groupi_n_11070 ,csa_tree_add_190_195_groupi_n_10342 ,csa_tree_add_190_195_groupi_n_10593);
  xnor csa_tree_add_190_195_groupi_g37941(csa_tree_add_190_195_groupi_n_11068 ,csa_tree_add_190_195_groupi_n_10591 ,csa_tree_add_190_195_groupi_n_10613);
  xnor csa_tree_add_190_195_groupi_g37942(csa_tree_add_190_195_groupi_n_11066 ,csa_tree_add_190_195_groupi_n_10068 ,csa_tree_add_190_195_groupi_n_10595);
  xnor csa_tree_add_190_195_groupi_g37943(csa_tree_add_190_195_groupi_n_11064 ,csa_tree_add_190_195_groupi_n_9322 ,csa_tree_add_190_195_groupi_n_10596);
  xnor csa_tree_add_190_195_groupi_g37944(csa_tree_add_190_195_groupi_n_11062 ,csa_tree_add_190_195_groupi_n_9941 ,csa_tree_add_190_195_groupi_n_10598);
  xnor csa_tree_add_190_195_groupi_g37945(csa_tree_add_190_195_groupi_n_11060 ,csa_tree_add_190_195_groupi_n_9896 ,csa_tree_add_190_195_groupi_n_10612);
  xnor csa_tree_add_190_195_groupi_g37946(csa_tree_add_190_195_groupi_n_11058 ,csa_tree_add_190_195_groupi_n_9757 ,csa_tree_add_190_195_groupi_n_149);
  and csa_tree_add_190_195_groupi_g37947(csa_tree_add_190_195_groupi_n_11057 ,csa_tree_add_190_195_groupi_n_10635 ,csa_tree_add_190_195_groupi_n_10835);
  or csa_tree_add_190_195_groupi_g37948(csa_tree_add_190_195_groupi_n_11055 ,csa_tree_add_190_195_groupi_n_10633 ,csa_tree_add_190_195_groupi_n_10907);
  xnor csa_tree_add_190_195_groupi_g37949(csa_tree_add_190_195_groupi_n_11052 ,csa_tree_add_190_195_groupi_n_9634 ,csa_tree_add_190_195_groupi_n_10609);
  xnor csa_tree_add_190_195_groupi_g37950(csa_tree_add_190_195_groupi_n_11051 ,csa_tree_add_190_195_groupi_n_10582 ,csa_tree_add_190_195_groupi_n_10608);
  xnor csa_tree_add_190_195_groupi_g37951(csa_tree_add_190_195_groupi_n_11049 ,csa_tree_add_190_195_groupi_n_10784 ,csa_tree_add_190_195_groupi_n_10616);
  xnor csa_tree_add_190_195_groupi_g37952(csa_tree_add_190_195_groupi_n_11047 ,csa_tree_add_190_195_groupi_n_10465 ,csa_tree_add_190_195_groupi_n_10604);
  xnor csa_tree_add_190_195_groupi_g37953(csa_tree_add_190_195_groupi_n_11045 ,csa_tree_add_190_195_groupi_n_10799 ,csa_tree_add_190_195_groupi_n_10610);
  xnor csa_tree_add_190_195_groupi_g37954(csa_tree_add_190_195_groupi_n_11043 ,csa_tree_add_190_195_groupi_n_10467 ,csa_tree_add_190_195_groupi_n_10611);
  xnor csa_tree_add_190_195_groupi_g37955(csa_tree_add_190_195_groupi_n_11041 ,csa_tree_add_190_195_groupi_n_10802 ,csa_tree_add_190_195_groupi_n_10105);
  xnor csa_tree_add_190_195_groupi_g37956(csa_tree_add_190_195_groupi_n_11039 ,csa_tree_add_190_195_groupi_n_9943 ,csa_tree_add_190_195_groupi_n_10607);
  xnor csa_tree_add_190_195_groupi_g37957(csa_tree_add_190_195_groupi_n_11037 ,csa_tree_add_190_195_groupi_n_10774 ,csa_tree_add_190_195_groupi_n_10357);
  and csa_tree_add_190_195_groupi_g37958(csa_tree_add_190_195_groupi_n_11035 ,csa_tree_add_190_195_groupi_n_10640 ,csa_tree_add_190_195_groupi_n_10926);
  xnor csa_tree_add_190_195_groupi_g37959(csa_tree_add_190_195_groupi_n_11033 ,csa_tree_add_190_195_groupi_n_10427 ,csa_tree_add_190_195_groupi_n_10619);
  xnor csa_tree_add_190_195_groupi_g37960(csa_tree_add_190_195_groupi_n_11031 ,csa_tree_add_190_195_groupi_n_10169 ,csa_tree_add_190_195_groupi_n_10621);
  xnor csa_tree_add_190_195_groupi_g37961(csa_tree_add_190_195_groupi_n_11029 ,csa_tree_add_190_195_groupi_n_10694 ,csa_tree_add_190_195_groupi_n_10624);
  xnor csa_tree_add_190_195_groupi_g37962(csa_tree_add_190_195_groupi_n_11028 ,csa_tree_add_190_195_groupi_n_10180 ,csa_tree_add_190_195_groupi_n_10623);
  xnor csa_tree_add_190_195_groupi_g37963(csa_tree_add_190_195_groupi_n_11027 ,csa_tree_add_190_195_groupi_n_9933 ,csa_tree_add_190_195_groupi_n_10605);
  xnor csa_tree_add_190_195_groupi_g37964(csa_tree_add_190_195_groupi_n_11025 ,csa_tree_add_190_195_groupi_n_10074 ,csa_tree_add_190_195_groupi_n_10622);
  xnor csa_tree_add_190_195_groupi_g37965(csa_tree_add_190_195_groupi_n_11023 ,csa_tree_add_190_195_groupi_n_9291 ,csa_tree_add_190_195_groupi_n_147);
  xnor csa_tree_add_190_195_groupi_g37966(csa_tree_add_190_195_groupi_n_11021 ,csa_tree_add_190_195_groupi_n_9894 ,csa_tree_add_190_195_groupi_n_10602);
  xnor csa_tree_add_190_195_groupi_g37967(csa_tree_add_190_195_groupi_n_11019 ,csa_tree_add_190_195_groupi_n_9314 ,csa_tree_add_190_195_groupi_n_134);
  not csa_tree_add_190_195_groupi_g37969(csa_tree_add_190_195_groupi_n_10981 ,csa_tree_add_190_195_groupi_n_10980);
  not csa_tree_add_190_195_groupi_g37973(csa_tree_add_190_195_groupi_n_10967 ,csa_tree_add_190_195_groupi_n_10968);
  not csa_tree_add_190_195_groupi_g37974(csa_tree_add_190_195_groupi_n_10966 ,csa_tree_add_190_195_groupi_n_10965);
  not csa_tree_add_190_195_groupi_g37975(csa_tree_add_190_195_groupi_n_10964 ,csa_tree_add_190_195_groupi_n_10963);
  not csa_tree_add_190_195_groupi_g37976(csa_tree_add_190_195_groupi_n_10960 ,csa_tree_add_190_195_groupi_n_10961);
  not csa_tree_add_190_195_groupi_g37977(csa_tree_add_190_195_groupi_n_10959 ,csa_tree_add_190_195_groupi_n_10958);
  not csa_tree_add_190_195_groupi_g37978(csa_tree_add_190_195_groupi_n_10957 ,csa_tree_add_190_195_groupi_n_10956);
  not csa_tree_add_190_195_groupi_g37979(csa_tree_add_190_195_groupi_n_10954 ,csa_tree_add_190_195_groupi_n_10955);
  not csa_tree_add_190_195_groupi_g37980(csa_tree_add_190_195_groupi_n_10952 ,csa_tree_add_190_195_groupi_n_10953);
  or csa_tree_add_190_195_groupi_g37981(csa_tree_add_190_195_groupi_n_10951 ,csa_tree_add_190_195_groupi_n_10779 ,csa_tree_add_190_195_groupi_n_10713);
  or csa_tree_add_190_195_groupi_g37982(csa_tree_add_190_195_groupi_n_10950 ,csa_tree_add_190_195_groupi_n_10067 ,csa_tree_add_190_195_groupi_n_10734);
  or csa_tree_add_190_195_groupi_g37983(csa_tree_add_190_195_groupi_n_10949 ,csa_tree_add_190_195_groupi_n_10468 ,csa_tree_add_190_195_groupi_n_10726);
  and csa_tree_add_190_195_groupi_g37984(csa_tree_add_190_195_groupi_n_10948 ,csa_tree_add_190_195_groupi_n_10305 ,csa_tree_add_190_195_groupi_n_10772);
  and csa_tree_add_190_195_groupi_g37985(csa_tree_add_190_195_groupi_n_10947 ,csa_tree_add_190_195_groupi_n_10583 ,csa_tree_add_190_195_groupi_n_10755);
  or csa_tree_add_190_195_groupi_g37986(csa_tree_add_190_195_groupi_n_10946 ,csa_tree_add_190_195_groupi_n_10777 ,csa_tree_add_190_195_groupi_n_10762);
  or csa_tree_add_190_195_groupi_g37987(csa_tree_add_190_195_groupi_n_10945 ,csa_tree_add_190_195_groupi_n_9851 ,csa_tree_add_190_195_groupi_n_10802);
  and csa_tree_add_190_195_groupi_g37988(csa_tree_add_190_195_groupi_n_10944 ,csa_tree_add_190_195_groupi_n_10636 ,csa_tree_add_190_195_groupi_n_10469);
  nor csa_tree_add_190_195_groupi_g37989(csa_tree_add_190_195_groupi_n_10943 ,csa_tree_add_190_195_groupi_n_9789 ,csa_tree_add_190_195_groupi_n_10756);
  or csa_tree_add_190_195_groupi_g37990(csa_tree_add_190_195_groupi_n_10942 ,csa_tree_add_190_195_groupi_n_10588 ,csa_tree_add_190_195_groupi_n_10731);
  nor csa_tree_add_190_195_groupi_g37991(csa_tree_add_190_195_groupi_n_10941 ,csa_tree_add_190_195_groupi_n_9957 ,csa_tree_add_190_195_groupi_n_10723);
  or csa_tree_add_190_195_groupi_g37992(csa_tree_add_190_195_groupi_n_10940 ,csa_tree_add_190_195_groupi_n_10647 ,csa_tree_add_190_195_groupi_n_135);
  nor csa_tree_add_190_195_groupi_g37993(csa_tree_add_190_195_groupi_n_10939 ,csa_tree_add_190_195_groupi_n_10646 ,csa_tree_add_190_195_groupi_n_10667);
  nor csa_tree_add_190_195_groupi_g37994(csa_tree_add_190_195_groupi_n_10938 ,csa_tree_add_190_195_groupi_n_10450 ,csa_tree_add_190_195_groupi_n_10679);
  nor csa_tree_add_190_195_groupi_g37995(csa_tree_add_190_195_groupi_n_10937 ,csa_tree_add_190_195_groupi_n_10460 ,csa_tree_add_190_195_groupi_n_10649);
  or csa_tree_add_190_195_groupi_g37996(csa_tree_add_190_195_groupi_n_10936 ,csa_tree_add_190_195_groupi_n_10240 ,csa_tree_add_190_195_groupi_n_10698);
  or csa_tree_add_190_195_groupi_g37997(csa_tree_add_190_195_groupi_n_10935 ,csa_tree_add_190_195_groupi_n_10577 ,csa_tree_add_190_195_groupi_n_10719);
  or csa_tree_add_190_195_groupi_g37998(csa_tree_add_190_195_groupi_n_10934 ,csa_tree_add_190_195_groupi_n_10449 ,csa_tree_add_190_195_groupi_n_10678);
  or csa_tree_add_190_195_groupi_g37999(csa_tree_add_190_195_groupi_n_10933 ,csa_tree_add_190_195_groupi_n_10701 ,csa_tree_add_190_195_groupi_n_10707);
  nor csa_tree_add_190_195_groupi_g38000(csa_tree_add_190_195_groupi_n_10932 ,csa_tree_add_190_195_groupi_n_10341 ,csa_tree_add_190_195_groupi_n_10733);
  or csa_tree_add_190_195_groupi_g38001(csa_tree_add_190_195_groupi_n_10931 ,csa_tree_add_190_195_groupi_n_10210 ,csa_tree_add_190_195_groupi_n_10672);
  nor csa_tree_add_190_195_groupi_g38002(csa_tree_add_190_195_groupi_n_10930 ,csa_tree_add_190_195_groupi_n_10211 ,csa_tree_add_190_195_groupi_n_10673);
  or csa_tree_add_190_195_groupi_g38003(csa_tree_add_190_195_groupi_n_10929 ,csa_tree_add_190_195_groupi_n_10482 ,csa_tree_add_190_195_groupi_n_10796);
  and csa_tree_add_190_195_groupi_g38004(csa_tree_add_190_195_groupi_n_10928 ,csa_tree_add_190_195_groupi_n_10487 ,csa_tree_add_190_195_groupi_n_10799);
  or csa_tree_add_190_195_groupi_g38005(csa_tree_add_190_195_groupi_n_10927 ,csa_tree_add_190_195_groupi_n_10549 ,csa_tree_add_190_195_groupi_n_10784);
  or csa_tree_add_190_195_groupi_g38006(csa_tree_add_190_195_groupi_n_10926 ,csa_tree_add_190_195_groupi_n_10704 ,csa_tree_add_190_195_groupi_n_10639);
  nor csa_tree_add_190_195_groupi_g38007(csa_tree_add_190_195_groupi_n_10925 ,csa_tree_add_190_195_groupi_n_10157 ,csa_tree_add_190_195_groupi_n_10683);
  or csa_tree_add_190_195_groupi_g38008(csa_tree_add_190_195_groupi_n_10924 ,csa_tree_add_190_195_groupi_n_10355 ,csa_tree_add_190_195_groupi_n_10746);
  and csa_tree_add_190_195_groupi_g38009(csa_tree_add_190_195_groupi_n_10923 ,csa_tree_add_190_195_groupi_n_10458 ,csa_tree_add_190_195_groupi_n_10687);
  nor csa_tree_add_190_195_groupi_g38010(csa_tree_add_190_195_groupi_n_10922 ,csa_tree_add_190_195_groupi_n_10590 ,csa_tree_add_190_195_groupi_n_10750);
  nor csa_tree_add_190_195_groupi_g38011(csa_tree_add_190_195_groupi_n_10921 ,csa_tree_add_190_195_groupi_n_10458 ,csa_tree_add_190_195_groupi_n_10687);
  nor csa_tree_add_190_195_groupi_g38012(csa_tree_add_190_195_groupi_n_10920 ,csa_tree_add_190_195_groupi_n_10660 ,csa_tree_add_190_195_groupi_n_10661);
  or csa_tree_add_190_195_groupi_g38013(csa_tree_add_190_195_groupi_n_10919 ,csa_tree_add_190_195_groupi_n_10659 ,csa_tree_add_190_195_groupi_n_10662);
  nor csa_tree_add_190_195_groupi_g38014(csa_tree_add_190_195_groupi_n_10918 ,csa_tree_add_190_195_groupi_n_10143 ,csa_tree_add_190_195_groupi_n_10774);
  or csa_tree_add_190_195_groupi_g38015(csa_tree_add_190_195_groupi_n_10917 ,csa_tree_add_190_195_groupi_n_10564 ,csa_tree_add_190_195_groupi_n_10688);
  or csa_tree_add_190_195_groupi_g38016(csa_tree_add_190_195_groupi_n_10916 ,csa_tree_add_190_195_groupi_n_10539 ,csa_tree_add_190_195_groupi_n_10695);
  nor csa_tree_add_190_195_groupi_g38017(csa_tree_add_190_195_groupi_n_10915 ,csa_tree_add_190_195_groupi_n_10563 ,csa_tree_add_190_195_groupi_n_10689);
  nor csa_tree_add_190_195_groupi_g38018(csa_tree_add_190_195_groupi_n_10914 ,csa_tree_add_190_195_groupi_n_10445 ,csa_tree_add_190_195_groupi_n_10684);
  or csa_tree_add_190_195_groupi_g38019(csa_tree_add_190_195_groupi_n_10913 ,csa_tree_add_190_195_groupi_n_10578 ,csa_tree_add_190_195_groupi_n_10759);
  or csa_tree_add_190_195_groupi_g38020(csa_tree_add_190_195_groupi_n_10912 ,csa_tree_add_190_195_groupi_n_10432 ,csa_tree_add_190_195_groupi_n_10663);
  nor csa_tree_add_190_195_groupi_g38021(csa_tree_add_190_195_groupi_n_10911 ,csa_tree_add_190_195_groupi_n_10433 ,csa_tree_add_190_195_groupi_n_10664);
  and csa_tree_add_190_195_groupi_g38022(csa_tree_add_190_195_groupi_n_10910 ,csa_tree_add_190_195_groupi_n_10761 ,csa_tree_add_190_195_groupi_n_10782);
  or csa_tree_add_190_195_groupi_g38023(csa_tree_add_190_195_groupi_n_10909 ,csa_tree_add_190_195_groupi_n_10766 ,csa_tree_add_190_195_groupi_n_10671);
  or csa_tree_add_190_195_groupi_g38024(csa_tree_add_190_195_groupi_n_10908 ,csa_tree_add_190_195_groupi_n_10444 ,csa_tree_add_190_195_groupi_n_10685);
  and csa_tree_add_190_195_groupi_g38025(csa_tree_add_190_195_groupi_n_10907 ,csa_tree_add_190_195_groupi_n_10632 ,csa_tree_add_190_195_groupi_n_10699);
  nor csa_tree_add_190_195_groupi_g38026(csa_tree_add_190_195_groupi_n_10906 ,csa_tree_add_190_195_groupi_n_9782 ,csa_tree_add_190_195_groupi_n_10681);
  or csa_tree_add_190_195_groupi_g38027(csa_tree_add_190_195_groupi_n_10905 ,csa_tree_add_190_195_groupi_n_10156 ,csa_tree_add_190_195_groupi_n_10682);
  or csa_tree_add_190_195_groupi_g38028(csa_tree_add_190_195_groupi_n_10904 ,csa_tree_add_190_195_groupi_n_10347 ,csa_tree_add_190_195_groupi_n_10641);
  and csa_tree_add_190_195_groupi_g38029(csa_tree_add_190_195_groupi_n_10986 ,csa_tree_add_190_195_groupi_n_10411 ,csa_tree_add_190_195_groupi_n_10643);
  and csa_tree_add_190_195_groupi_g38030(csa_tree_add_190_195_groupi_n_10985 ,csa_tree_add_190_195_groupi_n_10412 ,csa_tree_add_190_195_groupi_n_10712);
  and csa_tree_add_190_195_groupi_g38031(csa_tree_add_190_195_groupi_n_10984 ,csa_tree_add_190_195_groupi_n_10495 ,csa_tree_add_190_195_groupi_n_10716);
  and csa_tree_add_190_195_groupi_g38032(csa_tree_add_190_195_groupi_n_10983 ,csa_tree_add_190_195_groupi_n_10493 ,csa_tree_add_190_195_groupi_n_10715);
  or csa_tree_add_190_195_groupi_g38033(csa_tree_add_190_195_groupi_n_10982 ,csa_tree_add_190_195_groupi_n_10400 ,csa_tree_add_190_195_groupi_n_10725);
  or csa_tree_add_190_195_groupi_g38034(csa_tree_add_190_195_groupi_n_10980 ,csa_tree_add_190_195_groupi_n_10414 ,csa_tree_add_190_195_groupi_n_10637);
  and csa_tree_add_190_195_groupi_g38035(csa_tree_add_190_195_groupi_n_10979 ,csa_tree_add_190_195_groupi_n_10490 ,csa_tree_add_190_195_groupi_n_10711);
  and csa_tree_add_190_195_groupi_g38036(csa_tree_add_190_195_groupi_n_10978 ,csa_tree_add_190_195_groupi_n_10277 ,csa_tree_add_190_195_groupi_n_10708);
  and csa_tree_add_190_195_groupi_g38037(csa_tree_add_190_195_groupi_n_10977 ,csa_tree_add_190_195_groupi_n_10419 ,csa_tree_add_190_195_groupi_n_10744);
  and csa_tree_add_190_195_groupi_g38038(csa_tree_add_190_195_groupi_n_10976 ,csa_tree_add_190_195_groupi_n_10486 ,csa_tree_add_190_195_groupi_n_10738);
  and csa_tree_add_190_195_groupi_g38039(csa_tree_add_190_195_groupi_n_10975 ,csa_tree_add_190_195_groupi_n_10485 ,csa_tree_add_190_195_groupi_n_10706);
  and csa_tree_add_190_195_groupi_g38040(csa_tree_add_190_195_groupi_n_10974 ,csa_tree_add_190_195_groupi_n_10481 ,csa_tree_add_190_195_groupi_n_10722);
  and csa_tree_add_190_195_groupi_g38041(csa_tree_add_190_195_groupi_n_10973 ,csa_tree_add_190_195_groupi_n_10535 ,csa_tree_add_190_195_groupi_n_10752);
  and csa_tree_add_190_195_groupi_g38042(csa_tree_add_190_195_groupi_n_10972 ,csa_tree_add_190_195_groupi_n_10479 ,csa_tree_add_190_195_groupi_n_10729);
  and csa_tree_add_190_195_groupi_g38043(csa_tree_add_190_195_groupi_n_10971 ,csa_tree_add_190_195_groupi_n_10409 ,csa_tree_add_190_195_groupi_n_10627);
  and csa_tree_add_190_195_groupi_g38044(csa_tree_add_190_195_groupi_n_10970 ,csa_tree_add_190_195_groupi_n_10500 ,csa_tree_add_190_195_groupi_n_10737);
  and csa_tree_add_190_195_groupi_g38045(csa_tree_add_190_195_groupi_n_10969 ,csa_tree_add_190_195_groupi_n_10525 ,csa_tree_add_190_195_groupi_n_10751);
  and csa_tree_add_190_195_groupi_g38046(csa_tree_add_190_195_groupi_n_10968 ,csa_tree_add_190_195_groupi_n_10513 ,csa_tree_add_190_195_groupi_n_10742);
  or csa_tree_add_190_195_groupi_g38047(csa_tree_add_190_195_groupi_n_10965 ,csa_tree_add_190_195_groupi_n_10511 ,csa_tree_add_190_195_groupi_n_10739);
  and csa_tree_add_190_195_groupi_g38048(csa_tree_add_190_195_groupi_n_10963 ,csa_tree_add_190_195_groupi_n_10504 ,csa_tree_add_190_195_groupi_n_10736);
  and csa_tree_add_190_195_groupi_g38049(csa_tree_add_190_195_groupi_n_10962 ,csa_tree_add_190_195_groupi_n_10395 ,csa_tree_add_190_195_groupi_n_10634);
  or csa_tree_add_190_195_groupi_g38050(csa_tree_add_190_195_groupi_n_10961 ,csa_tree_add_190_195_groupi_n_10491 ,csa_tree_add_190_195_groupi_n_10710);
  and csa_tree_add_190_195_groupi_g38051(csa_tree_add_190_195_groupi_n_10958 ,csa_tree_add_190_195_groupi_n_10499 ,csa_tree_add_190_195_groupi_n_10763);
  and csa_tree_add_190_195_groupi_g38052(csa_tree_add_190_195_groupi_n_10956 ,csa_tree_add_190_195_groupi_n_10502 ,csa_tree_add_190_195_groupi_n_10721);
  or csa_tree_add_190_195_groupi_g38053(csa_tree_add_190_195_groupi_n_10955 ,csa_tree_add_190_195_groupi_n_10267 ,csa_tree_add_190_195_groupi_n_10747);
  and csa_tree_add_190_195_groupi_g38054(csa_tree_add_190_195_groupi_n_10953 ,csa_tree_add_190_195_groupi_n_10526 ,csa_tree_add_190_195_groupi_n_10748);
  not csa_tree_add_190_195_groupi_g38055(csa_tree_add_190_195_groupi_n_10901 ,csa_tree_add_190_195_groupi_n_10900);
  not csa_tree_add_190_195_groupi_g38056(csa_tree_add_190_195_groupi_n_10899 ,csa_tree_add_190_195_groupi_n_10898);
  not csa_tree_add_190_195_groupi_g38057(csa_tree_add_190_195_groupi_n_10897 ,csa_tree_add_190_195_groupi_n_10896);
  not csa_tree_add_190_195_groupi_g38058(csa_tree_add_190_195_groupi_n_10895 ,csa_tree_add_190_195_groupi_n_10894);
  not csa_tree_add_190_195_groupi_g38059(csa_tree_add_190_195_groupi_n_10893 ,csa_tree_add_190_195_groupi_n_10892);
  not csa_tree_add_190_195_groupi_g38060(csa_tree_add_190_195_groupi_n_10891 ,csa_tree_add_190_195_groupi_n_10890);
  not csa_tree_add_190_195_groupi_g38061(csa_tree_add_190_195_groupi_n_10889 ,csa_tree_add_190_195_groupi_n_10888);
  not csa_tree_add_190_195_groupi_g38062(csa_tree_add_190_195_groupi_n_10887 ,csa_tree_add_190_195_groupi_n_137);
  not csa_tree_add_190_195_groupi_g38063(csa_tree_add_190_195_groupi_n_10886 ,csa_tree_add_190_195_groupi_n_10885);
  not csa_tree_add_190_195_groupi_g38064(csa_tree_add_190_195_groupi_n_10884 ,csa_tree_add_190_195_groupi_n_10883);
  not csa_tree_add_190_195_groupi_g38065(csa_tree_add_190_195_groupi_n_10882 ,csa_tree_add_190_195_groupi_n_10881);
  not csa_tree_add_190_195_groupi_g38066(csa_tree_add_190_195_groupi_n_10880 ,csa_tree_add_190_195_groupi_n_10879);
  not csa_tree_add_190_195_groupi_g38067(csa_tree_add_190_195_groupi_n_10877 ,csa_tree_add_190_195_groupi_n_10876);
  not csa_tree_add_190_195_groupi_g38068(csa_tree_add_190_195_groupi_n_10875 ,csa_tree_add_190_195_groupi_n_10874);
  not csa_tree_add_190_195_groupi_g38069(csa_tree_add_190_195_groupi_n_10873 ,csa_tree_add_190_195_groupi_n_10872);
  not csa_tree_add_190_195_groupi_g38070(csa_tree_add_190_195_groupi_n_10871 ,csa_tree_add_190_195_groupi_n_10870);
  not csa_tree_add_190_195_groupi_g38071(csa_tree_add_190_195_groupi_n_10869 ,csa_tree_add_190_195_groupi_n_10868);
  not csa_tree_add_190_195_groupi_g38072(csa_tree_add_190_195_groupi_n_10867 ,csa_tree_add_190_195_groupi_n_144);
  not csa_tree_add_190_195_groupi_g38073(csa_tree_add_190_195_groupi_n_10866 ,csa_tree_add_190_195_groupi_n_10865);
  not csa_tree_add_190_195_groupi_g38074(csa_tree_add_190_195_groupi_n_10864 ,csa_tree_add_190_195_groupi_n_10863);
  not csa_tree_add_190_195_groupi_g38075(csa_tree_add_190_195_groupi_n_10862 ,csa_tree_add_190_195_groupi_n_10861);
  not csa_tree_add_190_195_groupi_g38076(csa_tree_add_190_195_groupi_n_10860 ,csa_tree_add_190_195_groupi_n_10859);
  not csa_tree_add_190_195_groupi_g38077(csa_tree_add_190_195_groupi_n_10858 ,csa_tree_add_190_195_groupi_n_10857);
  not csa_tree_add_190_195_groupi_g38078(csa_tree_add_190_195_groupi_n_10856 ,csa_tree_add_190_195_groupi_n_10855);
  not csa_tree_add_190_195_groupi_g38079(csa_tree_add_190_195_groupi_n_10854 ,csa_tree_add_190_195_groupi_n_10853);
  not csa_tree_add_190_195_groupi_g38080(csa_tree_add_190_195_groupi_n_10852 ,csa_tree_add_190_195_groupi_n_139);
  not csa_tree_add_190_195_groupi_g38081(csa_tree_add_190_195_groupi_n_10851 ,csa_tree_add_190_195_groupi_n_10850);
  not csa_tree_add_190_195_groupi_g38082(csa_tree_add_190_195_groupi_n_10849 ,csa_tree_add_190_195_groupi_n_10848);
  not csa_tree_add_190_195_groupi_g38083(csa_tree_add_190_195_groupi_n_10846 ,csa_tree_add_190_195_groupi_n_148);
  not csa_tree_add_190_195_groupi_g38084(csa_tree_add_190_195_groupi_n_10845 ,csa_tree_add_190_195_groupi_n_140);
  not csa_tree_add_190_195_groupi_g38085(csa_tree_add_190_195_groupi_n_10840 ,csa_tree_add_190_195_groupi_n_10839);
  not csa_tree_add_190_195_groupi_g38086(csa_tree_add_190_195_groupi_n_10837 ,csa_tree_add_190_195_groupi_n_10836);
  or csa_tree_add_190_195_groupi_g38087(csa_tree_add_190_195_groupi_n_10835 ,csa_tree_add_190_195_groupi_n_10344 ,csa_tree_add_190_195_groupi_n_10631);
  and csa_tree_add_190_195_groupi_g38088(csa_tree_add_190_195_groupi_n_10834 ,csa_tree_add_190_195_groupi_n_10800 ,csa_tree_add_190_195_groupi_n_10629);
  or csa_tree_add_190_195_groupi_g38089(csa_tree_add_190_195_groupi_n_10833 ,csa_tree_add_190_195_groupi_n_10696 ,csa_tree_add_190_195_groupi_n_10626);
  and csa_tree_add_190_195_groupi_g38090(csa_tree_add_190_195_groupi_n_10832 ,csa_tree_add_190_195_groupi_n_10766 ,csa_tree_add_190_195_groupi_n_10671);
  nor csa_tree_add_190_195_groupi_g38091(csa_tree_add_190_195_groupi_n_10831 ,csa_tree_add_190_195_groupi_n_10652 ,csa_tree_add_190_195_groupi_n_10658);
  and csa_tree_add_190_195_groupi_g38092(csa_tree_add_190_195_groupi_n_10830 ,csa_tree_add_190_195_groupi_n_10625 ,csa_tree_add_190_195_groupi_n_10350);
  or csa_tree_add_190_195_groupi_g38093(csa_tree_add_190_195_groupi_n_10829 ,csa_tree_add_190_195_groupi_n_10653 ,csa_tree_add_190_195_groupi_n_10657);
  or csa_tree_add_190_195_groupi_g38094(csa_tree_add_190_195_groupi_n_10828 ,csa_tree_add_190_195_groupi_n_10459 ,csa_tree_add_190_195_groupi_n_10648);
  or csa_tree_add_190_195_groupi_g38095(csa_tree_add_190_195_groupi_n_10827 ,csa_tree_add_190_195_groupi_n_9781 ,csa_tree_add_190_195_groupi_n_10680);
  xnor csa_tree_add_190_195_groupi_g38096(csa_tree_add_190_195_groupi_n_10826 ,csa_tree_add_190_195_groupi_n_10046 ,csa_tree_add_190_195_groupi_n_10559);
  xnor csa_tree_add_190_195_groupi_g38097(csa_tree_add_190_195_groupi_n_10825 ,csa_tree_add_190_195_groupi_n_10474 ,csa_tree_add_190_195_groupi_n_10206);
  xnor csa_tree_add_190_195_groupi_g38098(csa_tree_add_190_195_groupi_n_10824 ,csa_tree_add_190_195_groupi_n_10455 ,csa_tree_add_190_195_groupi_n_10190);
  xnor csa_tree_add_190_195_groupi_g38099(csa_tree_add_190_195_groupi_n_10823 ,csa_tree_add_190_195_groupi_n_10443 ,csa_tree_add_190_195_groupi_n_10343);
  xnor csa_tree_add_190_195_groupi_g38100(csa_tree_add_190_195_groupi_n_10822 ,csa_tree_add_190_195_groupi_n_10570 ,csa_tree_add_190_195_groupi_n_10209);
  xnor csa_tree_add_190_195_groupi_g38101(csa_tree_add_190_195_groupi_n_10821 ,csa_tree_add_190_195_groupi_n_10588 ,csa_tree_add_190_195_groupi_n_10422);
  xnor csa_tree_add_190_195_groupi_g38102(csa_tree_add_190_195_groupi_n_10820 ,csa_tree_add_190_195_groupi_n_10587 ,csa_tree_add_190_195_groupi_n_10450);
  xnor csa_tree_add_190_195_groupi_g38103(csa_tree_add_190_195_groupi_n_10819 ,csa_tree_add_190_195_groupi_n_10341 ,csa_tree_add_190_195_groupi_n_10423);
  xnor csa_tree_add_190_195_groupi_g38104(csa_tree_add_190_195_groupi_n_10818 ,csa_tree_add_190_195_groupi_n_10213 ,csa_tree_add_190_195_groupi_n_10578);
  xnor csa_tree_add_190_195_groupi_g38105(csa_tree_add_190_195_groupi_n_10817 ,csa_tree_add_190_195_groupi_n_9638 ,csa_tree_add_190_195_groupi_n_10568);
  xnor csa_tree_add_190_195_groupi_g38106(csa_tree_add_190_195_groupi_n_10816 ,csa_tree_add_190_195_groupi_n_10208 ,csa_tree_add_190_195_groupi_n_10431);
  xnor csa_tree_add_190_195_groupi_g38107(csa_tree_add_190_195_groupi_n_10815 ,csa_tree_add_190_195_groupi_n_10429 ,csa_tree_add_190_195_groupi_n_10161);
  xnor csa_tree_add_190_195_groupi_g38108(csa_tree_add_190_195_groupi_n_10814 ,csa_tree_add_190_195_groupi_n_10581 ,csa_tree_add_190_195_groupi_n_8505);
  xnor csa_tree_add_190_195_groupi_g38109(csa_tree_add_190_195_groupi_n_10813 ,csa_tree_add_190_195_groupi_n_10330 ,csa_tree_add_190_195_groupi_n_10555);
  xnor csa_tree_add_190_195_groupi_g38110(csa_tree_add_190_195_groupi_n_10812 ,csa_tree_add_190_195_groupi_n_10576 ,csa_tree_add_190_195_groupi_n_10447);
  xnor csa_tree_add_190_195_groupi_g38111(csa_tree_add_190_195_groupi_n_10811 ,csa_tree_add_190_195_groupi_n_10186 ,csa_tree_add_190_195_groupi_n_10452);
  xnor csa_tree_add_190_195_groupi_g38112(csa_tree_add_190_195_groupi_n_10810 ,csa_tree_add_190_195_groupi_n_10172 ,csa_tree_add_190_195_groupi_n_10439);
  xnor csa_tree_add_190_195_groupi_g38113(csa_tree_add_190_195_groupi_n_10809 ,csa_tree_add_190_195_groupi_n_10466 ,csa_tree_add_190_195_groupi_n_10590);
  xnor csa_tree_add_190_195_groupi_g38114(csa_tree_add_190_195_groupi_n_10808 ,csa_tree_add_190_195_groupi_n_10204 ,csa_tree_add_190_195_groupi_n_10470);
  xnor csa_tree_add_190_195_groupi_g38115(csa_tree_add_190_195_groupi_n_10807 ,csa_tree_add_190_195_groupi_n_10454 ,csa_tree_add_190_195_groupi_n_10557);
  xnor csa_tree_add_190_195_groupi_g38116(csa_tree_add_190_195_groupi_n_10806 ,csa_tree_add_190_195_groupi_n_10214 ,csa_tree_add_190_195_groupi_n_10579);
  xnor csa_tree_add_190_195_groupi_g38117(csa_tree_add_190_195_groupi_n_10805 ,csa_tree_add_190_195_groupi_n_10420 ,csa_tree_add_190_195_groupi_n_9776);
  xnor csa_tree_add_190_195_groupi_g38118(csa_tree_add_190_195_groupi_n_10804 ,csa_tree_add_190_195_groupi_n_10211 ,csa_tree_add_190_195_groupi_n_10589);
  xnor csa_tree_add_190_195_groupi_g38119(csa_tree_add_190_195_groupi_n_10803 ,csa_tree_add_190_195_groupi_n_10152 ,csa_tree_add_190_195_groupi_n_10565);
  xnor csa_tree_add_190_195_groupi_g38120(csa_tree_add_190_195_groupi_n_10903 ,csa_tree_add_190_195_groupi_n_10471 ,csa_tree_add_190_195_groupi_n_10375);
  xnor csa_tree_add_190_195_groupi_g38121(csa_tree_add_190_195_groupi_n_10902 ,csa_tree_add_190_195_groupi_n_9806 ,csa_tree_add_190_195_groupi_n_10376);
  xnor csa_tree_add_190_195_groupi_g38122(csa_tree_add_190_195_groupi_n_10900 ,csa_tree_add_190_195_groupi_n_9807 ,csa_tree_add_190_195_groupi_n_10373);
  xnor csa_tree_add_190_195_groupi_g38123(csa_tree_add_190_195_groupi_n_10898 ,csa_tree_add_190_195_groupi_n_9177 ,csa_tree_add_190_195_groupi_n_10372);
  xnor csa_tree_add_190_195_groupi_g38124(csa_tree_add_190_195_groupi_n_10896 ,csa_tree_add_190_195_groupi_n_9773 ,csa_tree_add_190_195_groupi_n_10377);
  xnor csa_tree_add_190_195_groupi_g38125(csa_tree_add_190_195_groupi_n_10894 ,csa_tree_add_190_195_groupi_n_10421 ,csa_tree_add_190_195_groupi_n_10370);
  xnor csa_tree_add_190_195_groupi_g38126(csa_tree_add_190_195_groupi_n_10892 ,csa_tree_add_190_195_groupi_n_10338 ,csa_tree_add_190_195_groupi_n_10378);
  xnor csa_tree_add_190_195_groupi_g38127(csa_tree_add_190_195_groupi_n_10890 ,csa_tree_add_190_195_groupi_n_9313 ,csa_tree_add_190_195_groupi_n_10358);
  xnor csa_tree_add_190_195_groupi_g38128(csa_tree_add_190_195_groupi_n_10888 ,csa_tree_add_190_195_groupi_n_8626 ,csa_tree_add_190_195_groupi_n_10380);
  xnor csa_tree_add_190_195_groupi_g38130(csa_tree_add_190_195_groupi_n_10885 ,csa_tree_add_190_195_groupi_n_10198 ,csa_tree_add_190_195_groupi_n_10381);
  xnor csa_tree_add_190_195_groupi_g38131(csa_tree_add_190_195_groupi_n_10883 ,csa_tree_add_190_195_groupi_n_9800 ,csa_tree_add_190_195_groupi_n_10366);
  xnor csa_tree_add_190_195_groupi_g38132(csa_tree_add_190_195_groupi_n_10881 ,csa_tree_add_190_195_groupi_n_9332 ,csa_tree_add_190_195_groupi_n_10365);
  xnor csa_tree_add_190_195_groupi_g38133(csa_tree_add_190_195_groupi_n_10879 ,csa_tree_add_190_195_groupi_n_10071 ,csa_tree_add_190_195_groupi_n_10364);
  xnor csa_tree_add_190_195_groupi_g38134(csa_tree_add_190_195_groupi_n_10878 ,csa_tree_add_190_195_groupi_n_9021 ,csa_tree_add_190_195_groupi_n_10382);
  xnor csa_tree_add_190_195_groupi_g38135(csa_tree_add_190_195_groupi_n_10876 ,csa_tree_add_190_195_groupi_n_10442 ,csa_tree_add_190_195_groupi_n_10363);
  xnor csa_tree_add_190_195_groupi_g38136(csa_tree_add_190_195_groupi_n_10874 ,csa_tree_add_190_195_groupi_n_10233 ,csa_tree_add_190_195_groupi_n_10379);
  xnor csa_tree_add_190_195_groupi_g38137(csa_tree_add_190_195_groupi_n_10872 ,csa_tree_add_190_195_groupi_n_9962 ,csa_tree_add_190_195_groupi_n_10362);
  xnor csa_tree_add_190_195_groupi_g38138(csa_tree_add_190_195_groupi_n_10870 ,csa_tree_add_190_195_groupi_n_10221 ,csa_tree_add_190_195_groupi_n_10386);
  xnor csa_tree_add_190_195_groupi_g38139(csa_tree_add_190_195_groupi_n_10868 ,csa_tree_add_190_195_groupi_n_9347 ,csa_tree_add_190_195_groupi_n_10387);
  xnor csa_tree_add_190_195_groupi_g38141(csa_tree_add_190_195_groupi_n_10865 ,csa_tree_add_190_195_groupi_n_10351 ,csa_tree_add_190_195_groupi_n_10369);
  xnor csa_tree_add_190_195_groupi_g38142(csa_tree_add_190_195_groupi_n_10863 ,csa_tree_add_190_195_groupi_n_9759 ,csa_tree_add_190_195_groupi_n_10360);
  xnor csa_tree_add_190_195_groupi_g38143(csa_tree_add_190_195_groupi_n_10861 ,csa_tree_add_190_195_groupi_n_10562 ,csa_tree_add_190_195_groupi_n_10359);
  xnor csa_tree_add_190_195_groupi_g38144(csa_tree_add_190_195_groupi_n_10859 ,csa_tree_add_190_195_groupi_n_9911 ,csa_tree_add_190_195_groupi_n_10374);
  xnor csa_tree_add_190_195_groupi_g38145(csa_tree_add_190_195_groupi_n_10857 ,csa_tree_add_190_195_groupi_n_10060 ,csa_tree_add_190_195_groupi_n_10388);
  xnor csa_tree_add_190_195_groupi_g38146(csa_tree_add_190_195_groupi_n_10855 ,csa_tree_add_190_195_groupi_n_9951 ,csa_tree_add_190_195_groupi_n_10356);
  xnor csa_tree_add_190_195_groupi_g38147(csa_tree_add_190_195_groupi_n_10853 ,csa_tree_add_190_195_groupi_n_9954 ,csa_tree_add_190_195_groupi_n_10385);
  xnor csa_tree_add_190_195_groupi_g38149(csa_tree_add_190_195_groupi_n_10850 ,csa_tree_add_190_195_groupi_n_8689 ,csa_tree_add_190_195_groupi_n_10389);
  xnor csa_tree_add_190_195_groupi_g38150(csa_tree_add_190_195_groupi_n_10848 ,csa_tree_add_190_195_groupi_n_9754 ,csa_tree_add_190_195_groupi_n_142);
  xnor csa_tree_add_190_195_groupi_g38151(csa_tree_add_190_195_groupi_n_10847 ,csa_tree_add_190_195_groupi_n_9901 ,csa_tree_add_190_195_groupi_n_10383);
  xnor csa_tree_add_190_195_groupi_g38154(csa_tree_add_190_195_groupi_n_10844 ,csa_tree_add_190_195_groupi_n_10339 ,csa_tree_add_190_195_groupi_n_10390);
  xnor csa_tree_add_190_195_groupi_g38155(csa_tree_add_190_195_groupi_n_10843 ,csa_tree_add_190_195_groupi_n_9490 ,csa_tree_add_190_195_groupi_n_136);
  xnor csa_tree_add_190_195_groupi_g38156(csa_tree_add_190_195_groupi_n_10842 ,csa_tree_add_190_195_groupi_n_7553 ,csa_tree_add_190_195_groupi_n_141);
  xnor csa_tree_add_190_195_groupi_g38157(csa_tree_add_190_195_groupi_n_10841 ,csa_tree_add_190_195_groupi_n_7631 ,csa_tree_add_190_195_groupi_n_10391);
  xnor csa_tree_add_190_195_groupi_g38158(csa_tree_add_190_195_groupi_n_10839 ,csa_tree_add_190_195_groupi_n_10585 ,csa_tree_add_190_195_groupi_n_10392);
  xnor csa_tree_add_190_195_groupi_g38159(csa_tree_add_190_195_groupi_n_10838 ,csa_tree_add_190_195_groupi_n_9798 ,csa_tree_add_190_195_groupi_n_10393);
  xnor csa_tree_add_190_195_groupi_g38160(csa_tree_add_190_195_groupi_n_10836 ,csa_tree_add_190_195_groupi_n_10314 ,csa_tree_add_190_195_groupi_n_10394);
  not csa_tree_add_190_195_groupi_g38162(csa_tree_add_190_195_groupi_n_10792 ,csa_tree_add_190_195_groupi_n_10791);
  not csa_tree_add_190_195_groupi_g38163(csa_tree_add_190_195_groupi_n_10790 ,csa_tree_add_190_195_groupi_n_10789);
  not csa_tree_add_190_195_groupi_g38166(csa_tree_add_190_195_groupi_n_10776 ,csa_tree_add_190_195_groupi_n_10775);
  not csa_tree_add_190_195_groupi_g38167(csa_tree_add_190_195_groupi_n_10770 ,csa_tree_add_190_195_groupi_n_10769);
  not csa_tree_add_190_195_groupi_g38168(csa_tree_add_190_195_groupi_n_10768 ,csa_tree_add_190_195_groupi_n_10767);
  not csa_tree_add_190_195_groupi_g38169(csa_tree_add_190_195_groupi_n_10765 ,csa_tree_add_190_195_groupi_n_10764);
  or csa_tree_add_190_195_groupi_g38170(csa_tree_add_190_195_groupi_n_10763 ,csa_tree_add_190_195_groupi_n_10497 ,csa_tree_add_190_195_groupi_n_10335);
  nor csa_tree_add_190_195_groupi_g38171(csa_tree_add_190_195_groupi_n_10762 ,csa_tree_add_190_195_groupi_n_10569 ,csa_tree_add_190_195_groupi_n_10209);
  or csa_tree_add_190_195_groupi_g38172(csa_tree_add_190_195_groupi_n_10761 ,csa_tree_add_190_195_groupi_n_10207 ,csa_tree_add_190_195_groupi_n_10431);
  nor csa_tree_add_190_195_groupi_g38173(csa_tree_add_190_195_groupi_n_10760 ,csa_tree_add_190_195_groupi_n_10208 ,csa_tree_add_190_195_groupi_n_10430);
  nor csa_tree_add_190_195_groupi_g38174(csa_tree_add_190_195_groupi_n_10759 ,csa_tree_add_190_195_groupi_n_10441 ,csa_tree_add_190_195_groupi_n_10213);
  or csa_tree_add_190_195_groupi_g38175(csa_tree_add_190_195_groupi_n_10758 ,csa_tree_add_190_195_groupi_n_10440 ,csa_tree_add_190_195_groupi_n_10212);
  nor csa_tree_add_190_195_groupi_g38176(csa_tree_add_190_195_groupi_n_10757 ,csa_tree_add_190_195_groupi_n_10330 ,csa_tree_add_190_195_groupi_n_10554);
  nor csa_tree_add_190_195_groupi_g38177(csa_tree_add_190_195_groupi_n_10756 ,csa_tree_add_190_195_groupi_n_9934 ,csa_tree_add_190_195_groupi_n_10442);
  or csa_tree_add_190_195_groupi_g38178(csa_tree_add_190_195_groupi_n_10755 ,csa_tree_add_190_195_groupi_n_10329 ,csa_tree_add_190_195_groupi_n_10555);
  or csa_tree_add_190_195_groupi_g38179(csa_tree_add_190_195_groupi_n_10754 ,csa_tree_add_190_195_groupi_n_10570 ,csa_tree_add_190_195_groupi_n_127);
  and csa_tree_add_190_195_groupi_g38180(csa_tree_add_190_195_groupi_n_10753 ,csa_tree_add_190_195_groupi_n_9934 ,csa_tree_add_190_195_groupi_n_10442);
  or csa_tree_add_190_195_groupi_g38181(csa_tree_add_190_195_groupi_n_10752 ,csa_tree_add_190_195_groupi_n_10068 ,csa_tree_add_190_195_groupi_n_10536);
  or csa_tree_add_190_195_groupi_g38182(csa_tree_add_190_195_groupi_n_10751 ,csa_tree_add_190_195_groupi_n_10582 ,csa_tree_add_190_195_groupi_n_10544);
  nor csa_tree_add_190_195_groupi_g38183(csa_tree_add_190_195_groupi_n_10750 ,csa_tree_add_190_195_groupi_n_10466 ,csa_tree_add_190_195_groupi_n_10463);
  nor csa_tree_add_190_195_groupi_g38184(csa_tree_add_190_195_groupi_n_10749 ,csa_tree_add_190_195_groupi_n_9638 ,csa_tree_add_190_195_groupi_n_10567);
  or csa_tree_add_190_195_groupi_g38185(csa_tree_add_190_195_groupi_n_10748 ,csa_tree_add_190_195_groupi_n_10078 ,csa_tree_add_190_195_groupi_n_10524);
  and csa_tree_add_190_195_groupi_g38186(csa_tree_add_190_195_groupi_n_10747 ,csa_tree_add_190_195_groupi_n_10266 ,csa_tree_add_190_195_groupi_n_10585);
  nor csa_tree_add_190_195_groupi_g38187(csa_tree_add_190_195_groupi_n_10746 ,csa_tree_add_190_195_groupi_n_10184 ,csa_tree_add_190_195_groupi_n_10427);
  or csa_tree_add_190_195_groupi_g38188(csa_tree_add_190_195_groupi_n_10745 ,csa_tree_add_190_195_groupi_n_10045 ,csa_tree_add_190_195_groupi_n_10559);
  or csa_tree_add_190_195_groupi_g38189(csa_tree_add_190_195_groupi_n_10744 ,csa_tree_add_190_195_groupi_n_10334 ,csa_tree_add_190_195_groupi_n_10406);
  and csa_tree_add_190_195_groupi_g38190(csa_tree_add_190_195_groupi_n_10743 ,csa_tree_add_190_195_groupi_n_10466 ,csa_tree_add_190_195_groupi_n_10463);
  or csa_tree_add_190_195_groupi_g38191(csa_tree_add_190_195_groupi_n_10742 ,csa_tree_add_190_195_groupi_n_10473 ,csa_tree_add_190_195_groupi_n_10514);
  or csa_tree_add_190_195_groupi_g38192(csa_tree_add_190_195_groupi_n_10741 ,csa_tree_add_190_195_groupi_n_10183 ,csa_tree_add_190_195_groupi_n_10426);
  nor csa_tree_add_190_195_groupi_g38193(csa_tree_add_190_195_groupi_n_10740 ,csa_tree_add_190_195_groupi_n_10046 ,csa_tree_add_190_195_groupi_n_10558);
  and csa_tree_add_190_195_groupi_g38194(csa_tree_add_190_195_groupi_n_10739 ,csa_tree_add_190_195_groupi_n_10342 ,csa_tree_add_190_195_groupi_n_10512);
  or csa_tree_add_190_195_groupi_g38195(csa_tree_add_190_195_groupi_n_10738 ,csa_tree_add_190_195_groupi_n_10475 ,csa_tree_add_190_195_groupi_n_10591);
  or csa_tree_add_190_195_groupi_g38196(csa_tree_add_190_195_groupi_n_10737 ,csa_tree_add_190_195_groupi_n_10074 ,csa_tree_add_190_195_groupi_n_10520);
  or csa_tree_add_190_195_groupi_g38197(csa_tree_add_190_195_groupi_n_10736 ,csa_tree_add_190_195_groupi_n_9662 ,csa_tree_add_190_195_groupi_n_10506);
  or csa_tree_add_190_195_groupi_g38198(csa_tree_add_190_195_groupi_n_10735 ,csa_tree_add_190_195_groupi_n_9640 ,csa_tree_add_190_195_groupi_n_10421);
  and csa_tree_add_190_195_groupi_g38199(csa_tree_add_190_195_groupi_n_10734 ,csa_tree_add_190_195_groupi_n_9640 ,csa_tree_add_190_195_groupi_n_10421);
  nor csa_tree_add_190_195_groupi_g38200(csa_tree_add_190_195_groupi_n_10733 ,csa_tree_add_190_195_groupi_n_9625 ,csa_tree_add_190_195_groupi_n_10423);
  or csa_tree_add_190_195_groupi_g38201(csa_tree_add_190_195_groupi_n_10732 ,csa_tree_add_190_195_groupi_n_9869 ,csa_tree_add_190_195_groupi_n_10422);
  and csa_tree_add_190_195_groupi_g38202(csa_tree_add_190_195_groupi_n_10731 ,csa_tree_add_190_195_groupi_n_9869 ,csa_tree_add_190_195_groupi_n_10422);
  nor csa_tree_add_190_195_groupi_g38203(csa_tree_add_190_195_groupi_n_10730 ,csa_tree_add_190_195_groupi_n_10571 ,csa_tree_add_190_195_groupi_n_10574);
  or csa_tree_add_190_195_groupi_g38204(csa_tree_add_190_195_groupi_n_10729 ,csa_tree_add_190_195_groupi_n_10230 ,csa_tree_add_190_195_groupi_n_10478);
  and csa_tree_add_190_195_groupi_g38205(csa_tree_add_190_195_groupi_n_10728 ,csa_tree_add_190_195_groupi_n_9625 ,csa_tree_add_190_195_groupi_n_10423);
  or csa_tree_add_190_195_groupi_g38206(csa_tree_add_190_195_groupi_n_10727 ,csa_tree_add_190_195_groupi_n_9776 ,csa_tree_add_190_195_groupi_n_10420);
  and csa_tree_add_190_195_groupi_g38207(csa_tree_add_190_195_groupi_n_10726 ,csa_tree_add_190_195_groupi_n_9776 ,csa_tree_add_190_195_groupi_n_10420);
  nor csa_tree_add_190_195_groupi_g38208(csa_tree_add_190_195_groupi_n_10725 ,csa_tree_add_190_195_groupi_n_10349 ,csa_tree_add_190_195_groupi_n_10399);
  and csa_tree_add_190_195_groupi_g38209(csa_tree_add_190_195_groupi_n_10724 ,csa_tree_add_190_195_groupi_n_9603 ,csa_tree_add_190_195_groupi_n_10562);
  nor csa_tree_add_190_195_groupi_g38210(csa_tree_add_190_195_groupi_n_10723 ,csa_tree_add_190_195_groupi_n_9603 ,csa_tree_add_190_195_groupi_n_10562);
  or csa_tree_add_190_195_groupi_g38211(csa_tree_add_190_195_groupi_n_10722 ,csa_tree_add_190_195_groupi_n_10229 ,csa_tree_add_190_195_groupi_n_10480);
  or csa_tree_add_190_195_groupi_g38212(csa_tree_add_190_195_groupi_n_10721 ,csa_tree_add_190_195_groupi_n_10086 ,csa_tree_add_190_195_groupi_n_10501);
  or csa_tree_add_190_195_groupi_g38213(csa_tree_add_190_195_groupi_n_10720 ,csa_tree_add_190_195_groupi_n_10576 ,csa_tree_add_190_195_groupi_n_10446);
  nor csa_tree_add_190_195_groupi_g38214(csa_tree_add_190_195_groupi_n_10719 ,csa_tree_add_190_195_groupi_n_10575 ,csa_tree_add_190_195_groupi_n_10447);
  and csa_tree_add_190_195_groupi_g38215(csa_tree_add_190_195_groupi_n_10718 ,csa_tree_add_190_195_groupi_n_10152 ,csa_tree_add_190_195_groupi_n_10566);
  or csa_tree_add_190_195_groupi_g38216(csa_tree_add_190_195_groupi_n_10717 ,csa_tree_add_190_195_groupi_n_10572 ,csa_tree_add_190_195_groupi_n_10573);
  or csa_tree_add_190_195_groupi_g38217(csa_tree_add_190_195_groupi_n_10716 ,csa_tree_add_190_195_groupi_n_9799 ,csa_tree_add_190_195_groupi_n_10494);
  or csa_tree_add_190_195_groupi_g38218(csa_tree_add_190_195_groupi_n_10715 ,csa_tree_add_190_195_groupi_n_10580 ,csa_tree_add_190_195_groupi_n_10492);
  or csa_tree_add_190_195_groupi_g38219(csa_tree_add_190_195_groupi_n_10714 ,csa_tree_add_190_195_groupi_n_10320 ,csa_tree_add_190_195_groupi_n_10462);
  nor csa_tree_add_190_195_groupi_g38220(csa_tree_add_190_195_groupi_n_10713 ,csa_tree_add_190_195_groupi_n_10321 ,csa_tree_add_190_195_groupi_n_10461);
  or csa_tree_add_190_195_groupi_g38221(csa_tree_add_190_195_groupi_n_10712 ,csa_tree_add_190_195_groupi_n_10226 ,csa_tree_add_190_195_groupi_n_10405);
  or csa_tree_add_190_195_groupi_g38222(csa_tree_add_190_195_groupi_n_10711 ,csa_tree_add_190_195_groupi_n_10340 ,csa_tree_add_190_195_groupi_n_10488);
  and csa_tree_add_190_195_groupi_g38223(csa_tree_add_190_195_groupi_n_10710 ,csa_tree_add_190_195_groupi_n_10470 ,csa_tree_add_190_195_groupi_n_10489);
  or csa_tree_add_190_195_groupi_g38224(csa_tree_add_190_195_groupi_n_10709 ,csa_tree_add_190_195_groupi_n_10454 ,csa_tree_add_190_195_groupi_n_10556);
  or csa_tree_add_190_195_groupi_g38225(csa_tree_add_190_195_groupi_n_10708 ,csa_tree_add_190_195_groupi_n_10285 ,csa_tree_add_190_195_groupi_n_10472);
  nor csa_tree_add_190_195_groupi_g38226(csa_tree_add_190_195_groupi_n_10707 ,csa_tree_add_190_195_groupi_n_10453 ,csa_tree_add_190_195_groupi_n_10557);
  or csa_tree_add_190_195_groupi_g38227(csa_tree_add_190_195_groupi_n_10706 ,csa_tree_add_190_195_groupi_n_10484 ,csa_tree_add_190_195_groupi_n_10354);
  nor csa_tree_add_190_195_groupi_g38228(csa_tree_add_190_195_groupi_n_10705 ,csa_tree_add_190_195_groupi_n_10152 ,csa_tree_add_190_195_groupi_n_10566);
  and csa_tree_add_190_195_groupi_g38229(csa_tree_add_190_195_groupi_n_10802 ,csa_tree_add_190_195_groupi_n_10264 ,csa_tree_add_190_195_groupi_n_10522);
  and csa_tree_add_190_195_groupi_g38230(csa_tree_add_190_195_groupi_n_10801 ,csa_tree_add_190_195_groupi_n_10256 ,csa_tree_add_190_195_groupi_n_10496);
  or csa_tree_add_190_195_groupi_g38231(csa_tree_add_190_195_groupi_n_10800 ,csa_tree_add_190_195_groupi_n_10260 ,csa_tree_add_190_195_groupi_n_10503);
  or csa_tree_add_190_195_groupi_g38232(csa_tree_add_190_195_groupi_n_10799 ,csa_tree_add_190_195_groupi_n_10238 ,csa_tree_add_190_195_groupi_n_10505);
  and csa_tree_add_190_195_groupi_g38233(csa_tree_add_190_195_groupi_n_10798 ,csa_tree_add_190_195_groupi_n_10128 ,csa_tree_add_190_195_groupi_n_10508);
  and csa_tree_add_190_195_groupi_g38234(csa_tree_add_190_195_groupi_n_10797 ,csa_tree_add_190_195_groupi_n_10243 ,csa_tree_add_190_195_groupi_n_10509);
  and csa_tree_add_190_195_groupi_g38235(csa_tree_add_190_195_groupi_n_10796 ,csa_tree_add_190_195_groupi_n_10296 ,csa_tree_add_190_195_groupi_n_10483);
  or csa_tree_add_190_195_groupi_g38236(csa_tree_add_190_195_groupi_n_10795 ,csa_tree_add_190_195_groupi_n_10245 ,csa_tree_add_190_195_groupi_n_10542);
  and csa_tree_add_190_195_groupi_g38237(csa_tree_add_190_195_groupi_n_10794 ,csa_tree_add_190_195_groupi_n_10249 ,csa_tree_add_190_195_groupi_n_10515);
  and csa_tree_add_190_195_groupi_g38238(csa_tree_add_190_195_groupi_n_10793 ,csa_tree_add_190_195_groupi_n_10302 ,csa_tree_add_190_195_groupi_n_10507);
  or csa_tree_add_190_195_groupi_g38239(csa_tree_add_190_195_groupi_n_10791 ,csa_tree_add_190_195_groupi_n_10253 ,csa_tree_add_190_195_groupi_n_10547);
  or csa_tree_add_190_195_groupi_g38240(csa_tree_add_190_195_groupi_n_10789 ,csa_tree_add_190_195_groupi_n_9844 ,csa_tree_add_190_195_groupi_n_10498);
  and csa_tree_add_190_195_groupi_g38241(csa_tree_add_190_195_groupi_n_10788 ,csa_tree_add_190_195_groupi_n_9848 ,csa_tree_add_190_195_groupi_n_10516);
  or csa_tree_add_190_195_groupi_g38242(csa_tree_add_190_195_groupi_n_10787 ,csa_tree_add_190_195_groupi_n_10234 ,csa_tree_add_190_195_groupi_n_10517);
  or csa_tree_add_190_195_groupi_g38243(csa_tree_add_190_195_groupi_n_10786 ,csa_tree_add_190_195_groupi_n_10126 ,csa_tree_add_190_195_groupi_n_10518);
  and csa_tree_add_190_195_groupi_g38244(csa_tree_add_190_195_groupi_n_10785 ,csa_tree_add_190_195_groupi_n_10004 ,csa_tree_add_190_195_groupi_n_10519);
  and csa_tree_add_190_195_groupi_g38245(csa_tree_add_190_195_groupi_n_10784 ,csa_tree_add_190_195_groupi_n_10255 ,csa_tree_add_190_195_groupi_n_10541);
  and csa_tree_add_190_195_groupi_g38246(csa_tree_add_190_195_groupi_n_10783 ,csa_tree_add_190_195_groupi_n_10270 ,csa_tree_add_190_195_groupi_n_10527);
  or csa_tree_add_190_195_groupi_g38247(csa_tree_add_190_195_groupi_n_10782 ,csa_tree_add_190_195_groupi_n_10286 ,csa_tree_add_190_195_groupi_n_10548);
  and csa_tree_add_190_195_groupi_g38248(csa_tree_add_190_195_groupi_n_10781 ,csa_tree_add_190_195_groupi_n_10012 ,csa_tree_add_190_195_groupi_n_10532);
  and csa_tree_add_190_195_groupi_g38249(csa_tree_add_190_195_groupi_n_10780 ,csa_tree_add_190_195_groupi_n_9096 ,csa_tree_add_190_195_groupi_n_10528);
  and csa_tree_add_190_195_groupi_g38250(csa_tree_add_190_195_groupi_n_10779 ,csa_tree_add_190_195_groupi_n_10259 ,csa_tree_add_190_195_groupi_n_10543);
  and csa_tree_add_190_195_groupi_g38251(csa_tree_add_190_195_groupi_n_10778 ,csa_tree_add_190_195_groupi_n_10142 ,csa_tree_add_190_195_groupi_n_10546);
  and csa_tree_add_190_195_groupi_g38252(csa_tree_add_190_195_groupi_n_10777 ,csa_tree_add_190_195_groupi_n_9587 ,csa_tree_add_190_195_groupi_n_10529);
  or csa_tree_add_190_195_groupi_g38253(csa_tree_add_190_195_groupi_n_10775 ,csa_tree_add_190_195_groupi_n_10281 ,csa_tree_add_190_195_groupi_n_10533);
  and csa_tree_add_190_195_groupi_g38254(csa_tree_add_190_195_groupi_n_10774 ,csa_tree_add_190_195_groupi_n_10282 ,csa_tree_add_190_195_groupi_n_10531);
  or csa_tree_add_190_195_groupi_g38255(csa_tree_add_190_195_groupi_n_10773 ,csa_tree_add_190_195_groupi_n_10114 ,csa_tree_add_190_195_groupi_n_10534);
  or csa_tree_add_190_195_groupi_g38256(csa_tree_add_190_195_groupi_n_10772 ,csa_tree_add_190_195_groupi_n_10289 ,csa_tree_add_190_195_groupi_n_10537);
  and csa_tree_add_190_195_groupi_g38257(csa_tree_add_190_195_groupi_n_10771 ,csa_tree_add_190_195_groupi_n_10293 ,csa_tree_add_190_195_groupi_n_10540);
  and csa_tree_add_190_195_groupi_g38258(csa_tree_add_190_195_groupi_n_10769 ,csa_tree_add_190_195_groupi_n_10303 ,csa_tree_add_190_195_groupi_n_10545);
  or csa_tree_add_190_195_groupi_g38259(csa_tree_add_190_195_groupi_n_10767 ,csa_tree_add_190_195_groupi_n_10307 ,csa_tree_add_190_195_groupi_n_10530);
  and csa_tree_add_190_195_groupi_g38260(csa_tree_add_190_195_groupi_n_10766 ,csa_tree_add_190_195_groupi_n_10274 ,csa_tree_add_190_195_groupi_n_10523);
  and csa_tree_add_190_195_groupi_g38261(csa_tree_add_190_195_groupi_n_10764 ,csa_tree_add_190_195_groupi_n_10247 ,csa_tree_add_190_195_groupi_n_10510);
  not csa_tree_add_190_195_groupi_g38262(csa_tree_add_190_195_groupi_n_10701 ,csa_tree_add_190_195_groupi_n_10700);
  not csa_tree_add_190_195_groupi_g38265(csa_tree_add_190_195_groupi_n_10695 ,csa_tree_add_190_195_groupi_n_10694);
  not csa_tree_add_190_195_groupi_g38266(csa_tree_add_190_195_groupi_n_10693 ,csa_tree_add_190_195_groupi_n_10692);
  not csa_tree_add_190_195_groupi_g38267(csa_tree_add_190_195_groupi_n_10691 ,csa_tree_add_190_195_groupi_n_10690);
  not csa_tree_add_190_195_groupi_g38268(csa_tree_add_190_195_groupi_n_10689 ,csa_tree_add_190_195_groupi_n_10688);
  not csa_tree_add_190_195_groupi_g38269(csa_tree_add_190_195_groupi_n_10687 ,csa_tree_add_190_195_groupi_n_10686);
  not csa_tree_add_190_195_groupi_g38270(csa_tree_add_190_195_groupi_n_10685 ,csa_tree_add_190_195_groupi_n_10684);
  not csa_tree_add_190_195_groupi_g38271(csa_tree_add_190_195_groupi_n_10683 ,csa_tree_add_190_195_groupi_n_10682);
  not csa_tree_add_190_195_groupi_g38272(csa_tree_add_190_195_groupi_n_10681 ,csa_tree_add_190_195_groupi_n_10680);
  not csa_tree_add_190_195_groupi_g38273(csa_tree_add_190_195_groupi_n_10679 ,csa_tree_add_190_195_groupi_n_10678);
  not csa_tree_add_190_195_groupi_g38274(csa_tree_add_190_195_groupi_n_10677 ,csa_tree_add_190_195_groupi_n_10676);
  not csa_tree_add_190_195_groupi_g38275(csa_tree_add_190_195_groupi_n_10675 ,csa_tree_add_190_195_groupi_n_10674);
  not csa_tree_add_190_195_groupi_g38276(csa_tree_add_190_195_groupi_n_10673 ,csa_tree_add_190_195_groupi_n_10672);
  not csa_tree_add_190_195_groupi_g38277(csa_tree_add_190_195_groupi_n_10671 ,csa_tree_add_190_195_groupi_n_10670);
  not csa_tree_add_190_195_groupi_g38278(csa_tree_add_190_195_groupi_n_10669 ,csa_tree_add_190_195_groupi_n_10668);
  not csa_tree_add_190_195_groupi_g38279(csa_tree_add_190_195_groupi_n_10667 ,csa_tree_add_190_195_groupi_n_135);
  not csa_tree_add_190_195_groupi_g38280(csa_tree_add_190_195_groupi_n_10666 ,csa_tree_add_190_195_groupi_n_10665);
  not csa_tree_add_190_195_groupi_g38281(csa_tree_add_190_195_groupi_n_10664 ,csa_tree_add_190_195_groupi_n_10663);
  not csa_tree_add_190_195_groupi_g38282(csa_tree_add_190_195_groupi_n_10662 ,csa_tree_add_190_195_groupi_n_10661);
  not csa_tree_add_190_195_groupi_g38283(csa_tree_add_190_195_groupi_n_10660 ,csa_tree_add_190_195_groupi_n_10659);
  not csa_tree_add_190_195_groupi_g38284(csa_tree_add_190_195_groupi_n_10657 ,csa_tree_add_190_195_groupi_n_10658);
  not csa_tree_add_190_195_groupi_g38285(csa_tree_add_190_195_groupi_n_10655 ,csa_tree_add_190_195_groupi_n_10654);
  not csa_tree_add_190_195_groupi_g38286(csa_tree_add_190_195_groupi_n_10653 ,csa_tree_add_190_195_groupi_n_10652);
  not csa_tree_add_190_195_groupi_g38287(csa_tree_add_190_195_groupi_n_10651 ,csa_tree_add_190_195_groupi_n_10650);
  not csa_tree_add_190_195_groupi_g38288(csa_tree_add_190_195_groupi_n_10649 ,csa_tree_add_190_195_groupi_n_10648);
  not csa_tree_add_190_195_groupi_g38289(csa_tree_add_190_195_groupi_n_10646 ,csa_tree_add_190_195_groupi_n_10647);
  not csa_tree_add_190_195_groupi_g38290(csa_tree_add_190_195_groupi_n_10645 ,csa_tree_add_190_195_groupi_n_10644);
  or csa_tree_add_190_195_groupi_g38291(csa_tree_add_190_195_groupi_n_10643 ,csa_tree_add_190_195_groupi_n_10231 ,csa_tree_add_190_195_groupi_n_10410);
  or csa_tree_add_190_195_groupi_g38292(csa_tree_add_190_195_groupi_n_10642 ,csa_tree_add_190_195_groupi_n_10201 ,csa_tree_add_190_195_groupi_n_10464);
  nor csa_tree_add_190_195_groupi_g38293(csa_tree_add_190_195_groupi_n_10641 ,csa_tree_add_190_195_groupi_n_10202 ,csa_tree_add_190_195_groupi_n_10465);
  or csa_tree_add_190_195_groupi_g38294(csa_tree_add_190_195_groupi_n_10640 ,csa_tree_add_190_195_groupi_n_10455 ,csa_tree_add_190_195_groupi_n_10189);
  nor csa_tree_add_190_195_groupi_g38295(csa_tree_add_190_195_groupi_n_10639 ,csa_tree_add_190_195_groupi_n_143 ,csa_tree_add_190_195_groupi_n_10190);
  nor csa_tree_add_190_195_groupi_g38296(csa_tree_add_190_195_groupi_n_10638 ,csa_tree_add_190_195_groupi_n_10186 ,csa_tree_add_190_195_groupi_n_10451);
  and csa_tree_add_190_195_groupi_g38297(csa_tree_add_190_195_groupi_n_10637 ,csa_tree_add_190_195_groupi_n_10467 ,csa_tree_add_190_195_groupi_n_10413);
  or csa_tree_add_190_195_groupi_g38298(csa_tree_add_190_195_groupi_n_10636 ,csa_tree_add_190_195_groupi_n_10185 ,csa_tree_add_190_195_groupi_n_10452);
  or csa_tree_add_190_195_groupi_g38299(csa_tree_add_190_195_groupi_n_10635 ,csa_tree_add_190_195_groupi_n_10047 ,csa_tree_add_190_195_groupi_n_10443);
  or csa_tree_add_190_195_groupi_g38300(csa_tree_add_190_195_groupi_n_10634 ,csa_tree_add_190_195_groupi_n_10474 ,csa_tree_add_190_195_groupi_n_10407);
  nor csa_tree_add_190_195_groupi_g38301(csa_tree_add_190_195_groupi_n_10633 ,csa_tree_add_190_195_groupi_n_10172 ,csa_tree_add_190_195_groupi_n_10438);
  or csa_tree_add_190_195_groupi_g38302(csa_tree_add_190_195_groupi_n_10632 ,csa_tree_add_190_195_groupi_n_10171 ,csa_tree_add_190_195_groupi_n_10439);
  and csa_tree_add_190_195_groupi_g38303(csa_tree_add_190_195_groupi_n_10631 ,csa_tree_add_190_195_groupi_n_10047 ,csa_tree_add_190_195_groupi_n_10443);
  nor csa_tree_add_190_195_groupi_g38304(csa_tree_add_190_195_groupi_n_10630 ,csa_tree_add_190_195_groupi_n_10437 ,csa_tree_add_190_195_groupi_n_10434);
  or csa_tree_add_190_195_groupi_g38305(csa_tree_add_190_195_groupi_n_10629 ,csa_tree_add_190_195_groupi_n_10436 ,csa_tree_add_190_195_groupi_n_10435);
  or csa_tree_add_190_195_groupi_g38306(csa_tree_add_190_195_groupi_n_10628 ,csa_tree_add_190_195_groupi_n_10429 ,csa_tree_add_190_195_groupi_n_10160);
  or csa_tree_add_190_195_groupi_g38307(csa_tree_add_190_195_groupi_n_10627 ,csa_tree_add_190_195_groupi_n_9661 ,csa_tree_add_190_195_groupi_n_10404);
  nor csa_tree_add_190_195_groupi_g38308(csa_tree_add_190_195_groupi_n_10626 ,csa_tree_add_190_195_groupi_n_10428 ,csa_tree_add_190_195_groupi_n_10161);
  or csa_tree_add_190_195_groupi_g38309(csa_tree_add_190_195_groupi_n_10625 ,csa_tree_add_190_195_groupi_n_9637 ,csa_tree_add_190_195_groupi_n_10568);
  xnor csa_tree_add_190_195_groupi_g38310(csa_tree_add_190_195_groupi_n_10624 ,csa_tree_add_190_195_groupi_n_10151 ,csa_tree_add_190_195_groupi_n_10149);
  xnor csa_tree_add_190_195_groupi_g38311(csa_tree_add_190_195_groupi_n_10623 ,csa_tree_add_190_195_groupi_n_10039 ,csa_tree_add_190_195_groupi_n_10226);
  xnor csa_tree_add_190_195_groupi_g38312(csa_tree_add_190_195_groupi_n_10622 ,csa_tree_add_190_195_groupi_n_9878 ,csa_tree_add_190_195_groupi_n_10192);
  xnor csa_tree_add_190_195_groupi_g38313(csa_tree_add_190_195_groupi_n_10621 ,csa_tree_add_190_195_groupi_n_9880 ,csa_tree_add_190_195_groupi_n_10334);
  xnor csa_tree_add_190_195_groupi_g38315(csa_tree_add_190_195_groupi_n_10620 ,csa_tree_add_190_195_groupi_n_9771 ,csa_tree_add_190_195_groupi_n_10170);
  xnor csa_tree_add_190_195_groupi_g38316(csa_tree_add_190_195_groupi_n_10619 ,csa_tree_add_190_195_groupi_n_10184 ,csa_tree_add_190_195_groupi_n_10355);
  xnor csa_tree_add_190_195_groupi_g38317(csa_tree_add_190_195_groupi_n_10618 ,csa_tree_add_190_195_groupi_n_9888 ,csa_tree_add_190_195_groupi_n_10178);
  xnor csa_tree_add_190_195_groupi_g38318(csa_tree_add_190_195_groupi_n_10617 ,csa_tree_add_190_195_groupi_n_7619 ,csa_tree_add_190_195_groupi_n_10218);
  xnor csa_tree_add_190_195_groupi_g38319(csa_tree_add_190_195_groupi_n_10616 ,csa_tree_add_190_195_groupi_n_10332 ,csa_tree_add_190_195_groupi_n_8630);
  xnor csa_tree_add_190_195_groupi_g38320(csa_tree_add_190_195_groupi_n_10615 ,csa_tree_add_190_195_groupi_n_9471 ,csa_tree_add_190_195_groupi_n_10219);
  xnor csa_tree_add_190_195_groupi_g38322(csa_tree_add_190_195_groupi_n_10614 ,csa_tree_add_190_195_groupi_n_10349 ,csa_tree_add_190_195_groupi_n_10154);
  xnor csa_tree_add_190_195_groupi_g38324(csa_tree_add_190_195_groupi_n_10613 ,csa_tree_add_190_195_groupi_n_9766 ,csa_tree_add_190_195_groupi_n_10174);
  xnor csa_tree_add_190_195_groupi_g38325(csa_tree_add_190_195_groupi_n_10612 ,csa_tree_add_190_195_groupi_n_10348 ,csa_tree_add_190_195_groupi_n_10058);
  xnor csa_tree_add_190_195_groupi_g38326(csa_tree_add_190_195_groupi_n_10611 ,csa_tree_add_190_195_groupi_n_10188 ,csa_tree_add_190_195_groupi_n_9899);
  xnor csa_tree_add_190_195_groupi_g38327(csa_tree_add_190_195_groupi_n_10610 ,csa_tree_add_190_195_groupi_n_10056 ,csa_tree_add_190_195_groupi_n_10194);
  xnor csa_tree_add_190_195_groupi_g38328(csa_tree_add_190_195_groupi_n_10609 ,csa_tree_add_190_195_groupi_n_9799 ,csa_tree_add_190_195_groupi_n_10217);
  xnor csa_tree_add_190_195_groupi_g38329(csa_tree_add_190_195_groupi_n_10608 ,csa_tree_add_190_195_groupi_n_10176 ,csa_tree_add_190_195_groupi_n_9945);
  xnor csa_tree_add_190_195_groupi_g38330(csa_tree_add_190_195_groupi_n_10607 ,csa_tree_add_190_195_groupi_n_10337 ,csa_tree_add_190_195_groupi_n_9928);
  xnor csa_tree_add_190_195_groupi_g38331(csa_tree_add_190_195_groupi_n_10606 ,csa_tree_add_190_195_groupi_n_9288 ,csa_tree_add_190_195_groupi_n_10335);
  xnor csa_tree_add_190_195_groupi_g38332(csa_tree_add_190_195_groupi_n_10605 ,csa_tree_add_190_195_groupi_n_10340 ,csa_tree_add_190_195_groupi_n_10200);
  xnor csa_tree_add_190_195_groupi_g38333(csa_tree_add_190_195_groupi_n_10604 ,csa_tree_add_190_195_groupi_n_10347 ,csa_tree_add_190_195_groupi_n_10202);
  xnor csa_tree_add_190_195_groupi_g38334(csa_tree_add_190_195_groupi_n_10603 ,csa_tree_add_190_195_groupi_n_10035 ,csa_tree_add_190_195_groupi_n_10225);
  xnor csa_tree_add_190_195_groupi_g38336(csa_tree_add_190_195_groupi_n_10602 ,csa_tree_add_190_195_groupi_n_10317 ,csa_tree_add_190_195_groupi_n_10230);
  xnor csa_tree_add_190_195_groupi_g38338(csa_tree_add_190_195_groupi_n_10601 ,csa_tree_add_190_195_groupi_n_10313 ,csa_tree_add_190_195_groupi_n_10354);
  xnor csa_tree_add_190_195_groupi_g38339(csa_tree_add_190_195_groupi_n_10600 ,csa_tree_add_190_195_groupi_n_8691 ,csa_tree_add_190_195_groupi_n_10322);
  xnor csa_tree_add_190_195_groupi_g38340(csa_tree_add_190_195_groupi_n_10599 ,csa_tree_add_190_195_groupi_n_9630 ,csa_tree_add_190_195_groupi_n_10147);
  xnor csa_tree_add_190_195_groupi_g38341(csa_tree_add_190_195_groupi_n_10598 ,csa_tree_add_190_195_groupi_n_10345 ,csa_tree_add_190_195_groupi_n_9939);
  xnor csa_tree_add_190_195_groupi_g38342(csa_tree_add_190_195_groupi_n_10597 ,csa_tree_add_190_195_groupi_n_9770 ,csa_tree_add_190_195_groupi_n_10333);
  xnor csa_tree_add_190_195_groupi_g38343(csa_tree_add_190_195_groupi_n_10596 ,csa_tree_add_190_195_groupi_n_9662 ,csa_tree_add_190_195_groupi_n_10324);
  xnor csa_tree_add_190_195_groupi_g38344(csa_tree_add_190_195_groupi_n_10595 ,csa_tree_add_190_195_groupi_n_9632 ,csa_tree_add_190_195_groupi_n_10159);
  xnor csa_tree_add_190_195_groupi_g38345(csa_tree_add_190_195_groupi_n_10594 ,csa_tree_add_190_195_groupi_n_9862 ,csa_tree_add_190_195_groupi_n_10182);
  xnor csa_tree_add_190_195_groupi_g38346(csa_tree_add_190_195_groupi_n_10593 ,csa_tree_add_190_195_groupi_n_10319 ,csa_tree_add_190_195_groupi_n_9868);
  xnor csa_tree_add_190_195_groupi_g38347(csa_tree_add_190_195_groupi_n_10592 ,csa_tree_add_190_195_groupi_n_9475 ,csa_tree_add_190_195_groupi_n_10163);
  and csa_tree_add_190_195_groupi_g38348(csa_tree_add_190_195_groupi_n_10704 ,csa_tree_add_190_195_groupi_n_10132 ,csa_tree_add_190_195_groupi_n_10416);
  or csa_tree_add_190_195_groupi_g38349(csa_tree_add_190_195_groupi_n_10703 ,csa_tree_add_190_195_groupi_n_10138 ,csa_tree_add_190_195_groupi_n_10396);
  xnor csa_tree_add_190_195_groupi_g38350(csa_tree_add_190_195_groupi_n_10702 ,csa_tree_add_190_195_groupi_n_8321 ,csa_tree_add_190_195_groupi_n_10090);
  xnor csa_tree_add_190_195_groupi_g38351(csa_tree_add_190_195_groupi_n_10700 ,csa_tree_add_190_195_groupi_n_10066 ,csa_tree_add_190_195_groupi_n_10109);
  xnor csa_tree_add_190_195_groupi_g38352(csa_tree_add_190_195_groupi_n_10699 ,csa_tree_add_190_195_groupi_n_10079 ,csa_tree_add_190_195_groupi_n_10111);
  xnor csa_tree_add_190_195_groupi_g38353(csa_tree_add_190_195_groupi_n_10698 ,csa_tree_add_190_195_groupi_n_9186 ,csa_tree_add_190_195_groupi_n_10113);
  and csa_tree_add_190_195_groupi_g38354(csa_tree_add_190_195_groupi_n_10697 ,csa_tree_add_190_195_groupi_n_10120 ,csa_tree_add_190_195_groupi_n_10398);
  and csa_tree_add_190_195_groupi_g38355(csa_tree_add_190_195_groupi_n_10696 ,csa_tree_add_190_195_groupi_n_10125 ,csa_tree_add_190_195_groupi_n_10401);
  xnor csa_tree_add_190_195_groupi_g38356(csa_tree_add_190_195_groupi_n_10694 ,csa_tree_add_190_195_groupi_n_9348 ,csa_tree_add_190_195_groupi_n_10096);
  xnor csa_tree_add_190_195_groupi_g38357(csa_tree_add_190_195_groupi_n_10692 ,csa_tree_add_190_195_groupi_n_9030 ,csa_tree_add_190_195_groupi_n_10100);
  xnor csa_tree_add_190_195_groupi_g38358(csa_tree_add_190_195_groupi_n_10690 ,csa_tree_add_190_195_groupi_n_8020 ,csa_tree_add_190_195_groupi_n_10091);
  xnor csa_tree_add_190_195_groupi_g38359(csa_tree_add_190_195_groupi_n_10688 ,csa_tree_add_190_195_groupi_n_9511 ,csa_tree_add_190_195_groupi_n_10095);
  xnor csa_tree_add_190_195_groupi_g38360(csa_tree_add_190_195_groupi_n_10686 ,csa_tree_add_190_195_groupi_n_9498 ,csa_tree_add_190_195_groupi_n_10089);
  xnor csa_tree_add_190_195_groupi_g38361(csa_tree_add_190_195_groupi_n_10684 ,csa_tree_add_190_195_groupi_n_9344 ,csa_tree_add_190_195_groupi_n_132);
  xnor csa_tree_add_190_195_groupi_g38362(csa_tree_add_190_195_groupi_n_10682 ,csa_tree_add_190_195_groupi_n_7354 ,csa_tree_add_190_195_groupi_n_10088);
  xnor csa_tree_add_190_195_groupi_g38363(csa_tree_add_190_195_groupi_n_10680 ,csa_tree_add_190_195_groupi_n_9482 ,csa_tree_add_190_195_groupi_n_10104);
  xnor csa_tree_add_190_195_groupi_g38364(csa_tree_add_190_195_groupi_n_10678 ,csa_tree_add_190_195_groupi_n_9035 ,csa_tree_add_190_195_groupi_n_10099);
  xnor csa_tree_add_190_195_groupi_g38365(csa_tree_add_190_195_groupi_n_10676 ,csa_tree_add_190_195_groupi_n_10220 ,csa_tree_add_190_195_groupi_n_9821);
  xnor csa_tree_add_190_195_groupi_g38366(csa_tree_add_190_195_groupi_n_10674 ,csa_tree_add_190_195_groupi_n_9796 ,csa_tree_add_190_195_groupi_n_10110);
  xnor csa_tree_add_190_195_groupi_g38367(csa_tree_add_190_195_groupi_n_10672 ,csa_tree_add_190_195_groupi_n_9480 ,csa_tree_add_190_195_groupi_n_10103);
  xnor csa_tree_add_190_195_groupi_g38368(csa_tree_add_190_195_groupi_n_10670 ,csa_tree_add_190_195_groupi_n_9318 ,csa_tree_add_190_195_groupi_n_10106);
  xnor csa_tree_add_190_195_groupi_g38369(csa_tree_add_190_195_groupi_n_10668 ,csa_tree_add_190_195_groupi_n_10087 ,csa_tree_add_190_195_groupi_n_10108);
  and csa_tree_add_190_195_groupi_g38371(csa_tree_add_190_195_groupi_n_10665 ,csa_tree_add_190_195_groupi_n_10135 ,csa_tree_add_190_195_groupi_n_10417);
  xnor csa_tree_add_190_195_groupi_g38372(csa_tree_add_190_195_groupi_n_10663 ,csa_tree_add_190_195_groupi_n_9790 ,csa_tree_add_190_195_groupi_n_10093);
  xnor csa_tree_add_190_195_groupi_g38373(csa_tree_add_190_195_groupi_n_10661 ,csa_tree_add_190_195_groupi_n_9311 ,csa_tree_add_190_195_groupi_n_10097);
  xnor csa_tree_add_190_195_groupi_g38374(csa_tree_add_190_195_groupi_n_10659 ,csa_tree_add_190_195_groupi_n_10232 ,csa_tree_add_190_195_groupi_n_10098);
  and csa_tree_add_190_195_groupi_g38375(csa_tree_add_190_195_groupi_n_10658 ,csa_tree_add_190_195_groupi_n_10123 ,csa_tree_add_190_195_groupi_n_10402);
  xnor csa_tree_add_190_195_groupi_g38376(csa_tree_add_190_195_groupi_n_10656 ,csa_tree_add_190_195_groupi_n_9793 ,csa_tree_add_190_195_groupi_n_10101);
  xnor csa_tree_add_190_195_groupi_g38377(csa_tree_add_190_195_groupi_n_10654 ,csa_tree_add_190_195_groupi_n_9920 ,csa_tree_add_190_195_groupi_n_10092);
  xnor csa_tree_add_190_195_groupi_g38378(csa_tree_add_190_195_groupi_n_10652 ,csa_tree_add_190_195_groupi_n_8027 ,csa_tree_add_190_195_groupi_n_133);
  and csa_tree_add_190_195_groupi_g38379(csa_tree_add_190_195_groupi_n_10650 ,csa_tree_add_190_195_groupi_n_10134 ,csa_tree_add_190_195_groupi_n_10418);
  xnor csa_tree_add_190_195_groupi_g38380(csa_tree_add_190_195_groupi_n_10648 ,csa_tree_add_190_195_groupi_n_7112 ,csa_tree_add_190_195_groupi_n_10102);
  xnor csa_tree_add_190_195_groupi_g38381(csa_tree_add_190_195_groupi_n_10647 ,csa_tree_add_190_195_groupi_n_9356 ,csa_tree_add_190_195_groupi_n_10112);
  xnor csa_tree_add_190_195_groupi_g38382(csa_tree_add_190_195_groupi_n_10644 ,csa_tree_add_190_195_groupi_n_7545 ,csa_tree_add_190_195_groupi_n_10094);
  not csa_tree_add_190_195_groupi_g38383(csa_tree_add_190_195_groupi_n_10580 ,csa_tree_add_190_195_groupi_n_10579);
  not csa_tree_add_190_195_groupi_g38385(csa_tree_add_190_195_groupi_n_10575 ,csa_tree_add_190_195_groupi_n_10576);
  not csa_tree_add_190_195_groupi_g38386(csa_tree_add_190_195_groupi_n_10573 ,csa_tree_add_190_195_groupi_n_10574);
  not csa_tree_add_190_195_groupi_g38387(csa_tree_add_190_195_groupi_n_10572 ,csa_tree_add_190_195_groupi_n_10571);
  not csa_tree_add_190_195_groupi_g38388(csa_tree_add_190_195_groupi_n_10569 ,csa_tree_add_190_195_groupi_n_10570);
  not csa_tree_add_190_195_groupi_g38389(csa_tree_add_190_195_groupi_n_10568 ,csa_tree_add_190_195_groupi_n_10567);
  not csa_tree_add_190_195_groupi_g38390(csa_tree_add_190_195_groupi_n_10566 ,csa_tree_add_190_195_groupi_n_10565);
  not csa_tree_add_190_195_groupi_g38391(csa_tree_add_190_195_groupi_n_10564 ,csa_tree_add_190_195_groupi_n_10563);
  not csa_tree_add_190_195_groupi_g38392(csa_tree_add_190_195_groupi_n_10560 ,csa_tree_add_190_195_groupi_n_10561);
  not csa_tree_add_190_195_groupi_g38393(csa_tree_add_190_195_groupi_n_10558 ,csa_tree_add_190_195_groupi_n_10559);
  not csa_tree_add_190_195_groupi_g38394(csa_tree_add_190_195_groupi_n_10557 ,csa_tree_add_190_195_groupi_n_10556);
  not csa_tree_add_190_195_groupi_g38395(csa_tree_add_190_195_groupi_n_10555 ,csa_tree_add_190_195_groupi_n_10554);
  not csa_tree_add_190_195_groupi_g38396(csa_tree_add_190_195_groupi_n_10553 ,csa_tree_add_190_195_groupi_n_10552);
  not csa_tree_add_190_195_groupi_g38397(csa_tree_add_190_195_groupi_n_10550 ,csa_tree_add_190_195_groupi_n_10551);
  nor csa_tree_add_190_195_groupi_g38398(csa_tree_add_190_195_groupi_n_10549 ,csa_tree_add_190_195_groupi_n_10331 ,csa_tree_add_190_195_groupi_n_8630);
  and csa_tree_add_190_195_groupi_g38399(csa_tree_add_190_195_groupi_n_10548 ,csa_tree_add_190_195_groupi_n_9962 ,csa_tree_add_190_195_groupi_n_10139);
  and csa_tree_add_190_195_groupi_g38400(csa_tree_add_190_195_groupi_n_10547 ,csa_tree_add_190_195_groupi_n_10309 ,csa_tree_add_190_195_groupi_n_10225);
  or csa_tree_add_190_195_groupi_g38401(csa_tree_add_190_195_groupi_n_10546 ,csa_tree_add_190_195_groupi_n_10073 ,csa_tree_add_190_195_groupi_n_10141);
  or csa_tree_add_190_195_groupi_g38402(csa_tree_add_190_195_groupi_n_10545 ,csa_tree_add_190_195_groupi_n_10337 ,csa_tree_add_190_195_groupi_n_10301);
  nor csa_tree_add_190_195_groupi_g38403(csa_tree_add_190_195_groupi_n_10544 ,csa_tree_add_190_195_groupi_n_10175 ,csa_tree_add_190_195_groupi_n_9945);
  or csa_tree_add_190_195_groupi_g38404(csa_tree_add_190_195_groupi_n_10543 ,csa_tree_add_190_195_groupi_n_9807 ,csa_tree_add_190_195_groupi_n_10271);
  and csa_tree_add_190_195_groupi_g38405(csa_tree_add_190_195_groupi_n_10542 ,csa_tree_add_190_195_groupi_n_10338 ,csa_tree_add_190_195_groupi_n_10244);
  or csa_tree_add_190_195_groupi_g38406(csa_tree_add_190_195_groupi_n_10541 ,csa_tree_add_190_195_groupi_n_10339 ,csa_tree_add_190_195_groupi_n_10283);
  or csa_tree_add_190_195_groupi_g38407(csa_tree_add_190_195_groupi_n_10540 ,csa_tree_add_190_195_groupi_n_10353 ,csa_tree_add_190_195_groupi_n_10292);
  nor csa_tree_add_190_195_groupi_g38408(csa_tree_add_190_195_groupi_n_10539 ,csa_tree_add_190_195_groupi_n_10150 ,csa_tree_add_190_195_groupi_n_10149);
  or csa_tree_add_190_195_groupi_g38409(csa_tree_add_190_195_groupi_n_10538 ,csa_tree_add_190_195_groupi_n_10151 ,csa_tree_add_190_195_groupi_n_10148);
  and csa_tree_add_190_195_groupi_g38410(csa_tree_add_190_195_groupi_n_10537 ,csa_tree_add_190_195_groupi_n_9798 ,csa_tree_add_190_195_groupi_n_10287);
  nor csa_tree_add_190_195_groupi_g38411(csa_tree_add_190_195_groupi_n_10536 ,csa_tree_add_190_195_groupi_n_9631 ,csa_tree_add_190_195_groupi_n_10159);
  or csa_tree_add_190_195_groupi_g38412(csa_tree_add_190_195_groupi_n_10535 ,csa_tree_add_190_195_groupi_n_9632 ,csa_tree_add_190_195_groupi_n_10158);
  and csa_tree_add_190_195_groupi_g38413(csa_tree_add_190_195_groupi_n_10534 ,csa_tree_add_190_195_groupi_n_10345 ,csa_tree_add_190_195_groupi_n_10129);
  nor csa_tree_add_190_195_groupi_g38414(csa_tree_add_190_195_groupi_n_10533 ,csa_tree_add_190_195_groupi_n_9800 ,csa_tree_add_190_195_groupi_n_10278);
  or csa_tree_add_190_195_groupi_g38415(csa_tree_add_190_195_groupi_n_10532 ,csa_tree_add_190_195_groupi_n_10015 ,csa_tree_add_190_195_groupi_n_10232);
  or csa_tree_add_190_195_groupi_g38416(csa_tree_add_190_195_groupi_n_10531 ,csa_tree_add_190_195_groupi_n_9955 ,csa_tree_add_190_195_groupi_n_10273);
  nor csa_tree_add_190_195_groupi_g38417(csa_tree_add_190_195_groupi_n_10530 ,csa_tree_add_190_195_groupi_n_10071 ,csa_tree_add_190_195_groupi_n_10311);
  or csa_tree_add_190_195_groupi_g38418(csa_tree_add_190_195_groupi_n_10529 ,csa_tree_add_190_195_groupi_n_9598 ,csa_tree_add_190_195_groupi_n_10220);
  or csa_tree_add_190_195_groupi_g38419(csa_tree_add_190_195_groupi_n_10528 ,csa_tree_add_190_195_groupi_n_9095 ,csa_tree_add_190_195_groupi_n_10218);
  or csa_tree_add_190_195_groupi_g38420(csa_tree_add_190_195_groupi_n_10527 ,csa_tree_add_190_195_groupi_n_9658 ,csa_tree_add_190_195_groupi_n_10269);
  or csa_tree_add_190_195_groupi_g38421(csa_tree_add_190_195_groupi_n_10526 ,csa_tree_add_190_195_groupi_n_9764 ,csa_tree_add_190_195_groupi_n_10314);
  or csa_tree_add_190_195_groupi_g38422(csa_tree_add_190_195_groupi_n_10525 ,csa_tree_add_190_195_groupi_n_10176 ,csa_tree_add_190_195_groupi_n_9944);
  and csa_tree_add_190_195_groupi_g38423(csa_tree_add_190_195_groupi_n_10524 ,csa_tree_add_190_195_groupi_n_9764 ,csa_tree_add_190_195_groupi_n_10314);
  or csa_tree_add_190_195_groupi_g38424(csa_tree_add_190_195_groupi_n_10523 ,csa_tree_add_190_195_groupi_n_10268 ,csa_tree_add_190_195_groupi_n_10233);
  or csa_tree_add_190_195_groupi_g38425(csa_tree_add_190_195_groupi_n_10522 ,csa_tree_add_190_195_groupi_n_9655 ,csa_tree_add_190_195_groupi_n_10263);
  or csa_tree_add_190_195_groupi_g38426(csa_tree_add_190_195_groupi_n_10521 ,csa_tree_add_190_195_groupi_n_9771 ,csa_tree_add_190_195_groupi_n_10170);
  nor csa_tree_add_190_195_groupi_g38427(csa_tree_add_190_195_groupi_n_10520 ,csa_tree_add_190_195_groupi_n_9877 ,csa_tree_add_190_195_groupi_n_10192);
  or csa_tree_add_190_195_groupi_g38428(csa_tree_add_190_195_groupi_n_10519 ,csa_tree_add_190_195_groupi_n_9995 ,csa_tree_add_190_195_groupi_n_10227);
  and csa_tree_add_190_195_groupi_g38429(csa_tree_add_190_195_groupi_n_10518 ,csa_tree_add_190_195_groupi_n_10348 ,csa_tree_add_190_195_groupi_n_10124);
  and csa_tree_add_190_195_groupi_g38430(csa_tree_add_190_195_groupi_n_10517 ,csa_tree_add_190_195_groupi_n_10119 ,csa_tree_add_190_195_groupi_n_10351);
  or csa_tree_add_190_195_groupi_g38431(csa_tree_add_190_195_groupi_n_10516 ,csa_tree_add_190_195_groupi_n_9847 ,csa_tree_add_190_195_groupi_n_10219);
  or csa_tree_add_190_195_groupi_g38432(csa_tree_add_190_195_groupi_n_10515 ,csa_tree_add_190_195_groupi_n_10333 ,csa_tree_add_190_195_groupi_n_10257);
  nor csa_tree_add_190_195_groupi_g38433(csa_tree_add_190_195_groupi_n_10514 ,csa_tree_add_190_195_groupi_n_9861 ,csa_tree_add_190_195_groupi_n_10182);
  or csa_tree_add_190_195_groupi_g38434(csa_tree_add_190_195_groupi_n_10513 ,csa_tree_add_190_195_groupi_n_9862 ,csa_tree_add_190_195_groupi_n_10181);
  or csa_tree_add_190_195_groupi_g38435(csa_tree_add_190_195_groupi_n_10512 ,csa_tree_add_190_195_groupi_n_10318 ,csa_tree_add_190_195_groupi_n_9868);
  nor csa_tree_add_190_195_groupi_g38436(csa_tree_add_190_195_groupi_n_10511 ,csa_tree_add_190_195_groupi_n_10319 ,csa_tree_add_190_195_groupi_n_9867);
  or csa_tree_add_190_195_groupi_g38437(csa_tree_add_190_195_groupi_n_10510 ,csa_tree_add_190_195_groupi_n_9954 ,csa_tree_add_190_195_groupi_n_10246);
  or csa_tree_add_190_195_groupi_g38438(csa_tree_add_190_195_groupi_n_10509 ,csa_tree_add_190_195_groupi_n_10077 ,csa_tree_add_190_195_groupi_n_10242);
  or csa_tree_add_190_195_groupi_g38439(csa_tree_add_190_195_groupi_n_10508 ,csa_tree_add_190_195_groupi_n_10083 ,csa_tree_add_190_195_groupi_n_10127);
  or csa_tree_add_190_195_groupi_g38440(csa_tree_add_190_195_groupi_n_10507 ,csa_tree_add_190_195_groupi_n_10070 ,csa_tree_add_190_195_groupi_n_10306);
  nor csa_tree_add_190_195_groupi_g38441(csa_tree_add_190_195_groupi_n_10506 ,csa_tree_add_190_195_groupi_n_9322 ,csa_tree_add_190_195_groupi_n_10324);
  and csa_tree_add_190_195_groupi_g38442(csa_tree_add_190_195_groupi_n_10505 ,csa_tree_add_190_195_groupi_n_9806 ,csa_tree_add_190_195_groupi_n_10237);
  or csa_tree_add_190_195_groupi_g38443(csa_tree_add_190_195_groupi_n_10504 ,csa_tree_add_190_195_groupi_n_9321 ,csa_tree_add_190_195_groupi_n_10323);
  nor csa_tree_add_190_195_groupi_g38444(csa_tree_add_190_195_groupi_n_10503 ,csa_tree_add_190_195_groupi_n_9667 ,csa_tree_add_190_195_groupi_n_10272);
  or csa_tree_add_190_195_groupi_g38445(csa_tree_add_190_195_groupi_n_10502 ,csa_tree_add_190_195_groupi_n_8659 ,csa_tree_add_190_195_groupi_n_10197);
  nor csa_tree_add_190_195_groupi_g38446(csa_tree_add_190_195_groupi_n_10501 ,csa_tree_add_190_195_groupi_n_8660 ,csa_tree_add_190_195_groupi_n_10198);
  or csa_tree_add_190_195_groupi_g38447(csa_tree_add_190_195_groupi_n_10500 ,csa_tree_add_190_195_groupi_n_9878 ,csa_tree_add_190_195_groupi_n_10191);
  or csa_tree_add_190_195_groupi_g38448(csa_tree_add_190_195_groupi_n_10499 ,csa_tree_add_190_195_groupi_n_9287 ,csa_tree_add_190_195_groupi_n_10166);
  and csa_tree_add_190_195_groupi_g38449(csa_tree_add_190_195_groupi_n_10498 ,csa_tree_add_190_195_groupi_n_10223 ,csa_tree_add_190_195_groupi_n_9966);
  nor csa_tree_add_190_195_groupi_g38450(csa_tree_add_190_195_groupi_n_10497 ,csa_tree_add_190_195_groupi_n_9288 ,csa_tree_add_190_195_groupi_n_10167);
  or csa_tree_add_190_195_groupi_g38451(csa_tree_add_190_195_groupi_n_10496 ,csa_tree_add_190_195_groupi_n_10336 ,csa_tree_add_190_195_groupi_n_10258);
  or csa_tree_add_190_195_groupi_g38452(csa_tree_add_190_195_groupi_n_10495 ,csa_tree_add_190_195_groupi_n_9633 ,csa_tree_add_190_195_groupi_n_10216);
  nor csa_tree_add_190_195_groupi_g38453(csa_tree_add_190_195_groupi_n_10494 ,csa_tree_add_190_195_groupi_n_9634 ,csa_tree_add_190_195_groupi_n_10217);
  or csa_tree_add_190_195_groupi_g38454(csa_tree_add_190_195_groupi_n_10493 ,csa_tree_add_190_195_groupi_n_10215 ,csa_tree_add_190_195_groupi_n_10214);
  and csa_tree_add_190_195_groupi_g38455(csa_tree_add_190_195_groupi_n_10492 ,csa_tree_add_190_195_groupi_n_10215 ,csa_tree_add_190_195_groupi_n_10214);
  nor csa_tree_add_190_195_groupi_g38456(csa_tree_add_190_195_groupi_n_10491 ,csa_tree_add_190_195_groupi_n_10325 ,csa_tree_add_190_195_groupi_n_10204);
  or csa_tree_add_190_195_groupi_g38457(csa_tree_add_190_195_groupi_n_10490 ,csa_tree_add_190_195_groupi_n_10199 ,csa_tree_add_190_195_groupi_n_9932);
  or csa_tree_add_190_195_groupi_g38458(csa_tree_add_190_195_groupi_n_10489 ,csa_tree_add_190_195_groupi_n_10326 ,csa_tree_add_190_195_groupi_n_10203);
  nor csa_tree_add_190_195_groupi_g38459(csa_tree_add_190_195_groupi_n_10488 ,csa_tree_add_190_195_groupi_n_10200 ,csa_tree_add_190_195_groupi_n_9933);
  or csa_tree_add_190_195_groupi_g38460(csa_tree_add_190_195_groupi_n_10487 ,csa_tree_add_190_195_groupi_n_10055 ,csa_tree_add_190_195_groupi_n_10194);
  or csa_tree_add_190_195_groupi_g38461(csa_tree_add_190_195_groupi_n_10486 ,csa_tree_add_190_195_groupi_n_9766 ,csa_tree_add_190_195_groupi_n_10173);
  or csa_tree_add_190_195_groupi_g38462(csa_tree_add_190_195_groupi_n_10485 ,csa_tree_add_190_195_groupi_n_9914 ,csa_tree_add_190_195_groupi_n_10312);
  nor csa_tree_add_190_195_groupi_g38463(csa_tree_add_190_195_groupi_n_10484 ,csa_tree_add_190_195_groupi_n_9915 ,csa_tree_add_190_195_groupi_n_10313);
  or csa_tree_add_190_195_groupi_g38464(csa_tree_add_190_195_groupi_n_10483 ,csa_tree_add_190_195_groupi_n_10069 ,csa_tree_add_190_195_groupi_n_10299);
  nor csa_tree_add_190_195_groupi_g38465(csa_tree_add_190_195_groupi_n_10482 ,csa_tree_add_190_195_groupi_n_10328 ,csa_tree_add_190_195_groupi_n_10195);
  or csa_tree_add_190_195_groupi_g38466(csa_tree_add_190_195_groupi_n_10481 ,csa_tree_add_190_195_groupi_n_9630 ,csa_tree_add_190_195_groupi_n_10146);
  nor csa_tree_add_190_195_groupi_g38467(csa_tree_add_190_195_groupi_n_10480 ,csa_tree_add_190_195_groupi_n_9629 ,csa_tree_add_190_195_groupi_n_10147);
  or csa_tree_add_190_195_groupi_g38468(csa_tree_add_190_195_groupi_n_10479 ,csa_tree_add_190_195_groupi_n_9894 ,csa_tree_add_190_195_groupi_n_10316);
  nor csa_tree_add_190_195_groupi_g38469(csa_tree_add_190_195_groupi_n_10478 ,csa_tree_add_190_195_groupi_n_9893 ,csa_tree_add_190_195_groupi_n_10317);
  nor csa_tree_add_190_195_groupi_g38470(csa_tree_add_190_195_groupi_n_10477 ,csa_tree_add_190_195_groupi_n_10056 ,csa_tree_add_190_195_groupi_n_10193);
  or csa_tree_add_190_195_groupi_g38471(csa_tree_add_190_195_groupi_n_10476 ,csa_tree_add_190_195_groupi_n_10327 ,csa_tree_add_190_195_groupi_n_10196);
  nor csa_tree_add_190_195_groupi_g38472(csa_tree_add_190_195_groupi_n_10475 ,csa_tree_add_190_195_groupi_n_9765 ,csa_tree_add_190_195_groupi_n_10174);
  and csa_tree_add_190_195_groupi_g38473(csa_tree_add_190_195_groupi_n_10591 ,csa_tree_add_190_195_groupi_n_8131 ,csa_tree_add_190_195_groupi_n_10298);
  and csa_tree_add_190_195_groupi_g38474(csa_tree_add_190_195_groupi_n_10590 ,csa_tree_add_190_195_groupi_n_9678 ,csa_tree_add_190_195_groupi_n_10235);
  and csa_tree_add_190_195_groupi_g38475(csa_tree_add_190_195_groupi_n_10589 ,csa_tree_add_190_195_groupi_n_9999 ,csa_tree_add_190_195_groupi_n_10239);
  and csa_tree_add_190_195_groupi_g38476(csa_tree_add_190_195_groupi_n_10588 ,csa_tree_add_190_195_groupi_n_9974 ,csa_tree_add_190_195_groupi_n_10241);
  and csa_tree_add_190_195_groupi_g38477(csa_tree_add_190_195_groupi_n_10587 ,csa_tree_add_190_195_groupi_n_9985 ,csa_tree_add_190_195_groupi_n_10251);
  and csa_tree_add_190_195_groupi_g38478(csa_tree_add_190_195_groupi_n_10586 ,csa_tree_add_190_195_groupi_n_9981 ,csa_tree_add_190_195_groupi_n_10262);
  or csa_tree_add_190_195_groupi_g38479(csa_tree_add_190_195_groupi_n_10585 ,csa_tree_add_190_195_groupi_n_9983 ,csa_tree_add_190_195_groupi_n_10265);
  and csa_tree_add_190_195_groupi_g38480(csa_tree_add_190_195_groupi_n_10584 ,csa_tree_add_190_195_groupi_n_9857 ,csa_tree_add_190_195_groupi_n_10275);
  or csa_tree_add_190_195_groupi_g38481(csa_tree_add_190_195_groupi_n_10583 ,csa_tree_add_190_195_groupi_n_10030 ,csa_tree_add_190_195_groupi_n_10115);
  and csa_tree_add_190_195_groupi_g38482(csa_tree_add_190_195_groupi_n_10582 ,csa_tree_add_190_195_groupi_n_9728 ,csa_tree_add_190_195_groupi_n_10280);
  and csa_tree_add_190_195_groupi_g38483(csa_tree_add_190_195_groupi_n_10581 ,csa_tree_add_190_195_groupi_n_9738 ,csa_tree_add_190_195_groupi_n_10291);
  or csa_tree_add_190_195_groupi_g38484(csa_tree_add_190_195_groupi_n_10579 ,csa_tree_add_190_195_groupi_n_10025 ,csa_tree_add_190_195_groupi_n_10300);
  and csa_tree_add_190_195_groupi_g38485(csa_tree_add_190_195_groupi_n_10578 ,csa_tree_add_190_195_groupi_n_9843 ,csa_tree_add_190_195_groupi_n_10140);
  and csa_tree_add_190_195_groupi_g38486(csa_tree_add_190_195_groupi_n_10577 ,csa_tree_add_190_195_groupi_n_9964 ,csa_tree_add_190_195_groupi_n_10254);
  and csa_tree_add_190_195_groupi_g38487(csa_tree_add_190_195_groupi_n_10576 ,csa_tree_add_190_195_groupi_n_10033 ,csa_tree_add_190_195_groupi_n_10310);
  or csa_tree_add_190_195_groupi_g38488(csa_tree_add_190_195_groupi_n_10574 ,csa_tree_add_190_195_groupi_n_9597 ,csa_tree_add_190_195_groupi_n_10295);
  or csa_tree_add_190_195_groupi_g38489(csa_tree_add_190_195_groupi_n_10571 ,csa_tree_add_190_195_groupi_n_9976 ,csa_tree_add_190_195_groupi_n_10294);
  and csa_tree_add_190_195_groupi_g38490(csa_tree_add_190_195_groupi_n_10570 ,csa_tree_add_190_195_groupi_n_8077 ,csa_tree_add_190_195_groupi_n_10276);
  and csa_tree_add_190_195_groupi_g38491(csa_tree_add_190_195_groupi_n_10567 ,csa_tree_add_190_195_groupi_n_9409 ,csa_tree_add_190_195_groupi_n_10279);
  or csa_tree_add_190_195_groupi_g38492(csa_tree_add_190_195_groupi_n_10565 ,csa_tree_add_190_195_groupi_n_9975 ,csa_tree_add_190_195_groupi_n_10288);
  or csa_tree_add_190_195_groupi_g38493(csa_tree_add_190_195_groupi_n_10563 ,csa_tree_add_190_195_groupi_n_10032 ,csa_tree_add_190_195_groupi_n_10144);
  or csa_tree_add_190_195_groupi_g38494(csa_tree_add_190_195_groupi_n_10562 ,csa_tree_add_190_195_groupi_n_9977 ,csa_tree_add_190_195_groupi_n_10248);
  or csa_tree_add_190_195_groupi_g38495(csa_tree_add_190_195_groupi_n_10561 ,csa_tree_add_190_195_groupi_n_10014 ,csa_tree_add_190_195_groupi_n_10290);
  and csa_tree_add_190_195_groupi_g38496(csa_tree_add_190_195_groupi_n_10559 ,csa_tree_add_190_195_groupi_n_9583 ,csa_tree_add_190_195_groupi_n_10250);
  and csa_tree_add_190_195_groupi_g38497(csa_tree_add_190_195_groupi_n_10556 ,csa_tree_add_190_195_groupi_n_9968 ,csa_tree_add_190_195_groupi_n_10284);
  and csa_tree_add_190_195_groupi_g38498(csa_tree_add_190_195_groupi_n_10554 ,csa_tree_add_190_195_groupi_n_9695 ,csa_tree_add_190_195_groupi_n_10252);
  or csa_tree_add_190_195_groupi_g38499(csa_tree_add_190_195_groupi_n_10552 ,csa_tree_add_190_195_groupi_n_9146 ,csa_tree_add_190_195_groupi_n_10304);
  and csa_tree_add_190_195_groupi_g38500(csa_tree_add_190_195_groupi_n_10551 ,csa_tree_add_190_195_groupi_n_10018 ,csa_tree_add_190_195_groupi_n_10261);
  not csa_tree_add_190_195_groupi_g38501(csa_tree_add_190_195_groupi_n_10472 ,csa_tree_add_190_195_groupi_n_10471);
  not csa_tree_add_190_195_groupi_g38502(csa_tree_add_190_195_groupi_n_10465 ,csa_tree_add_190_195_groupi_n_10464);
  not csa_tree_add_190_195_groupi_g38503(csa_tree_add_190_195_groupi_n_10462 ,csa_tree_add_190_195_groupi_n_10461);
  not csa_tree_add_190_195_groupi_g38504(csa_tree_add_190_195_groupi_n_10460 ,csa_tree_add_190_195_groupi_n_10459);
  not csa_tree_add_190_195_groupi_g38505(csa_tree_add_190_195_groupi_n_10457 ,csa_tree_add_190_195_groupi_n_10456);
  not csa_tree_add_190_195_groupi_g38506(csa_tree_add_190_195_groupi_n_10455 ,csa_tree_add_190_195_groupi_n_143);
  not csa_tree_add_190_195_groupi_g38507(csa_tree_add_190_195_groupi_n_10454 ,csa_tree_add_190_195_groupi_n_10453);
  not csa_tree_add_190_195_groupi_g38508(csa_tree_add_190_195_groupi_n_10452 ,csa_tree_add_190_195_groupi_n_10451);
  not csa_tree_add_190_195_groupi_g38509(csa_tree_add_190_195_groupi_n_10450 ,csa_tree_add_190_195_groupi_n_10449);
  not csa_tree_add_190_195_groupi_g38510(csa_tree_add_190_195_groupi_n_10448 ,csa_tree_add_190_195_groupi_n_138);
  not csa_tree_add_190_195_groupi_g38511(csa_tree_add_190_195_groupi_n_10447 ,csa_tree_add_190_195_groupi_n_10446);
  not csa_tree_add_190_195_groupi_g38512(csa_tree_add_190_195_groupi_n_10445 ,csa_tree_add_190_195_groupi_n_10444);
  not csa_tree_add_190_195_groupi_g38513(csa_tree_add_190_195_groupi_n_10441 ,csa_tree_add_190_195_groupi_n_10440);
  not csa_tree_add_190_195_groupi_g38514(csa_tree_add_190_195_groupi_n_10439 ,csa_tree_add_190_195_groupi_n_10438);
  not csa_tree_add_190_195_groupi_g38515(csa_tree_add_190_195_groupi_n_10437 ,csa_tree_add_190_195_groupi_n_10436);
  not csa_tree_add_190_195_groupi_g38516(csa_tree_add_190_195_groupi_n_10435 ,csa_tree_add_190_195_groupi_n_10434);
  not csa_tree_add_190_195_groupi_g38517(csa_tree_add_190_195_groupi_n_10433 ,csa_tree_add_190_195_groupi_n_10432);
  not csa_tree_add_190_195_groupi_g38518(csa_tree_add_190_195_groupi_n_10431 ,csa_tree_add_190_195_groupi_n_10430);
  not csa_tree_add_190_195_groupi_g38519(csa_tree_add_190_195_groupi_n_10429 ,csa_tree_add_190_195_groupi_n_10428);
  not csa_tree_add_190_195_groupi_g38520(csa_tree_add_190_195_groupi_n_10427 ,csa_tree_add_190_195_groupi_n_10426);
  not csa_tree_add_190_195_groupi_g38521(csa_tree_add_190_195_groupi_n_10425 ,csa_tree_add_190_195_groupi_n_10424);
  or csa_tree_add_190_195_groupi_g38522(csa_tree_add_190_195_groupi_n_10419 ,csa_tree_add_190_195_groupi_n_9879 ,csa_tree_add_190_195_groupi_n_10168);
  or csa_tree_add_190_195_groupi_g38523(csa_tree_add_190_195_groupi_n_10418 ,csa_tree_add_190_195_groupi_n_10085 ,csa_tree_add_190_195_groupi_n_10133);
  or csa_tree_add_190_195_groupi_g38524(csa_tree_add_190_195_groupi_n_10417 ,csa_tree_add_190_195_groupi_n_10075 ,csa_tree_add_190_195_groupi_n_10130);
  or csa_tree_add_190_195_groupi_g38525(csa_tree_add_190_195_groupi_n_10416 ,csa_tree_add_190_195_groupi_n_10082 ,csa_tree_add_190_195_groupi_n_10131);
  or csa_tree_add_190_195_groupi_g38526(csa_tree_add_190_195_groupi_n_10415 ,csa_tree_add_190_195_groupi_n_8691 ,csa_tree_add_190_195_groupi_n_10322);
  nor csa_tree_add_190_195_groupi_g38527(csa_tree_add_190_195_groupi_n_10414 ,csa_tree_add_190_195_groupi_n_10188 ,csa_tree_add_190_195_groupi_n_9898);
  or csa_tree_add_190_195_groupi_g38528(csa_tree_add_190_195_groupi_n_10413 ,csa_tree_add_190_195_groupi_n_10187 ,csa_tree_add_190_195_groupi_n_9899);
  or csa_tree_add_190_195_groupi_g38529(csa_tree_add_190_195_groupi_n_10412 ,csa_tree_add_190_195_groupi_n_10038 ,csa_tree_add_190_195_groupi_n_10180);
  or csa_tree_add_190_195_groupi_g38530(csa_tree_add_190_195_groupi_n_10411 ,csa_tree_add_190_195_groupi_n_9888 ,csa_tree_add_190_195_groupi_n_10177);
  nor csa_tree_add_190_195_groupi_g38531(csa_tree_add_190_195_groupi_n_10410 ,csa_tree_add_190_195_groupi_n_9887 ,csa_tree_add_190_195_groupi_n_10178);
  or csa_tree_add_190_195_groupi_g38532(csa_tree_add_190_195_groupi_n_10409 ,csa_tree_add_190_195_groupi_n_9475 ,csa_tree_add_190_195_groupi_n_10162);
  and csa_tree_add_190_195_groupi_g38533(csa_tree_add_190_195_groupi_n_10408 ,csa_tree_add_190_195_groupi_n_9771 ,csa_tree_add_190_195_groupi_n_10170);
  nor csa_tree_add_190_195_groupi_g38534(csa_tree_add_190_195_groupi_n_10407 ,csa_tree_add_190_195_groupi_n_9609 ,csa_tree_add_190_195_groupi_n_10206);
  nor csa_tree_add_190_195_groupi_g38535(csa_tree_add_190_195_groupi_n_10406 ,csa_tree_add_190_195_groupi_n_9880 ,csa_tree_add_190_195_groupi_n_10169);
  nor csa_tree_add_190_195_groupi_g38536(csa_tree_add_190_195_groupi_n_10405 ,csa_tree_add_190_195_groupi_n_10039 ,csa_tree_add_190_195_groupi_n_10179);
  nor csa_tree_add_190_195_groupi_g38537(csa_tree_add_190_195_groupi_n_10404 ,csa_tree_add_190_195_groupi_n_9474 ,csa_tree_add_190_195_groupi_n_10163);
  or csa_tree_add_190_195_groupi_g38538(csa_tree_add_190_195_groupi_n_10403 ,csa_tree_add_190_195_groupi_n_10332 ,csa_tree_add_190_195_groupi_n_8629);
  or csa_tree_add_190_195_groupi_g38539(csa_tree_add_190_195_groupi_n_10402 ,csa_tree_add_190_195_groupi_n_10222 ,csa_tree_add_190_195_groupi_n_10121);
  or csa_tree_add_190_195_groupi_g38540(csa_tree_add_190_195_groupi_n_10401 ,csa_tree_add_190_195_groupi_n_10122 ,csa_tree_add_190_195_groupi_n_10224);
  nor csa_tree_add_190_195_groupi_g38541(csa_tree_add_190_195_groupi_n_10400 ,csa_tree_add_190_195_groupi_n_9874 ,csa_tree_add_190_195_groupi_n_10155);
  and csa_tree_add_190_195_groupi_g38542(csa_tree_add_190_195_groupi_n_10399 ,csa_tree_add_190_195_groupi_n_9874 ,csa_tree_add_190_195_groupi_n_10155);
  or csa_tree_add_190_195_groupi_g38543(csa_tree_add_190_195_groupi_n_10398 ,csa_tree_add_190_195_groupi_n_10352 ,csa_tree_add_190_195_groupi_n_10117);
  and csa_tree_add_190_195_groupi_g38544(csa_tree_add_190_195_groupi_n_10397 ,csa_tree_add_190_195_groupi_n_8691 ,csa_tree_add_190_195_groupi_n_10322);
  nor csa_tree_add_190_195_groupi_g38545(csa_tree_add_190_195_groupi_n_10396 ,csa_tree_add_190_195_groupi_n_9794 ,csa_tree_add_190_195_groupi_n_10137);
  or csa_tree_add_190_195_groupi_g38546(csa_tree_add_190_195_groupi_n_10395 ,csa_tree_add_190_195_groupi_n_9608 ,csa_tree_add_190_195_groupi_n_10205);
  xor csa_tree_add_190_195_groupi_g38548(csa_tree_add_190_195_groupi_n_10394 ,csa_tree_add_190_195_groupi_n_10078 ,csa_tree_add_190_195_groupi_n_9764);
  xnor csa_tree_add_190_195_groupi_g38549(csa_tree_add_190_195_groupi_n_10393 ,csa_tree_add_190_195_groupi_n_8994 ,csa_tree_add_190_195_groupi_n_9866);
  xnor csa_tree_add_190_195_groupi_g38550(csa_tree_add_190_195_groupi_n_10392 ,csa_tree_add_190_195_groupi_n_9484 ,csa_tree_add_190_195_groupi_n_10041);
  xnor csa_tree_add_190_195_groupi_g38551(csa_tree_add_190_195_groupi_n_10391 ,csa_tree_add_190_195_groupi_n_9655 ,csa_tree_add_190_195_groupi_n_9864);
  xnor csa_tree_add_190_195_groupi_g38552(csa_tree_add_190_195_groupi_n_10390 ,csa_tree_add_190_195_groupi_n_9290 ,csa_tree_add_190_195_groupi_n_10044);
  xor csa_tree_add_190_195_groupi_g38554(csa_tree_add_190_195_groupi_n_10389 ,csa_tree_add_190_195_groupi_n_9931 ,csa_tree_add_190_195_groupi_n_9667);
  xnor csa_tree_add_190_195_groupi_g38555(csa_tree_add_190_195_groupi_n_10388 ,csa_tree_add_190_195_groupi_n_8488 ,csa_tree_add_190_195_groupi_n_9955);
  xnor csa_tree_add_190_195_groupi_g38556(csa_tree_add_190_195_groupi_n_10387 ,csa_tree_add_190_195_groupi_n_10080 ,csa_tree_add_190_195_groupi_n_9334);
  xnor csa_tree_add_190_195_groupi_g38557(csa_tree_add_190_195_groupi_n_10386 ,csa_tree_add_190_195_groupi_n_9619 ,csa_tree_add_190_195_groupi_n_10054);
  xnor csa_tree_add_190_195_groupi_g38559(csa_tree_add_190_195_groupi_n_10385 ,csa_tree_add_190_195_groupi_n_9892 ,csa_tree_add_190_195_groupi_n_9886);
  xnor csa_tree_add_190_195_groupi_g38560(csa_tree_add_190_195_groupi_n_10384 ,csa_tree_add_190_195_groupi_n_9494 ,csa_tree_add_190_195_groupi_n_9903);
  xnor csa_tree_add_190_195_groupi_g38561(csa_tree_add_190_195_groupi_n_10383 ,csa_tree_add_190_195_groupi_n_10082 ,csa_tree_add_190_195_groupi_n_8999);
  xnor csa_tree_add_190_195_groupi_g38562(csa_tree_add_190_195_groupi_n_10382 ,csa_tree_add_190_195_groupi_n_7129 ,csa_tree_add_190_195_groupi_n_9960);
  xnor csa_tree_add_190_195_groupi_g38563(csa_tree_add_190_195_groupi_n_10381 ,csa_tree_add_190_195_groupi_n_8660 ,csa_tree_add_190_195_groupi_n_10086);
  xnor csa_tree_add_190_195_groupi_g38564(csa_tree_add_190_195_groupi_n_10380 ,csa_tree_add_190_195_groupi_n_8693 ,csa_tree_add_190_195_groupi_n_10065);
  xnor csa_tree_add_190_195_groupi_g38565(csa_tree_add_190_195_groupi_n_10379 ,csa_tree_add_190_195_groupi_n_7551 ,csa_tree_add_190_195_groupi_n_10064);
  xnor csa_tree_add_190_195_groupi_g38566(csa_tree_add_190_195_groupi_n_10378 ,csa_tree_add_190_195_groupi_n_10042 ,csa_tree_add_190_195_groupi_n_9295);
  xnor csa_tree_add_190_195_groupi_g38567(csa_tree_add_190_195_groupi_n_10377 ,csa_tree_add_190_195_groupi_n_9961 ,csa_tree_add_190_195_groupi_n_9761);
  xnor csa_tree_add_190_195_groupi_g38568(csa_tree_add_190_195_groupi_n_10376 ,csa_tree_add_190_195_groupi_n_7591 ,csa_tree_add_190_195_groupi_n_9882);
  xnor csa_tree_add_190_195_groupi_g38569(csa_tree_add_190_195_groupi_n_10375 ,csa_tree_add_190_195_groupi_n_8504 ,csa_tree_add_190_195_groupi_n_9919);
  xnor csa_tree_add_190_195_groupi_g38570(csa_tree_add_190_195_groupi_n_10374 ,csa_tree_add_190_195_groupi_n_9658 ,csa_tree_add_190_195_groupi_n_9897);
  xnor csa_tree_add_190_195_groupi_g38571(csa_tree_add_190_195_groupi_n_10373 ,csa_tree_add_190_195_groupi_n_9294 ,csa_tree_add_190_195_groupi_n_9936);
  xnor csa_tree_add_190_195_groupi_g38572(csa_tree_add_190_195_groupi_n_10372 ,csa_tree_add_190_195_groupi_n_10069 ,csa_tree_add_190_195_groupi_n_9884);
  xnor csa_tree_add_190_195_groupi_g38573(csa_tree_add_190_195_groupi_n_10371 ,csa_tree_add_190_195_groupi_n_9873 ,csa_tree_add_190_195_groupi_n_10049);
  xnor csa_tree_add_190_195_groupi_g38574(csa_tree_add_190_195_groupi_n_10370 ,csa_tree_add_190_195_groupi_n_10067 ,csa_tree_add_190_195_groupi_n_9640);
  xnor csa_tree_add_190_195_groupi_g38575(csa_tree_add_190_195_groupi_n_10369 ,csa_tree_add_190_195_groupi_n_9477 ,csa_tree_add_190_195_groupi_n_9937);
  xnor csa_tree_add_190_195_groupi_g38576(csa_tree_add_190_195_groupi_n_10368 ,csa_tree_add_190_195_groupi_n_8964 ,csa_tree_add_190_195_groupi_n_9876);
  xnor csa_tree_add_190_195_groupi_g38577(csa_tree_add_190_195_groupi_n_10367 ,csa_tree_add_190_195_groupi_n_9909 ,csa_tree_add_190_195_groupi_n_9907);
  xnor csa_tree_add_190_195_groupi_g38578(csa_tree_add_190_195_groupi_n_10366 ,csa_tree_add_190_195_groupi_n_9501 ,csa_tree_add_190_195_groupi_n_9916);
  xnor csa_tree_add_190_195_groupi_g38579(csa_tree_add_190_195_groupi_n_10365 ,csa_tree_add_190_195_groupi_n_7070 ,csa_tree_add_190_195_groupi_n_9958);
  xnor csa_tree_add_190_195_groupi_g38580(csa_tree_add_190_195_groupi_n_10364 ,csa_tree_add_190_195_groupi_n_8945 ,csa_tree_add_190_195_groupi_n_9946);
  xnor csa_tree_add_190_195_groupi_g38581(csa_tree_add_190_195_groupi_n_10363 ,csa_tree_add_190_195_groupi_n_9934 ,csa_tree_add_190_195_groupi_n_9789);
  xnor csa_tree_add_190_195_groupi_g38582(csa_tree_add_190_195_groupi_n_10362 ,csa_tree_add_190_195_groupi_n_9926 ,csa_tree_add_190_195_groupi_n_9924);
  xnor csa_tree_add_190_195_groupi_g38583(csa_tree_add_190_195_groupi_n_10361 ,csa_tree_add_190_195_groupi_n_9622 ,csa_tree_add_190_195_groupi_n_10051);
  xnor csa_tree_add_190_195_groupi_g38584(csa_tree_add_190_195_groupi_n_10360 ,csa_tree_add_190_195_groupi_n_9905 ,csa_tree_add_190_195_groupi_n_10077);
  xnor csa_tree_add_190_195_groupi_g38585(csa_tree_add_190_195_groupi_n_10359 ,csa_tree_add_190_195_groupi_n_9603 ,csa_tree_add_190_195_groupi_n_9957);
  xnor csa_tree_add_190_195_groupi_g38586(csa_tree_add_190_195_groupi_n_10358 ,csa_tree_add_190_195_groupi_n_8840 ,csa_tree_add_190_195_groupi_n_9953);
  xnor csa_tree_add_190_195_groupi_g38587(csa_tree_add_190_195_groupi_n_10357 ,csa_tree_add_190_195_groupi_n_8617 ,csa_tree_add_190_195_groupi_n_10061);
  xnor csa_tree_add_190_195_groupi_g38588(csa_tree_add_190_195_groupi_n_10356 ,csa_tree_add_190_195_groupi_n_10083 ,csa_tree_add_190_195_groupi_n_9890);
  and csa_tree_add_190_195_groupi_g38589(csa_tree_add_190_195_groupi_n_10474 ,csa_tree_add_190_195_groupi_n_9855 ,csa_tree_add_190_195_groupi_n_10136);
  xnor csa_tree_add_190_195_groupi_g38590(csa_tree_add_190_195_groupi_n_10473 ,csa_tree_add_190_195_groupi_n_9301 ,csa_tree_add_190_195_groupi_n_9834);
  xnor csa_tree_add_190_195_groupi_g38591(csa_tree_add_190_195_groupi_n_10471 ,csa_tree_add_190_195_groupi_n_9011 ,csa_tree_add_190_195_groupi_n_9815);
  xnor csa_tree_add_190_195_groupi_g38592(csa_tree_add_190_195_groupi_n_10470 ,csa_tree_add_190_195_groupi_n_9358 ,csa_tree_add_190_195_groupi_n_131);
  xnor csa_tree_add_190_195_groupi_g38593(csa_tree_add_190_195_groupi_n_10469 ,csa_tree_add_190_195_groupi_n_7061 ,csa_tree_add_190_195_groupi_n_9814);
  xnor csa_tree_add_190_195_groupi_g38594(csa_tree_add_190_195_groupi_n_10468 ,csa_tree_add_190_195_groupi_n_9017 ,csa_tree_add_190_195_groupi_n_9812);
  xnor csa_tree_add_190_195_groupi_g38595(csa_tree_add_190_195_groupi_n_10467 ,csa_tree_add_190_195_groupi_n_9650 ,csa_tree_add_190_195_groupi_n_9824);
  xnor csa_tree_add_190_195_groupi_g38596(csa_tree_add_190_195_groupi_n_10466 ,csa_tree_add_190_195_groupi_n_9512 ,csa_tree_add_190_195_groupi_n_9833);
  xnor csa_tree_add_190_195_groupi_g38597(csa_tree_add_190_195_groupi_n_10464 ,csa_tree_add_190_195_groupi_n_9013 ,csa_tree_add_190_195_groupi_n_9826);
  xnor csa_tree_add_190_195_groupi_g38598(csa_tree_add_190_195_groupi_n_10463 ,csa_tree_add_190_195_groupi_n_9652 ,csa_tree_add_190_195_groupi_n_9832);
  xnor csa_tree_add_190_195_groupi_g38599(csa_tree_add_190_195_groupi_n_10461 ,csa_tree_add_190_195_groupi_n_7980 ,csa_tree_add_190_195_groupi_n_9836);
  and csa_tree_add_190_195_groupi_g38600(csa_tree_add_190_195_groupi_n_10459 ,csa_tree_add_190_195_groupi_n_9846 ,csa_tree_add_190_195_groupi_n_10118);
  xnor csa_tree_add_190_195_groupi_g38601(csa_tree_add_190_195_groupi_n_10458 ,csa_tree_add_190_195_groupi_n_9620 ,csa_tree_add_190_195_groupi_n_9825);
  and csa_tree_add_190_195_groupi_g38602(csa_tree_add_190_195_groupi_n_10456 ,csa_tree_add_190_195_groupi_n_10005 ,csa_tree_add_190_195_groupi_n_10145);
  xnor csa_tree_add_190_195_groupi_g38604(csa_tree_add_190_195_groupi_n_10453 ,csa_tree_add_190_195_groupi_n_8656 ,csa_tree_add_190_195_groupi_n_9840);
  xnor csa_tree_add_190_195_groupi_g38605(csa_tree_add_190_195_groupi_n_10451 ,csa_tree_add_190_195_groupi_n_7118 ,csa_tree_add_190_195_groupi_n_9823);
  xnor csa_tree_add_190_195_groupi_g38606(csa_tree_add_190_195_groupi_n_10449 ,csa_tree_add_190_195_groupi_n_7624 ,csa_tree_add_190_195_groupi_n_9822);
  xnor csa_tree_add_190_195_groupi_g38608(csa_tree_add_190_195_groupi_n_10446 ,csa_tree_add_190_195_groupi_n_9308 ,csa_tree_add_190_195_groupi_n_9813);
  xnor csa_tree_add_190_195_groupi_g38609(csa_tree_add_190_195_groupi_n_10444 ,csa_tree_add_190_195_groupi_n_7372 ,csa_tree_add_190_195_groupi_n_9831);
  xnor csa_tree_add_190_195_groupi_g38610(csa_tree_add_190_195_groupi_n_10443 ,csa_tree_add_190_195_groupi_n_9168 ,csa_tree_add_190_195_groupi_n_9820);
  xnor csa_tree_add_190_195_groupi_g38611(csa_tree_add_190_195_groupi_n_10442 ,csa_tree_add_190_195_groupi_n_8826 ,csa_tree_add_190_195_groupi_n_129);
  xnor csa_tree_add_190_195_groupi_g38612(csa_tree_add_190_195_groupi_n_10440 ,csa_tree_add_190_195_groupi_n_8637 ,csa_tree_add_190_195_groupi_n_9830);
  xnor csa_tree_add_190_195_groupi_g38613(csa_tree_add_190_195_groupi_n_10438 ,csa_tree_add_190_195_groupi_n_8649 ,csa_tree_add_190_195_groupi_n_9819);
  xnor csa_tree_add_190_195_groupi_g38614(csa_tree_add_190_195_groupi_n_10436 ,csa_tree_add_190_195_groupi_n_8639 ,csa_tree_add_190_195_groupi_n_130);
  xnor csa_tree_add_190_195_groupi_g38615(csa_tree_add_190_195_groupi_n_10434 ,csa_tree_add_190_195_groupi_n_8957 ,csa_tree_add_190_195_groupi_n_9818);
  xnor csa_tree_add_190_195_groupi_g38616(csa_tree_add_190_195_groupi_n_10432 ,csa_tree_add_190_195_groupi_n_9029 ,csa_tree_add_190_195_groupi_n_9829);
  xnor csa_tree_add_190_195_groupi_g38617(csa_tree_add_190_195_groupi_n_10430 ,csa_tree_add_190_195_groupi_n_8953 ,csa_tree_add_190_195_groupi_n_9828);
  xnor csa_tree_add_190_195_groupi_g38618(csa_tree_add_190_195_groupi_n_10428 ,csa_tree_add_190_195_groupi_n_8330 ,csa_tree_add_190_195_groupi_n_9817);
  xnor csa_tree_add_190_195_groupi_g38619(csa_tree_add_190_195_groupi_n_10426 ,csa_tree_add_190_195_groupi_n_9518 ,csa_tree_add_190_195_groupi_n_9835);
  xnor csa_tree_add_190_195_groupi_g38620(csa_tree_add_190_195_groupi_n_10424 ,csa_tree_add_190_195_groupi_n_9959 ,csa_tree_add_190_195_groupi_n_9827);
  xnor csa_tree_add_190_195_groupi_g38621(csa_tree_add_190_195_groupi_n_10423 ,csa_tree_add_190_195_groupi_n_9164 ,csa_tree_add_190_195_groupi_n_9837);
  xnor csa_tree_add_190_195_groupi_g38622(csa_tree_add_190_195_groupi_n_10422 ,csa_tree_add_190_195_groupi_n_9305 ,csa_tree_add_190_195_groupi_n_9841);
  xnor csa_tree_add_190_195_groupi_g38623(csa_tree_add_190_195_groupi_n_10421 ,csa_tree_add_190_195_groupi_n_7316 ,csa_tree_add_190_195_groupi_n_9816);
  xnor csa_tree_add_190_195_groupi_g38624(csa_tree_add_190_195_groupi_n_10420 ,csa_tree_add_190_195_groupi_n_9604 ,csa_tree_add_190_195_groupi_n_9838);
  not csa_tree_add_190_195_groupi_g38627(csa_tree_add_190_195_groupi_n_10344 ,csa_tree_add_190_195_groupi_n_10343);
  not csa_tree_add_190_195_groupi_g38629(csa_tree_add_190_195_groupi_n_10332 ,csa_tree_add_190_195_groupi_n_10331);
  not csa_tree_add_190_195_groupi_g38630(csa_tree_add_190_195_groupi_n_10329 ,csa_tree_add_190_195_groupi_n_10330);
  not csa_tree_add_190_195_groupi_g38631(csa_tree_add_190_195_groupi_n_10328 ,csa_tree_add_190_195_groupi_n_10327);
  not csa_tree_add_190_195_groupi_g38632(csa_tree_add_190_195_groupi_n_10326 ,csa_tree_add_190_195_groupi_n_10325);
  not csa_tree_add_190_195_groupi_g38633(csa_tree_add_190_195_groupi_n_10324 ,csa_tree_add_190_195_groupi_n_10323);
  not csa_tree_add_190_195_groupi_g38634(csa_tree_add_190_195_groupi_n_10321 ,csa_tree_add_190_195_groupi_n_10320);
  not csa_tree_add_190_195_groupi_g38635(csa_tree_add_190_195_groupi_n_10319 ,csa_tree_add_190_195_groupi_n_10318);
  not csa_tree_add_190_195_groupi_g38636(csa_tree_add_190_195_groupi_n_10317 ,csa_tree_add_190_195_groupi_n_10316);
  not csa_tree_add_190_195_groupi_g38637(csa_tree_add_190_195_groupi_n_10313 ,csa_tree_add_190_195_groupi_n_10312);
  and csa_tree_add_190_195_groupi_g38638(csa_tree_add_190_195_groupi_n_10311 ,csa_tree_add_190_195_groupi_n_8945 ,csa_tree_add_190_195_groupi_n_9947);
  or csa_tree_add_190_195_groupi_g38639(csa_tree_add_190_195_groupi_n_10310 ,csa_tree_add_190_195_groupi_n_10087 ,csa_tree_add_190_195_groupi_n_10031);
  or csa_tree_add_190_195_groupi_g38640(csa_tree_add_190_195_groupi_n_10309 ,csa_tree_add_190_195_groupi_n_7639 ,csa_tree_add_190_195_groupi_n_10035);
  nor csa_tree_add_190_195_groupi_g38641(csa_tree_add_190_195_groupi_n_10308 ,csa_tree_add_190_195_groupi_n_8617 ,csa_tree_add_190_195_groupi_n_10062);
  nor csa_tree_add_190_195_groupi_g38642(csa_tree_add_190_195_groupi_n_10307 ,csa_tree_add_190_195_groupi_n_8945 ,csa_tree_add_190_195_groupi_n_9947);
  nor csa_tree_add_190_195_groupi_g38643(csa_tree_add_190_195_groupi_n_10306 ,csa_tree_add_190_195_groupi_n_8963 ,csa_tree_add_190_195_groupi_n_9876);
  or csa_tree_add_190_195_groupi_g38644(csa_tree_add_190_195_groupi_n_10305 ,csa_tree_add_190_195_groupi_n_9768 ,csa_tree_add_190_195_groupi_n_10036);
  and csa_tree_add_190_195_groupi_g38645(csa_tree_add_190_195_groupi_n_10304 ,csa_tree_add_190_195_groupi_n_9144 ,csa_tree_add_190_195_groupi_n_10065);
  or csa_tree_add_190_195_groupi_g38646(csa_tree_add_190_195_groupi_n_10303 ,csa_tree_add_190_195_groupi_n_9943 ,csa_tree_add_190_195_groupi_n_9927);
  or csa_tree_add_190_195_groupi_g38647(csa_tree_add_190_195_groupi_n_10302 ,csa_tree_add_190_195_groupi_n_8964 ,csa_tree_add_190_195_groupi_n_9875);
  nor csa_tree_add_190_195_groupi_g38648(csa_tree_add_190_195_groupi_n_10301 ,csa_tree_add_190_195_groupi_n_9942 ,csa_tree_add_190_195_groupi_n_9928);
  nor csa_tree_add_190_195_groupi_g38649(csa_tree_add_190_195_groupi_n_10300 ,csa_tree_add_190_195_groupi_n_9666 ,csa_tree_add_190_195_groupi_n_10023);
  nor csa_tree_add_190_195_groupi_g38650(csa_tree_add_190_195_groupi_n_10299 ,csa_tree_add_190_195_groupi_n_9177 ,csa_tree_add_190_195_groupi_n_9884);
  or csa_tree_add_190_195_groupi_g38651(csa_tree_add_190_195_groupi_n_10298 ,csa_tree_add_190_195_groupi_n_8126 ,csa_tree_add_190_195_groupi_n_10076);
  nor csa_tree_add_190_195_groupi_g38652(csa_tree_add_190_195_groupi_n_10297 ,csa_tree_add_190_195_groupi_n_9767 ,csa_tree_add_190_195_groupi_n_10037);
  or csa_tree_add_190_195_groupi_g38653(csa_tree_add_190_195_groupi_n_10296 ,csa_tree_add_190_195_groupi_n_9176 ,csa_tree_add_190_195_groupi_n_9883);
  and csa_tree_add_190_195_groupi_g38654(csa_tree_add_190_195_groupi_n_10295 ,csa_tree_add_190_195_groupi_n_9596 ,csa_tree_add_190_195_groupi_n_9953);
  and csa_tree_add_190_195_groupi_g38655(csa_tree_add_190_195_groupi_n_10294 ,csa_tree_add_190_195_groupi_n_9793 ,csa_tree_add_190_195_groupi_n_9998);
  or csa_tree_add_190_195_groupi_g38656(csa_tree_add_190_195_groupi_n_10293 ,csa_tree_add_190_195_groupi_n_9756 ,csa_tree_add_190_195_groupi_n_9913);
  nor csa_tree_add_190_195_groupi_g38657(csa_tree_add_190_195_groupi_n_10292 ,csa_tree_add_190_195_groupi_n_9757 ,csa_tree_add_190_195_groupi_n_9912);
  or csa_tree_add_190_195_groupi_g38658(csa_tree_add_190_195_groupi_n_10291 ,csa_tree_add_190_195_groupi_n_9732 ,csa_tree_add_190_195_groupi_n_10072);
  nor csa_tree_add_190_195_groupi_g38659(csa_tree_add_190_195_groupi_n_10290 ,csa_tree_add_190_195_groupi_n_9511 ,csa_tree_add_190_195_groupi_n_10013);
  nor csa_tree_add_190_195_groupi_g38660(csa_tree_add_190_195_groupi_n_10289 ,csa_tree_add_190_195_groupi_n_8993 ,csa_tree_add_190_195_groupi_n_9866);
  nor csa_tree_add_190_195_groupi_g38661(csa_tree_add_190_195_groupi_n_10288 ,csa_tree_add_190_195_groupi_n_9656 ,csa_tree_add_190_195_groupi_n_9986);
  or csa_tree_add_190_195_groupi_g38662(csa_tree_add_190_195_groupi_n_10287 ,csa_tree_add_190_195_groupi_n_8994 ,csa_tree_add_190_195_groupi_n_9865);
  nor csa_tree_add_190_195_groupi_g38663(csa_tree_add_190_195_groupi_n_10286 ,csa_tree_add_190_195_groupi_n_9926 ,csa_tree_add_190_195_groupi_n_9923);
  nor csa_tree_add_190_195_groupi_g38664(csa_tree_add_190_195_groupi_n_10285 ,csa_tree_add_190_195_groupi_n_8503 ,csa_tree_add_190_195_groupi_n_9919);
  or csa_tree_add_190_195_groupi_g38665(csa_tree_add_190_195_groupi_n_10284 ,csa_tree_add_190_195_groupi_n_9961 ,csa_tree_add_190_195_groupi_n_9971);
  nor csa_tree_add_190_195_groupi_g38666(csa_tree_add_190_195_groupi_n_10283 ,csa_tree_add_190_195_groupi_n_9290 ,csa_tree_add_190_195_groupi_n_10044);
  or csa_tree_add_190_195_groupi_g38667(csa_tree_add_190_195_groupi_n_10282 ,csa_tree_add_190_195_groupi_n_8487 ,csa_tree_add_190_195_groupi_n_10059);
  nor csa_tree_add_190_195_groupi_g38668(csa_tree_add_190_195_groupi_n_10281 ,csa_tree_add_190_195_groupi_n_9501 ,csa_tree_add_190_195_groupi_n_9917);
  or csa_tree_add_190_195_groupi_g38669(csa_tree_add_190_195_groupi_n_10280 ,csa_tree_add_190_195_groupi_n_9725 ,csa_tree_add_190_195_groupi_n_9956);
  or csa_tree_add_190_195_groupi_g38670(csa_tree_add_190_195_groupi_n_10279 ,csa_tree_add_190_195_groupi_n_9403 ,csa_tree_add_190_195_groupi_n_9960);
  and csa_tree_add_190_195_groupi_g38671(csa_tree_add_190_195_groupi_n_10278 ,csa_tree_add_190_195_groupi_n_9501 ,csa_tree_add_190_195_groupi_n_9917);
  or csa_tree_add_190_195_groupi_g38672(csa_tree_add_190_195_groupi_n_10277 ,csa_tree_add_190_195_groupi_n_8504 ,csa_tree_add_190_195_groupi_n_9918);
  or csa_tree_add_190_195_groupi_g38673(csa_tree_add_190_195_groupi_n_10276 ,csa_tree_add_190_195_groupi_n_8076 ,csa_tree_add_190_195_groupi_n_10084);
  or csa_tree_add_190_195_groupi_g38674(csa_tree_add_190_195_groupi_n_10275 ,csa_tree_add_190_195_groupi_n_9795 ,csa_tree_add_190_195_groupi_n_9856);
  or csa_tree_add_190_195_groupi_g38675(csa_tree_add_190_195_groupi_n_10274 ,csa_tree_add_190_195_groupi_n_7550 ,csa_tree_add_190_195_groupi_n_10063);
  nor csa_tree_add_190_195_groupi_g38676(csa_tree_add_190_195_groupi_n_10273 ,csa_tree_add_190_195_groupi_n_8488 ,csa_tree_add_190_195_groupi_n_10060);
  and csa_tree_add_190_195_groupi_g38677(csa_tree_add_190_195_groupi_n_10272 ,csa_tree_add_190_195_groupi_n_8690 ,csa_tree_add_190_195_groupi_n_9931);
  nor csa_tree_add_190_195_groupi_g38678(csa_tree_add_190_195_groupi_n_10271 ,csa_tree_add_190_195_groupi_n_9294 ,csa_tree_add_190_195_groupi_n_9936);
  or csa_tree_add_190_195_groupi_g38679(csa_tree_add_190_195_groupi_n_10270 ,csa_tree_add_190_195_groupi_n_2405 ,csa_tree_add_190_195_groupi_n_9910);
  nor csa_tree_add_190_195_groupi_g38680(csa_tree_add_190_195_groupi_n_10269 ,csa_tree_add_190_195_groupi_n_1310 ,csa_tree_add_190_195_groupi_n_9911);
  nor csa_tree_add_190_195_groupi_g38681(csa_tree_add_190_195_groupi_n_10268 ,csa_tree_add_190_195_groupi_n_7551 ,csa_tree_add_190_195_groupi_n_10064);
  nor csa_tree_add_190_195_groupi_g38682(csa_tree_add_190_195_groupi_n_10267 ,csa_tree_add_190_195_groupi_n_9483 ,csa_tree_add_190_195_groupi_n_10041);
  or csa_tree_add_190_195_groupi_g38683(csa_tree_add_190_195_groupi_n_10266 ,csa_tree_add_190_195_groupi_n_9484 ,csa_tree_add_190_195_groupi_n_10040);
  and csa_tree_add_190_195_groupi_g38684(csa_tree_add_190_195_groupi_n_10265 ,csa_tree_add_190_195_groupi_n_9186 ,csa_tree_add_190_195_groupi_n_9982);
  or csa_tree_add_190_195_groupi_g38685(csa_tree_add_190_195_groupi_n_10264 ,csa_tree_add_190_195_groupi_n_7630 ,csa_tree_add_190_195_groupi_n_9863);
  nor csa_tree_add_190_195_groupi_g38686(csa_tree_add_190_195_groupi_n_10263 ,csa_tree_add_190_195_groupi_n_7631 ,csa_tree_add_190_195_groupi_n_9864);
  or csa_tree_add_190_195_groupi_g38687(csa_tree_add_190_195_groupi_n_10262 ,csa_tree_add_190_195_groupi_n_10079 ,csa_tree_add_190_195_groupi_n_9979);
  or csa_tree_add_190_195_groupi_g38688(csa_tree_add_190_195_groupi_n_10261 ,csa_tree_add_190_195_groupi_n_9796 ,csa_tree_add_190_195_groupi_n_9997);
  nor csa_tree_add_190_195_groupi_g38689(csa_tree_add_190_195_groupi_n_10260 ,csa_tree_add_190_195_groupi_n_8690 ,csa_tree_add_190_195_groupi_n_9931);
  or csa_tree_add_190_195_groupi_g38690(csa_tree_add_190_195_groupi_n_10259 ,csa_tree_add_190_195_groupi_n_9293 ,csa_tree_add_190_195_groupi_n_9935);
  and csa_tree_add_190_195_groupi_g38691(csa_tree_add_190_195_groupi_n_10258 ,csa_tree_add_190_195_groupi_n_9291 ,csa_tree_add_190_195_groupi_n_10052);
  nor csa_tree_add_190_195_groupi_g38692(csa_tree_add_190_195_groupi_n_10257 ,csa_tree_add_190_195_groupi_n_9770 ,csa_tree_add_190_195_groupi_n_9949);
  or csa_tree_add_190_195_groupi_g38693(csa_tree_add_190_195_groupi_n_10256 ,csa_tree_add_190_195_groupi_n_9291 ,csa_tree_add_190_195_groupi_n_10052);
  or csa_tree_add_190_195_groupi_g38694(csa_tree_add_190_195_groupi_n_10255 ,csa_tree_add_190_195_groupi_n_9289 ,csa_tree_add_190_195_groupi_n_10043);
  or csa_tree_add_190_195_groupi_g38695(csa_tree_add_190_195_groupi_n_10254 ,csa_tree_add_190_195_groupi_n_9963 ,csa_tree_add_190_195_groupi_n_10066);
  nor csa_tree_add_190_195_groupi_g38696(csa_tree_add_190_195_groupi_n_10253 ,csa_tree_add_190_195_groupi_n_7640 ,csa_tree_add_190_195_groupi_n_10034);
  or csa_tree_add_190_195_groupi_g38697(csa_tree_add_190_195_groupi_n_10252 ,csa_tree_add_190_195_groupi_n_9694 ,csa_tree_add_190_195_groupi_n_9958);
  or csa_tree_add_190_195_groupi_g38698(csa_tree_add_190_195_groupi_n_10251 ,csa_tree_add_190_195_groupi_n_9356 ,csa_tree_add_190_195_groupi_n_9984);
  or csa_tree_add_190_195_groupi_g38699(csa_tree_add_190_195_groupi_n_10250 ,csa_tree_add_190_195_groupi_n_10080 ,csa_tree_add_190_195_groupi_n_9576);
  or csa_tree_add_190_195_groupi_g38700(csa_tree_add_190_195_groupi_n_10249 ,csa_tree_add_190_195_groupi_n_9769 ,csa_tree_add_190_195_groupi_n_9948);
  and csa_tree_add_190_195_groupi_g38701(csa_tree_add_190_195_groupi_n_10248 ,csa_tree_add_190_195_groupi_n_9035 ,csa_tree_add_190_195_groupi_n_9978);
  or csa_tree_add_190_195_groupi_g38702(csa_tree_add_190_195_groupi_n_10247 ,csa_tree_add_190_195_groupi_n_9891 ,csa_tree_add_190_195_groupi_n_9885);
  nor csa_tree_add_190_195_groupi_g38703(csa_tree_add_190_195_groupi_n_10246 ,csa_tree_add_190_195_groupi_n_9892 ,csa_tree_add_190_195_groupi_n_9886);
  and csa_tree_add_190_195_groupi_g38704(csa_tree_add_190_195_groupi_n_10245 ,csa_tree_add_190_195_groupi_n_10042 ,csa_tree_add_190_195_groupi_n_9295);
  or csa_tree_add_190_195_groupi_g38705(csa_tree_add_190_195_groupi_n_10244 ,csa_tree_add_190_195_groupi_n_10042 ,csa_tree_add_190_195_groupi_n_9295);
  or csa_tree_add_190_195_groupi_g38706(csa_tree_add_190_195_groupi_n_10243 ,csa_tree_add_190_195_groupi_n_9758 ,csa_tree_add_190_195_groupi_n_9905);
  nor csa_tree_add_190_195_groupi_g38707(csa_tree_add_190_195_groupi_n_10242 ,csa_tree_add_190_195_groupi_n_9759 ,csa_tree_add_190_195_groupi_n_9904);
  or csa_tree_add_190_195_groupi_g38708(csa_tree_add_190_195_groupi_n_10241 ,csa_tree_add_190_195_groupi_n_9791 ,csa_tree_add_190_195_groupi_n_9973);
  and csa_tree_add_190_195_groupi_g38709(csa_tree_add_190_195_groupi_n_10240 ,csa_tree_add_190_195_groupi_n_9860 ,csa_tree_add_190_195_groupi_n_9952);
  or csa_tree_add_190_195_groupi_g38710(csa_tree_add_190_195_groupi_n_10239 ,csa_tree_add_190_195_groupi_n_9803 ,csa_tree_add_190_195_groupi_n_10001);
  nor csa_tree_add_190_195_groupi_g38711(csa_tree_add_190_195_groupi_n_10238 ,csa_tree_add_190_195_groupi_n_7590 ,csa_tree_add_190_195_groupi_n_9882);
  or csa_tree_add_190_195_groupi_g38712(csa_tree_add_190_195_groupi_n_10237 ,csa_tree_add_190_195_groupi_n_7591 ,csa_tree_add_190_195_groupi_n_9881);
  or csa_tree_add_190_195_groupi_g38713(csa_tree_add_190_195_groupi_n_10236 ,csa_tree_add_190_195_groupi_n_9860 ,csa_tree_add_190_195_groupi_n_9952);
  or csa_tree_add_190_195_groupi_g38714(csa_tree_add_190_195_groupi_n_10235 ,csa_tree_add_190_195_groupi_n_9677 ,csa_tree_add_190_195_groupi_n_9959);
  and csa_tree_add_190_195_groupi_g38715(csa_tree_add_190_195_groupi_n_10234 ,csa_tree_add_190_195_groupi_n_9477 ,csa_tree_add_190_195_groupi_n_9937);
  and csa_tree_add_190_195_groupi_g38716(csa_tree_add_190_195_groupi_n_10355 ,csa_tree_add_190_195_groupi_n_9731 ,csa_tree_add_190_195_groupi_n_10008);
  and csa_tree_add_190_195_groupi_g38717(csa_tree_add_190_195_groupi_n_10354 ,csa_tree_add_190_195_groupi_n_9680 ,csa_tree_add_190_195_groupi_n_9970);
  and csa_tree_add_190_195_groupi_g38718(csa_tree_add_190_195_groupi_n_10353 ,csa_tree_add_190_195_groupi_n_9686 ,csa_tree_add_190_195_groupi_n_9972);
  and csa_tree_add_190_195_groupi_g38719(csa_tree_add_190_195_groupi_n_10352 ,csa_tree_add_190_195_groupi_n_9700 ,csa_tree_add_190_195_groupi_n_9988);
  or csa_tree_add_190_195_groupi_g38720(csa_tree_add_190_195_groupi_n_10351 ,csa_tree_add_190_195_groupi_n_9704 ,csa_tree_add_190_195_groupi_n_9990);
  or csa_tree_add_190_195_groupi_g38721(csa_tree_add_190_195_groupi_n_10350 ,csa_tree_add_190_195_groupi_n_9703 ,csa_tree_add_190_195_groupi_n_9987);
  and csa_tree_add_190_195_groupi_g38722(csa_tree_add_190_195_groupi_n_10349 ,csa_tree_add_190_195_groupi_n_9693 ,csa_tree_add_190_195_groupi_n_9991);
  or csa_tree_add_190_195_groupi_g38723(csa_tree_add_190_195_groupi_n_10348 ,csa_tree_add_190_195_groupi_n_9707 ,csa_tree_add_190_195_groupi_n_9993);
  and csa_tree_add_190_195_groupi_g38724(csa_tree_add_190_195_groupi_n_10347 ,csa_tree_add_190_195_groupi_n_9720 ,csa_tree_add_190_195_groupi_n_10002);
  or csa_tree_add_190_195_groupi_g38725(csa_tree_add_190_195_groupi_n_10346 ,csa_tree_add_190_195_groupi_n_9722 ,csa_tree_add_190_195_groupi_n_10003);
  or csa_tree_add_190_195_groupi_g38726(csa_tree_add_190_195_groupi_n_10345 ,csa_tree_add_190_195_groupi_n_9589 ,csa_tree_add_190_195_groupi_n_10006);
  or csa_tree_add_190_195_groupi_g38727(csa_tree_add_190_195_groupi_n_10343 ,csa_tree_add_190_195_groupi_n_9682 ,csa_tree_add_190_195_groupi_n_9969);
  or csa_tree_add_190_195_groupi_g38728(csa_tree_add_190_195_groupi_n_10342 ,csa_tree_add_190_195_groupi_n_9733 ,csa_tree_add_190_195_groupi_n_10009);
  and csa_tree_add_190_195_groupi_g38729(csa_tree_add_190_195_groupi_n_10341 ,csa_tree_add_190_195_groupi_n_8312 ,csa_tree_add_190_195_groupi_n_10000);
  and csa_tree_add_190_195_groupi_g38730(csa_tree_add_190_195_groupi_n_10340 ,csa_tree_add_190_195_groupi_n_9136 ,csa_tree_add_190_195_groupi_n_10019);
  and csa_tree_add_190_195_groupi_g38731(csa_tree_add_190_195_groupi_n_10339 ,csa_tree_add_190_195_groupi_n_9698 ,csa_tree_add_190_195_groupi_n_10020);
  or csa_tree_add_190_195_groupi_g38732(csa_tree_add_190_195_groupi_n_10338 ,csa_tree_add_190_195_groupi_n_9600 ,csa_tree_add_190_195_groupi_n_10021);
  and csa_tree_add_190_195_groupi_g38733(csa_tree_add_190_195_groupi_n_10337 ,csa_tree_add_190_195_groupi_n_9745 ,csa_tree_add_190_195_groupi_n_10026);
  and csa_tree_add_190_195_groupi_g38734(csa_tree_add_190_195_groupi_n_10336 ,csa_tree_add_190_195_groupi_n_8802 ,csa_tree_add_190_195_groupi_n_10024);
  and csa_tree_add_190_195_groupi_g38735(csa_tree_add_190_195_groupi_n_10335 ,csa_tree_add_190_195_groupi_n_9454 ,csa_tree_add_190_195_groupi_n_10028);
  and csa_tree_add_190_195_groupi_g38736(csa_tree_add_190_195_groupi_n_10334 ,csa_tree_add_190_195_groupi_n_9578 ,csa_tree_add_190_195_groupi_n_9996);
  and csa_tree_add_190_195_groupi_g38737(csa_tree_add_190_195_groupi_n_10333 ,csa_tree_add_190_195_groupi_n_9458 ,csa_tree_add_190_195_groupi_n_10027);
  or csa_tree_add_190_195_groupi_g38738(csa_tree_add_190_195_groupi_n_10331 ,csa_tree_add_190_195_groupi_n_7688 ,csa_tree_add_190_195_groupi_n_9992);
  and csa_tree_add_190_195_groupi_g38739(csa_tree_add_190_195_groupi_n_10330 ,csa_tree_add_190_195_groupi_n_8097 ,csa_tree_add_190_195_groupi_n_10007);
  and csa_tree_add_190_195_groupi_g38740(csa_tree_add_190_195_groupi_n_10327 ,csa_tree_add_190_195_groupi_n_9675 ,csa_tree_add_190_195_groupi_n_9967);
  and csa_tree_add_190_195_groupi_g38741(csa_tree_add_190_195_groupi_n_10325 ,csa_tree_add_190_195_groupi_n_9138 ,csa_tree_add_190_195_groupi_n_10022);
  and csa_tree_add_190_195_groupi_g38742(csa_tree_add_190_195_groupi_n_10323 ,csa_tree_add_190_195_groupi_n_9594 ,csa_tree_add_190_195_groupi_n_10010);
  or csa_tree_add_190_195_groupi_g38743(csa_tree_add_190_195_groupi_n_10322 ,csa_tree_add_190_195_groupi_n_8742 ,csa_tree_add_190_195_groupi_n_9989);
  and csa_tree_add_190_195_groupi_g38744(csa_tree_add_190_195_groupi_n_10320 ,csa_tree_add_190_195_groupi_n_9670 ,csa_tree_add_190_195_groupi_n_9965);
  or csa_tree_add_190_195_groupi_g38745(csa_tree_add_190_195_groupi_n_10318 ,csa_tree_add_190_195_groupi_n_9418 ,csa_tree_add_190_195_groupi_n_10011);
  and csa_tree_add_190_195_groupi_g38746(csa_tree_add_190_195_groupi_n_10316 ,csa_tree_add_190_195_groupi_n_9283 ,csa_tree_add_190_195_groupi_n_9994);
  and csa_tree_add_190_195_groupi_g38747(csa_tree_add_190_195_groupi_n_10315 ,csa_tree_add_190_195_groupi_n_9749 ,csa_tree_add_190_195_groupi_n_10029);
  and csa_tree_add_190_195_groupi_g38748(csa_tree_add_190_195_groupi_n_10314 ,csa_tree_add_190_195_groupi_n_9582 ,csa_tree_add_190_195_groupi_n_9980);
  and csa_tree_add_190_195_groupi_g38749(csa_tree_add_190_195_groupi_n_10312 ,csa_tree_add_190_195_groupi_n_9740 ,csa_tree_add_190_195_groupi_n_10016);
  not csa_tree_add_190_195_groupi_g38750(csa_tree_add_190_195_groupi_n_10229 ,csa_tree_add_190_195_groupi_n_10228);
  not csa_tree_add_190_195_groupi_g38753(csa_tree_add_190_195_groupi_n_10222 ,csa_tree_add_190_195_groupi_n_10221);
  not csa_tree_add_190_195_groupi_g38754(csa_tree_add_190_195_groupi_n_10217 ,csa_tree_add_190_195_groupi_n_10216);
  not csa_tree_add_190_195_groupi_g38755(csa_tree_add_190_195_groupi_n_10213 ,csa_tree_add_190_195_groupi_n_10212);
  not csa_tree_add_190_195_groupi_g38756(csa_tree_add_190_195_groupi_n_10211 ,csa_tree_add_190_195_groupi_n_10210);
  not csa_tree_add_190_195_groupi_g38757(csa_tree_add_190_195_groupi_n_10209 ,csa_tree_add_190_195_groupi_n_127);
  not csa_tree_add_190_195_groupi_g38758(csa_tree_add_190_195_groupi_n_10208 ,csa_tree_add_190_195_groupi_n_10207);
  not csa_tree_add_190_195_groupi_g38759(csa_tree_add_190_195_groupi_n_10206 ,csa_tree_add_190_195_groupi_n_10205);
  not csa_tree_add_190_195_groupi_g38760(csa_tree_add_190_195_groupi_n_10204 ,csa_tree_add_190_195_groupi_n_10203);
  not csa_tree_add_190_195_groupi_g38761(csa_tree_add_190_195_groupi_n_10202 ,csa_tree_add_190_195_groupi_n_10201);
  not csa_tree_add_190_195_groupi_g38762(csa_tree_add_190_195_groupi_n_10200 ,csa_tree_add_190_195_groupi_n_10199);
  not csa_tree_add_190_195_groupi_g38763(csa_tree_add_190_195_groupi_n_10198 ,csa_tree_add_190_195_groupi_n_10197);
  not csa_tree_add_190_195_groupi_g38764(csa_tree_add_190_195_groupi_n_10196 ,csa_tree_add_190_195_groupi_n_10195);
  not csa_tree_add_190_195_groupi_g38765(csa_tree_add_190_195_groupi_n_10194 ,csa_tree_add_190_195_groupi_n_10193);
  not csa_tree_add_190_195_groupi_g38766(csa_tree_add_190_195_groupi_n_10192 ,csa_tree_add_190_195_groupi_n_10191);
  not csa_tree_add_190_195_groupi_g38767(csa_tree_add_190_195_groupi_n_10190 ,csa_tree_add_190_195_groupi_n_10189);
  not csa_tree_add_190_195_groupi_g38768(csa_tree_add_190_195_groupi_n_10188 ,csa_tree_add_190_195_groupi_n_10187);
  not csa_tree_add_190_195_groupi_g38769(csa_tree_add_190_195_groupi_n_10186 ,csa_tree_add_190_195_groupi_n_10185);
  not csa_tree_add_190_195_groupi_g38770(csa_tree_add_190_195_groupi_n_10184 ,csa_tree_add_190_195_groupi_n_10183);
  not csa_tree_add_190_195_groupi_g38771(csa_tree_add_190_195_groupi_n_10182 ,csa_tree_add_190_195_groupi_n_10181);
  not csa_tree_add_190_195_groupi_g38772(csa_tree_add_190_195_groupi_n_10180 ,csa_tree_add_190_195_groupi_n_10179);
  not csa_tree_add_190_195_groupi_g38773(csa_tree_add_190_195_groupi_n_10178 ,csa_tree_add_190_195_groupi_n_10177);
  not csa_tree_add_190_195_groupi_g38774(csa_tree_add_190_195_groupi_n_10176 ,csa_tree_add_190_195_groupi_n_10175);
  not csa_tree_add_190_195_groupi_g38775(csa_tree_add_190_195_groupi_n_10174 ,csa_tree_add_190_195_groupi_n_10173);
  not csa_tree_add_190_195_groupi_g38776(csa_tree_add_190_195_groupi_n_10172 ,csa_tree_add_190_195_groupi_n_10171);
  not csa_tree_add_190_195_groupi_g38777(csa_tree_add_190_195_groupi_n_10169 ,csa_tree_add_190_195_groupi_n_10168);
  not csa_tree_add_190_195_groupi_g38778(csa_tree_add_190_195_groupi_n_10167 ,csa_tree_add_190_195_groupi_n_10166);
  not csa_tree_add_190_195_groupi_g38779(csa_tree_add_190_195_groupi_n_10165 ,csa_tree_add_190_195_groupi_n_10164);
  not csa_tree_add_190_195_groupi_g38780(csa_tree_add_190_195_groupi_n_10163 ,csa_tree_add_190_195_groupi_n_10162);
  not csa_tree_add_190_195_groupi_g38781(csa_tree_add_190_195_groupi_n_10161 ,csa_tree_add_190_195_groupi_n_10160);
  not csa_tree_add_190_195_groupi_g38782(csa_tree_add_190_195_groupi_n_10159 ,csa_tree_add_190_195_groupi_n_10158);
  not csa_tree_add_190_195_groupi_g38783(csa_tree_add_190_195_groupi_n_10157 ,csa_tree_add_190_195_groupi_n_10156);
  not csa_tree_add_190_195_groupi_g38784(csa_tree_add_190_195_groupi_n_10155 ,csa_tree_add_190_195_groupi_n_10154);
  not csa_tree_add_190_195_groupi_g38785(csa_tree_add_190_195_groupi_n_10151 ,csa_tree_add_190_195_groupi_n_10150);
  not csa_tree_add_190_195_groupi_g38786(csa_tree_add_190_195_groupi_n_10149 ,csa_tree_add_190_195_groupi_n_10148);
  not csa_tree_add_190_195_groupi_g38787(csa_tree_add_190_195_groupi_n_10147 ,csa_tree_add_190_195_groupi_n_10146);
  or csa_tree_add_190_195_groupi_g38788(csa_tree_add_190_195_groupi_n_10145 ,csa_tree_add_190_195_groupi_n_9797 ,csa_tree_add_190_195_groupi_n_10017);
  and csa_tree_add_190_195_groupi_g38789(csa_tree_add_190_195_groupi_n_10144 ,csa_tree_add_190_195_groupi_n_9790 ,csa_tree_add_190_195_groupi_n_9842);
  and csa_tree_add_190_195_groupi_g38790(csa_tree_add_190_195_groupi_n_10143 ,csa_tree_add_190_195_groupi_n_8617 ,csa_tree_add_190_195_groupi_n_10062);
  or csa_tree_add_190_195_groupi_g38791(csa_tree_add_190_195_groupi_n_10142 ,csa_tree_add_190_195_groupi_n_9622 ,csa_tree_add_190_195_groupi_n_10050);
  nor csa_tree_add_190_195_groupi_g38792(csa_tree_add_190_195_groupi_n_10141 ,csa_tree_add_190_195_groupi_n_9621 ,csa_tree_add_190_195_groupi_n_10051);
  or csa_tree_add_190_195_groupi_g38793(csa_tree_add_190_195_groupi_n_10140 ,csa_tree_add_190_195_groupi_n_9504 ,csa_tree_add_190_195_groupi_n_9858);
  or csa_tree_add_190_195_groupi_g38794(csa_tree_add_190_195_groupi_n_10139 ,csa_tree_add_190_195_groupi_n_9925 ,csa_tree_add_190_195_groupi_n_9924);
  and csa_tree_add_190_195_groupi_g38795(csa_tree_add_190_195_groupi_n_10138 ,csa_tree_add_190_195_groupi_n_9639 ,csa_tree_add_190_195_groupi_n_9920);
  nor csa_tree_add_190_195_groupi_g38796(csa_tree_add_190_195_groupi_n_10137 ,csa_tree_add_190_195_groupi_n_9639 ,csa_tree_add_190_195_groupi_n_9920);
  or csa_tree_add_190_195_groupi_g38797(csa_tree_add_190_195_groupi_n_10136 ,csa_tree_add_190_195_groupi_n_9355 ,csa_tree_add_190_195_groupi_n_9854);
  or csa_tree_add_190_195_groupi_g38798(csa_tree_add_190_195_groupi_n_10135 ,csa_tree_add_190_195_groupi_n_9494 ,csa_tree_add_190_195_groupi_n_9902);
  or csa_tree_add_190_195_groupi_g38799(csa_tree_add_190_195_groupi_n_10134 ,csa_tree_add_190_195_groupi_n_9909 ,csa_tree_add_190_195_groupi_n_9906);
  nor csa_tree_add_190_195_groupi_g38800(csa_tree_add_190_195_groupi_n_10133 ,csa_tree_add_190_195_groupi_n_9908 ,csa_tree_add_190_195_groupi_n_9907);
  or csa_tree_add_190_195_groupi_g38801(csa_tree_add_190_195_groupi_n_10132 ,csa_tree_add_190_195_groupi_n_9901 ,csa_tree_add_190_195_groupi_n_8998);
  nor csa_tree_add_190_195_groupi_g38802(csa_tree_add_190_195_groupi_n_10131 ,csa_tree_add_190_195_groupi_n_9900 ,csa_tree_add_190_195_groupi_n_8999);
  nor csa_tree_add_190_195_groupi_g38803(csa_tree_add_190_195_groupi_n_10130 ,csa_tree_add_190_195_groupi_n_9493 ,csa_tree_add_190_195_groupi_n_9903);
  or csa_tree_add_190_195_groupi_g38804(csa_tree_add_190_195_groupi_n_10129 ,csa_tree_add_190_195_groupi_n_9941 ,csa_tree_add_190_195_groupi_n_9938);
  or csa_tree_add_190_195_groupi_g38805(csa_tree_add_190_195_groupi_n_10128 ,csa_tree_add_190_195_groupi_n_9889 ,csa_tree_add_190_195_groupi_n_9950);
  nor csa_tree_add_190_195_groupi_g38806(csa_tree_add_190_195_groupi_n_10127 ,csa_tree_add_190_195_groupi_n_9890 ,csa_tree_add_190_195_groupi_n_9951);
  nor csa_tree_add_190_195_groupi_g38807(csa_tree_add_190_195_groupi_n_10126 ,csa_tree_add_190_195_groupi_n_9895 ,csa_tree_add_190_195_groupi_n_10058);
  or csa_tree_add_190_195_groupi_g38808(csa_tree_add_190_195_groupi_n_10125 ,csa_tree_add_190_195_groupi_n_9502 ,csa_tree_add_190_195_groupi_n_9922);
  or csa_tree_add_190_195_groupi_g38809(csa_tree_add_190_195_groupi_n_10124 ,csa_tree_add_190_195_groupi_n_9896 ,csa_tree_add_190_195_groupi_n_10057);
  or csa_tree_add_190_195_groupi_g38810(csa_tree_add_190_195_groupi_n_10123 ,csa_tree_add_190_195_groupi_n_9619 ,csa_tree_add_190_195_groupi_n_10053);
  nor csa_tree_add_190_195_groupi_g38811(csa_tree_add_190_195_groupi_n_10122 ,csa_tree_add_190_195_groupi_n_9503 ,csa_tree_add_190_195_groupi_n_9921);
  nor csa_tree_add_190_195_groupi_g38812(csa_tree_add_190_195_groupi_n_10121 ,csa_tree_add_190_195_groupi_n_9618 ,csa_tree_add_190_195_groupi_n_10054);
  or csa_tree_add_190_195_groupi_g38813(csa_tree_add_190_195_groupi_n_10120 ,csa_tree_add_190_195_groupi_n_9873 ,csa_tree_add_190_195_groupi_n_10048);
  or csa_tree_add_190_195_groupi_g38814(csa_tree_add_190_195_groupi_n_10119 ,csa_tree_add_190_195_groupi_n_9477 ,csa_tree_add_190_195_groupi_n_9937);
  or csa_tree_add_190_195_groupi_g38815(csa_tree_add_190_195_groupi_n_10118 ,csa_tree_add_190_195_groupi_n_9845 ,csa_tree_add_190_195_groupi_n_10081);
  nor csa_tree_add_190_195_groupi_g38816(csa_tree_add_190_195_groupi_n_10117 ,csa_tree_add_190_195_groupi_n_9872 ,csa_tree_add_190_195_groupi_n_10049);
  xnor csa_tree_add_190_195_groupi_g38817(out1[1] ,csa_tree_add_190_195_groupi_n_8501 ,csa_tree_add_190_195_groupi_n_9535);
  nor csa_tree_add_190_195_groupi_g38818(csa_tree_add_190_195_groupi_n_10115 ,csa_tree_add_190_195_groupi_n_9203 ,csa_tree_add_190_195_groupi_n_9859);
  nor csa_tree_add_190_195_groupi_g38819(csa_tree_add_190_195_groupi_n_10114 ,csa_tree_add_190_195_groupi_n_9940 ,csa_tree_add_190_195_groupi_n_9939);
  xnor csa_tree_add_190_195_groupi_g38821(csa_tree_add_190_195_groupi_n_10113 ,csa_tree_add_190_195_groupi_n_7072 ,csa_tree_add_190_195_groupi_n_9643);
  xnor csa_tree_add_190_195_groupi_g38822(csa_tree_add_190_195_groupi_n_10112 ,csa_tree_add_190_195_groupi_n_8992 ,csa_tree_add_190_195_groupi_n_9763);
  xnor csa_tree_add_190_195_groupi_g38823(csa_tree_add_190_195_groupi_n_10111 ,csa_tree_add_190_195_groupi_n_9784 ,csa_tree_add_190_195_groupi_n_9636);
  xnor csa_tree_add_190_195_groupi_g38824(csa_tree_add_190_195_groupi_n_10110 ,csa_tree_add_190_195_groupi_n_9606 ,csa_tree_add_190_195_groupi_n_9340);
  xnor csa_tree_add_190_195_groupi_g38825(csa_tree_add_190_195_groupi_n_10109 ,csa_tree_add_190_195_groupi_n_9160 ,csa_tree_add_190_195_groupi_n_9647);
  xnor csa_tree_add_190_195_groupi_g38826(csa_tree_add_190_195_groupi_n_10108 ,csa_tree_add_190_195_groupi_n_9473 ,csa_tree_add_190_195_groupi_n_9649);
  xnor csa_tree_add_190_195_groupi_g38827(csa_tree_add_190_195_groupi_n_10107 ,csa_tree_add_190_195_groupi_n_9342 ,csa_tree_add_190_195_groupi_n_9641);
  xnor csa_tree_add_190_195_groupi_g38828(csa_tree_add_190_195_groupi_n_10106 ,csa_tree_add_190_195_groupi_n_8627 ,csa_tree_add_190_195_groupi_n_9669);
  xnor csa_tree_add_190_195_groupi_g38829(csa_tree_add_190_195_groupi_n_10105 ,csa_tree_add_190_195_groupi_n_9751 ,csa_tree_add_190_195_groupi_n_8666);
  xnor csa_tree_add_190_195_groupi_g38830(csa_tree_add_190_195_groupi_n_10104 ,csa_tree_add_190_195_groupi_n_7574 ,csa_tree_add_190_195_groupi_n_9804);
  xnor csa_tree_add_190_195_groupi_g38831(csa_tree_add_190_195_groupi_n_10103 ,csa_tree_add_190_195_groupi_n_8966 ,csa_tree_add_190_195_groupi_n_9786);
  xnor csa_tree_add_190_195_groupi_g38832(csa_tree_add_190_195_groupi_n_10102 ,csa_tree_add_190_195_groupi_n_9791 ,csa_tree_add_190_195_groupi_n_9624);
  xnor csa_tree_add_190_195_groupi_g38833(csa_tree_add_190_195_groupi_n_10101 ,csa_tree_add_190_195_groupi_n_9645 ,csa_tree_add_190_195_groupi_n_9310);
  xnor csa_tree_add_190_195_groupi_g38834(csa_tree_add_190_195_groupi_n_10100 ,csa_tree_add_190_195_groupi_n_9777 ,csa_tree_add_190_195_groupi_n_9656);
  xnor csa_tree_add_190_195_groupi_g38835(csa_tree_add_190_195_groupi_n_10099 ,csa_tree_add_190_195_groupi_n_9602 ,csa_tree_add_190_195_groupi_n_9307);
  xnor csa_tree_add_190_195_groupi_g38836(csa_tree_add_190_195_groupi_n_10098 ,csa_tree_add_190_195_groupi_n_9753 ,csa_tree_add_190_195_groupi_n_9329);
  xnor csa_tree_add_190_195_groupi_g38837(csa_tree_add_190_195_groupi_n_10097 ,csa_tree_add_190_195_groupi_n_9617 ,csa_tree_add_190_195_groupi_n_9803);
  xnor csa_tree_add_190_195_groupi_g38838(csa_tree_add_190_195_groupi_n_10096 ,csa_tree_add_190_195_groupi_n_7497 ,csa_tree_add_190_195_groupi_n_9801);
  xnor csa_tree_add_190_195_groupi_g38839(csa_tree_add_190_195_groupi_n_10095 ,csa_tree_add_190_195_groupi_n_9755 ,csa_tree_add_190_195_groupi_n_9780);
  xnor csa_tree_add_190_195_groupi_g38840(csa_tree_add_190_195_groupi_n_10094 ,csa_tree_add_190_195_groupi_n_9607 ,csa_tree_add_190_195_groupi_n_9666);
  xnor csa_tree_add_190_195_groupi_g38842(csa_tree_add_190_195_groupi_n_10093 ,csa_tree_add_190_195_groupi_n_9338 ,csa_tree_add_190_195_groupi_n_9613);
  xnor csa_tree_add_190_195_groupi_g38843(csa_tree_add_190_195_groupi_n_10092 ,csa_tree_add_190_195_groupi_n_9794 ,csa_tree_add_190_195_groupi_n_9639);
  xnor csa_tree_add_190_195_groupi_g38844(csa_tree_add_190_195_groupi_n_10091 ,csa_tree_add_190_195_groupi_n_8197 ,csa_tree_add_190_195_groupi_n_9810);
  xnor csa_tree_add_190_195_groupi_g38845(csa_tree_add_190_195_groupi_n_10090 ,csa_tree_add_190_195_groupi_n_9203 ,csa_tree_add_190_195_groupi_n_9626);
  xnor csa_tree_add_190_195_groupi_g38846(csa_tree_add_190_195_groupi_n_10089 ,csa_tree_add_190_195_groupi_n_9795 ,csa_tree_add_190_195_groupi_n_9615);
  xnor csa_tree_add_190_195_groupi_g38847(csa_tree_add_190_195_groupi_n_10088 ,csa_tree_add_190_195_groupi_n_9651 ,csa_tree_add_190_195_groupi_n_7632);
  and csa_tree_add_190_195_groupi_g38848(csa_tree_add_190_195_groupi_n_10233 ,csa_tree_add_190_195_groupi_n_9580 ,csa_tree_add_190_195_groupi_n_9850);
  xnor csa_tree_add_190_195_groupi_g38849(csa_tree_add_190_195_groupi_n_10232 ,csa_tree_add_190_195_groupi_n_8377 ,csa_tree_add_190_195_groupi_n_9551);
  xnor csa_tree_add_190_195_groupi_g38850(csa_tree_add_190_195_groupi_n_10231 ,csa_tree_add_190_195_groupi_n_9316 ,csa_tree_add_190_195_groupi_n_9540);
  xnor csa_tree_add_190_195_groupi_g38851(csa_tree_add_190_195_groupi_n_10230 ,csa_tree_add_190_195_groupi_n_9657 ,csa_tree_add_190_195_groupi_n_9229);
  xnor csa_tree_add_190_195_groupi_g38852(csa_tree_add_190_195_groupi_n_10228 ,csa_tree_add_190_195_groupi_n_8876 ,csa_tree_add_190_195_groupi_n_9558);
  xnor csa_tree_add_190_195_groupi_g38853(csa_tree_add_190_195_groupi_n_10227 ,csa_tree_add_190_195_groupi_n_9336 ,csa_tree_add_190_195_groupi_n_9536);
  xnor csa_tree_add_190_195_groupi_g38854(csa_tree_add_190_195_groupi_n_10226 ,csa_tree_add_190_195_groupi_n_8211 ,csa_tree_add_190_195_groupi_n_9537);
  xnor csa_tree_add_190_195_groupi_g38855(csa_tree_add_190_195_groupi_n_10225 ,csa_tree_add_190_195_groupi_n_5333 ,csa_tree_add_190_195_groupi_n_9564);
  xnor csa_tree_add_190_195_groupi_g38856(csa_tree_add_190_195_groupi_n_10224 ,csa_tree_add_190_195_groupi_n_6760 ,csa_tree_add_190_195_groupi_n_9533);
  xnor csa_tree_add_190_195_groupi_g38857(csa_tree_add_190_195_groupi_n_10223 ,csa_tree_add_190_195_groupi_n_5433 ,csa_tree_add_190_195_groupi_n_9528);
  or csa_tree_add_190_195_groupi_g38858(csa_tree_add_190_195_groupi_n_10221 ,csa_tree_add_190_195_groupi_n_9574 ,csa_tree_add_190_195_groupi_n_9849);
  xnor csa_tree_add_190_195_groupi_g38859(csa_tree_add_190_195_groupi_n_10220 ,csa_tree_add_190_195_groupi_n_7596 ,csa_tree_add_190_195_groupi_n_9569);
  xnor csa_tree_add_190_195_groupi_g38860(csa_tree_add_190_195_groupi_n_10219 ,csa_tree_add_190_195_groupi_n_8201 ,csa_tree_add_190_195_groupi_n_9559);
  xnor csa_tree_add_190_195_groupi_g38861(csa_tree_add_190_195_groupi_n_10218 ,csa_tree_add_190_195_groupi_n_7083 ,csa_tree_add_190_195_groupi_n_9568);
  xnor csa_tree_add_190_195_groupi_g38862(csa_tree_add_190_195_groupi_n_10216 ,csa_tree_add_190_195_groupi_n_9194 ,csa_tree_add_190_195_groupi_n_9561);
  xnor csa_tree_add_190_195_groupi_g38863(csa_tree_add_190_195_groupi_n_10215 ,csa_tree_add_190_195_groupi_n_9175 ,csa_tree_add_190_195_groupi_n_9560);
  xnor csa_tree_add_190_195_groupi_g38864(csa_tree_add_190_195_groupi_n_10214 ,csa_tree_add_190_195_groupi_n_7626 ,csa_tree_add_190_195_groupi_n_125);
  xnor csa_tree_add_190_195_groupi_g38865(csa_tree_add_190_195_groupi_n_10212 ,csa_tree_add_190_195_groupi_n_8713 ,csa_tree_add_190_195_groupi_n_9529);
  xnor csa_tree_add_190_195_groupi_g38866(csa_tree_add_190_195_groupi_n_10210 ,csa_tree_add_190_195_groupi_n_9808 ,csa_tree_add_190_195_groupi_n_9557);
  xnor csa_tree_add_190_195_groupi_g38868(csa_tree_add_190_195_groupi_n_10207 ,csa_tree_add_190_195_groupi_n_9659 ,csa_tree_add_190_195_groupi_n_9545);
  xnor csa_tree_add_190_195_groupi_g38869(csa_tree_add_190_195_groupi_n_10205 ,csa_tree_add_190_195_groupi_n_9527 ,csa_tree_add_190_195_groupi_n_9544);
  xnor csa_tree_add_190_195_groupi_g38870(csa_tree_add_190_195_groupi_n_10203 ,csa_tree_add_190_195_groupi_n_8699 ,csa_tree_add_190_195_groupi_n_9566);
  xnor csa_tree_add_190_195_groupi_g38871(csa_tree_add_190_195_groupi_n_10201 ,csa_tree_add_190_195_groupi_n_7601 ,csa_tree_add_190_195_groupi_n_124);
  xnor csa_tree_add_190_195_groupi_g38872(csa_tree_add_190_195_groupi_n_10199 ,csa_tree_add_190_195_groupi_n_9327 ,csa_tree_add_190_195_groupi_n_9567);
  xnor csa_tree_add_190_195_groupi_g38873(csa_tree_add_190_195_groupi_n_10197 ,csa_tree_add_190_195_groupi_n_8391 ,csa_tree_add_190_195_groupi_n_9565);
  xnor csa_tree_add_190_195_groupi_g38874(csa_tree_add_190_195_groupi_n_10195 ,csa_tree_add_190_195_groupi_n_9043 ,csa_tree_add_190_195_groupi_n_9555);
  xnor csa_tree_add_190_195_groupi_g38875(csa_tree_add_190_195_groupi_n_10193 ,csa_tree_add_190_195_groupi_n_9792 ,csa_tree_add_190_195_groupi_n_8896);
  xnor csa_tree_add_190_195_groupi_g38876(csa_tree_add_190_195_groupi_n_10191 ,csa_tree_add_190_195_groupi_n_9663 ,csa_tree_add_190_195_groupi_n_9223);
  xnor csa_tree_add_190_195_groupi_g38877(csa_tree_add_190_195_groupi_n_10189 ,csa_tree_add_190_195_groupi_n_8853 ,csa_tree_add_190_195_groupi_n_9543);
  xnor csa_tree_add_190_195_groupi_g38878(csa_tree_add_190_195_groupi_n_10187 ,csa_tree_add_190_195_groupi_n_8679 ,csa_tree_add_190_195_groupi_n_9542);
  xnor csa_tree_add_190_195_groupi_g38879(csa_tree_add_190_195_groupi_n_10185 ,csa_tree_add_190_195_groupi_n_7097 ,csa_tree_add_190_195_groupi_n_9563);
  xnor csa_tree_add_190_195_groupi_g38880(csa_tree_add_190_195_groupi_n_10183 ,csa_tree_add_190_195_groupi_n_8369 ,csa_tree_add_190_195_groupi_n_9553);
  xnor csa_tree_add_190_195_groupi_g38881(csa_tree_add_190_195_groupi_n_10181 ,csa_tree_add_190_195_groupi_n_8032 ,csa_tree_add_190_195_groupi_n_9552);
  xnor csa_tree_add_190_195_groupi_g38882(csa_tree_add_190_195_groupi_n_10179 ,csa_tree_add_190_195_groupi_n_6960 ,csa_tree_add_190_195_groupi_n_9554);
  xnor csa_tree_add_190_195_groupi_g38883(csa_tree_add_190_195_groupi_n_10177 ,csa_tree_add_190_195_groupi_n_8704 ,csa_tree_add_190_195_groupi_n_9541);
  xnor csa_tree_add_190_195_groupi_g38884(csa_tree_add_190_195_groupi_n_10175 ,csa_tree_add_190_195_groupi_n_9785 ,csa_tree_add_190_195_groupi_n_7887);
  xnor csa_tree_add_190_195_groupi_g38885(csa_tree_add_190_195_groupi_n_10173 ,csa_tree_add_190_195_groupi_n_8822 ,csa_tree_add_190_195_groupi_n_9556);
  xnor csa_tree_add_190_195_groupi_g38886(csa_tree_add_190_195_groupi_n_10171 ,csa_tree_add_190_195_groupi_n_8848 ,csa_tree_add_190_195_groupi_n_9539);
  xnor csa_tree_add_190_195_groupi_g38887(csa_tree_add_190_195_groupi_n_10170 ,csa_tree_add_190_195_groupi_n_9665 ,csa_tree_add_190_195_groupi_n_8894);
  xnor csa_tree_add_190_195_groupi_g38888(csa_tree_add_190_195_groupi_n_10168 ,csa_tree_add_190_195_groupi_n_9524 ,csa_tree_add_190_195_groupi_n_9538);
  xnor csa_tree_add_190_195_groupi_g38889(csa_tree_add_190_195_groupi_n_10166 ,csa_tree_add_190_195_groupi_n_8025 ,csa_tree_add_190_195_groupi_n_9562);
  xnor csa_tree_add_190_195_groupi_g38890(csa_tree_add_190_195_groupi_n_10164 ,csa_tree_add_190_195_groupi_n_9788 ,csa_tree_add_190_195_groupi_n_9550);
  xnor csa_tree_add_190_195_groupi_g38891(csa_tree_add_190_195_groupi_n_10162 ,csa_tree_add_190_195_groupi_n_9171 ,csa_tree_add_190_195_groupi_n_128);
  xnor csa_tree_add_190_195_groupi_g38892(csa_tree_add_190_195_groupi_n_10160 ,csa_tree_add_190_195_groupi_n_9352 ,csa_tree_add_190_195_groupi_n_9534);
  xnor csa_tree_add_190_195_groupi_g38893(csa_tree_add_190_195_groupi_n_10158 ,csa_tree_add_190_195_groupi_n_8835 ,csa_tree_add_190_195_groupi_n_9549);
  and csa_tree_add_190_195_groupi_g38894(csa_tree_add_190_195_groupi_n_10156 ,csa_tree_add_190_195_groupi_n_9265 ,csa_tree_add_190_195_groupi_n_9853);
  xnor csa_tree_add_190_195_groupi_g38895(csa_tree_add_190_195_groupi_n_10154 ,csa_tree_add_190_195_groupi_n_7614 ,csa_tree_add_190_195_groupi_n_9532);
  xnor csa_tree_add_190_195_groupi_g38896(csa_tree_add_190_195_groupi_n_10153 ,csa_tree_add_190_195_groupi_n_7582 ,csa_tree_add_190_195_groupi_n_9531);
  xnor csa_tree_add_190_195_groupi_g38897(csa_tree_add_190_195_groupi_n_10152 ,csa_tree_add_190_195_groupi_n_9330 ,csa_tree_add_190_195_groupi_n_9530);
  xnor csa_tree_add_190_195_groupi_g38898(csa_tree_add_190_195_groupi_n_10150 ,csa_tree_add_190_195_groupi_n_7569 ,csa_tree_add_190_195_groupi_n_9548);
  xnor csa_tree_add_190_195_groupi_g38899(csa_tree_add_190_195_groupi_n_10148 ,csa_tree_add_190_195_groupi_n_9654 ,csa_tree_add_190_195_groupi_n_9547);
  xnor csa_tree_add_190_195_groupi_g38900(csa_tree_add_190_195_groupi_n_10146 ,csa_tree_add_190_195_groupi_n_8372 ,csa_tree_add_190_195_groupi_n_126);
  not csa_tree_add_190_195_groupi_g38909(csa_tree_add_190_195_groupi_n_10064 ,csa_tree_add_190_195_groupi_n_10063);
  not csa_tree_add_190_195_groupi_g38910(csa_tree_add_190_195_groupi_n_10062 ,csa_tree_add_190_195_groupi_n_10061);
  not csa_tree_add_190_195_groupi_g38911(csa_tree_add_190_195_groupi_n_10059 ,csa_tree_add_190_195_groupi_n_10060);
  not csa_tree_add_190_195_groupi_g38912(csa_tree_add_190_195_groupi_n_10058 ,csa_tree_add_190_195_groupi_n_10057);
  not csa_tree_add_190_195_groupi_g38913(csa_tree_add_190_195_groupi_n_10056 ,csa_tree_add_190_195_groupi_n_10055);
  not csa_tree_add_190_195_groupi_g38914(csa_tree_add_190_195_groupi_n_10054 ,csa_tree_add_190_195_groupi_n_10053);
  not csa_tree_add_190_195_groupi_g38915(csa_tree_add_190_195_groupi_n_10051 ,csa_tree_add_190_195_groupi_n_10050);
  not csa_tree_add_190_195_groupi_g38916(csa_tree_add_190_195_groupi_n_10049 ,csa_tree_add_190_195_groupi_n_10048);
  not csa_tree_add_190_195_groupi_g38917(csa_tree_add_190_195_groupi_n_10045 ,csa_tree_add_190_195_groupi_n_10046);
  not csa_tree_add_190_195_groupi_g38918(csa_tree_add_190_195_groupi_n_10043 ,csa_tree_add_190_195_groupi_n_10044);
  not csa_tree_add_190_195_groupi_g38919(csa_tree_add_190_195_groupi_n_10040 ,csa_tree_add_190_195_groupi_n_10041);
  not csa_tree_add_190_195_groupi_g38920(csa_tree_add_190_195_groupi_n_10039 ,csa_tree_add_190_195_groupi_n_10038);
  not csa_tree_add_190_195_groupi_g38921(csa_tree_add_190_195_groupi_n_10037 ,csa_tree_add_190_195_groupi_n_10036);
  not csa_tree_add_190_195_groupi_g38922(csa_tree_add_190_195_groupi_n_10034 ,csa_tree_add_190_195_groupi_n_10035);
  or csa_tree_add_190_195_groupi_g38923(csa_tree_add_190_195_groupi_n_10033 ,csa_tree_add_190_195_groupi_n_9473 ,csa_tree_add_190_195_groupi_n_9648);
  nor csa_tree_add_190_195_groupi_g38924(csa_tree_add_190_195_groupi_n_10032 ,csa_tree_add_190_195_groupi_n_9338 ,csa_tree_add_190_195_groupi_n_9612);
  nor csa_tree_add_190_195_groupi_g38925(csa_tree_add_190_195_groupi_n_10031 ,csa_tree_add_190_195_groupi_n_9472 ,csa_tree_add_190_195_groupi_n_9649);
  and csa_tree_add_190_195_groupi_g38926(csa_tree_add_190_195_groupi_n_10030 ,csa_tree_add_190_195_groupi_n_8321 ,csa_tree_add_190_195_groupi_n_9626);
  or csa_tree_add_190_195_groupi_g38927(csa_tree_add_190_195_groupi_n_10029 ,csa_tree_add_190_195_groupi_n_9805 ,csa_tree_add_190_195_groupi_n_9748);
  or csa_tree_add_190_195_groupi_g38928(csa_tree_add_190_195_groupi_n_10028 ,csa_tree_add_190_195_groupi_n_9452 ,csa_tree_add_190_195_groupi_n_9809);
  or csa_tree_add_190_195_groupi_g38929(csa_tree_add_190_195_groupi_n_10027 ,csa_tree_add_190_195_groupi_n_9450 ,csa_tree_add_190_195_groupi_n_9654);
  or csa_tree_add_190_195_groupi_g38930(csa_tree_add_190_195_groupi_n_10026 ,csa_tree_add_190_195_groupi_n_8871 ,csa_tree_add_190_195_groupi_n_9744);
  nor csa_tree_add_190_195_groupi_g38931(csa_tree_add_190_195_groupi_n_10025 ,csa_tree_add_190_195_groupi_n_7546 ,csa_tree_add_190_195_groupi_n_9607);
  or csa_tree_add_190_195_groupi_g38932(csa_tree_add_190_195_groupi_n_10024 ,csa_tree_add_190_195_groupi_n_8797 ,csa_tree_add_190_195_groupi_n_9792);
  and csa_tree_add_190_195_groupi_g38933(csa_tree_add_190_195_groupi_n_10023 ,csa_tree_add_190_195_groupi_n_7546 ,csa_tree_add_190_195_groupi_n_9607);
  or csa_tree_add_190_195_groupi_g38934(csa_tree_add_190_195_groupi_n_10022 ,csa_tree_add_190_195_groupi_n_9137 ,csa_tree_add_190_195_groupi_n_9664);
  and csa_tree_add_190_195_groupi_g38935(csa_tree_add_190_195_groupi_n_10021 ,csa_tree_add_190_195_groupi_n_9599 ,csa_tree_add_190_195_groupi_n_9518);
  or csa_tree_add_190_195_groupi_g38936(csa_tree_add_190_195_groupi_n_10020 ,csa_tree_add_190_195_groupi_n_9362 ,csa_tree_add_190_195_groupi_n_9697);
  or csa_tree_add_190_195_groupi_g38937(csa_tree_add_190_195_groupi_n_10019 ,csa_tree_add_190_195_groupi_n_9134 ,csa_tree_add_190_195_groupi_n_9657);
  or csa_tree_add_190_195_groupi_g38938(csa_tree_add_190_195_groupi_n_10018 ,csa_tree_add_190_195_groupi_n_9605 ,csa_tree_add_190_195_groupi_n_9340);
  nor csa_tree_add_190_195_groupi_g38939(csa_tree_add_190_195_groupi_n_10017 ,csa_tree_add_190_195_groupi_n_9341 ,csa_tree_add_190_195_groupi_n_9641);
  or csa_tree_add_190_195_groupi_g38940(csa_tree_add_190_195_groupi_n_10016 ,csa_tree_add_190_195_groupi_n_9354 ,csa_tree_add_190_195_groupi_n_9739);
  nor csa_tree_add_190_195_groupi_g38941(csa_tree_add_190_195_groupi_n_10015 ,csa_tree_add_190_195_groupi_n_9752 ,csa_tree_add_190_195_groupi_n_9329);
  and csa_tree_add_190_195_groupi_g38942(csa_tree_add_190_195_groupi_n_10014 ,csa_tree_add_190_195_groupi_n_9755 ,csa_tree_add_190_195_groupi_n_9780);
  nor csa_tree_add_190_195_groupi_g38943(csa_tree_add_190_195_groupi_n_10013 ,csa_tree_add_190_195_groupi_n_9755 ,csa_tree_add_190_195_groupi_n_9780);
  or csa_tree_add_190_195_groupi_g38944(csa_tree_add_190_195_groupi_n_10012 ,csa_tree_add_190_195_groupi_n_9753 ,csa_tree_add_190_195_groupi_n_9328);
  nor csa_tree_add_190_195_groupi_g38945(csa_tree_add_190_195_groupi_n_10011 ,csa_tree_add_190_195_groupi_n_9416 ,csa_tree_add_190_195_groupi_n_9659);
  or csa_tree_add_190_195_groupi_g38946(csa_tree_add_190_195_groupi_n_10010 ,csa_tree_add_190_195_groupi_n_8390 ,csa_tree_add_190_195_groupi_n_9593);
  and csa_tree_add_190_195_groupi_g38947(csa_tree_add_190_195_groupi_n_10009 ,csa_tree_add_190_195_groupi_n_9515 ,csa_tree_add_190_195_groupi_n_9730);
  or csa_tree_add_190_195_groupi_g38948(csa_tree_add_190_195_groupi_n_10008 ,csa_tree_add_190_195_groupi_n_9196 ,csa_tree_add_190_195_groupi_n_9729);
  or csa_tree_add_190_195_groupi_g38949(csa_tree_add_190_195_groupi_n_10007 ,csa_tree_add_190_195_groupi_n_8094 ,csa_tree_add_190_195_groupi_n_9651);
  and csa_tree_add_190_195_groupi_g38950(csa_tree_add_190_195_groupi_n_10006 ,csa_tree_add_190_195_groupi_n_9184 ,csa_tree_add_190_195_groupi_n_9588);
  or csa_tree_add_190_195_groupi_g38951(csa_tree_add_190_195_groupi_n_10005 ,csa_tree_add_190_195_groupi_n_9342 ,csa_tree_add_190_195_groupi_n_117);
  or csa_tree_add_190_195_groupi_g38952(csa_tree_add_190_195_groupi_n_10004 ,csa_tree_add_190_195_groupi_n_9774 ,csa_tree_add_190_195_groupi_n_9627);
  nor csa_tree_add_190_195_groupi_g38953(csa_tree_add_190_195_groupi_n_10003 ,csa_tree_add_190_195_groupi_n_9721 ,csa_tree_add_190_195_groupi_n_9358);
  or csa_tree_add_190_195_groupi_g38954(csa_tree_add_190_195_groupi_n_10002 ,csa_tree_add_190_195_groupi_n_9719 ,csa_tree_add_190_195_groupi_n_9650);
  nor csa_tree_add_190_195_groupi_g38955(csa_tree_add_190_195_groupi_n_10001 ,csa_tree_add_190_195_groupi_n_9311 ,csa_tree_add_190_195_groupi_n_9617);
  or csa_tree_add_190_195_groupi_g38956(csa_tree_add_190_195_groupi_n_10000 ,csa_tree_add_190_195_groupi_n_8298 ,csa_tree_add_190_195_groupi_n_9811);
  or csa_tree_add_190_195_groupi_g38957(csa_tree_add_190_195_groupi_n_9999 ,csa_tree_add_190_195_groupi_n_119 ,csa_tree_add_190_195_groupi_n_9616);
  or csa_tree_add_190_195_groupi_g38958(csa_tree_add_190_195_groupi_n_9998 ,csa_tree_add_190_195_groupi_n_9644 ,csa_tree_add_190_195_groupi_n_9310);
  nor csa_tree_add_190_195_groupi_g38959(csa_tree_add_190_195_groupi_n_9997 ,csa_tree_add_190_195_groupi_n_9606 ,csa_tree_add_190_195_groupi_n_9339);
  or csa_tree_add_190_195_groupi_g38960(csa_tree_add_190_195_groupi_n_9996 ,csa_tree_add_190_195_groupi_n_8842 ,csa_tree_add_190_195_groupi_n_9577);
  nor csa_tree_add_190_195_groupi_g38961(csa_tree_add_190_195_groupi_n_9995 ,csa_tree_add_190_195_groupi_n_9775 ,csa_tree_add_190_195_groupi_n_9628);
  or csa_tree_add_190_195_groupi_g38962(csa_tree_add_190_195_groupi_n_9994 ,csa_tree_add_190_195_groupi_n_9788 ,csa_tree_add_190_195_groupi_n_9281);
  nor csa_tree_add_190_195_groupi_g38963(csa_tree_add_190_195_groupi_n_9993 ,csa_tree_add_190_195_groupi_n_9188 ,csa_tree_add_190_195_groupi_n_9706);
  and csa_tree_add_190_195_groupi_g38964(csa_tree_add_190_195_groupi_n_9992 ,csa_tree_add_190_195_groupi_n_7685 ,csa_tree_add_190_195_groupi_n_9785);
  or csa_tree_add_190_195_groupi_g38965(csa_tree_add_190_195_groupi_n_9991 ,csa_tree_add_190_195_groupi_n_9201 ,csa_tree_add_190_195_groupi_n_9692);
  nor csa_tree_add_190_195_groupi_g38966(csa_tree_add_190_195_groupi_n_9990 ,csa_tree_add_190_195_groupi_n_9522 ,csa_tree_add_190_195_groupi_n_9701);
  nor csa_tree_add_190_195_groupi_g38967(csa_tree_add_190_195_groupi_n_9989 ,csa_tree_add_190_195_groupi_n_8766 ,csa_tree_add_190_195_groupi_n_9665);
  or csa_tree_add_190_195_groupi_g38968(csa_tree_add_190_195_groupi_n_9988 ,csa_tree_add_190_195_groupi_n_9802 ,csa_tree_add_190_195_groupi_n_9699);
  nor csa_tree_add_190_195_groupi_g38969(csa_tree_add_190_195_groupi_n_9987 ,csa_tree_add_190_195_groupi_n_9669 ,csa_tree_add_190_195_groupi_n_9743);
  and csa_tree_add_190_195_groupi_g38970(csa_tree_add_190_195_groupi_n_9986 ,csa_tree_add_190_195_groupi_n_9030 ,csa_tree_add_190_195_groupi_n_9778);
  or csa_tree_add_190_195_groupi_g38971(csa_tree_add_190_195_groupi_n_9985 ,csa_tree_add_190_195_groupi_n_8991 ,csa_tree_add_190_195_groupi_n_9762);
  nor csa_tree_add_190_195_groupi_g38972(csa_tree_add_190_195_groupi_n_9984 ,csa_tree_add_190_195_groupi_n_8992 ,csa_tree_add_190_195_groupi_n_9763);
  nor csa_tree_add_190_195_groupi_g38973(csa_tree_add_190_195_groupi_n_9983 ,csa_tree_add_190_195_groupi_n_7071 ,csa_tree_add_190_195_groupi_n_9643);
  or csa_tree_add_190_195_groupi_g38974(csa_tree_add_190_195_groupi_n_9982 ,csa_tree_add_190_195_groupi_n_7072 ,csa_tree_add_190_195_groupi_n_9642);
  or csa_tree_add_190_195_groupi_g38975(csa_tree_add_190_195_groupi_n_9981 ,csa_tree_add_190_195_groupi_n_9784 ,csa_tree_add_190_195_groupi_n_9635);
  or csa_tree_add_190_195_groupi_g38976(csa_tree_add_190_195_groupi_n_9980 ,csa_tree_add_190_195_groupi_n_9183 ,csa_tree_add_190_195_groupi_n_9581);
  nor csa_tree_add_190_195_groupi_g38977(csa_tree_add_190_195_groupi_n_9979 ,csa_tree_add_190_195_groupi_n_9783 ,csa_tree_add_190_195_groupi_n_9636);
  or csa_tree_add_190_195_groupi_g38978(csa_tree_add_190_195_groupi_n_9978 ,csa_tree_add_190_195_groupi_n_9602 ,csa_tree_add_190_195_groupi_n_9306);
  nor csa_tree_add_190_195_groupi_g38979(csa_tree_add_190_195_groupi_n_9977 ,csa_tree_add_190_195_groupi_n_9601 ,csa_tree_add_190_195_groupi_n_9307);
  nor csa_tree_add_190_195_groupi_g38980(csa_tree_add_190_195_groupi_n_9976 ,csa_tree_add_190_195_groupi_n_9645 ,csa_tree_add_190_195_groupi_n_9309);
  nor csa_tree_add_190_195_groupi_g38981(csa_tree_add_190_195_groupi_n_9975 ,csa_tree_add_190_195_groupi_n_9030 ,csa_tree_add_190_195_groupi_n_9778);
  or csa_tree_add_190_195_groupi_g38982(csa_tree_add_190_195_groupi_n_9974 ,csa_tree_add_190_195_groupi_n_7111 ,csa_tree_add_190_195_groupi_n_9623);
  nor csa_tree_add_190_195_groupi_g38983(csa_tree_add_190_195_groupi_n_9973 ,csa_tree_add_190_195_groupi_n_7112 ,csa_tree_add_190_195_groupi_n_9624);
  or csa_tree_add_190_195_groupi_g38984(csa_tree_add_190_195_groupi_n_9972 ,csa_tree_add_190_195_groupi_n_9507 ,csa_tree_add_190_195_groupi_n_9685);
  nor csa_tree_add_190_195_groupi_g38985(csa_tree_add_190_195_groupi_n_9971 ,csa_tree_add_190_195_groupi_n_9761 ,csa_tree_add_190_195_groupi_n_9773);
  or csa_tree_add_190_195_groupi_g38986(csa_tree_add_190_195_groupi_n_9970 ,csa_tree_add_190_195_groupi_n_9679 ,csa_tree_add_190_195_groupi_n_9652);
  nor csa_tree_add_190_195_groupi_g38987(csa_tree_add_190_195_groupi_n_9969 ,csa_tree_add_190_195_groupi_n_9506 ,csa_tree_add_190_195_groupi_n_9681);
  or csa_tree_add_190_195_groupi_g38988(csa_tree_add_190_195_groupi_n_9968 ,csa_tree_add_190_195_groupi_n_9760 ,csa_tree_add_190_195_groupi_n_9772);
  or csa_tree_add_190_195_groupi_g38989(csa_tree_add_190_195_groupi_n_9967 ,csa_tree_add_190_195_groupi_n_9512 ,csa_tree_add_190_195_groupi_n_9674);
  or csa_tree_add_190_195_groupi_g38990(csa_tree_add_190_195_groupi_n_9966 ,csa_tree_add_190_195_groupi_n_9314 ,csa_tree_add_190_195_groupi_n_9779);
  or csa_tree_add_190_195_groupi_g38991(csa_tree_add_190_195_groupi_n_9965 ,csa_tree_add_190_195_groupi_n_9787 ,csa_tree_add_190_195_groupi_n_9570);
  or csa_tree_add_190_195_groupi_g38992(csa_tree_add_190_195_groupi_n_9964 ,csa_tree_add_190_195_groupi_n_9160 ,csa_tree_add_190_195_groupi_n_9646);
  nor csa_tree_add_190_195_groupi_g38993(csa_tree_add_190_195_groupi_n_9963 ,csa_tree_add_190_195_groupi_n_9159 ,csa_tree_add_190_195_groupi_n_9647);
  and csa_tree_add_190_195_groupi_g38994(csa_tree_add_190_195_groupi_n_10087 ,csa_tree_add_190_195_groupi_n_9461 ,csa_tree_add_190_195_groupi_n_9712);
  and csa_tree_add_190_195_groupi_g38995(csa_tree_add_190_195_groupi_n_10086 ,csa_tree_add_190_195_groupi_n_8937 ,csa_tree_add_190_195_groupi_n_9672);
  and csa_tree_add_190_195_groupi_g38996(csa_tree_add_190_195_groupi_n_10085 ,csa_tree_add_190_195_groupi_n_9413 ,csa_tree_add_190_195_groupi_n_9676);
  and csa_tree_add_190_195_groupi_g38997(csa_tree_add_190_195_groupi_n_10084 ,csa_tree_add_190_195_groupi_n_9399 ,csa_tree_add_190_195_groupi_n_9684);
  and csa_tree_add_190_195_groupi_g38998(csa_tree_add_190_195_groupi_n_10083 ,csa_tree_add_190_195_groupi_n_9257 ,csa_tree_add_190_195_groupi_n_9689);
  and csa_tree_add_190_195_groupi_g38999(csa_tree_add_190_195_groupi_n_10082 ,csa_tree_add_190_195_groupi_n_8060 ,csa_tree_add_190_195_groupi_n_9691);
  and csa_tree_add_190_195_groupi_g39000(csa_tree_add_190_195_groupi_n_10081 ,csa_tree_add_190_195_groupi_n_9387 ,csa_tree_add_190_195_groupi_n_9696);
  and csa_tree_add_190_195_groupi_g39001(csa_tree_add_190_195_groupi_n_10080 ,csa_tree_add_190_195_groupi_n_7703 ,csa_tree_add_190_195_groupi_n_9709);
  and csa_tree_add_190_195_groupi_g39002(csa_tree_add_190_195_groupi_n_10079 ,csa_tree_add_190_195_groupi_n_9255 ,csa_tree_add_190_195_groupi_n_9711);
  and csa_tree_add_190_195_groupi_g39003(csa_tree_add_190_195_groupi_n_10078 ,csa_tree_add_190_195_groupi_n_9261 ,csa_tree_add_190_195_groupi_n_9715);
  and csa_tree_add_190_195_groupi_g39004(csa_tree_add_190_195_groupi_n_10077 ,csa_tree_add_190_195_groupi_n_9393 ,csa_tree_add_190_195_groupi_n_9717);
  and csa_tree_add_190_195_groupi_g39005(csa_tree_add_190_195_groupi_n_10076 ,csa_tree_add_190_195_groupi_n_9429 ,csa_tree_add_190_195_groupi_n_9595);
  and csa_tree_add_190_195_groupi_g39006(csa_tree_add_190_195_groupi_n_10075 ,csa_tree_add_190_195_groupi_n_9391 ,csa_tree_add_190_195_groupi_n_9716);
  and csa_tree_add_190_195_groupi_g39007(csa_tree_add_190_195_groupi_n_10074 ,csa_tree_add_190_195_groupi_n_9279 ,csa_tree_add_190_195_groupi_n_9592);
  and csa_tree_add_190_195_groupi_g39008(csa_tree_add_190_195_groupi_n_10073 ,csa_tree_add_190_195_groupi_n_9402 ,csa_tree_add_190_195_groupi_n_9723);
  and csa_tree_add_190_195_groupi_g39009(csa_tree_add_190_195_groupi_n_10072 ,csa_tree_add_190_195_groupi_n_9417 ,csa_tree_add_190_195_groupi_n_9726);
  and csa_tree_add_190_195_groupi_g39010(csa_tree_add_190_195_groupi_n_10071 ,csa_tree_add_190_195_groupi_n_9277 ,csa_tree_add_190_195_groupi_n_9591);
  and csa_tree_add_190_195_groupi_g39011(csa_tree_add_190_195_groupi_n_10070 ,csa_tree_add_190_195_groupi_n_9422 ,csa_tree_add_190_195_groupi_n_9734);
  and csa_tree_add_190_195_groupi_g39012(csa_tree_add_190_195_groupi_n_10069 ,csa_tree_add_190_195_groupi_n_9430 ,csa_tree_add_190_195_groupi_n_9736);
  and csa_tree_add_190_195_groupi_g39013(csa_tree_add_190_195_groupi_n_10068 ,csa_tree_add_190_195_groupi_n_8927 ,csa_tree_add_190_195_groupi_n_9590);
  and csa_tree_add_190_195_groupi_g39014(csa_tree_add_190_195_groupi_n_10067 ,csa_tree_add_190_195_groupi_n_9462 ,csa_tree_add_190_195_groupi_n_9741);
  and csa_tree_add_190_195_groupi_g39015(csa_tree_add_190_195_groupi_n_10066 ,csa_tree_add_190_195_groupi_n_9457 ,csa_tree_add_190_195_groupi_n_9747);
  or csa_tree_add_190_195_groupi_g39016(csa_tree_add_190_195_groupi_n_10065 ,csa_tree_add_190_195_groupi_n_9419 ,csa_tree_add_190_195_groupi_n_9671);
  and csa_tree_add_190_195_groupi_g39017(csa_tree_add_190_195_groupi_n_10063 ,csa_tree_add_190_195_groupi_n_7721 ,csa_tree_add_190_195_groupi_n_9718);
  or csa_tree_add_190_195_groupi_g39018(csa_tree_add_190_195_groupi_n_10061 ,csa_tree_add_190_195_groupi_n_8760 ,csa_tree_add_190_195_groupi_n_9727);
  or csa_tree_add_190_195_groupi_g39019(csa_tree_add_190_195_groupi_n_10060 ,csa_tree_add_190_195_groupi_n_9272 ,csa_tree_add_190_195_groupi_n_9683);
  or csa_tree_add_190_195_groupi_g39020(csa_tree_add_190_195_groupi_n_10057 ,csa_tree_add_190_195_groupi_n_9072 ,csa_tree_add_190_195_groupi_n_9708);
  or csa_tree_add_190_195_groupi_g39021(csa_tree_add_190_195_groupi_n_10055 ,csa_tree_add_190_195_groupi_n_9432 ,csa_tree_add_190_195_groupi_n_9737);
  and csa_tree_add_190_195_groupi_g39022(csa_tree_add_190_195_groupi_n_10053 ,csa_tree_add_190_195_groupi_n_9068 ,csa_tree_add_190_195_groupi_n_9705);
  and csa_tree_add_190_195_groupi_g39023(csa_tree_add_190_195_groupi_n_10052 ,csa_tree_add_190_195_groupi_n_9149 ,csa_tree_add_190_195_groupi_n_9746);
  and csa_tree_add_190_195_groupi_g39024(csa_tree_add_190_195_groupi_n_10050 ,csa_tree_add_190_195_groupi_n_9107 ,csa_tree_add_190_195_groupi_n_9724);
  and csa_tree_add_190_195_groupi_g39025(csa_tree_add_190_195_groupi_n_10048 ,csa_tree_add_190_195_groupi_n_9372 ,csa_tree_add_190_195_groupi_n_9702);
  and csa_tree_add_190_195_groupi_g39026(csa_tree_add_190_195_groupi_n_10047 ,csa_tree_add_190_195_groupi_n_9382 ,csa_tree_add_190_195_groupi_n_9713);
  or csa_tree_add_190_195_groupi_g39027(csa_tree_add_190_195_groupi_n_10046 ,csa_tree_add_190_195_groupi_n_9379 ,csa_tree_add_190_195_groupi_n_9710);
  or csa_tree_add_190_195_groupi_g39028(csa_tree_add_190_195_groupi_n_10044 ,csa_tree_add_190_195_groupi_n_9453 ,csa_tree_add_190_195_groupi_n_9690);
  or csa_tree_add_190_195_groupi_g39029(csa_tree_add_190_195_groupi_n_10042 ,csa_tree_add_190_195_groupi_n_8796 ,csa_tree_add_190_195_groupi_n_9742);
  and csa_tree_add_190_195_groupi_g39030(csa_tree_add_190_195_groupi_n_10041 ,csa_tree_add_190_195_groupi_n_9260 ,csa_tree_add_190_195_groupi_n_9688);
  and csa_tree_add_190_195_groupi_g39031(csa_tree_add_190_195_groupi_n_10038 ,csa_tree_add_190_195_groupi_n_9122 ,csa_tree_add_190_195_groupi_n_9687);
  or csa_tree_add_190_195_groupi_g39032(csa_tree_add_190_195_groupi_n_10036 ,csa_tree_add_190_195_groupi_n_9426 ,csa_tree_add_190_195_groupi_n_9735);
  or csa_tree_add_190_195_groupi_g39033(csa_tree_add_190_195_groupi_n_10035 ,csa_tree_add_190_195_groupi_n_9466 ,csa_tree_add_190_195_groupi_n_9714);
  not csa_tree_add_190_195_groupi_g39035(csa_tree_add_190_195_groupi_n_9951 ,csa_tree_add_190_195_groupi_n_9950);
  not csa_tree_add_190_195_groupi_g39036(csa_tree_add_190_195_groupi_n_9949 ,csa_tree_add_190_195_groupi_n_9948);
  not csa_tree_add_190_195_groupi_g39037(csa_tree_add_190_195_groupi_n_9947 ,csa_tree_add_190_195_groupi_n_9946);
  not csa_tree_add_190_195_groupi_g39038(csa_tree_add_190_195_groupi_n_9945 ,csa_tree_add_190_195_groupi_n_9944);
  not csa_tree_add_190_195_groupi_g39039(csa_tree_add_190_195_groupi_n_9943 ,csa_tree_add_190_195_groupi_n_9942);
  not csa_tree_add_190_195_groupi_g39040(csa_tree_add_190_195_groupi_n_9941 ,csa_tree_add_190_195_groupi_n_9940);
  not csa_tree_add_190_195_groupi_g39041(csa_tree_add_190_195_groupi_n_9939 ,csa_tree_add_190_195_groupi_n_9938);
  not csa_tree_add_190_195_groupi_g39042(csa_tree_add_190_195_groupi_n_9936 ,csa_tree_add_190_195_groupi_n_9935);
  not csa_tree_add_190_195_groupi_g39043(csa_tree_add_190_195_groupi_n_9933 ,csa_tree_add_190_195_groupi_n_9932);
  not csa_tree_add_190_195_groupi_g39044(csa_tree_add_190_195_groupi_n_9930 ,csa_tree_add_190_195_groupi_n_9929);
  not csa_tree_add_190_195_groupi_g39045(csa_tree_add_190_195_groupi_n_9927 ,csa_tree_add_190_195_groupi_n_9928);
  not csa_tree_add_190_195_groupi_g39046(csa_tree_add_190_195_groupi_n_9926 ,csa_tree_add_190_195_groupi_n_9925);
  not csa_tree_add_190_195_groupi_g39047(csa_tree_add_190_195_groupi_n_9924 ,csa_tree_add_190_195_groupi_n_9923);
  not csa_tree_add_190_195_groupi_g39048(csa_tree_add_190_195_groupi_n_9922 ,csa_tree_add_190_195_groupi_n_9921);
  not csa_tree_add_190_195_groupi_g39049(csa_tree_add_190_195_groupi_n_9919 ,csa_tree_add_190_195_groupi_n_9918);
  not csa_tree_add_190_195_groupi_g39050(csa_tree_add_190_195_groupi_n_9917 ,csa_tree_add_190_195_groupi_n_9916);
  not csa_tree_add_190_195_groupi_g39051(csa_tree_add_190_195_groupi_n_9915 ,csa_tree_add_190_195_groupi_n_9914);
  not csa_tree_add_190_195_groupi_g39052(csa_tree_add_190_195_groupi_n_9913 ,csa_tree_add_190_195_groupi_n_9912);
  not csa_tree_add_190_195_groupi_g39053(csa_tree_add_190_195_groupi_n_9911 ,csa_tree_add_190_195_groupi_n_9910);
  not csa_tree_add_190_195_groupi_g39054(csa_tree_add_190_195_groupi_n_9909 ,csa_tree_add_190_195_groupi_n_9908);
  not csa_tree_add_190_195_groupi_g39055(csa_tree_add_190_195_groupi_n_9907 ,csa_tree_add_190_195_groupi_n_9906);
  not csa_tree_add_190_195_groupi_g39056(csa_tree_add_190_195_groupi_n_9905 ,csa_tree_add_190_195_groupi_n_9904);
  not csa_tree_add_190_195_groupi_g39057(csa_tree_add_190_195_groupi_n_9903 ,csa_tree_add_190_195_groupi_n_9902);
  not csa_tree_add_190_195_groupi_g39058(csa_tree_add_190_195_groupi_n_9901 ,csa_tree_add_190_195_groupi_n_9900);
  not csa_tree_add_190_195_groupi_g39059(csa_tree_add_190_195_groupi_n_9899 ,csa_tree_add_190_195_groupi_n_9898);
  not csa_tree_add_190_195_groupi_g39061(csa_tree_add_190_195_groupi_n_9896 ,csa_tree_add_190_195_groupi_n_9895);
  not csa_tree_add_190_195_groupi_g39062(csa_tree_add_190_195_groupi_n_9894 ,csa_tree_add_190_195_groupi_n_9893);
  not csa_tree_add_190_195_groupi_g39063(csa_tree_add_190_195_groupi_n_9891 ,csa_tree_add_190_195_groupi_n_9892);
  not csa_tree_add_190_195_groupi_g39064(csa_tree_add_190_195_groupi_n_9890 ,csa_tree_add_190_195_groupi_n_9889);
  not csa_tree_add_190_195_groupi_g39065(csa_tree_add_190_195_groupi_n_9888 ,csa_tree_add_190_195_groupi_n_9887);
  not csa_tree_add_190_195_groupi_g39066(csa_tree_add_190_195_groupi_n_9885 ,csa_tree_add_190_195_groupi_n_9886);
  not csa_tree_add_190_195_groupi_g39067(csa_tree_add_190_195_groupi_n_9884 ,csa_tree_add_190_195_groupi_n_9883);
  not csa_tree_add_190_195_groupi_g39068(csa_tree_add_190_195_groupi_n_9882 ,csa_tree_add_190_195_groupi_n_9881);
  not csa_tree_add_190_195_groupi_g39069(csa_tree_add_190_195_groupi_n_9880 ,csa_tree_add_190_195_groupi_n_9879);
  not csa_tree_add_190_195_groupi_g39070(csa_tree_add_190_195_groupi_n_9878 ,csa_tree_add_190_195_groupi_n_9877);
  not csa_tree_add_190_195_groupi_g39071(csa_tree_add_190_195_groupi_n_9876 ,csa_tree_add_190_195_groupi_n_9875);
  not csa_tree_add_190_195_groupi_g39072(csa_tree_add_190_195_groupi_n_9873 ,csa_tree_add_190_195_groupi_n_9872);
  not csa_tree_add_190_195_groupi_g39073(csa_tree_add_190_195_groupi_n_9871 ,csa_tree_add_190_195_groupi_n_9870);
  not csa_tree_add_190_195_groupi_g39074(csa_tree_add_190_195_groupi_n_9868 ,csa_tree_add_190_195_groupi_n_9867);
  not csa_tree_add_190_195_groupi_g39075(csa_tree_add_190_195_groupi_n_9865 ,csa_tree_add_190_195_groupi_n_9866);
  not csa_tree_add_190_195_groupi_g39076(csa_tree_add_190_195_groupi_n_9863 ,csa_tree_add_190_195_groupi_n_9864);
  not csa_tree_add_190_195_groupi_g39077(csa_tree_add_190_195_groupi_n_9862 ,csa_tree_add_190_195_groupi_n_9861);
  nor csa_tree_add_190_195_groupi_g39078(csa_tree_add_190_195_groupi_n_9859 ,csa_tree_add_190_195_groupi_n_8321 ,csa_tree_add_190_195_groupi_n_9626);
  nor csa_tree_add_190_195_groupi_g39079(csa_tree_add_190_195_groupi_n_9858 ,csa_tree_add_190_195_groupi_n_9620 ,csa_tree_add_190_195_groupi_n_9346);
  or csa_tree_add_190_195_groupi_g39080(csa_tree_add_190_195_groupi_n_9857 ,csa_tree_add_190_195_groupi_n_9498 ,csa_tree_add_190_195_groupi_n_9614);
  nor csa_tree_add_190_195_groupi_g39081(csa_tree_add_190_195_groupi_n_9856 ,csa_tree_add_190_195_groupi_n_9497 ,csa_tree_add_190_195_groupi_n_9615);
  or csa_tree_add_190_195_groupi_g39082(csa_tree_add_190_195_groupi_n_9855 ,csa_tree_add_190_195_groupi_n_7138 ,csa_tree_add_190_195_groupi_n_9604);
  and csa_tree_add_190_195_groupi_g39083(csa_tree_add_190_195_groupi_n_9854 ,csa_tree_add_190_195_groupi_n_7138 ,csa_tree_add_190_195_groupi_n_9604);
  or csa_tree_add_190_195_groupi_g39084(csa_tree_add_190_195_groupi_n_9853 ,csa_tree_add_190_195_groupi_n_9668 ,csa_tree_add_190_195_groupi_n_9263);
  or csa_tree_add_190_195_groupi_g39085(csa_tree_add_190_195_groupi_n_9852 ,csa_tree_add_190_195_groupi_n_9750 ,csa_tree_add_190_195_groupi_n_8665);
  nor csa_tree_add_190_195_groupi_g39086(csa_tree_add_190_195_groupi_n_9851 ,csa_tree_add_190_195_groupi_n_9751 ,csa_tree_add_190_195_groupi_n_8666);
  or csa_tree_add_190_195_groupi_g39087(csa_tree_add_190_195_groupi_n_9850 ,csa_tree_add_190_195_groupi_n_9571 ,csa_tree_add_190_195_groupi_n_9653);
  nor csa_tree_add_190_195_groupi_g39088(csa_tree_add_190_195_groupi_n_9849 ,csa_tree_add_190_195_groupi_n_9526 ,csa_tree_add_190_195_groupi_n_9573);
  or csa_tree_add_190_195_groupi_g39089(csa_tree_add_190_195_groupi_n_9848 ,csa_tree_add_190_195_groupi_n_9470 ,csa_tree_add_190_195_groupi_n_9611);
  nor csa_tree_add_190_195_groupi_g39090(csa_tree_add_190_195_groupi_n_9847 ,csa_tree_add_190_195_groupi_n_9471 ,csa_tree_add_190_195_groupi_n_9610);
  or csa_tree_add_190_195_groupi_g39091(csa_tree_add_190_195_groupi_n_9846 ,csa_tree_add_190_195_groupi_n_9317 ,csa_tree_add_190_195_groupi_n_9754);
  and csa_tree_add_190_195_groupi_g39092(csa_tree_add_190_195_groupi_n_9845 ,csa_tree_add_190_195_groupi_n_9317 ,csa_tree_add_190_195_groupi_n_9754);
  and csa_tree_add_190_195_groupi_g39093(csa_tree_add_190_195_groupi_n_9844 ,csa_tree_add_190_195_groupi_n_9314 ,csa_tree_add_190_195_groupi_n_9779);
  or csa_tree_add_190_195_groupi_g39094(csa_tree_add_190_195_groupi_n_9843 ,csa_tree_add_190_195_groupi_n_110 ,csa_tree_add_190_195_groupi_n_9345);
  or csa_tree_add_190_195_groupi_g39095(csa_tree_add_190_195_groupi_n_9842 ,csa_tree_add_190_195_groupi_n_9337 ,csa_tree_add_190_195_groupi_n_9613);
  xnor csa_tree_add_190_195_groupi_g39096(csa_tree_add_190_195_groupi_n_9841 ,csa_tree_add_190_195_groupi_n_7168 ,csa_tree_add_190_195_groupi_n_9507);
  xnor csa_tree_add_190_195_groupi_g39097(csa_tree_add_190_195_groupi_n_9840 ,csa_tree_add_190_195_groupi_n_8818 ,csa_tree_add_190_195_groupi_n_9349);
  xnor csa_tree_add_190_195_groupi_g39098(csa_tree_add_190_195_groupi_n_9839 ,csa_tree_add_190_195_groupi_n_7593 ,csa_tree_add_190_195_groupi_n_9479);
  xnor csa_tree_add_190_195_groupi_g39099(csa_tree_add_190_195_groupi_n_9838 ,csa_tree_add_190_195_groupi_n_9355 ,csa_tree_add_190_195_groupi_n_7138);
  xnor csa_tree_add_190_195_groupi_g39100(csa_tree_add_190_195_groupi_n_9837 ,csa_tree_add_190_195_groupi_n_8955 ,csa_tree_add_190_195_groupi_n_9523);
  xnor csa_tree_add_190_195_groupi_g39101(csa_tree_add_190_195_groupi_n_9836 ,csa_tree_add_190_195_groupi_n_9526 ,csa_tree_add_190_195_groupi_n_9468);
  xnor csa_tree_add_190_195_groupi_g39102(csa_tree_add_190_195_groupi_n_9835 ,csa_tree_add_190_195_groupi_n_9025 ,csa_tree_add_190_195_groupi_n_9297);
  xor csa_tree_add_190_195_groupi_g39103(csa_tree_add_190_195_groupi_n_9834 ,csa_tree_add_190_195_groupi_n_9354 ,csa_tree_add_190_195_groupi_n_7562);
  xnor csa_tree_add_190_195_groupi_g39104(csa_tree_add_190_195_groupi_n_9833 ,csa_tree_add_190_195_groupi_n_9009 ,csa_tree_add_190_195_groupi_n_9320);
  xnor csa_tree_add_190_195_groupi_g39105(csa_tree_add_190_195_groupi_n_9832 ,csa_tree_add_190_195_groupi_n_9166 ,csa_tree_add_190_195_groupi_n_9303);
  xnor csa_tree_add_190_195_groupi_g39106(csa_tree_add_190_195_groupi_n_9831 ,csa_tree_add_190_195_groupi_n_7144 ,csa_tree_add_190_195_groupi_n_9350);
  xnor csa_tree_add_190_195_groupi_g39108(csa_tree_add_190_195_groupi_n_9830 ,csa_tree_add_190_195_groupi_n_8390 ,csa_tree_add_190_195_groupi_n_9324);
  xnor csa_tree_add_190_195_groupi_g39109(csa_tree_add_190_195_groupi_n_9829 ,csa_tree_add_190_195_groupi_n_9184 ,csa_tree_add_190_195_groupi_n_9285);
  xnor csa_tree_add_190_195_groupi_g39110(csa_tree_add_190_195_groupi_n_9828 ,csa_tree_add_190_195_groupi_n_9326 ,csa_tree_add_190_195_groupi_n_9515);
  xnor csa_tree_add_190_195_groupi_g39111(csa_tree_add_190_195_groupi_n_9827 ,csa_tree_add_190_195_groupi_n_9486 ,csa_tree_add_190_195_groupi_n_9500);
  xnor csa_tree_add_190_195_groupi_g39113(csa_tree_add_190_195_groupi_n_9826 ,csa_tree_add_190_195_groupi_n_9505 ,csa_tree_add_190_195_groupi_n_9012);
  xnor csa_tree_add_190_195_groupi_g39114(csa_tree_add_190_195_groupi_n_9825 ,csa_tree_add_190_195_groupi_n_9504 ,csa_tree_add_190_195_groupi_n_9346);
  xnor csa_tree_add_190_195_groupi_g39115(csa_tree_add_190_195_groupi_n_9824 ,csa_tree_add_190_195_groupi_n_8609 ,csa_tree_add_190_195_groupi_n_9496);
  xnor csa_tree_add_190_195_groupi_g39116(csa_tree_add_190_195_groupi_n_9823 ,csa_tree_add_190_195_groupi_n_7116 ,csa_tree_add_190_195_groupi_n_9360);
  xnor csa_tree_add_190_195_groupi_g39117(csa_tree_add_190_195_groupi_n_9822 ,csa_tree_add_190_195_groupi_n_9508 ,csa_tree_add_190_195_groupi_n_9001);
  xnor csa_tree_add_190_195_groupi_g39118(csa_tree_add_190_195_groupi_n_9821 ,csa_tree_add_190_195_groupi_n_9492 ,csa_tree_add_190_195_groupi_n_9015);
  xnor csa_tree_add_190_195_groupi_g39119(csa_tree_add_190_195_groupi_n_9820 ,csa_tree_add_190_195_groupi_n_7172 ,csa_tree_add_190_195_groupi_n_9359);
  xnor csa_tree_add_190_195_groupi_g39120(csa_tree_add_190_195_groupi_n_9819 ,csa_tree_add_190_195_groupi_n_9519 ,csa_tree_add_190_195_groupi_n_8990);
  xor csa_tree_add_190_195_groupi_g39122(csa_tree_add_190_195_groupi_n_9818 ,csa_tree_add_190_195_groupi_n_9196 ,csa_tree_add_190_195_groupi_n_9488);
  xnor csa_tree_add_190_195_groupi_g39123(csa_tree_add_190_195_groupi_n_9817 ,csa_tree_add_190_195_groupi_n_9169 ,csa_tree_add_190_195_groupi_n_9516);
  xnor csa_tree_add_190_195_groupi_g39124(csa_tree_add_190_195_groupi_n_9816 ,csa_tree_add_190_195_groupi_n_9521 ,csa_tree_add_190_195_groupi_n_5417);
  xnor csa_tree_add_190_195_groupi_g39125(csa_tree_add_190_195_groupi_n_9815 ,csa_tree_add_190_195_groupi_n_9299 ,csa_tree_add_190_195_groupi_n_9362);
  xor csa_tree_add_190_195_groupi_g39126(csa_tree_add_190_195_groupi_n_9814 ,csa_tree_add_190_195_groupi_n_9522 ,csa_tree_add_190_195_groupi_n_9286);
  xnor csa_tree_add_190_195_groupi_g39127(csa_tree_add_190_195_groupi_n_9813 ,csa_tree_add_190_195_groupi_n_9476 ,csa_tree_add_190_195_groupi_n_9506);
  xnor csa_tree_add_190_195_groupi_g39128(csa_tree_add_190_195_groupi_n_9812 ,csa_tree_add_190_195_groupi_n_7515 ,csa_tree_add_190_195_groupi_n_9520);
  or csa_tree_add_190_195_groupi_g39129(csa_tree_add_190_195_groupi_n_9962 ,csa_tree_add_190_195_groupi_n_9268 ,csa_tree_add_190_195_groupi_n_9584);
  xnor csa_tree_add_190_195_groupi_g39130(csa_tree_add_190_195_groupi_n_9961 ,csa_tree_add_190_195_groupi_n_75 ,csa_tree_add_190_195_groupi_n_9237);
  and csa_tree_add_190_195_groupi_g39131(csa_tree_add_190_195_groupi_n_9960 ,csa_tree_add_190_195_groupi_n_9271 ,csa_tree_add_190_195_groupi_n_9585);
  xnor csa_tree_add_190_195_groupi_g39132(csa_tree_add_190_195_groupi_n_9959 ,csa_tree_add_190_195_groupi_n_8207 ,csa_tree_add_190_195_groupi_n_9217);
  xnor csa_tree_add_190_195_groupi_g39133(csa_tree_add_190_195_groupi_n_9958 ,csa_tree_add_190_195_groupi_n_5393 ,csa_tree_add_190_195_groupi_n_9244);
  xnor csa_tree_add_190_195_groupi_g39134(csa_tree_add_190_195_groupi_n_9957 ,csa_tree_add_190_195_groupi_n_8846 ,csa_tree_add_190_195_groupi_n_9222);
  xnor csa_tree_add_190_195_groupi_g39135(csa_tree_add_190_195_groupi_n_9956 ,csa_tree_add_190_195_groupi_n_5435 ,csa_tree_add_190_195_groupi_n_9212);
  and csa_tree_add_190_195_groupi_g39136(csa_tree_add_190_195_groupi_n_9955 ,csa_tree_add_190_195_groupi_n_7958 ,csa_tree_add_190_195_groupi_n_9586);
  and csa_tree_add_190_195_groupi_g39137(csa_tree_add_190_195_groupi_n_9954 ,csa_tree_add_190_195_groupi_n_9253 ,csa_tree_add_190_195_groupi_n_9579);
  xnor csa_tree_add_190_195_groupi_g39138(csa_tree_add_190_195_groupi_n_9953 ,csa_tree_add_190_195_groupi_n_9368 ,csa_tree_add_190_195_groupi_n_9245);
  xnor csa_tree_add_190_195_groupi_g39139(csa_tree_add_190_195_groupi_n_9952 ,csa_tree_add_190_195_groupi_n_9363 ,csa_tree_add_190_195_groupi_n_9248);
  and csa_tree_add_190_195_groupi_g39140(csa_tree_add_190_195_groupi_n_9950 ,csa_tree_add_190_195_groupi_n_9282 ,csa_tree_add_190_195_groupi_n_9673);
  xnor csa_tree_add_190_195_groupi_g39141(csa_tree_add_190_195_groupi_n_9948 ,csa_tree_add_190_195_groupi_n_9357 ,csa_tree_add_190_195_groupi_n_8258);
  xnor csa_tree_add_190_195_groupi_g39142(csa_tree_add_190_195_groupi_n_9946 ,csa_tree_add_190_195_groupi_n_9367 ,csa_tree_add_190_195_groupi_n_9216);
  xnor csa_tree_add_190_195_groupi_g39143(csa_tree_add_190_195_groupi_n_9944 ,csa_tree_add_190_195_groupi_n_7607 ,csa_tree_add_190_195_groupi_n_9215);
  xnor csa_tree_add_190_195_groupi_g39144(csa_tree_add_190_195_groupi_n_9942 ,csa_tree_add_190_195_groupi_n_8030 ,csa_tree_add_190_195_groupi_n_121);
  xnor csa_tree_add_190_195_groupi_g39145(csa_tree_add_190_195_groupi_n_9940 ,csa_tree_add_190_195_groupi_n_8622 ,csa_tree_add_190_195_groupi_n_9252);
  xnor csa_tree_add_190_195_groupi_g39146(csa_tree_add_190_195_groupi_n_9938 ,csa_tree_add_190_195_groupi_n_9187 ,csa_tree_add_190_195_groupi_n_9213);
  or csa_tree_add_190_195_groupi_g39147(csa_tree_add_190_195_groupi_n_9937 ,csa_tree_add_190_195_groupi_n_7478 ,csa_tree_add_190_195_groupi_n_9572);
  xnor csa_tree_add_190_195_groupi_g39148(csa_tree_add_190_195_groupi_n_9935 ,csa_tree_add_190_195_groupi_n_8357 ,csa_tree_add_190_195_groupi_n_9242);
  xnor csa_tree_add_190_195_groupi_g39149(csa_tree_add_190_195_groupi_n_9934 ,csa_tree_add_190_195_groupi_n_7565 ,csa_tree_add_190_195_groupi_n_9211);
  xnor csa_tree_add_190_195_groupi_g39150(csa_tree_add_190_195_groupi_n_9932 ,csa_tree_add_190_195_groupi_n_9365 ,csa_tree_add_190_195_groupi_n_9239);
  xnor csa_tree_add_190_195_groupi_g39151(csa_tree_add_190_195_groupi_n_9931 ,csa_tree_add_190_195_groupi_n_5321 ,csa_tree_add_190_195_groupi_n_9251);
  xnor csa_tree_add_190_195_groupi_g39152(csa_tree_add_190_195_groupi_n_9929 ,csa_tree_add_190_195_groupi_n_8867 ,csa_tree_add_190_195_groupi_n_9238);
  xnor csa_tree_add_190_195_groupi_g39153(csa_tree_add_190_195_groupi_n_9928 ,csa_tree_add_190_195_groupi_n_8519 ,csa_tree_add_190_195_groupi_n_9241);
  xnor csa_tree_add_190_195_groupi_g39154(csa_tree_add_190_195_groupi_n_9925 ,csa_tree_add_190_195_groupi_n_8521 ,csa_tree_add_190_195_groupi_n_9209);
  xnor csa_tree_add_190_195_groupi_g39155(csa_tree_add_190_195_groupi_n_9923 ,csa_tree_add_190_195_groupi_n_8524 ,csa_tree_add_190_195_groupi_n_9208);
  or csa_tree_add_190_195_groupi_g39156(csa_tree_add_190_195_groupi_n_9921 ,csa_tree_add_190_195_groupi_n_9270 ,csa_tree_add_190_195_groupi_n_9575);
  xnor csa_tree_add_190_195_groupi_g39157(csa_tree_add_190_195_groupi_n_9920 ,csa_tree_add_190_195_groupi_n_7166 ,csa_tree_add_190_195_groupi_n_9224);
  xnor csa_tree_add_190_195_groupi_g39158(csa_tree_add_190_195_groupi_n_9918 ,csa_tree_add_190_195_groupi_n_8841 ,csa_tree_add_190_195_groupi_n_9240);
  xnor csa_tree_add_190_195_groupi_g39159(csa_tree_add_190_195_groupi_n_9916 ,csa_tree_add_190_195_groupi_n_7826 ,csa_tree_add_190_195_groupi_n_9246);
  xnor csa_tree_add_190_195_groupi_g39160(csa_tree_add_190_195_groupi_n_9914 ,csa_tree_add_190_195_groupi_n_7583 ,csa_tree_add_190_195_groupi_n_9236);
  xnor csa_tree_add_190_195_groupi_g39161(csa_tree_add_190_195_groupi_n_9912 ,csa_tree_add_190_195_groupi_n_8974 ,csa_tree_add_190_195_groupi_n_9233);
  xnor csa_tree_add_190_195_groupi_g39162(csa_tree_add_190_195_groupi_n_9910 ,csa_tree_add_190_195_groupi_n_8021 ,csa_tree_add_190_195_groupi_n_9204);
  xnor csa_tree_add_190_195_groupi_g39163(csa_tree_add_190_195_groupi_n_9908 ,csa_tree_add_190_195_groupi_n_8611 ,csa_tree_add_190_195_groupi_n_122);
  xnor csa_tree_add_190_195_groupi_g39164(csa_tree_add_190_195_groupi_n_9906 ,csa_tree_add_190_195_groupi_n_8323 ,csa_tree_add_190_195_groupi_n_9207);
  xnor csa_tree_add_190_195_groupi_g39165(csa_tree_add_190_195_groupi_n_9904 ,csa_tree_add_190_195_groupi_n_8858 ,csa_tree_add_190_195_groupi_n_9228);
  xnor csa_tree_add_190_195_groupi_g39166(csa_tree_add_190_195_groupi_n_9902 ,csa_tree_add_190_195_groupi_n_8492 ,csa_tree_add_190_195_groupi_n_9206);
  xnor csa_tree_add_190_195_groupi_g39167(csa_tree_add_190_195_groupi_n_9900 ,csa_tree_add_190_195_groupi_n_7308 ,csa_tree_add_190_195_groupi_n_9205);
  xnor csa_tree_add_190_195_groupi_g39168(csa_tree_add_190_195_groupi_n_9898 ,csa_tree_add_190_195_groupi_n_9003 ,csa_tree_add_190_195_groupi_n_9210);
  xnor csa_tree_add_190_195_groupi_g39169(csa_tree_add_190_195_groupi_n_9897 ,csa_tree_add_190_195_groupi_n_7833 ,csa_tree_add_190_195_groupi_n_9247);
  xnor csa_tree_add_190_195_groupi_g39170(csa_tree_add_190_195_groupi_n_9895 ,csa_tree_add_190_195_groupi_n_9509 ,csa_tree_add_190_195_groupi_n_8262);
  xnor csa_tree_add_190_195_groupi_g39171(csa_tree_add_190_195_groupi_n_9893 ,csa_tree_add_190_195_groupi_n_9292 ,csa_tree_add_190_195_groupi_n_9230);
  xnor csa_tree_add_190_195_groupi_g39172(csa_tree_add_190_195_groupi_n_9892 ,csa_tree_add_190_195_groupi_n_8533 ,csa_tree_add_190_195_groupi_n_9234);
  xnor csa_tree_add_190_195_groupi_g39173(csa_tree_add_190_195_groupi_n_9889 ,csa_tree_add_190_195_groupi_n_8342 ,csa_tree_add_190_195_groupi_n_123);
  xnor csa_tree_add_190_195_groupi_g39174(csa_tree_add_190_195_groupi_n_9887 ,csa_tree_add_190_195_groupi_n_8677 ,csa_tree_add_190_195_groupi_n_9243);
  xnor csa_tree_add_190_195_groupi_g39175(csa_tree_add_190_195_groupi_n_9886 ,csa_tree_add_190_195_groupi_n_9049 ,csa_tree_add_190_195_groupi_n_9232);
  xnor csa_tree_add_190_195_groupi_g39176(csa_tree_add_190_195_groupi_n_9883 ,csa_tree_add_190_195_groupi_n_8875 ,csa_tree_add_190_195_groupi_n_9226);
  xnor csa_tree_add_190_195_groupi_g39177(csa_tree_add_190_195_groupi_n_9881 ,csa_tree_add_190_195_groupi_n_5454 ,csa_tree_add_190_195_groupi_n_9225);
  xnor csa_tree_add_190_195_groupi_g39178(csa_tree_add_190_195_groupi_n_9879 ,csa_tree_add_190_195_groupi_n_8983 ,csa_tree_add_190_195_groupi_n_9214);
  xnor csa_tree_add_190_195_groupi_g39179(csa_tree_add_190_195_groupi_n_9877 ,csa_tree_add_190_195_groupi_n_9192 ,csa_tree_add_190_195_groupi_n_9235);
  xnor csa_tree_add_190_195_groupi_g39180(csa_tree_add_190_195_groupi_n_9875 ,csa_tree_add_190_195_groupi_n_8352 ,csa_tree_add_190_195_groupi_n_9221);
  xnor csa_tree_add_190_195_groupi_g39181(csa_tree_add_190_195_groupi_n_9874 ,csa_tree_add_190_195_groupi_n_7617 ,csa_tree_add_190_195_groupi_n_9219);
  xnor csa_tree_add_190_195_groupi_g39182(csa_tree_add_190_195_groupi_n_9872 ,csa_tree_add_190_195_groupi_n_7366 ,csa_tree_add_190_195_groupi_n_9227);
  xnor csa_tree_add_190_195_groupi_g39183(csa_tree_add_190_195_groupi_n_9870 ,csa_tree_add_190_195_groupi_n_9514 ,csa_tree_add_190_195_groupi_n_8882);
  xnor csa_tree_add_190_195_groupi_g39184(csa_tree_add_190_195_groupi_n_9869 ,csa_tree_add_190_195_groupi_n_9513 ,csa_tree_add_190_195_groupi_n_8909);
  xnor csa_tree_add_190_195_groupi_g39185(csa_tree_add_190_195_groupi_n_9867 ,csa_tree_add_190_195_groupi_n_8620 ,csa_tree_add_190_195_groupi_n_9220);
  xnor csa_tree_add_190_195_groupi_g39186(csa_tree_add_190_195_groupi_n_9866 ,csa_tree_add_190_195_groupi_n_5926 ,csa_tree_add_190_195_groupi_n_9250);
  xnor csa_tree_add_190_195_groupi_g39187(csa_tree_add_190_195_groupi_n_9864 ,csa_tree_add_190_195_groupi_n_4611 ,csa_tree_add_190_195_groupi_n_9231);
  xnor csa_tree_add_190_195_groupi_g39188(csa_tree_add_190_195_groupi_n_9861 ,csa_tree_add_190_195_groupi_n_8661 ,csa_tree_add_190_195_groupi_n_9218);
  xnor csa_tree_add_190_195_groupi_g39189(csa_tree_add_190_195_groupi_n_9860 ,csa_tree_add_190_195_groupi_n_9181 ,csa_tree_add_190_195_groupi_n_9249);
  not csa_tree_add_190_195_groupi_g39190(csa_tree_add_190_195_groupi_n_9811 ,csa_tree_add_190_195_groupi_n_9810);
  not csa_tree_add_190_195_groupi_g39191(csa_tree_add_190_195_groupi_n_9809 ,csa_tree_add_190_195_groupi_n_9808);
  not csa_tree_add_190_195_groupi_g39192(csa_tree_add_190_195_groupi_n_9805 ,csa_tree_add_190_195_groupi_n_9804);
  not csa_tree_add_190_195_groupi_g39193(csa_tree_add_190_195_groupi_n_9802 ,csa_tree_add_190_195_groupi_n_9801);
  not csa_tree_add_190_195_groupi_g39195(csa_tree_add_190_195_groupi_n_9787 ,csa_tree_add_190_195_groupi_n_9786);
  not csa_tree_add_190_195_groupi_g39196(csa_tree_add_190_195_groupi_n_9784 ,csa_tree_add_190_195_groupi_n_9783);
  not csa_tree_add_190_195_groupi_g39197(csa_tree_add_190_195_groupi_n_9782 ,csa_tree_add_190_195_groupi_n_9781);
  not csa_tree_add_190_195_groupi_g39199(csa_tree_add_190_195_groupi_n_9778 ,csa_tree_add_190_195_groupi_n_9777);
  not csa_tree_add_190_195_groupi_g39200(csa_tree_add_190_195_groupi_n_9774 ,csa_tree_add_190_195_groupi_n_9775);
  not csa_tree_add_190_195_groupi_g39201(csa_tree_add_190_195_groupi_n_9773 ,csa_tree_add_190_195_groupi_n_9772);
  not csa_tree_add_190_195_groupi_g39202(csa_tree_add_190_195_groupi_n_9770 ,csa_tree_add_190_195_groupi_n_9769);
  not csa_tree_add_190_195_groupi_g39203(csa_tree_add_190_195_groupi_n_9767 ,csa_tree_add_190_195_groupi_n_9768);
  not csa_tree_add_190_195_groupi_g39204(csa_tree_add_190_195_groupi_n_9766 ,csa_tree_add_190_195_groupi_n_9765);
  not csa_tree_add_190_195_groupi_g39205(csa_tree_add_190_195_groupi_n_9762 ,csa_tree_add_190_195_groupi_n_9763);
  not csa_tree_add_190_195_groupi_g39206(csa_tree_add_190_195_groupi_n_9761 ,csa_tree_add_190_195_groupi_n_9760);
  not csa_tree_add_190_195_groupi_g39207(csa_tree_add_190_195_groupi_n_9758 ,csa_tree_add_190_195_groupi_n_9759);
  not csa_tree_add_190_195_groupi_g39208(csa_tree_add_190_195_groupi_n_9756 ,csa_tree_add_190_195_groupi_n_9757);
  not csa_tree_add_190_195_groupi_g39209(csa_tree_add_190_195_groupi_n_9752 ,csa_tree_add_190_195_groupi_n_9753);
  not csa_tree_add_190_195_groupi_g39210(csa_tree_add_190_195_groupi_n_9751 ,csa_tree_add_190_195_groupi_n_9750);
  or csa_tree_add_190_195_groupi_g39211(csa_tree_add_190_195_groupi_n_9749 ,csa_tree_add_190_195_groupi_n_7574 ,csa_tree_add_190_195_groupi_n_9482);
  and csa_tree_add_190_195_groupi_g39212(csa_tree_add_190_195_groupi_n_9748 ,csa_tree_add_190_195_groupi_n_7574 ,csa_tree_add_190_195_groupi_n_9482);
  or csa_tree_add_190_195_groupi_g39213(csa_tree_add_190_195_groupi_n_9747 ,csa_tree_add_190_195_groupi_n_9043 ,csa_tree_add_190_195_groupi_n_9456);
  or csa_tree_add_190_195_groupi_g39214(csa_tree_add_190_195_groupi_n_9746 ,csa_tree_add_190_195_groupi_n_9145 ,csa_tree_add_190_195_groupi_n_9369);
  or csa_tree_add_190_195_groupi_g39215(csa_tree_add_190_195_groupi_n_9745 ,csa_tree_add_190_195_groupi_n_8339 ,csa_tree_add_190_195_groupi_n_9292);
  and csa_tree_add_190_195_groupi_g39216(csa_tree_add_190_195_groupi_n_9744 ,csa_tree_add_190_195_groupi_n_8339 ,csa_tree_add_190_195_groupi_n_9292);
  and csa_tree_add_190_195_groupi_g39217(csa_tree_add_190_195_groupi_n_9743 ,csa_tree_add_190_195_groupi_n_8628 ,csa_tree_add_190_195_groupi_n_9318);
  and csa_tree_add_190_195_groupi_g39218(csa_tree_add_190_195_groupi_n_9742 ,csa_tree_add_190_195_groupi_n_8795 ,csa_tree_add_190_195_groupi_n_9513);
  or csa_tree_add_190_195_groupi_g39219(csa_tree_add_190_195_groupi_n_9741 ,csa_tree_add_190_195_groupi_n_8843 ,csa_tree_add_190_195_groupi_n_9464);
  or csa_tree_add_190_195_groupi_g39220(csa_tree_add_190_195_groupi_n_9740 ,csa_tree_add_190_195_groupi_n_7562 ,csa_tree_add_190_195_groupi_n_9300);
  nor csa_tree_add_190_195_groupi_g39221(csa_tree_add_190_195_groupi_n_9739 ,csa_tree_add_190_195_groupi_n_7561 ,csa_tree_add_190_195_groupi_n_9301);
  or csa_tree_add_190_195_groupi_g39222(csa_tree_add_190_195_groupi_n_9738 ,csa_tree_add_190_195_groupi_n_7592 ,csa_tree_add_190_195_groupi_n_9479);
  and csa_tree_add_190_195_groupi_g39223(csa_tree_add_190_195_groupi_n_9737 ,csa_tree_add_190_195_groupi_n_9431 ,csa_tree_add_190_195_groupi_n_9352);
  or csa_tree_add_190_195_groupi_g39224(csa_tree_add_190_195_groupi_n_9736 ,csa_tree_add_190_195_groupi_n_8845 ,csa_tree_add_190_195_groupi_n_9428);
  and csa_tree_add_190_195_groupi_g39225(csa_tree_add_190_195_groupi_n_9735 ,csa_tree_add_190_195_groupi_n_9359 ,csa_tree_add_190_195_groupi_n_9423);
  or csa_tree_add_190_195_groupi_g39226(csa_tree_add_190_195_groupi_n_9734 ,csa_tree_add_190_195_groupi_n_8713 ,csa_tree_add_190_195_groupi_n_9421);
  nor csa_tree_add_190_195_groupi_g39227(csa_tree_add_190_195_groupi_n_9733 ,csa_tree_add_190_195_groupi_n_8953 ,csa_tree_add_190_195_groupi_n_9325);
  nor csa_tree_add_190_195_groupi_g39228(csa_tree_add_190_195_groupi_n_9732 ,csa_tree_add_190_195_groupi_n_7593 ,csa_tree_add_190_195_groupi_n_9478);
  or csa_tree_add_190_195_groupi_g39229(csa_tree_add_190_195_groupi_n_9731 ,csa_tree_add_190_195_groupi_n_8956 ,csa_tree_add_190_195_groupi_n_9488);
  or csa_tree_add_190_195_groupi_g39230(csa_tree_add_190_195_groupi_n_9730 ,csa_tree_add_190_195_groupi_n_8952 ,csa_tree_add_190_195_groupi_n_9326);
  nor csa_tree_add_190_195_groupi_g39231(csa_tree_add_190_195_groupi_n_9729 ,csa_tree_add_190_195_groupi_n_8957 ,csa_tree_add_190_195_groupi_n_9487);
  or csa_tree_add_190_195_groupi_g39232(csa_tree_add_190_195_groupi_n_9728 ,csa_tree_add_190_195_groupi_n_7162 ,csa_tree_add_190_195_groupi_n_9489);
  nor csa_tree_add_190_195_groupi_g39233(csa_tree_add_190_195_groupi_n_9727 ,csa_tree_add_190_195_groupi_n_9514 ,csa_tree_add_190_195_groupi_n_8751);
  or csa_tree_add_190_195_groupi_g39234(csa_tree_add_190_195_groupi_n_9726 ,csa_tree_add_190_195_groupi_n_8389 ,csa_tree_add_190_195_groupi_n_9396);
  nor csa_tree_add_190_195_groupi_g39235(csa_tree_add_190_195_groupi_n_9725 ,csa_tree_add_190_195_groupi_n_7161 ,csa_tree_add_190_195_groupi_n_9490);
  or csa_tree_add_190_195_groupi_g39236(csa_tree_add_190_195_groupi_n_9724 ,csa_tree_add_190_195_groupi_n_9103 ,csa_tree_add_190_195_groupi_n_9361);
  or csa_tree_add_190_195_groupi_g39237(csa_tree_add_190_195_groupi_n_9723 ,csa_tree_add_190_195_groupi_n_8212 ,csa_tree_add_190_195_groupi_n_9401);
  nor csa_tree_add_190_195_groupi_g39238(csa_tree_add_190_195_groupi_n_9722 ,csa_tree_add_190_195_groupi_n_6956 ,csa_tree_add_190_195_groupi_n_9467);
  and csa_tree_add_190_195_groupi_g39239(csa_tree_add_190_195_groupi_n_9721 ,csa_tree_add_190_195_groupi_n_6956 ,csa_tree_add_190_195_groupi_n_9467);
  or csa_tree_add_190_195_groupi_g39240(csa_tree_add_190_195_groupi_n_9720 ,csa_tree_add_190_195_groupi_n_8608 ,csa_tree_add_190_195_groupi_n_9496);
  nor csa_tree_add_190_195_groupi_g39241(csa_tree_add_190_195_groupi_n_9719 ,csa_tree_add_190_195_groupi_n_8609 ,csa_tree_add_190_195_groupi_n_9495);
  or csa_tree_add_190_195_groupi_g39242(csa_tree_add_190_195_groupi_n_9718 ,csa_tree_add_190_195_groupi_n_7714 ,csa_tree_add_190_195_groupi_n_9351);
  or csa_tree_add_190_195_groupi_g39243(csa_tree_add_190_195_groupi_n_9717 ,csa_tree_add_190_195_groupi_n_9508 ,csa_tree_add_190_195_groupi_n_9370);
  or csa_tree_add_190_195_groupi_g39244(csa_tree_add_190_195_groupi_n_9716 ,csa_tree_add_190_195_groupi_n_9037 ,csa_tree_add_190_195_groupi_n_9386);
  or csa_tree_add_190_195_groupi_g39245(csa_tree_add_190_195_groupi_n_9715 ,csa_tree_add_190_195_groupi_n_8704 ,csa_tree_add_190_195_groupi_n_9269);
  and csa_tree_add_190_195_groupi_g39246(csa_tree_add_190_195_groupi_n_9714 ,csa_tree_add_190_195_groupi_n_9527 ,csa_tree_add_190_195_groupi_n_9463);
  or csa_tree_add_190_195_groupi_g39247(csa_tree_add_190_195_groupi_n_9713 ,csa_tree_add_190_195_groupi_n_8874 ,csa_tree_add_190_195_groupi_n_9381);
  or csa_tree_add_190_195_groupi_g39248(csa_tree_add_190_195_groupi_n_9712 ,csa_tree_add_190_195_groupi_n_8876 ,csa_tree_add_190_195_groupi_n_9459);
  or csa_tree_add_190_195_groupi_g39249(csa_tree_add_190_195_groupi_n_9711 ,csa_tree_add_190_195_groupi_n_8872 ,csa_tree_add_190_195_groupi_n_9254);
  and csa_tree_add_190_195_groupi_g39250(csa_tree_add_190_195_groupi_n_9710 ,csa_tree_add_190_195_groupi_n_9375 ,csa_tree_add_190_195_groupi_n_9520);
  or csa_tree_add_190_195_groupi_g39251(csa_tree_add_190_195_groupi_n_9709 ,csa_tree_add_190_195_groupi_n_7693 ,csa_tree_add_190_195_groupi_n_9521);
  and csa_tree_add_190_195_groupi_g39252(csa_tree_add_190_195_groupi_n_9708 ,csa_tree_add_190_195_groupi_n_9071 ,csa_tree_add_190_195_groupi_n_9349);
  nor csa_tree_add_190_195_groupi_g39253(csa_tree_add_190_195_groupi_n_9707 ,csa_tree_add_190_195_groupi_n_7622 ,csa_tree_add_190_195_groupi_n_9330);
  and csa_tree_add_190_195_groupi_g39254(csa_tree_add_190_195_groupi_n_9706 ,csa_tree_add_190_195_groupi_n_7622 ,csa_tree_add_190_195_groupi_n_9330);
  or csa_tree_add_190_195_groupi_g39255(csa_tree_add_190_195_groupi_n_9705 ,csa_tree_add_190_195_groupi_n_9366 ,csa_tree_add_190_195_groupi_n_9067);
  and csa_tree_add_190_195_groupi_g39256(csa_tree_add_190_195_groupi_n_9704 ,csa_tree_add_190_195_groupi_n_7061 ,csa_tree_add_190_195_groupi_n_9286);
  nor csa_tree_add_190_195_groupi_g39257(csa_tree_add_190_195_groupi_n_9703 ,csa_tree_add_190_195_groupi_n_8628 ,csa_tree_add_190_195_groupi_n_9318);
  or csa_tree_add_190_195_groupi_g39258(csa_tree_add_190_195_groupi_n_9702 ,csa_tree_add_190_195_groupi_n_9197 ,csa_tree_add_190_195_groupi_n_9377);
  nor csa_tree_add_190_195_groupi_g39259(csa_tree_add_190_195_groupi_n_9701 ,csa_tree_add_190_195_groupi_n_7061 ,csa_tree_add_190_195_groupi_n_9286);
  or csa_tree_add_190_195_groupi_g39260(csa_tree_add_190_195_groupi_n_9700 ,csa_tree_add_190_195_groupi_n_7497 ,csa_tree_add_190_195_groupi_n_9348);
  and csa_tree_add_190_195_groupi_g39261(csa_tree_add_190_195_groupi_n_9699 ,csa_tree_add_190_195_groupi_n_7497 ,csa_tree_add_190_195_groupi_n_9348);
  or csa_tree_add_190_195_groupi_g39262(csa_tree_add_190_195_groupi_n_9698 ,csa_tree_add_190_195_groupi_n_9010 ,csa_tree_add_190_195_groupi_n_9299);
  nor csa_tree_add_190_195_groupi_g39263(csa_tree_add_190_195_groupi_n_9697 ,csa_tree_add_190_195_groupi_n_9011 ,csa_tree_add_190_195_groupi_n_9298);
  or csa_tree_add_190_195_groupi_g39264(csa_tree_add_190_195_groupi_n_9696 ,csa_tree_add_190_195_groupi_n_9195 ,csa_tree_add_190_195_groupi_n_9388);
  or csa_tree_add_190_195_groupi_g39265(csa_tree_add_190_195_groupi_n_9695 ,csa_tree_add_190_195_groupi_n_7069 ,csa_tree_add_190_195_groupi_n_9331);
  nor csa_tree_add_190_195_groupi_g39266(csa_tree_add_190_195_groupi_n_9694 ,csa_tree_add_190_195_groupi_n_7070 ,csa_tree_add_190_195_groupi_n_9332);
  or csa_tree_add_190_195_groupi_g39267(csa_tree_add_190_195_groupi_n_9693 ,csa_tree_add_190_195_groupi_n_7098 ,csa_tree_add_190_195_groupi_n_111);
  nor csa_tree_add_190_195_groupi_g39268(csa_tree_add_190_195_groupi_n_9692 ,csa_tree_add_190_195_groupi_n_7099 ,csa_tree_add_190_195_groupi_n_9327);
  or csa_tree_add_190_195_groupi_g39269(csa_tree_add_190_195_groupi_n_9691 ,csa_tree_add_190_195_groupi_n_8067 ,csa_tree_add_190_195_groupi_n_9510);
  nor csa_tree_add_190_195_groupi_g39270(csa_tree_add_190_195_groupi_n_9690 ,csa_tree_add_190_195_groupi_n_8699 ,csa_tree_add_190_195_groupi_n_9443);
  or csa_tree_add_190_195_groupi_g39271(csa_tree_add_190_195_groupi_n_9689 ,csa_tree_add_190_195_groupi_n_8849 ,csa_tree_add_190_195_groupi_n_9256);
  or csa_tree_add_190_195_groupi_g39272(csa_tree_add_190_195_groupi_n_9688 ,csa_tree_add_190_195_groupi_n_8723 ,csa_tree_add_190_195_groupi_n_9259);
  or csa_tree_add_190_195_groupi_g39273(csa_tree_add_190_195_groupi_n_9687 ,csa_tree_add_190_195_groupi_n_9127 ,csa_tree_add_190_195_groupi_n_9364);
  or csa_tree_add_190_195_groupi_g39274(csa_tree_add_190_195_groupi_n_9686 ,csa_tree_add_190_195_groupi_n_7167 ,csa_tree_add_190_195_groupi_n_9304);
  nor csa_tree_add_190_195_groupi_g39275(csa_tree_add_190_195_groupi_n_9685 ,csa_tree_add_190_195_groupi_n_7168 ,csa_tree_add_190_195_groupi_n_9305);
  or csa_tree_add_190_195_groupi_g39276(csa_tree_add_190_195_groupi_n_9684 ,csa_tree_add_190_195_groupi_n_8865 ,csa_tree_add_190_195_groupi_n_9400);
  and csa_tree_add_190_195_groupi_g39277(csa_tree_add_190_195_groupi_n_9683 ,csa_tree_add_190_195_groupi_n_8391 ,csa_tree_add_190_195_groupi_n_9280);
  nor csa_tree_add_190_195_groupi_g39278(csa_tree_add_190_195_groupi_n_9682 ,csa_tree_add_190_195_groupi_n_9308 ,csa_tree_add_190_195_groupi_n_9476);
  and csa_tree_add_190_195_groupi_g39279(csa_tree_add_190_195_groupi_n_9681 ,csa_tree_add_190_195_groupi_n_9308 ,csa_tree_add_190_195_groupi_n_9476);
  or csa_tree_add_190_195_groupi_g39280(csa_tree_add_190_195_groupi_n_9680 ,csa_tree_add_190_195_groupi_n_9165 ,csa_tree_add_190_195_groupi_n_9303);
  nor csa_tree_add_190_195_groupi_g39281(csa_tree_add_190_195_groupi_n_9679 ,csa_tree_add_190_195_groupi_n_9166 ,csa_tree_add_190_195_groupi_n_9302);
  or csa_tree_add_190_195_groupi_g39282(csa_tree_add_190_195_groupi_n_9678 ,csa_tree_add_190_195_groupi_n_9485 ,csa_tree_add_190_195_groupi_n_9500);
  nor csa_tree_add_190_195_groupi_g39283(csa_tree_add_190_195_groupi_n_9677 ,csa_tree_add_190_195_groupi_n_9486 ,csa_tree_add_190_195_groupi_n_9499);
  or csa_tree_add_190_195_groupi_g39284(csa_tree_add_190_195_groupi_n_9676 ,csa_tree_add_190_195_groupi_n_8515 ,csa_tree_add_190_195_groupi_n_9414);
  or csa_tree_add_190_195_groupi_g39285(csa_tree_add_190_195_groupi_n_9675 ,csa_tree_add_190_195_groupi_n_9009 ,csa_tree_add_190_195_groupi_n_9319);
  nor csa_tree_add_190_195_groupi_g39286(csa_tree_add_190_195_groupi_n_9674 ,csa_tree_add_190_195_groupi_n_9008 ,csa_tree_add_190_195_groupi_n_9320);
  or csa_tree_add_190_195_groupi_g39287(csa_tree_add_190_195_groupi_n_9673 ,csa_tree_add_190_195_groupi_n_9519 ,csa_tree_add_190_195_groupi_n_9258);
  or csa_tree_add_190_195_groupi_g39288(csa_tree_add_190_195_groupi_n_9672 ,csa_tree_add_190_195_groupi_n_9367 ,csa_tree_add_190_195_groupi_n_8936);
  and csa_tree_add_190_195_groupi_g39289(csa_tree_add_190_195_groupi_n_9671 ,csa_tree_add_190_195_groupi_n_9523 ,csa_tree_add_190_195_groupi_n_9434);
  or csa_tree_add_190_195_groupi_g39290(csa_tree_add_190_195_groupi_n_9670 ,csa_tree_add_190_195_groupi_n_8966 ,csa_tree_add_190_195_groupi_n_9481);
  or csa_tree_add_190_195_groupi_g39291(csa_tree_add_190_195_groupi_n_9810 ,csa_tree_add_190_195_groupi_n_7769 ,csa_tree_add_190_195_groupi_n_9433);
  or csa_tree_add_190_195_groupi_g39292(csa_tree_add_190_195_groupi_n_9808 ,csa_tree_add_190_195_groupi_n_9148 ,csa_tree_add_190_195_groupi_n_9451);
  and csa_tree_add_190_195_groupi_g39293(csa_tree_add_190_195_groupi_n_9807 ,csa_tree_add_190_195_groupi_n_8597 ,csa_tree_add_190_195_groupi_n_9444);
  or csa_tree_add_190_195_groupi_g39294(csa_tree_add_190_195_groupi_n_9806 ,csa_tree_add_190_195_groupi_n_7275 ,csa_tree_add_190_195_groupi_n_9427);
  or csa_tree_add_190_195_groupi_g39295(csa_tree_add_190_195_groupi_n_9804 ,csa_tree_add_190_195_groupi_n_7241 ,csa_tree_add_190_195_groupi_n_9380);
  and csa_tree_add_190_195_groupi_g39296(csa_tree_add_190_195_groupi_n_9803 ,csa_tree_add_190_195_groupi_n_8929 ,csa_tree_add_190_195_groupi_n_9407);
  or csa_tree_add_190_195_groupi_g39297(csa_tree_add_190_195_groupi_n_9801 ,csa_tree_add_190_195_groupi_n_6098 ,csa_tree_add_190_195_groupi_n_9378);
  and csa_tree_add_190_195_groupi_g39298(csa_tree_add_190_195_groupi_n_9800 ,csa_tree_add_190_195_groupi_n_9106 ,csa_tree_add_190_195_groupi_n_9406);
  and csa_tree_add_190_195_groupi_g39299(csa_tree_add_190_195_groupi_n_9799 ,csa_tree_add_190_195_groupi_n_8803 ,csa_tree_add_190_195_groupi_n_9449);
  or csa_tree_add_190_195_groupi_g39300(csa_tree_add_190_195_groupi_n_9798 ,csa_tree_add_190_195_groupi_n_8427 ,csa_tree_add_190_195_groupi_n_9415);
  and csa_tree_add_190_195_groupi_g39301(csa_tree_add_190_195_groupi_n_9797 ,csa_tree_add_190_195_groupi_n_9086 ,csa_tree_add_190_195_groupi_n_9383);
  and csa_tree_add_190_195_groupi_g39302(csa_tree_add_190_195_groupi_n_9796 ,csa_tree_add_190_195_groupi_n_9076 ,csa_tree_add_190_195_groupi_n_9374);
  and csa_tree_add_190_195_groupi_g39303(csa_tree_add_190_195_groupi_n_9795 ,csa_tree_add_190_195_groupi_n_9099 ,csa_tree_add_190_195_groupi_n_9397);
  and csa_tree_add_190_195_groupi_g39304(csa_tree_add_190_195_groupi_n_9794 ,csa_tree_add_190_195_groupi_n_9153 ,csa_tree_add_190_195_groupi_n_9410);
  or csa_tree_add_190_195_groupi_g39305(csa_tree_add_190_195_groupi_n_9793 ,csa_tree_add_190_195_groupi_n_7779 ,csa_tree_add_190_195_groupi_n_9411);
  and csa_tree_add_190_195_groupi_g39306(csa_tree_add_190_195_groupi_n_9792 ,csa_tree_add_190_195_groupi_n_9142 ,csa_tree_add_190_195_groupi_n_9447);
  and csa_tree_add_190_195_groupi_g39307(csa_tree_add_190_195_groupi_n_9791 ,csa_tree_add_190_195_groupi_n_6244 ,csa_tree_add_190_195_groupi_n_9405);
  or csa_tree_add_190_195_groupi_g39308(csa_tree_add_190_195_groupi_n_9790 ,csa_tree_add_190_195_groupi_n_9060 ,csa_tree_add_190_195_groupi_n_9392);
  and csa_tree_add_190_195_groupi_g39309(csa_tree_add_190_195_groupi_n_9789 ,csa_tree_add_190_195_groupi_n_8917 ,csa_tree_add_190_195_groupi_n_9394);
  and csa_tree_add_190_195_groupi_g39310(csa_tree_add_190_195_groupi_n_9788 ,csa_tree_add_190_195_groupi_n_9126 ,csa_tree_add_190_195_groupi_n_9435);
  or csa_tree_add_190_195_groupi_g39311(csa_tree_add_190_195_groupi_n_9786 ,csa_tree_add_190_195_groupi_n_9141 ,csa_tree_add_190_195_groupi_n_9446);
  or csa_tree_add_190_195_groupi_g39312(csa_tree_add_190_195_groupi_n_9785 ,csa_tree_add_190_195_groupi_n_8941 ,csa_tree_add_190_195_groupi_n_9455);
  or csa_tree_add_190_195_groupi_g39313(csa_tree_add_190_195_groupi_n_9783 ,csa_tree_add_190_195_groupi_n_9104 ,csa_tree_add_190_195_groupi_n_9371);
  or csa_tree_add_190_195_groupi_g39314(csa_tree_add_190_195_groupi_n_9781 ,csa_tree_add_190_195_groupi_n_9151 ,csa_tree_add_190_195_groupi_n_9404);
  or csa_tree_add_190_195_groupi_g39315(csa_tree_add_190_195_groupi_n_9780 ,csa_tree_add_190_195_groupi_n_9121 ,csa_tree_add_190_195_groupi_n_9424);
  or csa_tree_add_190_195_groupi_g39316(csa_tree_add_190_195_groupi_n_9779 ,csa_tree_add_190_195_groupi_n_8461 ,csa_tree_add_190_195_groupi_n_9385);
  or csa_tree_add_190_195_groupi_g39317(csa_tree_add_190_195_groupi_n_9777 ,csa_tree_add_190_195_groupi_n_8447 ,csa_tree_add_190_195_groupi_n_9437);
  and csa_tree_add_190_195_groupi_g39318(csa_tree_add_190_195_groupi_n_9776 ,csa_tree_add_190_195_groupi_n_7957 ,csa_tree_add_190_195_groupi_n_9408);
  or csa_tree_add_190_195_groupi_g39319(csa_tree_add_190_195_groupi_n_9775 ,csa_tree_add_190_195_groupi_n_8921 ,csa_tree_add_190_195_groupi_n_9373);
  and csa_tree_add_190_195_groupi_g39320(csa_tree_add_190_195_groupi_n_9772 ,csa_tree_add_190_195_groupi_n_9130 ,csa_tree_add_190_195_groupi_n_9439);
  or csa_tree_add_190_195_groupi_g39321(csa_tree_add_190_195_groupi_n_9771 ,csa_tree_add_190_195_groupi_n_9074 ,csa_tree_add_190_195_groupi_n_9441);
  and csa_tree_add_190_195_groupi_g39322(csa_tree_add_190_195_groupi_n_9769 ,csa_tree_add_190_195_groupi_n_9154 ,csa_tree_add_190_195_groupi_n_9460);
  or csa_tree_add_190_195_groupi_g39323(csa_tree_add_190_195_groupi_n_9768 ,csa_tree_add_190_195_groupi_n_9059 ,csa_tree_add_190_195_groupi_n_9390);
  or csa_tree_add_190_195_groupi_g39324(csa_tree_add_190_195_groupi_n_9765 ,csa_tree_add_190_195_groupi_n_9128 ,csa_tree_add_190_195_groupi_n_9436);
  and csa_tree_add_190_195_groupi_g39325(csa_tree_add_190_195_groupi_n_9764 ,csa_tree_add_190_195_groupi_n_9090 ,csa_tree_add_190_195_groupi_n_9389);
  or csa_tree_add_190_195_groupi_g39326(csa_tree_add_190_195_groupi_n_9763 ,csa_tree_add_190_195_groupi_n_9084 ,csa_tree_add_190_195_groupi_n_9384);
  and csa_tree_add_190_195_groupi_g39327(csa_tree_add_190_195_groupi_n_9760 ,csa_tree_add_190_195_groupi_n_9132 ,csa_tree_add_190_195_groupi_n_9440);
  or csa_tree_add_190_195_groupi_g39328(csa_tree_add_190_195_groupi_n_9759 ,csa_tree_add_190_195_groupi_n_8918 ,csa_tree_add_190_195_groupi_n_9398);
  or csa_tree_add_190_195_groupi_g39329(csa_tree_add_190_195_groupi_n_9757 ,csa_tree_add_190_195_groupi_n_8142 ,csa_tree_add_190_195_groupi_n_9438);
  or csa_tree_add_190_195_groupi_g39330(csa_tree_add_190_195_groupi_n_9755 ,csa_tree_add_190_195_groupi_n_9055 ,csa_tree_add_190_195_groupi_n_9425);
  and csa_tree_add_190_195_groupi_g39331(csa_tree_add_190_195_groupi_n_9754 ,csa_tree_add_190_195_groupi_n_9063 ,csa_tree_add_190_195_groupi_n_9376);
  and csa_tree_add_190_195_groupi_g39332(csa_tree_add_190_195_groupi_n_9753 ,csa_tree_add_190_195_groupi_n_9113 ,csa_tree_add_190_195_groupi_n_9412);
  and csa_tree_add_190_195_groupi_g39333(csa_tree_add_190_195_groupi_n_9750 ,csa_tree_add_190_195_groupi_n_8143 ,csa_tree_add_190_195_groupi_n_9395);
  not csa_tree_add_190_195_groupi_g39335(csa_tree_add_190_195_groupi_n_9664 ,csa_tree_add_190_195_groupi_n_9663);
  not csa_tree_add_190_195_groupi_g39336(csa_tree_add_190_195_groupi_n_9661 ,csa_tree_add_190_195_groupi_n_9660);
  not csa_tree_add_190_195_groupi_g39338(csa_tree_add_190_195_groupi_n_9649 ,csa_tree_add_190_195_groupi_n_9648);
  not csa_tree_add_190_195_groupi_g39339(csa_tree_add_190_195_groupi_n_9647 ,csa_tree_add_190_195_groupi_n_9646);
  not csa_tree_add_190_195_groupi_g39340(csa_tree_add_190_195_groupi_n_9645 ,csa_tree_add_190_195_groupi_n_9644);
  not csa_tree_add_190_195_groupi_g39341(csa_tree_add_190_195_groupi_n_9643 ,csa_tree_add_190_195_groupi_n_9642);
  not csa_tree_add_190_195_groupi_g39342(csa_tree_add_190_195_groupi_n_9641 ,csa_tree_add_190_195_groupi_n_117);
  not csa_tree_add_190_195_groupi_g39343(csa_tree_add_190_195_groupi_n_9638 ,csa_tree_add_190_195_groupi_n_9637);
  not csa_tree_add_190_195_groupi_g39344(csa_tree_add_190_195_groupi_n_9635 ,csa_tree_add_190_195_groupi_n_9636);
  not csa_tree_add_190_195_groupi_g39345(csa_tree_add_190_195_groupi_n_9634 ,csa_tree_add_190_195_groupi_n_9633);
  not csa_tree_add_190_195_groupi_g39346(csa_tree_add_190_195_groupi_n_9632 ,csa_tree_add_190_195_groupi_n_9631);
  not csa_tree_add_190_195_groupi_g39347(csa_tree_add_190_195_groupi_n_9630 ,csa_tree_add_190_195_groupi_n_9629);
  not csa_tree_add_190_195_groupi_g39348(csa_tree_add_190_195_groupi_n_9628 ,csa_tree_add_190_195_groupi_n_9627);
  not csa_tree_add_190_195_groupi_g39349(csa_tree_add_190_195_groupi_n_9623 ,csa_tree_add_190_195_groupi_n_9624);
  not csa_tree_add_190_195_groupi_g39350(csa_tree_add_190_195_groupi_n_9622 ,csa_tree_add_190_195_groupi_n_9621);
  not csa_tree_add_190_195_groupi_g39351(csa_tree_add_190_195_groupi_n_9620 ,csa_tree_add_190_195_groupi_n_110);
  not csa_tree_add_190_195_groupi_g39352(csa_tree_add_190_195_groupi_n_9619 ,csa_tree_add_190_195_groupi_n_9618);
  not csa_tree_add_190_195_groupi_g39353(csa_tree_add_190_195_groupi_n_9617 ,csa_tree_add_190_195_groupi_n_9616);
  not csa_tree_add_190_195_groupi_g39354(csa_tree_add_190_195_groupi_n_9615 ,csa_tree_add_190_195_groupi_n_9614);
  not csa_tree_add_190_195_groupi_g39355(csa_tree_add_190_195_groupi_n_9613 ,csa_tree_add_190_195_groupi_n_9612);
  not csa_tree_add_190_195_groupi_g39356(csa_tree_add_190_195_groupi_n_9611 ,csa_tree_add_190_195_groupi_n_9610);
  not csa_tree_add_190_195_groupi_g39357(csa_tree_add_190_195_groupi_n_9609 ,csa_tree_add_190_195_groupi_n_9608);
  not csa_tree_add_190_195_groupi_g39358(csa_tree_add_190_195_groupi_n_9605 ,csa_tree_add_190_195_groupi_n_9606);
  not csa_tree_add_190_195_groupi_g39359(csa_tree_add_190_195_groupi_n_9602 ,csa_tree_add_190_195_groupi_n_9601);
  nor csa_tree_add_190_195_groupi_g39360(csa_tree_add_190_195_groupi_n_9600 ,csa_tree_add_190_195_groupi_n_9025 ,csa_tree_add_190_195_groupi_n_9296);
  or csa_tree_add_190_195_groupi_g39361(csa_tree_add_190_195_groupi_n_9599 ,csa_tree_add_190_195_groupi_n_9024 ,csa_tree_add_190_195_groupi_n_9297);
  nor csa_tree_add_190_195_groupi_g39362(csa_tree_add_190_195_groupi_n_9598 ,csa_tree_add_190_195_groupi_n_9491 ,csa_tree_add_190_195_groupi_n_9015);
  nor csa_tree_add_190_195_groupi_g39363(csa_tree_add_190_195_groupi_n_9597 ,csa_tree_add_190_195_groupi_n_8840 ,csa_tree_add_190_195_groupi_n_9313);
  or csa_tree_add_190_195_groupi_g39364(csa_tree_add_190_195_groupi_n_9596 ,csa_tree_add_190_195_groupi_n_8839 ,csa_tree_add_190_195_groupi_n_9312);
  or csa_tree_add_190_195_groupi_g39365(csa_tree_add_190_195_groupi_n_9595 ,csa_tree_add_190_195_groupi_n_8518 ,csa_tree_add_190_195_groupi_n_9420);
  or csa_tree_add_190_195_groupi_g39366(csa_tree_add_190_195_groupi_n_9594 ,csa_tree_add_190_195_groupi_n_8636 ,csa_tree_add_190_195_groupi_n_9323);
  nor csa_tree_add_190_195_groupi_g39367(csa_tree_add_190_195_groupi_n_9593 ,csa_tree_add_190_195_groupi_n_8637 ,csa_tree_add_190_195_groupi_n_9324);
  or csa_tree_add_190_195_groupi_g39368(csa_tree_add_190_195_groupi_n_9592 ,csa_tree_add_190_195_groupi_n_9517 ,csa_tree_add_190_195_groupi_n_9278);
  or csa_tree_add_190_195_groupi_g39369(csa_tree_add_190_195_groupi_n_9591 ,csa_tree_add_190_195_groupi_n_8854 ,csa_tree_add_190_195_groupi_n_9276);
  or csa_tree_add_190_195_groupi_g39370(csa_tree_add_190_195_groupi_n_9590 ,csa_tree_add_190_195_groupi_n_9353 ,csa_tree_add_190_195_groupi_n_8925);
  nor csa_tree_add_190_195_groupi_g39371(csa_tree_add_190_195_groupi_n_9589 ,csa_tree_add_190_195_groupi_n_9285 ,csa_tree_add_190_195_groupi_n_9028);
  or csa_tree_add_190_195_groupi_g39372(csa_tree_add_190_195_groupi_n_9588 ,csa_tree_add_190_195_groupi_n_9284 ,csa_tree_add_190_195_groupi_n_9029);
  or csa_tree_add_190_195_groupi_g39373(csa_tree_add_190_195_groupi_n_9587 ,csa_tree_add_190_195_groupi_n_9492 ,csa_tree_add_190_195_groupi_n_9014);
  or csa_tree_add_190_195_groupi_g39374(csa_tree_add_190_195_groupi_n_9586 ,csa_tree_add_190_195_groupi_n_7949 ,csa_tree_add_190_195_groupi_n_9357);
  or csa_tree_add_190_195_groupi_g39375(csa_tree_add_190_195_groupi_n_9585 ,csa_tree_add_190_195_groupi_n_9198 ,csa_tree_add_190_195_groupi_n_9275);
  nor csa_tree_add_190_195_groupi_g39376(csa_tree_add_190_195_groupi_n_9584 ,csa_tree_add_190_195_groupi_n_9505 ,csa_tree_add_190_195_groupi_n_9267);
  or csa_tree_add_190_195_groupi_g39377(csa_tree_add_190_195_groupi_n_9583 ,csa_tree_add_190_195_groupi_n_9347 ,csa_tree_add_190_195_groupi_n_9333);
  or csa_tree_add_190_195_groupi_g39378(csa_tree_add_190_195_groupi_n_9582 ,csa_tree_add_190_195_groupi_n_8816 ,csa_tree_add_190_195_groupi_n_9315);
  nor csa_tree_add_190_195_groupi_g39379(csa_tree_add_190_195_groupi_n_9581 ,csa_tree_add_190_195_groupi_n_8817 ,csa_tree_add_190_195_groupi_n_9316);
  or csa_tree_add_190_195_groupi_g39380(csa_tree_add_190_195_groupi_n_9580 ,csa_tree_add_190_195_groupi_n_6909 ,csa_tree_add_190_195_groupi_n_9343);
  or csa_tree_add_190_195_groupi_g39381(csa_tree_add_190_195_groupi_n_9579 ,csa_tree_add_190_195_groupi_n_9525 ,csa_tree_add_190_195_groupi_n_9262);
  or csa_tree_add_190_195_groupi_g39382(csa_tree_add_190_195_groupi_n_9578 ,csa_tree_add_190_195_groupi_n_8978 ,csa_tree_add_190_195_groupi_n_9335);
  nor csa_tree_add_190_195_groupi_g39383(csa_tree_add_190_195_groupi_n_9577 ,csa_tree_add_190_195_groupi_n_8979 ,csa_tree_add_190_195_groupi_n_9336);
  nor csa_tree_add_190_195_groupi_g39384(csa_tree_add_190_195_groupi_n_9576 ,csa_tree_add_190_195_groupi_n_120 ,csa_tree_add_190_195_groupi_n_9334);
  nor csa_tree_add_190_195_groupi_g39385(csa_tree_add_190_195_groupi_n_9575 ,csa_tree_add_190_195_groupi_n_8862 ,csa_tree_add_190_195_groupi_n_9274);
  nor csa_tree_add_190_195_groupi_g39386(csa_tree_add_190_195_groupi_n_9574 ,csa_tree_add_190_195_groupi_n_7980 ,csa_tree_add_190_195_groupi_n_9469);
  and csa_tree_add_190_195_groupi_g39387(csa_tree_add_190_195_groupi_n_9573 ,csa_tree_add_190_195_groupi_n_7980 ,csa_tree_add_190_195_groupi_n_9469);
  and csa_tree_add_190_195_groupi_g39388(csa_tree_add_190_195_groupi_n_9572 ,csa_tree_add_190_195_groupi_n_7477 ,csa_tree_add_190_195_groupi_n_9360);
  nor csa_tree_add_190_195_groupi_g39389(csa_tree_add_190_195_groupi_n_9571 ,csa_tree_add_190_195_groupi_n_6908 ,csa_tree_add_190_195_groupi_n_9344);
  and csa_tree_add_190_195_groupi_g39390(csa_tree_add_190_195_groupi_n_9570 ,csa_tree_add_190_195_groupi_n_8966 ,csa_tree_add_190_195_groupi_n_9481);
  xnor csa_tree_add_190_195_groupi_g39391(csa_tree_add_190_195_groupi_n_9569 ,csa_tree_add_190_195_groupi_n_7560 ,csa_tree_add_190_195_groupi_n_9042);
  xnor csa_tree_add_190_195_groupi_g39392(csa_tree_add_190_195_groupi_n_9568 ,csa_tree_add_190_195_groupi_n_7352 ,csa_tree_add_190_195_groupi_n_9038);
  xnor csa_tree_add_190_195_groupi_g39393(csa_tree_add_190_195_groupi_n_9567 ,csa_tree_add_190_195_groupi_n_7099 ,csa_tree_add_190_195_groupi_n_9201);
  xnor csa_tree_add_190_195_groupi_g39394(csa_tree_add_190_195_groupi_n_9566 ,csa_tree_add_190_195_groupi_n_8484 ,csa_tree_add_190_195_groupi_n_8965);
  xnor csa_tree_add_190_195_groupi_g39395(csa_tree_add_190_195_groupi_n_9565 ,csa_tree_add_190_195_groupi_n_8825 ,csa_tree_add_190_195_groupi_n_9023);
  xnor csa_tree_add_190_195_groupi_g39396(csa_tree_add_190_195_groupi_n_9564 ,csa_tree_add_190_195_groupi_n_8518 ,csa_tree_add_190_195_groupi_n_9005);
  xnor csa_tree_add_190_195_groupi_g39397(csa_tree_add_190_195_groupi_n_9563 ,csa_tree_add_190_195_groupi_n_7376 ,csa_tree_add_190_195_groupi_n_9199);
  xnor csa_tree_add_190_195_groupi_g39398(csa_tree_add_190_195_groupi_n_9562 ,csa_tree_add_190_195_groupi_n_7496 ,csa_tree_add_190_195_groupi_n_9193);
  xnor csa_tree_add_190_195_groupi_g39399(csa_tree_add_190_195_groupi_n_9561 ,csa_tree_add_190_195_groupi_n_7983 ,csa_tree_add_190_195_groupi_n_8962);
  xnor csa_tree_add_190_195_groupi_g39400(csa_tree_add_190_195_groupi_n_9560 ,csa_tree_add_190_195_groupi_n_9179 ,csa_tree_add_190_195_groupi_n_9037);
  xnor csa_tree_add_190_195_groupi_g39402(csa_tree_add_190_195_groupi_n_9559 ,csa_tree_add_190_195_groupi_n_5964 ,csa_tree_add_190_195_groupi_n_9048);
  xnor csa_tree_add_190_195_groupi_g39404(csa_tree_add_190_195_groupi_n_9558 ,csa_tree_add_190_195_groupi_n_8366 ,csa_tree_add_190_195_groupi_n_9158);
  xnor csa_tree_add_190_195_groupi_g39405(csa_tree_add_190_195_groupi_n_9557 ,csa_tree_add_190_195_groupi_n_9162 ,csa_tree_add_190_195_groupi_n_8959);
  xnor csa_tree_add_190_195_groupi_g39406(csa_tree_add_190_195_groupi_n_9556 ,csa_tree_add_190_195_groupi_n_8389 ,csa_tree_add_190_195_groupi_n_9173);
  xnor csa_tree_add_190_195_groupi_g39407(csa_tree_add_190_195_groupi_n_9555 ,csa_tree_add_190_195_groupi_n_8011 ,csa_tree_add_190_195_groupi_n_8971);
  xnor csa_tree_add_190_195_groupi_g39408(csa_tree_add_190_195_groupi_n_9554 ,csa_tree_add_190_195_groupi_n_8865 ,csa_tree_add_190_195_groupi_n_8949);
  xnor csa_tree_add_190_195_groupi_g39409(csa_tree_add_190_195_groupi_n_9553 ,csa_tree_add_190_195_groupi_n_8843 ,csa_tree_add_190_195_groupi_n_8968);
  xnor csa_tree_add_190_195_groupi_g39410(csa_tree_add_190_195_groupi_n_9552 ,csa_tree_add_190_195_groupi_n_8004 ,csa_tree_add_190_195_groupi_n_9200);
  xnor csa_tree_add_190_195_groupi_g39411(csa_tree_add_190_195_groupi_n_9551 ,csa_tree_add_190_195_groupi_n_7189 ,csa_tree_add_190_195_groupi_n_9039);
  xnor csa_tree_add_190_195_groupi_g39412(csa_tree_add_190_195_groupi_n_9550 ,csa_tree_add_190_195_groupi_n_8987 ,csa_tree_add_190_195_groupi_n_9027);
  xnor csa_tree_add_190_195_groupi_g39413(csa_tree_add_190_195_groupi_n_9549 ,csa_tree_add_190_195_groupi_n_8969 ,csa_tree_add_190_195_groupi_n_8845);
  xnor csa_tree_add_190_195_groupi_g39414(csa_tree_add_190_195_groupi_n_9548 ,csa_tree_add_190_195_groupi_n_7512 ,csa_tree_add_190_195_groupi_n_9044);
  xnor csa_tree_add_190_195_groupi_g39415(csa_tree_add_190_195_groupi_n_9547 ,csa_tree_add_190_195_groupi_n_8975 ,csa_tree_add_190_195_groupi_n_7353);
  xnor csa_tree_add_190_195_groupi_g39416(csa_tree_add_190_195_groupi_n_9546 ,csa_tree_add_190_195_groupi_n_8332 ,csa_tree_add_190_195_groupi_n_8947);
  xnor csa_tree_add_190_195_groupi_g39417(csa_tree_add_190_195_groupi_n_9545 ,csa_tree_add_190_195_groupi_n_7984 ,csa_tree_add_190_195_groupi_n_8960);
  xnor csa_tree_add_190_195_groupi_g39418(csa_tree_add_190_195_groupi_n_9544 ,csa_tree_add_190_195_groupi_n_8334 ,csa_tree_add_190_195_groupi_n_8977);
  xnor csa_tree_add_190_195_groupi_g39420(csa_tree_add_190_195_groupi_n_9543 ,csa_tree_add_190_195_groupi_n_9034 ,csa_tree_add_190_195_groupi_n_9032);
  xnor csa_tree_add_190_195_groupi_g39421(csa_tree_add_190_195_groupi_n_9542 ,csa_tree_add_190_195_groupi_n_8681 ,csa_tree_add_190_195_groupi_n_9182);
  xnor csa_tree_add_190_195_groupi_g39422(csa_tree_add_190_195_groupi_n_9541 ,csa_tree_add_190_195_groupi_n_8813 ,csa_tree_add_190_195_groupi_n_8995);
  xnor csa_tree_add_190_195_groupi_g39423(csa_tree_add_190_195_groupi_n_9540 ,csa_tree_add_190_195_groupi_n_8817 ,csa_tree_add_190_195_groupi_n_9183);
  xnor csa_tree_add_190_195_groupi_g39424(csa_tree_add_190_195_groupi_n_9539 ,csa_tree_add_190_195_groupi_n_8815 ,csa_tree_add_190_195_groupi_n_8988);
  xnor csa_tree_add_190_195_groupi_g39425(csa_tree_add_190_195_groupi_n_9538 ,csa_tree_add_190_195_groupi_n_8668 ,csa_tree_add_190_195_groupi_n_8981);
  xnor csa_tree_add_190_195_groupi_g39426(csa_tree_add_190_195_groupi_n_9537 ,csa_tree_add_190_195_groupi_n_9019 ,csa_tree_add_190_195_groupi_n_8951);
  xnor csa_tree_add_190_195_groupi_g39427(csa_tree_add_190_195_groupi_n_9536 ,csa_tree_add_190_195_groupi_n_8842 ,csa_tree_add_190_195_groupi_n_8979);
  xnor csa_tree_add_190_195_groupi_g39429(csa_tree_add_190_195_groupi_n_9535 ,csa_tree_add_190_195_groupi_n_8658 ,csa_tree_add_190_195_groupi_n_9052);
  xnor csa_tree_add_190_195_groupi_g39430(csa_tree_add_190_195_groupi_n_9534 ,csa_tree_add_190_195_groupi_n_7589 ,csa_tree_add_190_195_groupi_n_8973);
  xnor csa_tree_add_190_195_groupi_g39431(csa_tree_add_190_195_groupi_n_9533 ,csa_tree_add_190_195_groupi_n_5193 ,csa_tree_add_190_195_groupi_n_9045);
  xnor csa_tree_add_190_195_groupi_g39432(csa_tree_add_190_195_groupi_n_9532 ,csa_tree_add_190_195_groupi_n_8723 ,csa_tree_add_190_195_groupi_n_8997);
  xnor csa_tree_add_190_195_groupi_g39433(csa_tree_add_190_195_groupi_n_9531 ,csa_tree_add_190_195_groupi_n_8834 ,csa_tree_add_190_195_groupi_n_9191);
  xnor csa_tree_add_190_195_groupi_g39434(csa_tree_add_190_195_groupi_n_9530 ,csa_tree_add_190_195_groupi_n_9188 ,csa_tree_add_190_195_groupi_n_7622);
  xnor csa_tree_add_190_195_groupi_g39435(csa_tree_add_190_195_groupi_n_9529 ,csa_tree_add_190_195_groupi_n_8336 ,csa_tree_add_190_195_groupi_n_8985);
  xnor csa_tree_add_190_195_groupi_g39436(csa_tree_add_190_195_groupi_n_9528 ,csa_tree_add_190_195_groupi_n_5253 ,csa_tree_add_190_195_groupi_n_25);
  and csa_tree_add_190_195_groupi_g39437(csa_tree_add_190_195_groupi_n_9669 ,csa_tree_add_190_195_groupi_n_7476 ,csa_tree_add_190_195_groupi_n_9442);
  and csa_tree_add_190_195_groupi_g39438(csa_tree_add_190_195_groupi_n_9668 ,csa_tree_add_190_195_groupi_n_7959 ,csa_tree_add_190_195_groupi_n_9264);
  xnor csa_tree_add_190_195_groupi_g39439(csa_tree_add_190_195_groupi_n_9667 ,csa_tree_add_190_195_groupi_n_64 ,csa_tree_add_190_195_groupi_n_8885);
  xnor csa_tree_add_190_195_groupi_g39440(csa_tree_add_190_195_groupi_n_9666 ,csa_tree_add_190_195_groupi_n_5301 ,csa_tree_add_190_195_groupi_n_8904);
  and csa_tree_add_190_195_groupi_g39441(csa_tree_add_190_195_groupi_n_9665 ,csa_tree_add_190_195_groupi_n_7747 ,csa_tree_add_190_195_groupi_n_9445);
  xnor csa_tree_add_190_195_groupi_g39442(csa_tree_add_190_195_groupi_n_9663 ,csa_tree_add_190_195_groupi_n_8543 ,csa_tree_add_190_195_groupi_n_8903);
  xnor csa_tree_add_190_195_groupi_g39443(csa_tree_add_190_195_groupi_n_9662 ,csa_tree_add_190_195_groupi_n_7612 ,csa_tree_add_190_195_groupi_n_116);
  xnor csa_tree_add_190_195_groupi_g39444(csa_tree_add_190_195_groupi_n_9660 ,csa_tree_add_190_195_groupi_n_9040 ,csa_tree_add_190_195_groupi_n_7916);
  xnor csa_tree_add_190_195_groupi_g39445(csa_tree_add_190_195_groupi_n_9659 ,csa_tree_add_190_195_groupi_n_7979 ,csa_tree_add_190_195_groupi_n_8895);
  xnor csa_tree_add_190_195_groupi_g39446(csa_tree_add_190_195_groupi_n_9658 ,csa_tree_add_190_195_groupi_n_8714 ,csa_tree_add_190_195_groupi_n_8888);
  xnor csa_tree_add_190_195_groupi_g39447(csa_tree_add_190_195_groupi_n_9657 ,csa_tree_add_190_195_groupi_n_5200 ,csa_tree_add_190_195_groupi_n_8902);
  xnor csa_tree_add_190_195_groupi_g39448(csa_tree_add_190_195_groupi_n_9656 ,csa_tree_add_190_195_groupi_n_7362 ,csa_tree_add_190_195_groupi_n_8900);
  xnor csa_tree_add_190_195_groupi_g39449(csa_tree_add_190_195_groupi_n_9655 ,csa_tree_add_190_195_groupi_n_4994 ,csa_tree_add_190_195_groupi_n_8908);
  xnor csa_tree_add_190_195_groupi_g39450(csa_tree_add_190_195_groupi_n_9654 ,csa_tree_add_190_195_groupi_n_4625 ,csa_tree_add_190_195_groupi_n_8879);
  xnor csa_tree_add_190_195_groupi_g39451(csa_tree_add_190_195_groupi_n_9653 ,csa_tree_add_190_195_groupi_n_7841 ,csa_tree_add_190_195_groupi_n_115);
  and csa_tree_add_190_195_groupi_g39452(csa_tree_add_190_195_groupi_n_9652 ,csa_tree_add_190_195_groupi_n_8932 ,csa_tree_add_190_195_groupi_n_9465);
  xnor csa_tree_add_190_195_groupi_g39453(csa_tree_add_190_195_groupi_n_9651 ,csa_tree_add_190_195_groupi_n_9036 ,csa_tree_add_190_195_groupi_n_6613);
  and csa_tree_add_190_195_groupi_g39454(csa_tree_add_190_195_groupi_n_9650 ,csa_tree_add_190_195_groupi_n_8919 ,csa_tree_add_190_195_groupi_n_9266);
  xnor csa_tree_add_190_195_groupi_g39455(csa_tree_add_190_195_groupi_n_9648 ,csa_tree_add_190_195_groupi_n_7096 ,csa_tree_add_190_195_groupi_n_8907);
  xnor csa_tree_add_190_195_groupi_g39456(csa_tree_add_190_195_groupi_n_9646 ,csa_tree_add_190_195_groupi_n_7336 ,csa_tree_add_190_195_groupi_n_8878);
  xnor csa_tree_add_190_195_groupi_g39457(csa_tree_add_190_195_groupi_n_9644 ,csa_tree_add_190_195_groupi_n_9185 ,csa_tree_add_190_195_groupi_n_7461);
  xnor csa_tree_add_190_195_groupi_g39458(csa_tree_add_190_195_groupi_n_9642 ,csa_tree_add_190_195_groupi_n_7090 ,csa_tree_add_190_195_groupi_n_8887);
  and csa_tree_add_190_195_groupi_g39460(csa_tree_add_190_195_groupi_n_9640 ,csa_tree_add_190_195_groupi_n_8934 ,csa_tree_add_190_195_groupi_n_9448);
  xnor csa_tree_add_190_195_groupi_g39461(csa_tree_add_190_195_groupi_n_9639 ,csa_tree_add_190_195_groupi_n_8387 ,csa_tree_add_190_195_groupi_n_8891);
  xnor csa_tree_add_190_195_groupi_g39462(csa_tree_add_190_195_groupi_n_9637 ,csa_tree_add_190_195_groupi_n_9202 ,csa_tree_add_190_195_groupi_n_7917);
  xnor csa_tree_add_190_195_groupi_g39463(csa_tree_add_190_195_groupi_n_9636 ,csa_tree_add_190_195_groupi_n_7520 ,csa_tree_add_190_195_groupi_n_8910);
  xnor csa_tree_add_190_195_groupi_g39464(csa_tree_add_190_195_groupi_n_9633 ,csa_tree_add_190_195_groupi_n_8494 ,csa_tree_add_190_195_groupi_n_8906);
  xnor csa_tree_add_190_195_groupi_g39465(csa_tree_add_190_195_groupi_n_9631 ,csa_tree_add_190_195_groupi_n_8319 ,csa_tree_add_190_195_groupi_n_8893);
  xnor csa_tree_add_190_195_groupi_g39466(csa_tree_add_190_195_groupi_n_9629 ,csa_tree_add_190_195_groupi_n_7839 ,csa_tree_add_190_195_groupi_n_8899);
  xnor csa_tree_add_190_195_groupi_g39467(csa_tree_add_190_195_groupi_n_9627 ,csa_tree_add_190_195_groupi_n_8662 ,csa_tree_add_190_195_groupi_n_8884);
  xnor csa_tree_add_190_195_groupi_g39468(csa_tree_add_190_195_groupi_n_9626 ,csa_tree_add_190_195_groupi_n_6767 ,csa_tree_add_190_195_groupi_n_8912);
  xnor csa_tree_add_190_195_groupi_g39469(csa_tree_add_190_195_groupi_n_9625 ,csa_tree_add_190_195_groupi_n_8632 ,csa_tree_add_190_195_groupi_n_8898);
  xnor csa_tree_add_190_195_groupi_g39470(csa_tree_add_190_195_groupi_n_9624 ,csa_tree_add_190_195_groupi_n_8523 ,csa_tree_add_190_195_groupi_n_8880);
  xnor csa_tree_add_190_195_groupi_g39471(csa_tree_add_190_195_groupi_n_9621 ,csa_tree_add_190_195_groupi_n_8823 ,csa_tree_add_190_195_groupi_n_99);
  xnor csa_tree_add_190_195_groupi_g39473(csa_tree_add_190_195_groupi_n_9618 ,csa_tree_add_190_195_groupi_n_9190 ,csa_tree_add_190_195_groupi_n_8266);
  xnor csa_tree_add_190_195_groupi_g39474(csa_tree_add_190_195_groupi_n_9616 ,csa_tree_add_190_195_groupi_n_8374 ,csa_tree_add_190_195_groupi_n_118);
  xnor csa_tree_add_190_195_groupi_g39475(csa_tree_add_190_195_groupi_n_9614 ,csa_tree_add_190_195_groupi_n_8023 ,csa_tree_add_190_195_groupi_n_8890);
  and csa_tree_add_190_195_groupi_g39476(csa_tree_add_190_195_groupi_n_9612 ,csa_tree_add_190_195_groupi_n_8923 ,csa_tree_add_190_195_groupi_n_9273);
  xnor csa_tree_add_190_195_groupi_g39477(csa_tree_add_190_195_groupi_n_9610 ,csa_tree_add_190_195_groupi_n_8019 ,csa_tree_add_190_195_groupi_n_8883);
  xnor csa_tree_add_190_195_groupi_g39478(csa_tree_add_190_195_groupi_n_9608 ,csa_tree_add_190_195_groupi_n_6936 ,csa_tree_add_190_195_groupi_n_8889);
  xnor csa_tree_add_190_195_groupi_g39479(csa_tree_add_190_195_groupi_n_9607 ,csa_tree_add_190_195_groupi_n_8383 ,csa_tree_add_190_195_groupi_n_8905);
  xnor csa_tree_add_190_195_groupi_g39480(csa_tree_add_190_195_groupi_n_9606 ,csa_tree_add_190_195_groupi_n_7517 ,csa_tree_add_190_195_groupi_n_8901);
  xnor csa_tree_add_190_195_groupi_g39481(csa_tree_add_190_195_groupi_n_9604 ,csa_tree_add_190_195_groupi_n_8040 ,csa_tree_add_190_195_groupi_n_8892);
  xnor csa_tree_add_190_195_groupi_g39482(csa_tree_add_190_195_groupi_n_9603 ,csa_tree_add_190_195_groupi_n_8697 ,csa_tree_add_190_195_groupi_n_8881);
  xnor csa_tree_add_190_195_groupi_g39483(csa_tree_add_190_195_groupi_n_9601 ,csa_tree_add_190_195_groupi_n_7995 ,csa_tree_add_190_195_groupi_n_8897);
  not csa_tree_add_190_195_groupi_g39484(csa_tree_add_190_195_groupi_n_9525 ,csa_tree_add_190_195_groupi_n_9524);
  not csa_tree_add_190_195_groupi_g39485(csa_tree_add_190_195_groupi_n_9517 ,csa_tree_add_190_195_groupi_n_9516);
  not csa_tree_add_190_195_groupi_g39486(csa_tree_add_190_195_groupi_n_9510 ,csa_tree_add_190_195_groupi_n_9509);
  not csa_tree_add_190_195_groupi_g39487(csa_tree_add_190_195_groupi_n_9503 ,csa_tree_add_190_195_groupi_n_9502);
  not csa_tree_add_190_195_groupi_g39488(csa_tree_add_190_195_groupi_n_9499 ,csa_tree_add_190_195_groupi_n_9500);
  not csa_tree_add_190_195_groupi_g39489(csa_tree_add_190_195_groupi_n_9498 ,csa_tree_add_190_195_groupi_n_9497);
  not csa_tree_add_190_195_groupi_g39490(csa_tree_add_190_195_groupi_n_9495 ,csa_tree_add_190_195_groupi_n_9496);
  not csa_tree_add_190_195_groupi_g39491(csa_tree_add_190_195_groupi_n_9494 ,csa_tree_add_190_195_groupi_n_9493);
  not csa_tree_add_190_195_groupi_g39492(csa_tree_add_190_195_groupi_n_9492 ,csa_tree_add_190_195_groupi_n_9491);
  not csa_tree_add_190_195_groupi_g39493(csa_tree_add_190_195_groupi_n_9489 ,csa_tree_add_190_195_groupi_n_9490);
  not csa_tree_add_190_195_groupi_g39494(csa_tree_add_190_195_groupi_n_9487 ,csa_tree_add_190_195_groupi_n_9488);
  not csa_tree_add_190_195_groupi_g39495(csa_tree_add_190_195_groupi_n_9485 ,csa_tree_add_190_195_groupi_n_9486);
  not csa_tree_add_190_195_groupi_g39496(csa_tree_add_190_195_groupi_n_9483 ,csa_tree_add_190_195_groupi_n_9484);
  not csa_tree_add_190_195_groupi_g39497(csa_tree_add_190_195_groupi_n_9481 ,csa_tree_add_190_195_groupi_n_9480);
  not csa_tree_add_190_195_groupi_g39498(csa_tree_add_190_195_groupi_n_9479 ,csa_tree_add_190_195_groupi_n_9478);
  not csa_tree_add_190_195_groupi_g39499(csa_tree_add_190_195_groupi_n_9475 ,csa_tree_add_190_195_groupi_n_9474);
  not csa_tree_add_190_195_groupi_g39500(csa_tree_add_190_195_groupi_n_9472 ,csa_tree_add_190_195_groupi_n_9473);
  not csa_tree_add_190_195_groupi_g39501(csa_tree_add_190_195_groupi_n_9471 ,csa_tree_add_190_195_groupi_n_9470);
  not csa_tree_add_190_195_groupi_g39502(csa_tree_add_190_195_groupi_n_9469 ,csa_tree_add_190_195_groupi_n_9468);
  nor csa_tree_add_190_195_groupi_g39504(csa_tree_add_190_195_groupi_n_9466 ,csa_tree_add_190_195_groupi_n_8333 ,csa_tree_add_190_195_groupi_n_8977);
  or csa_tree_add_190_195_groupi_g39505(csa_tree_add_190_195_groupi_n_9465 ,csa_tree_add_190_195_groupi_n_8507 ,csa_tree_add_190_195_groupi_n_8931);
  nor csa_tree_add_190_195_groupi_g39506(csa_tree_add_190_195_groupi_n_9464 ,csa_tree_add_190_195_groupi_n_8369 ,csa_tree_add_190_195_groupi_n_8968);
  or csa_tree_add_190_195_groupi_g39507(csa_tree_add_190_195_groupi_n_9463 ,csa_tree_add_190_195_groupi_n_8334 ,csa_tree_add_190_195_groupi_n_8976);
  or csa_tree_add_190_195_groupi_g39508(csa_tree_add_190_195_groupi_n_9462 ,csa_tree_add_190_195_groupi_n_8368 ,csa_tree_add_190_195_groupi_n_8967);
  or csa_tree_add_190_195_groupi_g39509(csa_tree_add_190_195_groupi_n_9461 ,csa_tree_add_190_195_groupi_n_8365 ,csa_tree_add_190_195_groupi_n_9158);
  or csa_tree_add_190_195_groupi_g39510(csa_tree_add_190_195_groupi_n_9460 ,csa_tree_add_190_195_groupi_n_8542 ,csa_tree_add_190_195_groupi_n_9152);
  nor csa_tree_add_190_195_groupi_g39511(csa_tree_add_190_195_groupi_n_9459 ,csa_tree_add_190_195_groupi_n_8366 ,csa_tree_add_190_195_groupi_n_9157);
  or csa_tree_add_190_195_groupi_g39512(csa_tree_add_190_195_groupi_n_9458 ,csa_tree_add_190_195_groupi_n_7353 ,csa_tree_add_190_195_groupi_n_8975);
  or csa_tree_add_190_195_groupi_g39513(csa_tree_add_190_195_groupi_n_9457 ,csa_tree_add_190_195_groupi_n_8011 ,csa_tree_add_190_195_groupi_n_8970);
  nor csa_tree_add_190_195_groupi_g39514(csa_tree_add_190_195_groupi_n_9456 ,csa_tree_add_190_195_groupi_n_8010 ,csa_tree_add_190_195_groupi_n_8971);
  and csa_tree_add_190_195_groupi_g39515(csa_tree_add_190_195_groupi_n_9455 ,csa_tree_add_190_195_groupi_n_8215 ,csa_tree_add_190_195_groupi_n_8942);
  or csa_tree_add_190_195_groupi_g39516(csa_tree_add_190_195_groupi_n_9454 ,csa_tree_add_190_195_groupi_n_9161 ,csa_tree_add_190_195_groupi_n_8959);
  nor csa_tree_add_190_195_groupi_g39517(csa_tree_add_190_195_groupi_n_9453 ,csa_tree_add_190_195_groupi_n_8485 ,csa_tree_add_190_195_groupi_n_8965);
  nor csa_tree_add_190_195_groupi_g39518(csa_tree_add_190_195_groupi_n_9452 ,csa_tree_add_190_195_groupi_n_9162 ,csa_tree_add_190_195_groupi_n_8958);
  and csa_tree_add_190_195_groupi_g39519(csa_tree_add_190_195_groupi_n_9451 ,csa_tree_add_190_195_groupi_n_9147 ,csa_tree_add_190_195_groupi_n_8875);
  and csa_tree_add_190_195_groupi_g39520(csa_tree_add_190_195_groupi_n_9450 ,csa_tree_add_190_195_groupi_n_7353 ,csa_tree_add_190_195_groupi_n_8975);
  or csa_tree_add_190_195_groupi_g39521(csa_tree_add_190_195_groupi_n_9449 ,csa_tree_add_190_195_groupi_n_8801 ,csa_tree_add_190_195_groupi_n_9189);
  or csa_tree_add_190_195_groupi_g39522(csa_tree_add_190_195_groupi_n_9448 ,csa_tree_add_190_195_groupi_n_8511 ,csa_tree_add_190_195_groupi_n_8933);
  or csa_tree_add_190_195_groupi_g39523(csa_tree_add_190_195_groupi_n_9447 ,csa_tree_add_190_195_groupi_n_8525 ,csa_tree_add_190_195_groupi_n_9140);
  and csa_tree_add_190_195_groupi_g39524(csa_tree_add_190_195_groupi_n_9446 ,csa_tree_add_190_195_groupi_n_8219 ,csa_tree_add_190_195_groupi_n_9139);
  or csa_tree_add_190_195_groupi_g39525(csa_tree_add_190_195_groupi_n_9445 ,csa_tree_add_190_195_groupi_n_7775 ,csa_tree_add_190_195_groupi_n_9202);
  or csa_tree_add_190_195_groupi_g39526(csa_tree_add_190_195_groupi_n_9444 ,csa_tree_add_190_195_groupi_n_8596 ,csa_tree_add_190_195_groupi_n_9039);
  and csa_tree_add_190_195_groupi_g39527(csa_tree_add_190_195_groupi_n_9443 ,csa_tree_add_190_195_groupi_n_8485 ,csa_tree_add_190_195_groupi_n_8965);
  or csa_tree_add_190_195_groupi_g39528(csa_tree_add_190_195_groupi_n_9442 ,csa_tree_add_190_195_groupi_n_7489 ,csa_tree_add_190_195_groupi_n_9041);
  nor csa_tree_add_190_195_groupi_g39529(csa_tree_add_190_195_groupi_n_9441 ,csa_tree_add_190_195_groupi_n_8867 ,csa_tree_add_190_195_groupi_n_9117);
  or csa_tree_add_190_195_groupi_g39530(csa_tree_add_190_195_groupi_n_9440 ,csa_tree_add_190_195_groupi_n_8855 ,csa_tree_add_190_195_groupi_n_9131);
  or csa_tree_add_190_195_groupi_g39531(csa_tree_add_190_195_groupi_n_9439 ,csa_tree_add_190_195_groupi_n_8850 ,csa_tree_add_190_195_groupi_n_9129);
  and csa_tree_add_190_195_groupi_g39532(csa_tree_add_190_195_groupi_n_9438 ,csa_tree_add_190_195_groupi_n_8141 ,csa_tree_add_190_195_groupi_n_9042);
  and csa_tree_add_190_195_groupi_g39533(csa_tree_add_190_195_groupi_n_9437 ,csa_tree_add_190_195_groupi_n_8446 ,csa_tree_add_190_195_groupi_n_9200);
  nor csa_tree_add_190_195_groupi_g39534(csa_tree_add_190_195_groupi_n_9436 ,csa_tree_add_190_195_groupi_n_8841 ,csa_tree_add_190_195_groupi_n_9124);
  or csa_tree_add_190_195_groupi_g39535(csa_tree_add_190_195_groupi_n_9435 ,csa_tree_add_190_195_groupi_n_8385 ,csa_tree_add_190_195_groupi_n_9125);
  or csa_tree_add_190_195_groupi_g39536(csa_tree_add_190_195_groupi_n_9434 ,csa_tree_add_190_195_groupi_n_9163 ,csa_tree_add_190_195_groupi_n_8954);
  nor csa_tree_add_190_195_groupi_g39537(csa_tree_add_190_195_groupi_n_9433 ,csa_tree_add_190_195_groupi_n_7767 ,csa_tree_add_190_195_groupi_n_9038);
  nor csa_tree_add_190_195_groupi_g39538(csa_tree_add_190_195_groupi_n_9432 ,csa_tree_add_190_195_groupi_n_7588 ,csa_tree_add_190_195_groupi_n_8973);
  or csa_tree_add_190_195_groupi_g39539(csa_tree_add_190_195_groupi_n_9431 ,csa_tree_add_190_195_groupi_n_7589 ,csa_tree_add_190_195_groupi_n_8972);
  or csa_tree_add_190_195_groupi_g39540(csa_tree_add_190_195_groupi_n_9430 ,csa_tree_add_190_195_groupi_n_8835 ,csa_tree_add_190_195_groupi_n_8969);
  or csa_tree_add_190_195_groupi_g39541(csa_tree_add_190_195_groupi_n_9429 ,csa_tree_add_190_195_groupi_n_5333 ,csa_tree_add_190_195_groupi_n_9004);
  and csa_tree_add_190_195_groupi_g39542(csa_tree_add_190_195_groupi_n_9428 ,csa_tree_add_190_195_groupi_n_8835 ,csa_tree_add_190_195_groupi_n_8969);
  and csa_tree_add_190_195_groupi_g39543(csa_tree_add_190_195_groupi_n_9427 ,csa_tree_add_190_195_groupi_n_7274 ,csa_tree_add_190_195_groupi_n_9045);
  nor csa_tree_add_190_195_groupi_g39544(csa_tree_add_190_195_groupi_n_9426 ,csa_tree_add_190_195_groupi_n_7172 ,csa_tree_add_190_195_groupi_n_9167);
  and csa_tree_add_190_195_groupi_g39545(csa_tree_add_190_195_groupi_n_9425 ,csa_tree_add_190_195_groupi_n_8521 ,csa_tree_add_190_195_groupi_n_9054);
  and csa_tree_add_190_195_groupi_g39546(csa_tree_add_190_195_groupi_n_9424 ,csa_tree_add_190_195_groupi_n_8524 ,csa_tree_add_190_195_groupi_n_9120);
  or csa_tree_add_190_195_groupi_g39547(csa_tree_add_190_195_groupi_n_9423 ,csa_tree_add_190_195_groupi_n_7171 ,csa_tree_add_190_195_groupi_n_9168);
  or csa_tree_add_190_195_groupi_g39548(csa_tree_add_190_195_groupi_n_9422 ,csa_tree_add_190_195_groupi_n_8335 ,csa_tree_add_190_195_groupi_n_8984);
  nor csa_tree_add_190_195_groupi_g39549(csa_tree_add_190_195_groupi_n_9421 ,csa_tree_add_190_195_groupi_n_8336 ,csa_tree_add_190_195_groupi_n_8985);
  nor csa_tree_add_190_195_groupi_g39550(csa_tree_add_190_195_groupi_n_9420 ,csa_tree_add_190_195_groupi_n_5332 ,csa_tree_add_190_195_groupi_n_9005);
  nor csa_tree_add_190_195_groupi_g39551(csa_tree_add_190_195_groupi_n_9419 ,csa_tree_add_190_195_groupi_n_9164 ,csa_tree_add_190_195_groupi_n_8955);
  nor csa_tree_add_190_195_groupi_g39552(csa_tree_add_190_195_groupi_n_9418 ,csa_tree_add_190_195_groupi_n_7985 ,csa_tree_add_190_195_groupi_n_8960);
  or csa_tree_add_190_195_groupi_g39553(csa_tree_add_190_195_groupi_n_9417 ,csa_tree_add_190_195_groupi_n_8821 ,csa_tree_add_190_195_groupi_n_9172);
  and csa_tree_add_190_195_groupi_g39554(csa_tree_add_190_195_groupi_n_9416 ,csa_tree_add_190_195_groupi_n_7985 ,csa_tree_add_190_195_groupi_n_8960);
  and csa_tree_add_190_195_groupi_g39555(csa_tree_add_190_195_groupi_n_9415 ,csa_tree_add_190_195_groupi_n_8425 ,csa_tree_add_190_195_groupi_n_9048);
  nor csa_tree_add_190_195_groupi_g39556(csa_tree_add_190_195_groupi_n_9414 ,csa_tree_add_190_195_groupi_n_9003 ,csa_tree_add_190_195_groupi_n_8644);
  or csa_tree_add_190_195_groupi_g39557(csa_tree_add_190_195_groupi_n_9413 ,csa_tree_add_190_195_groupi_n_9002 ,csa_tree_add_190_195_groupi_n_8643);
  or csa_tree_add_190_195_groupi_g39558(csa_tree_add_190_195_groupi_n_9412 ,csa_tree_add_190_195_groupi_n_8707 ,csa_tree_add_190_195_groupi_n_9112);
  nor csa_tree_add_190_195_groupi_g39559(csa_tree_add_190_195_groupi_n_9411 ,csa_tree_add_190_195_groupi_n_9199 ,csa_tree_add_190_195_groupi_n_7771);
  or csa_tree_add_190_195_groupi_g39560(csa_tree_add_190_195_groupi_n_9410 ,csa_tree_add_190_195_groupi_n_9150 ,csa_tree_add_190_195_groupi_n_9046);
  or csa_tree_add_190_195_groupi_g39561(csa_tree_add_190_195_groupi_n_9409 ,csa_tree_add_190_195_groupi_n_7128 ,csa_tree_add_190_195_groupi_n_9020);
  or csa_tree_add_190_195_groupi_g39562(csa_tree_add_190_195_groupi_n_9408 ,csa_tree_add_190_195_groupi_n_7956 ,csa_tree_add_190_195_groupi_n_9044);
  or csa_tree_add_190_195_groupi_g39563(csa_tree_add_190_195_groupi_n_9407 ,csa_tree_add_190_195_groupi_n_9187 ,csa_tree_add_190_195_groupi_n_8928);
  or csa_tree_add_190_195_groupi_g39564(csa_tree_add_190_195_groupi_n_9406 ,csa_tree_add_190_195_groupi_n_8536 ,csa_tree_add_190_195_groupi_n_9105);
  or csa_tree_add_190_195_groupi_g39565(csa_tree_add_190_195_groupi_n_9405 ,csa_tree_add_190_195_groupi_n_6250 ,csa_tree_add_190_195_groupi_n_9047);
  and csa_tree_add_190_195_groupi_g39566(csa_tree_add_190_195_groupi_n_9404 ,csa_tree_add_190_195_groupi_n_9192 ,csa_tree_add_190_195_groupi_n_9088);
  nor csa_tree_add_190_195_groupi_g39567(csa_tree_add_190_195_groupi_n_9403 ,csa_tree_add_190_195_groupi_n_7129 ,csa_tree_add_190_195_groupi_n_9021);
  or csa_tree_add_190_195_groupi_g39568(csa_tree_add_190_195_groupi_n_9402 ,csa_tree_add_190_195_groupi_n_9018 ,csa_tree_add_190_195_groupi_n_8951);
  nor csa_tree_add_190_195_groupi_g39569(csa_tree_add_190_195_groupi_n_9401 ,csa_tree_add_190_195_groupi_n_9019 ,csa_tree_add_190_195_groupi_n_8950);
  nor csa_tree_add_190_195_groupi_g39570(csa_tree_add_190_195_groupi_n_9400 ,csa_tree_add_190_195_groupi_n_6959 ,csa_tree_add_190_195_groupi_n_8949);
  or csa_tree_add_190_195_groupi_g39571(csa_tree_add_190_195_groupi_n_9399 ,csa_tree_add_190_195_groupi_n_6960 ,csa_tree_add_190_195_groupi_n_8948);
  and csa_tree_add_190_195_groupi_g39572(csa_tree_add_190_195_groupi_n_9398 ,csa_tree_add_190_195_groupi_n_9182 ,csa_tree_add_190_195_groupi_n_8913);
  or csa_tree_add_190_195_groupi_g39573(csa_tree_add_190_195_groupi_n_9397 ,csa_tree_add_190_195_groupi_n_8509 ,csa_tree_add_190_195_groupi_n_9098);
  nor csa_tree_add_190_195_groupi_g39574(csa_tree_add_190_195_groupi_n_9396 ,csa_tree_add_190_195_groupi_n_8822 ,csa_tree_add_190_195_groupi_n_9173);
  or csa_tree_add_190_195_groupi_g39575(csa_tree_add_190_195_groupi_n_9395 ,csa_tree_add_190_195_groupi_n_8133 ,csa_tree_add_190_195_groupi_n_9051);
  or csa_tree_add_190_195_groupi_g39576(csa_tree_add_190_195_groupi_n_9394 ,csa_tree_add_190_195_groupi_n_8847 ,csa_tree_add_190_195_groupi_n_8944);
  or csa_tree_add_190_195_groupi_g39577(csa_tree_add_190_195_groupi_n_9393 ,csa_tree_add_190_195_groupi_n_7623 ,csa_tree_add_190_195_groupi_n_9000);
  nor csa_tree_add_190_195_groupi_g39578(csa_tree_add_190_195_groupi_n_9392 ,csa_tree_add_190_195_groupi_n_8858 ,csa_tree_add_190_195_groupi_n_9092);
  or csa_tree_add_190_195_groupi_g39579(csa_tree_add_190_195_groupi_n_9391 ,csa_tree_add_190_195_groupi_n_9178 ,csa_tree_add_190_195_groupi_n_9174);
  and csa_tree_add_190_195_groupi_g39580(csa_tree_add_190_195_groupi_n_9390 ,csa_tree_add_190_195_groupi_n_9058 ,csa_tree_add_190_195_groupi_n_9191);
  or csa_tree_add_190_195_groupi_g39581(csa_tree_add_190_195_groupi_n_9389 ,csa_tree_add_190_195_groupi_n_8870 ,csa_tree_add_190_195_groupi_n_9089);
  nor csa_tree_add_190_195_groupi_g39582(csa_tree_add_190_195_groupi_n_9388 ,csa_tree_add_190_195_groupi_n_7983 ,csa_tree_add_190_195_groupi_n_8961);
  or csa_tree_add_190_195_groupi_g39583(csa_tree_add_190_195_groupi_n_9387 ,csa_tree_add_190_195_groupi_n_7982 ,csa_tree_add_190_195_groupi_n_8962);
  nor csa_tree_add_190_195_groupi_g39584(csa_tree_add_190_195_groupi_n_9386 ,csa_tree_add_190_195_groupi_n_9179 ,csa_tree_add_190_195_groupi_n_9175);
  and csa_tree_add_190_195_groupi_g39585(csa_tree_add_190_195_groupi_n_9385 ,csa_tree_add_190_195_groupi_n_9193 ,csa_tree_add_190_195_groupi_n_8477);
  and csa_tree_add_190_195_groupi_g39586(csa_tree_add_190_195_groupi_n_9384 ,csa_tree_add_190_195_groupi_n_8533 ,csa_tree_add_190_195_groupi_n_9083);
  or csa_tree_add_190_195_groupi_g39587(csa_tree_add_190_195_groupi_n_9383 ,csa_tree_add_190_195_groupi_n_9082 ,csa_tree_add_190_195_groupi_n_9050);
  or csa_tree_add_190_195_groupi_g39588(csa_tree_add_190_195_groupi_n_9382 ,csa_tree_add_190_195_groupi_n_7326 ,csa_tree_add_190_195_groupi_n_9180);
  nor csa_tree_add_190_195_groupi_g39589(csa_tree_add_190_195_groupi_n_9381 ,csa_tree_add_190_195_groupi_n_7327 ,csa_tree_add_190_195_groupi_n_9181);
  and csa_tree_add_190_195_groupi_g39590(csa_tree_add_190_195_groupi_n_9380 ,csa_tree_add_190_195_groupi_n_7239 ,csa_tree_add_190_195_groupi_n_9185);
  nor csa_tree_add_190_195_groupi_g39591(csa_tree_add_190_195_groupi_n_9379 ,csa_tree_add_190_195_groupi_n_7515 ,csa_tree_add_190_195_groupi_n_9016);
  nor csa_tree_add_190_195_groupi_g39592(csa_tree_add_190_195_groupi_n_9378 ,csa_tree_add_190_195_groupi_n_6096 ,csa_tree_add_190_195_groupi_n_9036);
  nor csa_tree_add_190_195_groupi_g39593(csa_tree_add_190_195_groupi_n_9377 ,csa_tree_add_190_195_groupi_n_8332 ,csa_tree_add_190_195_groupi_n_8946);
  or csa_tree_add_190_195_groupi_g39594(csa_tree_add_190_195_groupi_n_9376 ,csa_tree_add_190_195_groupi_n_8520 ,csa_tree_add_190_195_groupi_n_9061);
  or csa_tree_add_190_195_groupi_g39595(csa_tree_add_190_195_groupi_n_9375 ,csa_tree_add_190_195_groupi_n_7514 ,csa_tree_add_190_195_groupi_n_9017);
  or csa_tree_add_190_195_groupi_g39596(csa_tree_add_190_195_groupi_n_9374 ,csa_tree_add_190_195_groupi_n_8522 ,csa_tree_add_190_195_groupi_n_9133);
  and csa_tree_add_190_195_groupi_g39597(csa_tree_add_190_195_groupi_n_9373 ,csa_tree_add_190_195_groupi_n_8930 ,csa_tree_add_190_195_groupi_n_9052);
  or csa_tree_add_190_195_groupi_g39598(csa_tree_add_190_195_groupi_n_9372 ,csa_tree_add_190_195_groupi_n_8331 ,csa_tree_add_190_195_groupi_n_8947);
  and csa_tree_add_190_195_groupi_g39599(csa_tree_add_190_195_groupi_n_9371 ,csa_tree_add_190_195_groupi_n_8210 ,csa_tree_add_190_195_groupi_n_9080);
  nor csa_tree_add_190_195_groupi_g39600(csa_tree_add_190_195_groupi_n_9370 ,csa_tree_add_190_195_groupi_n_7624 ,csa_tree_add_190_195_groupi_n_9001);
  or csa_tree_add_190_195_groupi_g39601(csa_tree_add_190_195_groupi_n_9527 ,csa_tree_add_190_195_groupi_n_8810 ,csa_tree_add_190_195_groupi_n_9097);
  and csa_tree_add_190_195_groupi_g39602(csa_tree_add_190_195_groupi_n_9526 ,csa_tree_add_190_195_groupi_n_8753 ,csa_tree_add_190_195_groupi_n_9065);
  or csa_tree_add_190_195_groupi_g39603(csa_tree_add_190_195_groupi_n_9524 ,csa_tree_add_190_195_groupi_n_8736 ,csa_tree_add_190_195_groupi_n_9078);
  or csa_tree_add_190_195_groupi_g39604(csa_tree_add_190_195_groupi_n_9523 ,csa_tree_add_190_195_groupi_n_6523 ,csa_tree_add_190_195_groupi_n_9143);
  and csa_tree_add_190_195_groupi_g39605(csa_tree_add_190_195_groupi_n_9522 ,csa_tree_add_190_195_groupi_n_8457 ,csa_tree_add_190_195_groupi_n_9062);
  and csa_tree_add_190_195_groupi_g39606(csa_tree_add_190_195_groupi_n_9521 ,csa_tree_add_190_195_groupi_n_8778 ,csa_tree_add_190_195_groupi_n_9073);
  or csa_tree_add_190_195_groupi_g39607(csa_tree_add_190_195_groupi_n_9520 ,csa_tree_add_190_195_groupi_n_8601 ,csa_tree_add_190_195_groupi_n_9075);
  and csa_tree_add_190_195_groupi_g39608(csa_tree_add_190_195_groupi_n_9519 ,csa_tree_add_190_195_groupi_n_8727 ,csa_tree_add_190_195_groupi_n_9081);
  or csa_tree_add_190_195_groupi_g39609(csa_tree_add_190_195_groupi_n_9518 ,csa_tree_add_190_195_groupi_n_8792 ,csa_tree_add_190_195_groupi_n_9135);
  or csa_tree_add_190_195_groupi_g39610(csa_tree_add_190_195_groupi_n_9516 ,csa_tree_add_190_195_groupi_n_7750 ,csa_tree_add_190_195_groupi_n_9116);
  or csa_tree_add_190_195_groupi_g39611(csa_tree_add_190_195_groupi_n_9515 ,csa_tree_add_190_195_groupi_n_8112 ,csa_tree_add_190_195_groupi_n_9115);
  and csa_tree_add_190_195_groupi_g39612(csa_tree_add_190_195_groupi_n_9514 ,csa_tree_add_190_195_groupi_n_6190 ,csa_tree_add_190_195_groupi_n_9110);
  or csa_tree_add_190_195_groupi_g39613(csa_tree_add_190_195_groupi_n_9513 ,csa_tree_add_190_195_groupi_n_8794 ,csa_tree_add_190_195_groupi_n_9057);
  and csa_tree_add_190_195_groupi_g39614(csa_tree_add_190_195_groupi_n_9512 ,csa_tree_add_190_195_groupi_n_8775 ,csa_tree_add_190_195_groupi_n_9056);
  and csa_tree_add_190_195_groupi_g39615(csa_tree_add_190_195_groupi_n_9511 ,csa_tree_add_190_195_groupi_n_8790 ,csa_tree_add_190_195_groupi_n_9053);
  or csa_tree_add_190_195_groupi_g39616(csa_tree_add_190_195_groupi_n_9509 ,csa_tree_add_190_195_groupi_n_7705 ,csa_tree_add_190_195_groupi_n_9091);
  and csa_tree_add_190_195_groupi_g39617(csa_tree_add_190_195_groupi_n_9508 ,csa_tree_add_190_195_groupi_n_8732 ,csa_tree_add_190_195_groupi_n_9093);
  and csa_tree_add_190_195_groupi_g39618(csa_tree_add_190_195_groupi_n_9507 ,csa_tree_add_190_195_groupi_n_6452 ,csa_tree_add_190_195_groupi_n_8940);
  and csa_tree_add_190_195_groupi_g39619(csa_tree_add_190_195_groupi_n_9506 ,csa_tree_add_190_195_groupi_n_8804 ,csa_tree_add_190_195_groupi_n_8943);
  and csa_tree_add_190_195_groupi_g39620(csa_tree_add_190_195_groupi_n_9505 ,csa_tree_add_190_195_groupi_n_8786 ,csa_tree_add_190_195_groupi_n_9119);
  and csa_tree_add_190_195_groupi_g39621(csa_tree_add_190_195_groupi_n_9504 ,csa_tree_add_190_195_groupi_n_8745 ,csa_tree_add_190_195_groupi_n_9102);
  and csa_tree_add_190_195_groupi_g39622(csa_tree_add_190_195_groupi_n_9502 ,csa_tree_add_190_195_groupi_n_7976 ,csa_tree_add_190_195_groupi_n_9069);
  and csa_tree_add_190_195_groupi_g39623(csa_tree_add_190_195_groupi_n_9501 ,csa_tree_add_190_195_groupi_n_8750 ,csa_tree_add_190_195_groupi_n_9108);
  and csa_tree_add_190_195_groupi_g39624(csa_tree_add_190_195_groupi_n_9500 ,csa_tree_add_190_195_groupi_n_8592 ,csa_tree_add_190_195_groupi_n_9155);
  or csa_tree_add_190_195_groupi_g39625(csa_tree_add_190_195_groupi_n_9497 ,csa_tree_add_190_195_groupi_n_8811 ,csa_tree_add_190_195_groupi_n_9100);
  and csa_tree_add_190_195_groupi_g39626(csa_tree_add_190_195_groupi_n_9496 ,csa_tree_add_190_195_groupi_n_8738 ,csa_tree_add_190_195_groupi_n_9118);
  or csa_tree_add_190_195_groupi_g39627(csa_tree_add_190_195_groupi_n_9493 ,csa_tree_add_190_195_groupi_n_8737 ,csa_tree_add_190_195_groupi_n_9094);
  or csa_tree_add_190_195_groupi_g39628(csa_tree_add_190_195_groupi_n_9491 ,csa_tree_add_190_195_groupi_n_7738 ,csa_tree_add_190_195_groupi_n_9111);
  or csa_tree_add_190_195_groupi_g39629(csa_tree_add_190_195_groupi_n_9490 ,csa_tree_add_190_195_groupi_n_7264 ,csa_tree_add_190_195_groupi_n_9109);
  and csa_tree_add_190_195_groupi_g39630(csa_tree_add_190_195_groupi_n_9488 ,csa_tree_add_190_195_groupi_n_6847 ,csa_tree_add_190_195_groupi_n_9114);
  or csa_tree_add_190_195_groupi_g39631(csa_tree_add_190_195_groupi_n_9486 ,csa_tree_add_190_195_groupi_n_8607 ,csa_tree_add_190_195_groupi_n_8938);
  or csa_tree_add_190_195_groupi_g39632(csa_tree_add_190_195_groupi_n_9484 ,csa_tree_add_190_195_groupi_n_7947 ,csa_tree_add_190_195_groupi_n_9087);
  and csa_tree_add_190_195_groupi_g39633(csa_tree_add_190_195_groupi_n_9482 ,csa_tree_add_190_195_groupi_n_7704 ,csa_tree_add_190_195_groupi_n_9085);
  or csa_tree_add_190_195_groupi_g39634(csa_tree_add_190_195_groupi_n_9480 ,csa_tree_add_190_195_groupi_n_8599 ,csa_tree_add_190_195_groupi_n_8935);
  or csa_tree_add_190_195_groupi_g39635(csa_tree_add_190_195_groupi_n_9478 ,csa_tree_add_190_195_groupi_n_6408 ,csa_tree_add_190_195_groupi_n_9123);
  or csa_tree_add_190_195_groupi_g39636(csa_tree_add_190_195_groupi_n_9477 ,csa_tree_add_190_195_groupi_n_8725 ,csa_tree_add_190_195_groupi_n_9070);
  and csa_tree_add_190_195_groupi_g39637(csa_tree_add_190_195_groupi_n_9476 ,csa_tree_add_190_195_groupi_n_8770 ,csa_tree_add_190_195_groupi_n_9079);
  or csa_tree_add_190_195_groupi_g39638(csa_tree_add_190_195_groupi_n_9474 ,csa_tree_add_190_195_groupi_n_8145 ,csa_tree_add_190_195_groupi_n_9077);
  and csa_tree_add_190_195_groupi_g39639(csa_tree_add_190_195_groupi_n_9473 ,csa_tree_add_190_195_groupi_n_7968 ,csa_tree_add_190_195_groupi_n_9156);
  and csa_tree_add_190_195_groupi_g39640(csa_tree_add_190_195_groupi_n_9470 ,csa_tree_add_190_195_groupi_n_8454 ,csa_tree_add_190_195_groupi_n_9064);
  or csa_tree_add_190_195_groupi_g39641(csa_tree_add_190_195_groupi_n_9468 ,csa_tree_add_190_195_groupi_n_8749 ,csa_tree_add_190_195_groupi_n_9066);
  and csa_tree_add_190_195_groupi_g39642(csa_tree_add_190_195_groupi_n_9467 ,csa_tree_add_190_195_groupi_n_8746 ,csa_tree_add_190_195_groupi_n_9101);
  not csa_tree_add_190_195_groupi_g39643(csa_tree_add_190_195_groupi_n_9369 ,csa_tree_add_190_195_groupi_n_9368);
  not csa_tree_add_190_195_groupi_g39644(csa_tree_add_190_195_groupi_n_9366 ,csa_tree_add_190_195_groupi_n_9365);
  not csa_tree_add_190_195_groupi_g39645(csa_tree_add_190_195_groupi_n_9364 ,csa_tree_add_190_195_groupi_n_9363);
  not csa_tree_add_190_195_groupi_g39648(csa_tree_add_190_195_groupi_n_9351 ,csa_tree_add_190_195_groupi_n_9350);
  not csa_tree_add_190_195_groupi_g39649(csa_tree_add_190_195_groupi_n_9347 ,csa_tree_add_190_195_groupi_n_120);
  not csa_tree_add_190_195_groupi_g39650(csa_tree_add_190_195_groupi_n_9346 ,csa_tree_add_190_195_groupi_n_9345);
  not csa_tree_add_190_195_groupi_g39651(csa_tree_add_190_195_groupi_n_9344 ,csa_tree_add_190_195_groupi_n_9343);
  not csa_tree_add_190_195_groupi_g39652(csa_tree_add_190_195_groupi_n_9342 ,csa_tree_add_190_195_groupi_n_9341);
  not csa_tree_add_190_195_groupi_g39653(csa_tree_add_190_195_groupi_n_9340 ,csa_tree_add_190_195_groupi_n_9339);
  not csa_tree_add_190_195_groupi_g39654(csa_tree_add_190_195_groupi_n_9338 ,csa_tree_add_190_195_groupi_n_9337);
  not csa_tree_add_190_195_groupi_g39655(csa_tree_add_190_195_groupi_n_9336 ,csa_tree_add_190_195_groupi_n_9335);
  not csa_tree_add_190_195_groupi_g39656(csa_tree_add_190_195_groupi_n_9334 ,csa_tree_add_190_195_groupi_n_9333);
  not csa_tree_add_190_195_groupi_g39657(csa_tree_add_190_195_groupi_n_9332 ,csa_tree_add_190_195_groupi_n_9331);
  not csa_tree_add_190_195_groupi_g39658(csa_tree_add_190_195_groupi_n_9329 ,csa_tree_add_190_195_groupi_n_9328);
  not csa_tree_add_190_195_groupi_g39659(csa_tree_add_190_195_groupi_n_9327 ,csa_tree_add_190_195_groupi_n_111);
  not csa_tree_add_190_195_groupi_g39660(csa_tree_add_190_195_groupi_n_9326 ,csa_tree_add_190_195_groupi_n_9325);
  not csa_tree_add_190_195_groupi_g39661(csa_tree_add_190_195_groupi_n_9324 ,csa_tree_add_190_195_groupi_n_9323);
  not csa_tree_add_190_195_groupi_g39662(csa_tree_add_190_195_groupi_n_9322 ,csa_tree_add_190_195_groupi_n_9321);
  not csa_tree_add_190_195_groupi_g39663(csa_tree_add_190_195_groupi_n_9320 ,csa_tree_add_190_195_groupi_n_9319);
  not csa_tree_add_190_195_groupi_g39664(csa_tree_add_190_195_groupi_n_9316 ,csa_tree_add_190_195_groupi_n_9315);
  not csa_tree_add_190_195_groupi_g39665(csa_tree_add_190_195_groupi_n_9313 ,csa_tree_add_190_195_groupi_n_9312);
  not csa_tree_add_190_195_groupi_g39666(csa_tree_add_190_195_groupi_n_9311 ,csa_tree_add_190_195_groupi_n_119);
  not csa_tree_add_190_195_groupi_g39667(csa_tree_add_190_195_groupi_n_9310 ,csa_tree_add_190_195_groupi_n_9309);
  not csa_tree_add_190_195_groupi_g39668(csa_tree_add_190_195_groupi_n_9306 ,csa_tree_add_190_195_groupi_n_9307);
  not csa_tree_add_190_195_groupi_g39669(csa_tree_add_190_195_groupi_n_9305 ,csa_tree_add_190_195_groupi_n_9304);
  not csa_tree_add_190_195_groupi_g39670(csa_tree_add_190_195_groupi_n_9303 ,csa_tree_add_190_195_groupi_n_9302);
  not csa_tree_add_190_195_groupi_g39671(csa_tree_add_190_195_groupi_n_9301 ,csa_tree_add_190_195_groupi_n_9300);
  not csa_tree_add_190_195_groupi_g39672(csa_tree_add_190_195_groupi_n_9298 ,csa_tree_add_190_195_groupi_n_9299);
  not csa_tree_add_190_195_groupi_g39673(csa_tree_add_190_195_groupi_n_9297 ,csa_tree_add_190_195_groupi_n_9296);
  not csa_tree_add_190_195_groupi_g39674(csa_tree_add_190_195_groupi_n_9294 ,csa_tree_add_190_195_groupi_n_9293);
  not csa_tree_add_190_195_groupi_g39675(csa_tree_add_190_195_groupi_n_9290 ,csa_tree_add_190_195_groupi_n_9289);
  not csa_tree_add_190_195_groupi_g39676(csa_tree_add_190_195_groupi_n_9288 ,csa_tree_add_190_195_groupi_n_9287);
  not csa_tree_add_190_195_groupi_g39677(csa_tree_add_190_195_groupi_n_9285 ,csa_tree_add_190_195_groupi_n_9284);
  or csa_tree_add_190_195_groupi_g39678(csa_tree_add_190_195_groupi_n_9283 ,csa_tree_add_190_195_groupi_n_8987 ,csa_tree_add_190_195_groupi_n_9026);
  or csa_tree_add_190_195_groupi_g39679(csa_tree_add_190_195_groupi_n_9282 ,csa_tree_add_190_195_groupi_n_8648 ,csa_tree_add_190_195_groupi_n_8989);
  nor csa_tree_add_190_195_groupi_g39680(csa_tree_add_190_195_groupi_n_9281 ,csa_tree_add_190_195_groupi_n_8986 ,csa_tree_add_190_195_groupi_n_9027);
  or csa_tree_add_190_195_groupi_g39681(csa_tree_add_190_195_groupi_n_9280 ,csa_tree_add_190_195_groupi_n_8824 ,csa_tree_add_190_195_groupi_n_9023);
  or csa_tree_add_190_195_groupi_g39682(csa_tree_add_190_195_groupi_n_9279 ,csa_tree_add_190_195_groupi_n_9169 ,csa_tree_add_190_195_groupi_n_8330);
  and csa_tree_add_190_195_groupi_g39683(csa_tree_add_190_195_groupi_n_9278 ,csa_tree_add_190_195_groupi_n_9169 ,csa_tree_add_190_195_groupi_n_8330);
  or csa_tree_add_190_195_groupi_g39684(csa_tree_add_190_195_groupi_n_9277 ,csa_tree_add_190_195_groupi_n_9034 ,csa_tree_add_190_195_groupi_n_9031);
  nor csa_tree_add_190_195_groupi_g39685(csa_tree_add_190_195_groupi_n_9276 ,csa_tree_add_190_195_groupi_n_9033 ,csa_tree_add_190_195_groupi_n_9032);
  nor csa_tree_add_190_195_groupi_g39686(csa_tree_add_190_195_groupi_n_9275 ,csa_tree_add_190_195_groupi_n_6954 ,csa_tree_add_190_195_groupi_n_9171);
  and csa_tree_add_190_195_groupi_g39687(csa_tree_add_190_195_groupi_n_9274 ,csa_tree_add_190_195_groupi_n_7123 ,csa_tree_add_190_195_groupi_n_8974);
  or csa_tree_add_190_195_groupi_g39688(csa_tree_add_190_195_groupi_n_9273 ,csa_tree_add_190_195_groupi_n_8857 ,csa_tree_add_190_195_groupi_n_8922);
  nor csa_tree_add_190_195_groupi_g39689(csa_tree_add_190_195_groupi_n_9272 ,csa_tree_add_190_195_groupi_n_8825 ,csa_tree_add_190_195_groupi_n_9022);
  or csa_tree_add_190_195_groupi_g39690(csa_tree_add_190_195_groupi_n_9271 ,csa_tree_add_190_195_groupi_n_6955 ,csa_tree_add_190_195_groupi_n_9170);
  nor csa_tree_add_190_195_groupi_g39691(csa_tree_add_190_195_groupi_n_9270 ,csa_tree_add_190_195_groupi_n_7123 ,csa_tree_add_190_195_groupi_n_8974);
  nor csa_tree_add_190_195_groupi_g39692(csa_tree_add_190_195_groupi_n_9269 ,csa_tree_add_190_195_groupi_n_8813 ,csa_tree_add_190_195_groupi_n_8995);
  and csa_tree_add_190_195_groupi_g39693(csa_tree_add_190_195_groupi_n_9268 ,csa_tree_add_190_195_groupi_n_9013 ,csa_tree_add_190_195_groupi_n_9012);
  nor csa_tree_add_190_195_groupi_g39694(csa_tree_add_190_195_groupi_n_9267 ,csa_tree_add_190_195_groupi_n_9013 ,csa_tree_add_190_195_groupi_n_9012);
  or csa_tree_add_190_195_groupi_g39695(csa_tree_add_190_195_groupi_n_9266 ,csa_tree_add_190_195_groupi_n_8868 ,csa_tree_add_190_195_groupi_n_8915);
  or csa_tree_add_190_195_groupi_g39696(csa_tree_add_190_195_groupi_n_9265 ,csa_tree_add_190_195_groupi_n_8026 ,csa_tree_add_190_195_groupi_n_9007);
  or csa_tree_add_190_195_groupi_g39697(csa_tree_add_190_195_groupi_n_9264 ,csa_tree_add_190_195_groupi_n_7952 ,csa_tree_add_190_195_groupi_n_9190);
  nor csa_tree_add_190_195_groupi_g39698(csa_tree_add_190_195_groupi_n_9263 ,csa_tree_add_190_195_groupi_n_8027 ,csa_tree_add_190_195_groupi_n_9006);
  nor csa_tree_add_190_195_groupi_g39699(csa_tree_add_190_195_groupi_n_9262 ,csa_tree_add_190_195_groupi_n_8667 ,csa_tree_add_190_195_groupi_n_8981);
  or csa_tree_add_190_195_groupi_g39700(csa_tree_add_190_195_groupi_n_9261 ,csa_tree_add_190_195_groupi_n_8812 ,csa_tree_add_190_195_groupi_n_105);
  or csa_tree_add_190_195_groupi_g39701(csa_tree_add_190_195_groupi_n_9260 ,csa_tree_add_190_195_groupi_n_7614 ,csa_tree_add_190_195_groupi_n_8996);
  nor csa_tree_add_190_195_groupi_g39702(csa_tree_add_190_195_groupi_n_9259 ,csa_tree_add_190_195_groupi_n_7613 ,csa_tree_add_190_195_groupi_n_8997);
  nor csa_tree_add_190_195_groupi_g39703(csa_tree_add_190_195_groupi_n_9258 ,csa_tree_add_190_195_groupi_n_8649 ,csa_tree_add_190_195_groupi_n_8990);
  or csa_tree_add_190_195_groupi_g39704(csa_tree_add_190_195_groupi_n_9257 ,csa_tree_add_190_195_groupi_n_8814 ,csa_tree_add_190_195_groupi_n_103);
  nor csa_tree_add_190_195_groupi_g39705(csa_tree_add_190_195_groupi_n_9256 ,csa_tree_add_190_195_groupi_n_8815 ,csa_tree_add_190_195_groupi_n_8988);
  or csa_tree_add_190_195_groupi_g39706(csa_tree_add_190_195_groupi_n_9255 ,csa_tree_add_190_195_groupi_n_8829 ,csa_tree_add_190_195_groupi_n_8982);
  nor csa_tree_add_190_195_groupi_g39707(csa_tree_add_190_195_groupi_n_9254 ,csa_tree_add_190_195_groupi_n_8830 ,csa_tree_add_190_195_groupi_n_8983);
  or csa_tree_add_190_195_groupi_g39708(csa_tree_add_190_195_groupi_n_9253 ,csa_tree_add_190_195_groupi_n_8668 ,csa_tree_add_190_195_groupi_n_8980);
  xnor csa_tree_add_190_195_groupi_g39709(csa_tree_add_190_195_groupi_n_9252 ,csa_tree_add_190_195_groupi_n_7637 ,csa_tree_add_190_195_groupi_n_8707);
  xnor csa_tree_add_190_195_groupi_g39710(csa_tree_add_190_195_groupi_n_9251 ,csa_tree_add_190_195_groupi_n_8705 ,csa_tree_add_190_195_groupi_n_6275);
  xnor csa_tree_add_190_195_groupi_g39711(csa_tree_add_190_195_groupi_n_9250 ,csa_tree_add_190_195_groupi_n_8338 ,csa_tree_add_190_195_groupi_n_8706);
  xnor csa_tree_add_190_195_groupi_g39712(csa_tree_add_190_195_groupi_n_9249 ,csa_tree_add_190_195_groupi_n_7327 ,csa_tree_add_190_195_groupi_n_8874);
  xnor csa_tree_add_190_195_groupi_g39713(csa_tree_add_190_195_groupi_n_9248 ,csa_tree_add_190_195_groupi_n_7131 ,csa_tree_add_190_195_groupi_n_8832);
  xnor csa_tree_add_190_195_groupi_g39714(csa_tree_add_190_195_groupi_n_9247 ,csa_tree_add_190_195_groupi_n_8616 ,csa_tree_add_190_195_groupi_n_8509);
  xnor csa_tree_add_190_195_groupi_g39715(csa_tree_add_190_195_groupi_n_9246 ,csa_tree_add_190_195_groupi_n_7825 ,csa_tree_add_190_195_groupi_n_8851);
  xnor csa_tree_add_190_195_groupi_g39716(csa_tree_add_190_195_groupi_n_9245 ,csa_tree_add_190_195_groupi_n_7323 ,csa_tree_add_190_195_groupi_n_8687);
  xnor csa_tree_add_190_195_groupi_g39717(csa_tree_add_190_195_groupi_n_9244 ,csa_tree_add_190_195_groupi_n_8709 ,csa_tree_add_190_195_groupi_n_5392);
  xor csa_tree_add_190_195_groupi_g39719(csa_tree_add_190_195_groupi_n_9243 ,csa_tree_add_190_195_groupi_n_7508 ,csa_tree_add_190_195_groupi_n_8870);
  xnor csa_tree_add_190_195_groupi_g39720(csa_tree_add_190_195_groupi_n_9242 ,csa_tree_add_190_195_groupi_n_6259 ,csa_tree_add_190_195_groupi_n_8722);
  xnor csa_tree_add_190_195_groupi_g39721(csa_tree_add_190_195_groupi_n_9241 ,csa_tree_add_190_195_groupi_n_8610 ,csa_tree_add_190_195_groupi_n_7498);
  xnor csa_tree_add_190_195_groupi_g39722(csa_tree_add_190_195_groupi_n_9240 ,csa_tree_add_190_195_groupi_n_7313 ,csa_tree_add_190_195_groupi_n_8838);
  xnor csa_tree_add_190_195_groupi_g39723(csa_tree_add_190_195_groupi_n_9239 ,csa_tree_add_190_195_groupi_n_7504 ,csa_tree_add_190_195_groupi_n_8655);
  xnor csa_tree_add_190_195_groupi_g39724(csa_tree_add_190_195_groupi_n_9238 ,csa_tree_add_190_195_groupi_n_8497 ,csa_tree_add_190_195_groupi_n_8688);
  xnor csa_tree_add_190_195_groupi_g39725(csa_tree_add_190_195_groupi_n_9237 ,csa_tree_add_190_195_groupi_n_77 ,csa_tree_add_190_195_groupi_n_72);
  xnor csa_tree_add_190_195_groupi_g39726(csa_tree_add_190_195_groupi_n_9236 ,csa_tree_add_190_195_groupi_n_8708 ,csa_tree_add_190_195_groupi_n_7179);
  xnor csa_tree_add_190_195_groupi_g39727(csa_tree_add_190_195_groupi_n_9235 ,csa_tree_add_190_195_groupi_n_7598 ,csa_tree_add_190_195_groupi_n_8633);
  xnor csa_tree_add_190_195_groupi_g39728(csa_tree_add_190_195_groupi_n_9234 ,csa_tree_add_190_195_groupi_n_8663 ,csa_tree_add_190_195_groupi_n_8489);
  xnor csa_tree_add_190_195_groupi_g39729(csa_tree_add_190_195_groupi_n_9233 ,csa_tree_add_190_195_groupi_n_7122 ,csa_tree_add_190_195_groupi_n_8862);
  xnor csa_tree_add_190_195_groupi_g39730(csa_tree_add_190_195_groupi_n_9232 ,csa_tree_add_190_195_groupi_n_8635 ,csa_tree_add_190_195_groupi_n_7991);
  xnor csa_tree_add_190_195_groupi_g39731(csa_tree_add_190_195_groupi_n_9231 ,csa_tree_add_190_195_groupi_n_8000 ,csa_tree_add_190_195_groupi_n_8702);
  xor csa_tree_add_190_195_groupi_g39732(csa_tree_add_190_195_groupi_n_9230 ,csa_tree_add_190_195_groupi_n_8339 ,csa_tree_add_190_195_groupi_n_8871);
  xnor csa_tree_add_190_195_groupi_g39734(csa_tree_add_190_195_groupi_n_9229 ,csa_tree_add_190_195_groupi_n_8828 ,csa_tree_add_190_195_groupi_n_8672);
  xnor csa_tree_add_190_195_groupi_g39735(csa_tree_add_190_195_groupi_n_9228 ,csa_tree_add_190_195_groupi_n_8358 ,csa_tree_add_190_195_groupi_n_8698);
  xnor csa_tree_add_190_195_groupi_g39736(csa_tree_add_190_195_groupi_n_9227 ,csa_tree_add_190_195_groupi_n_8327 ,csa_tree_add_190_195_groupi_n_8861);
  xnor csa_tree_add_190_195_groupi_g39737(csa_tree_add_190_195_groupi_n_9226 ,csa_tree_add_190_195_groupi_n_7819 ,csa_tree_add_190_195_groupi_n_8613);
  xnor csa_tree_add_190_195_groupi_g39738(csa_tree_add_190_195_groupi_n_9225 ,csa_tree_add_190_195_groupi_n_8675 ,csa_tree_add_190_195_groupi_n_8525);
  xnor csa_tree_add_190_195_groupi_g39739(csa_tree_add_190_195_groupi_n_9224 ,csa_tree_add_190_195_groupi_n_8712 ,csa_tree_add_190_195_groupi_n_8317);
  xnor csa_tree_add_190_195_groupi_g39740(csa_tree_add_190_195_groupi_n_9223 ,csa_tree_add_190_195_groupi_n_8670 ,csa_tree_add_190_195_groupi_n_8624);
  xnor csa_tree_add_190_195_groupi_g39741(csa_tree_add_190_195_groupi_n_9222 ,csa_tree_add_190_195_groupi_n_8483 ,csa_tree_add_190_195_groupi_n_8695);
  xnor csa_tree_add_190_195_groupi_g39742(csa_tree_add_190_195_groupi_n_9221 ,csa_tree_add_190_195_groupi_n_8507 ,csa_tree_add_190_195_groupi_n_8651);
  xnor csa_tree_add_190_195_groupi_g39743(csa_tree_add_190_195_groupi_n_9220 ,csa_tree_add_190_195_groupi_n_8855 ,csa_tree_add_190_195_groupi_n_8370);
  xnor csa_tree_add_190_195_groupi_g39744(csa_tree_add_190_195_groupi_n_9219 ,csa_tree_add_190_195_groupi_n_7348 ,csa_tree_add_190_195_groupi_n_8873);
  xnor csa_tree_add_190_195_groupi_g39745(csa_tree_add_190_195_groupi_n_9218 ,csa_tree_add_190_195_groupi_n_7603 ,csa_tree_add_190_195_groupi_n_8850);
  xor csa_tree_add_190_195_groupi_g39746(csa_tree_add_190_195_groupi_n_9217 ,csa_tree_add_190_195_groupi_n_8385 ,csa_tree_add_190_195_groupi_n_8619);
  xnor csa_tree_add_190_195_groupi_g39747(csa_tree_add_190_195_groupi_n_9216 ,csa_tree_add_190_195_groupi_n_7585 ,csa_tree_add_190_195_groupi_n_8634);
  xnor csa_tree_add_190_195_groupi_g39748(csa_tree_add_190_195_groupi_n_9215 ,csa_tree_add_190_195_groupi_n_7638 ,csa_tree_add_190_195_groupi_n_8869);
  xnor csa_tree_add_190_195_groupi_g39749(csa_tree_add_190_195_groupi_n_9214 ,csa_tree_add_190_195_groupi_n_8830 ,csa_tree_add_190_195_groupi_n_8872);
  xnor csa_tree_add_190_195_groupi_g39750(csa_tree_add_190_195_groupi_n_9213 ,csa_tree_add_190_195_groupi_n_8646 ,csa_tree_add_190_195_groupi_n_8837);
  xnor csa_tree_add_190_195_groupi_g39751(csa_tree_add_190_195_groupi_n_9212 ,csa_tree_add_190_195_groupi_n_5533 ,csa_tree_add_190_195_groupi_n_8721);
  xnor csa_tree_add_190_195_groupi_g39752(csa_tree_add_190_195_groupi_n_9211 ,csa_tree_add_190_195_groupi_n_8315 ,csa_tree_add_190_195_groupi_n_8852);
  xnor csa_tree_add_190_195_groupi_g39753(csa_tree_add_190_195_groupi_n_9210 ,csa_tree_add_190_195_groupi_n_8515 ,csa_tree_add_190_195_groupi_n_8644);
  xnor csa_tree_add_190_195_groupi_g39754(csa_tree_add_190_195_groupi_n_9209 ,csa_tree_add_190_195_groupi_n_7824 ,csa_tree_add_190_195_groupi_n_8642);
  xnor csa_tree_add_190_195_groupi_g39755(csa_tree_add_190_195_groupi_n_9208 ,csa_tree_add_190_195_groupi_n_7549 ,csa_tree_add_190_195_groupi_n_8641);
  xnor csa_tree_add_190_195_groupi_g39757(csa_tree_add_190_195_groupi_n_9207 ,csa_tree_add_190_195_groupi_n_8017 ,csa_tree_add_190_195_groupi_n_8859);
  xnor csa_tree_add_190_195_groupi_g39758(csa_tree_add_190_195_groupi_n_9206 ,csa_tree_add_190_195_groupi_n_6964 ,csa_tree_add_190_195_groupi_n_8864);
  xnor csa_tree_add_190_195_groupi_g39759(csa_tree_add_190_195_groupi_n_9205 ,csa_tree_add_190_195_groupi_n_7066 ,csa_tree_add_190_195_groupi_n_8866);
  xnor csa_tree_add_190_195_groupi_g39760(csa_tree_add_190_195_groupi_n_9204 ,csa_tree_add_190_195_groupi_n_8481 ,csa_tree_add_190_195_groupi_n_8700);
  xnor csa_tree_add_190_195_groupi_g39761(csa_tree_add_190_195_groupi_n_9368 ,csa_tree_add_190_195_groupi_n_4601 ,csa_tree_add_190_195_groupi_n_8574);
  xnor csa_tree_add_190_195_groupi_g39762(csa_tree_add_190_195_groupi_n_9367 ,csa_tree_add_190_195_groupi_n_4716 ,csa_tree_add_190_195_groupi_n_8576);
  or csa_tree_add_190_195_groupi_g39763(csa_tree_add_190_195_groupi_n_9365 ,csa_tree_add_190_195_groupi_n_6393 ,csa_tree_add_190_195_groupi_n_8914);
  xnor csa_tree_add_190_195_groupi_g39764(csa_tree_add_190_195_groupi_n_9363 ,csa_tree_add_190_195_groupi_n_6927 ,csa_tree_add_190_195_groupi_n_8550);
  xnor csa_tree_add_190_195_groupi_g39765(csa_tree_add_190_195_groupi_n_9362 ,csa_tree_add_190_195_groupi_n_4704 ,csa_tree_add_190_195_groupi_n_8582);
  xnor csa_tree_add_190_195_groupi_g39766(csa_tree_add_190_195_groupi_n_9361 ,csa_tree_add_190_195_groupi_n_8710 ,csa_tree_add_190_195_groupi_n_6641);
  xnor csa_tree_add_190_195_groupi_g39767(csa_tree_add_190_195_groupi_n_9360 ,csa_tree_add_190_195_groupi_n_5072 ,csa_tree_add_190_195_groupi_n_8555);
  xnor csa_tree_add_190_195_groupi_g39768(csa_tree_add_190_195_groupi_n_9359 ,csa_tree_add_190_195_groupi_n_6573 ,csa_tree_add_190_195_groupi_n_8561);
  xnor csa_tree_add_190_195_groupi_g39769(csa_tree_add_190_195_groupi_n_9358 ,csa_tree_add_190_195_groupi_n_4925 ,csa_tree_add_190_195_groupi_n_8587);
  and csa_tree_add_190_195_groupi_g39770(csa_tree_add_190_195_groupi_n_9357 ,csa_tree_add_190_195_groupi_n_6569 ,csa_tree_add_190_195_groupi_n_8920);
  xnor csa_tree_add_190_195_groupi_g39771(csa_tree_add_190_195_groupi_n_9356 ,csa_tree_add_190_195_groupi_n_8187 ,csa_tree_add_190_195_groupi_n_8577);
  xnor csa_tree_add_190_195_groupi_g39772(csa_tree_add_190_195_groupi_n_9355 ,csa_tree_add_190_195_groupi_n_5069 ,csa_tree_add_190_195_groupi_n_8554);
  xnor csa_tree_add_190_195_groupi_g39773(csa_tree_add_190_195_groupi_n_9354 ,csa_tree_add_190_195_groupi_n_5388 ,csa_tree_add_190_195_groupi_n_8568);
  and csa_tree_add_190_195_groupi_g39774(csa_tree_add_190_195_groupi_n_9353 ,csa_tree_add_190_195_groupi_n_8758 ,csa_tree_add_190_195_groupi_n_8926);
  xnor csa_tree_add_190_195_groupi_g39775(csa_tree_add_190_195_groupi_n_9352 ,csa_tree_add_190_195_groupi_n_5272 ,csa_tree_add_190_195_groupi_n_8566);
  or csa_tree_add_190_195_groupi_g39776(csa_tree_add_190_195_groupi_n_9350 ,csa_tree_add_190_195_groupi_n_6164 ,csa_tree_add_190_195_groupi_n_8916);
  xnor csa_tree_add_190_195_groupi_g39777(csa_tree_add_190_195_groupi_n_9349 ,csa_tree_add_190_195_groupi_n_8720 ,csa_tree_add_190_195_groupi_n_7918);
  xnor csa_tree_add_190_195_groupi_g39778(csa_tree_add_190_195_groupi_n_9348 ,csa_tree_add_190_195_groupi_n_8718 ,csa_tree_add_190_195_groupi_n_6642);
  xnor csa_tree_add_190_195_groupi_g39780(csa_tree_add_190_195_groupi_n_9345 ,csa_tree_add_190_195_groupi_n_8340 ,csa_tree_add_190_195_groupi_n_8558);
  xnor csa_tree_add_190_195_groupi_g39781(csa_tree_add_190_195_groupi_n_9343 ,csa_tree_add_190_195_groupi_n_8044 ,csa_tree_add_190_195_groupi_n_8560);
  xnor csa_tree_add_190_195_groupi_g39782(csa_tree_add_190_195_groupi_n_9341 ,csa_tree_add_190_195_groupi_n_8354 ,csa_tree_add_190_195_groupi_n_8585);
  xnor csa_tree_add_190_195_groupi_g39783(csa_tree_add_190_195_groupi_n_9339 ,csa_tree_add_190_195_groupi_n_8664 ,csa_tree_add_190_195_groupi_n_8549);
  xnor csa_tree_add_190_195_groupi_g39784(csa_tree_add_190_195_groupi_n_9337 ,csa_tree_add_190_195_groupi_n_8395 ,csa_tree_add_190_195_groupi_n_8548);
  xnor csa_tree_add_190_195_groupi_g39785(csa_tree_add_190_195_groupi_n_9335 ,csa_tree_add_190_195_groupi_n_8346 ,csa_tree_add_190_195_groupi_n_8547);
  xnor csa_tree_add_190_195_groupi_g39786(csa_tree_add_190_195_groupi_n_9333 ,csa_tree_add_190_195_groupi_n_8877 ,csa_tree_add_190_195_groupi_n_7910);
  xnor csa_tree_add_190_195_groupi_g39787(csa_tree_add_190_195_groupi_n_9331 ,csa_tree_add_190_195_groupi_n_5506 ,csa_tree_add_190_195_groupi_n_8559);
  xnor csa_tree_add_190_195_groupi_g39788(csa_tree_add_190_195_groupi_n_9330 ,csa_tree_add_190_195_groupi_n_5436 ,csa_tree_add_190_195_groupi_n_8552);
  xnor csa_tree_add_190_195_groupi_g39789(csa_tree_add_190_195_groupi_n_9328 ,csa_tree_add_190_195_groupi_n_8673 ,csa_tree_add_190_195_groupi_n_8583);
  xnor csa_tree_add_190_195_groupi_g39791(csa_tree_add_190_195_groupi_n_9325 ,csa_tree_add_190_195_groupi_n_7329 ,csa_tree_add_190_195_groupi_n_8562);
  xnor csa_tree_add_190_195_groupi_g39792(csa_tree_add_190_195_groupi_n_9323 ,csa_tree_add_190_195_groupi_n_5544 ,csa_tree_add_190_195_groupi_n_8564);
  xnor csa_tree_add_190_195_groupi_g39793(csa_tree_add_190_195_groupi_n_9321 ,csa_tree_add_190_195_groupi_n_8015 ,csa_tree_add_190_195_groupi_n_8565);
  xnor csa_tree_add_190_195_groupi_g39794(csa_tree_add_190_195_groupi_n_9319 ,csa_tree_add_190_195_groupi_n_7194 ,csa_tree_add_190_195_groupi_n_8556);
  xnor csa_tree_add_190_195_groupi_g39795(csa_tree_add_190_195_groupi_n_9318 ,csa_tree_add_190_195_groupi_n_7375 ,csa_tree_add_190_195_groupi_n_8563);
  xnor csa_tree_add_190_195_groupi_g39796(csa_tree_add_190_195_groupi_n_9317 ,csa_tree_add_190_195_groupi_n_8191 ,csa_tree_add_190_195_groupi_n_8557);
  xnor csa_tree_add_190_195_groupi_g39797(csa_tree_add_190_195_groupi_n_9315 ,csa_tree_add_190_195_groupi_n_7599 ,csa_tree_add_190_195_groupi_n_8551);
  xnor csa_tree_add_190_195_groupi_g39798(csa_tree_add_190_195_groupi_n_9314 ,csa_tree_add_190_195_groupi_n_5382 ,csa_tree_add_190_195_groupi_n_113);
  xnor csa_tree_add_190_195_groupi_g39799(csa_tree_add_190_195_groupi_n_9312 ,csa_tree_add_190_195_groupi_n_8701 ,csa_tree_add_190_195_groupi_n_7893);
  xnor csa_tree_add_190_195_groupi_g39801(csa_tree_add_190_195_groupi_n_9309 ,csa_tree_add_190_195_groupi_n_8856 ,csa_tree_add_190_195_groupi_n_7460);
  xnor csa_tree_add_190_195_groupi_g39802(csa_tree_add_190_195_groupi_n_9308 ,csa_tree_add_190_195_groupi_n_5291 ,csa_tree_add_190_195_groupi_n_8573);
  xnor csa_tree_add_190_195_groupi_g39803(csa_tree_add_190_195_groupi_n_9307 ,csa_tree_add_190_195_groupi_n_7332 ,csa_tree_add_190_195_groupi_n_8579);
  xnor csa_tree_add_190_195_groupi_g39804(csa_tree_add_190_195_groupi_n_9304 ,csa_tree_add_190_195_groupi_n_8362 ,csa_tree_add_190_195_groupi_n_8580);
  xnor csa_tree_add_190_195_groupi_g39805(csa_tree_add_190_195_groupi_n_9302 ,csa_tree_add_190_195_groupi_n_7578 ,csa_tree_add_190_195_groupi_n_8567);
  xnor csa_tree_add_190_195_groupi_g39806(csa_tree_add_190_195_groupi_n_9300 ,csa_tree_add_190_195_groupi_n_8213 ,csa_tree_add_190_195_groupi_n_8569);
  xnor csa_tree_add_190_195_groupi_g39807(csa_tree_add_190_195_groupi_n_9299 ,csa_tree_add_190_195_groupi_n_4930 ,csa_tree_add_190_195_groupi_n_8581);
  xnor csa_tree_add_190_195_groupi_g39808(csa_tree_add_190_195_groupi_n_9296 ,csa_tree_add_190_195_groupi_n_5497 ,csa_tree_add_190_195_groupi_n_8570);
  xnor csa_tree_add_190_195_groupi_g39809(csa_tree_add_190_195_groupi_n_9295 ,csa_tree_add_190_195_groupi_n_8863 ,csa_tree_add_190_195_groupi_n_8249);
  xnor csa_tree_add_190_195_groupi_g39810(csa_tree_add_190_195_groupi_n_9293 ,csa_tree_add_190_195_groupi_n_7856 ,csa_tree_add_190_195_groupi_n_8571);
  xnor csa_tree_add_190_195_groupi_g39811(csa_tree_add_190_195_groupi_n_9292 ,csa_tree_add_190_195_groupi_n_7848 ,csa_tree_add_190_195_groupi_n_8572);
  xnor csa_tree_add_190_195_groupi_g39812(csa_tree_add_190_195_groupi_n_9291 ,csa_tree_add_190_195_groupi_n_8647 ,csa_tree_add_190_195_groupi_n_8578);
  xnor csa_tree_add_190_195_groupi_g39813(csa_tree_add_190_195_groupi_n_9289 ,csa_tree_add_190_195_groupi_n_8844 ,csa_tree_add_190_195_groupi_n_6616);
  xnor csa_tree_add_190_195_groupi_g39814(csa_tree_add_190_195_groupi_n_9287 ,csa_tree_add_190_195_groupi_n_7334 ,csa_tree_add_190_195_groupi_n_8575);
  xnor csa_tree_add_190_195_groupi_g39815(csa_tree_add_190_195_groupi_n_9286 ,csa_tree_add_190_195_groupi_n_4700 ,csa_tree_add_190_195_groupi_n_8586);
  or csa_tree_add_190_195_groupi_g39816(csa_tree_add_190_195_groupi_n_9284 ,csa_tree_add_190_195_groupi_n_8593 ,csa_tree_add_190_195_groupi_n_8924);
  not csa_tree_add_190_195_groupi_g39819(csa_tree_add_190_195_groupi_n_9195 ,csa_tree_add_190_195_groupi_n_9194);
  not csa_tree_add_190_195_groupi_g39821(csa_tree_add_190_195_groupi_n_9181 ,csa_tree_add_190_195_groupi_n_9180);
  not csa_tree_add_190_195_groupi_g39822(csa_tree_add_190_195_groupi_n_9178 ,csa_tree_add_190_195_groupi_n_9179);
  not csa_tree_add_190_195_groupi_g39823(csa_tree_add_190_195_groupi_n_9177 ,csa_tree_add_190_195_groupi_n_9176);
  not csa_tree_add_190_195_groupi_g39824(csa_tree_add_190_195_groupi_n_9174 ,csa_tree_add_190_195_groupi_n_9175);
  not csa_tree_add_190_195_groupi_g39825(csa_tree_add_190_195_groupi_n_9172 ,csa_tree_add_190_195_groupi_n_9173);
  not csa_tree_add_190_195_groupi_g39826(csa_tree_add_190_195_groupi_n_9171 ,csa_tree_add_190_195_groupi_n_9170);
  not csa_tree_add_190_195_groupi_g39827(csa_tree_add_190_195_groupi_n_9167 ,csa_tree_add_190_195_groupi_n_9168);
  not csa_tree_add_190_195_groupi_g39828(csa_tree_add_190_195_groupi_n_9165 ,csa_tree_add_190_195_groupi_n_9166);
  not csa_tree_add_190_195_groupi_g39829(csa_tree_add_190_195_groupi_n_9164 ,csa_tree_add_190_195_groupi_n_9163);
  not csa_tree_add_190_195_groupi_g39830(csa_tree_add_190_195_groupi_n_9161 ,csa_tree_add_190_195_groupi_n_9162);
  not csa_tree_add_190_195_groupi_g39831(csa_tree_add_190_195_groupi_n_9160 ,csa_tree_add_190_195_groupi_n_9159);
  not csa_tree_add_190_195_groupi_g39832(csa_tree_add_190_195_groupi_n_9157 ,csa_tree_add_190_195_groupi_n_9158);
  or csa_tree_add_190_195_groupi_g39833(csa_tree_add_190_195_groupi_n_9156 ,csa_tree_add_190_195_groupi_n_7967 ,csa_tree_add_190_195_groupi_n_8708);
  or csa_tree_add_190_195_groupi_g39834(csa_tree_add_190_195_groupi_n_9155 ,csa_tree_add_190_195_groupi_n_8712 ,csa_tree_add_190_195_groupi_n_8591);
  or csa_tree_add_190_195_groupi_g39835(csa_tree_add_190_195_groupi_n_9154 ,csa_tree_add_190_195_groupi_n_7093 ,csa_tree_add_190_195_groupi_n_8631);
  or csa_tree_add_190_195_groupi_g39836(csa_tree_add_190_195_groupi_n_9153 ,csa_tree_add_190_195_groupi_n_7601 ,csa_tree_add_190_195_groupi_n_8652);
  nor csa_tree_add_190_195_groupi_g39837(csa_tree_add_190_195_groupi_n_9152 ,csa_tree_add_190_195_groupi_n_7092 ,csa_tree_add_190_195_groupi_n_8632);
  and csa_tree_add_190_195_groupi_g39838(csa_tree_add_190_195_groupi_n_9151 ,csa_tree_add_190_195_groupi_n_7598 ,csa_tree_add_190_195_groupi_n_8633);
  nor csa_tree_add_190_195_groupi_g39839(csa_tree_add_190_195_groupi_n_9150 ,csa_tree_add_190_195_groupi_n_7600 ,csa_tree_add_190_195_groupi_n_8653);
  or csa_tree_add_190_195_groupi_g39840(csa_tree_add_190_195_groupi_n_9149 ,csa_tree_add_190_195_groupi_n_7322 ,csa_tree_add_190_195_groupi_n_8686);
  nor csa_tree_add_190_195_groupi_g39841(csa_tree_add_190_195_groupi_n_9148 ,csa_tree_add_190_195_groupi_n_7818 ,csa_tree_add_190_195_groupi_n_8613);
  or csa_tree_add_190_195_groupi_g39842(csa_tree_add_190_195_groupi_n_9147 ,csa_tree_add_190_195_groupi_n_7819 ,csa_tree_add_190_195_groupi_n_8612);
  nor csa_tree_add_190_195_groupi_g39843(csa_tree_add_190_195_groupi_n_9146 ,csa_tree_add_190_195_groupi_n_8693 ,csa_tree_add_190_195_groupi_n_8626);
  nor csa_tree_add_190_195_groupi_g39844(csa_tree_add_190_195_groupi_n_9145 ,csa_tree_add_190_195_groupi_n_7323 ,csa_tree_add_190_195_groupi_n_8687);
  or csa_tree_add_190_195_groupi_g39845(csa_tree_add_190_195_groupi_n_9144 ,csa_tree_add_190_195_groupi_n_8692 ,csa_tree_add_190_195_groupi_n_8625);
  nor csa_tree_add_190_195_groupi_g39846(csa_tree_add_190_195_groupi_n_9143 ,csa_tree_add_190_195_groupi_n_6521 ,csa_tree_add_190_195_groupi_n_8709);
  or csa_tree_add_190_195_groupi_g39847(csa_tree_add_190_195_groupi_n_9142 ,csa_tree_add_190_195_groupi_n_5453 ,csa_tree_add_190_195_groupi_n_8675);
  and csa_tree_add_190_195_groupi_g39848(csa_tree_add_190_195_groupi_n_9141 ,csa_tree_add_190_195_groupi_n_7378 ,csa_tree_add_190_195_groupi_n_8673);
  nor csa_tree_add_190_195_groupi_g39849(csa_tree_add_190_195_groupi_n_9140 ,csa_tree_add_190_195_groupi_n_5454 ,csa_tree_add_190_195_groupi_n_8674);
  or csa_tree_add_190_195_groupi_g39850(csa_tree_add_190_195_groupi_n_9139 ,csa_tree_add_190_195_groupi_n_7378 ,csa_tree_add_190_195_groupi_n_8673);
  or csa_tree_add_190_195_groupi_g39851(csa_tree_add_190_195_groupi_n_9138 ,csa_tree_add_190_195_groupi_n_8669 ,csa_tree_add_190_195_groupi_n_8624);
  nor csa_tree_add_190_195_groupi_g39852(csa_tree_add_190_195_groupi_n_9137 ,csa_tree_add_190_195_groupi_n_8670 ,csa_tree_add_190_195_groupi_n_8623);
  or csa_tree_add_190_195_groupi_g39853(csa_tree_add_190_195_groupi_n_9136 ,csa_tree_add_190_195_groupi_n_8827 ,csa_tree_add_190_195_groupi_n_8671);
  and csa_tree_add_190_195_groupi_g39854(csa_tree_add_190_195_groupi_n_9135 ,csa_tree_add_190_195_groupi_n_8523 ,csa_tree_add_190_195_groupi_n_8788);
  nor csa_tree_add_190_195_groupi_g39855(csa_tree_add_190_195_groupi_n_9134 ,csa_tree_add_190_195_groupi_n_8828 ,csa_tree_add_190_195_groupi_n_8672);
  and csa_tree_add_190_195_groupi_g39856(csa_tree_add_190_195_groupi_n_9133 ,csa_tree_add_190_195_groupi_n_7988 ,csa_tree_add_190_195_groupi_n_8662);
  or csa_tree_add_190_195_groupi_g39857(csa_tree_add_190_195_groupi_n_9132 ,csa_tree_add_190_195_groupi_n_8370 ,csa_tree_add_190_195_groupi_n_8620);
  and csa_tree_add_190_195_groupi_g39858(csa_tree_add_190_195_groupi_n_9131 ,csa_tree_add_190_195_groupi_n_8370 ,csa_tree_add_190_195_groupi_n_8620);
  or csa_tree_add_190_195_groupi_g39859(csa_tree_add_190_195_groupi_n_9130 ,csa_tree_add_190_195_groupi_n_7602 ,csa_tree_add_190_195_groupi_n_8661);
  nor csa_tree_add_190_195_groupi_g39860(csa_tree_add_190_195_groupi_n_9129 ,csa_tree_add_190_195_groupi_n_7603 ,csa_tree_add_190_195_groupi_n_112);
  and csa_tree_add_190_195_groupi_g39861(csa_tree_add_190_195_groupi_n_9128 ,csa_tree_add_190_195_groupi_n_7313 ,csa_tree_add_190_195_groupi_n_8838);
  nor csa_tree_add_190_195_groupi_g39862(csa_tree_add_190_195_groupi_n_9127 ,csa_tree_add_190_195_groupi_n_7130 ,csa_tree_add_190_195_groupi_n_8832);
  or csa_tree_add_190_195_groupi_g39863(csa_tree_add_190_195_groupi_n_9126 ,csa_tree_add_190_195_groupi_n_8206 ,csa_tree_add_190_195_groupi_n_8619);
  nor csa_tree_add_190_195_groupi_g39864(csa_tree_add_190_195_groupi_n_9125 ,csa_tree_add_190_195_groupi_n_8207 ,csa_tree_add_190_195_groupi_n_8618);
  nor csa_tree_add_190_195_groupi_g39865(csa_tree_add_190_195_groupi_n_9124 ,csa_tree_add_190_195_groupi_n_7313 ,csa_tree_add_190_195_groupi_n_8838);
  nor csa_tree_add_190_195_groupi_g39866(csa_tree_add_190_195_groupi_n_9123 ,csa_tree_add_190_195_groupi_n_6395 ,csa_tree_add_190_195_groupi_n_8844);
  or csa_tree_add_190_195_groupi_g39867(csa_tree_add_190_195_groupi_n_9122 ,csa_tree_add_190_195_groupi_n_7131 ,csa_tree_add_190_195_groupi_n_8831);
  nor csa_tree_add_190_195_groupi_g39868(csa_tree_add_190_195_groupi_n_9121 ,csa_tree_add_190_195_groupi_n_7549 ,csa_tree_add_190_195_groupi_n_8640);
  or csa_tree_add_190_195_groupi_g39869(csa_tree_add_190_195_groupi_n_9120 ,csa_tree_add_190_195_groupi_n_7548 ,csa_tree_add_190_195_groupi_n_8641);
  or csa_tree_add_190_195_groupi_g39870(csa_tree_add_190_195_groupi_n_9119 ,csa_tree_add_190_195_groupi_n_8233 ,csa_tree_add_190_195_groupi_n_8787);
  or csa_tree_add_190_195_groupi_g39871(csa_tree_add_190_195_groupi_n_9118 ,csa_tree_add_190_195_groupi_n_7657 ,csa_tree_add_190_195_groupi_n_8773);
  and csa_tree_add_190_195_groupi_g39872(csa_tree_add_190_195_groupi_n_9117 ,csa_tree_add_190_195_groupi_n_8498 ,csa_tree_add_190_195_groupi_n_8688);
  nor csa_tree_add_190_195_groupi_g39873(csa_tree_add_190_195_groupi_n_9116 ,csa_tree_add_190_195_groupi_n_7817 ,csa_tree_add_190_195_groupi_n_8877);
  and csa_tree_add_190_195_groupi_g39874(csa_tree_add_190_195_groupi_n_9115 ,csa_tree_add_190_195_groupi_n_8110 ,csa_tree_add_190_195_groupi_n_8851);
  or csa_tree_add_190_195_groupi_g39875(csa_tree_add_190_195_groupi_n_9114 ,csa_tree_add_190_195_groupi_n_6845 ,csa_tree_add_190_195_groupi_n_8705);
  or csa_tree_add_190_195_groupi_g39876(csa_tree_add_190_195_groupi_n_9113 ,csa_tree_add_190_195_groupi_n_7636 ,csa_tree_add_190_195_groupi_n_8621);
  nor csa_tree_add_190_195_groupi_g39877(csa_tree_add_190_195_groupi_n_9112 ,csa_tree_add_190_195_groupi_n_7637 ,csa_tree_add_190_195_groupi_n_8622);
  nor csa_tree_add_190_195_groupi_g39878(csa_tree_add_190_195_groupi_n_9111 ,csa_tree_add_190_195_groupi_n_7748 ,csa_tree_add_190_195_groupi_n_8866);
  or csa_tree_add_190_195_groupi_g39879(csa_tree_add_190_195_groupi_n_9110 ,csa_tree_add_190_195_groupi_n_6325 ,csa_tree_add_190_195_groupi_n_8716);
  and csa_tree_add_190_195_groupi_g39880(csa_tree_add_190_195_groupi_n_9109 ,csa_tree_add_190_195_groupi_n_7262 ,csa_tree_add_190_195_groupi_n_8856);
  or csa_tree_add_190_195_groupi_g39881(csa_tree_add_190_195_groupi_n_9108 ,csa_tree_add_190_195_groupi_n_8860 ,csa_tree_add_190_195_groupi_n_8748);
  or csa_tree_add_190_195_groupi_g39882(csa_tree_add_190_195_groupi_n_9107 ,csa_tree_add_190_195_groupi_n_8819 ,csa_tree_add_190_195_groupi_n_8638);
  or csa_tree_add_190_195_groupi_g39883(csa_tree_add_190_195_groupi_n_9106 ,csa_tree_add_190_195_groupi_n_7358 ,csa_tree_add_190_195_groupi_n_8696);
  nor csa_tree_add_190_195_groupi_g39884(csa_tree_add_190_195_groupi_n_9105 ,csa_tree_add_190_195_groupi_n_7357 ,csa_tree_add_190_195_groupi_n_8697);
  and csa_tree_add_190_195_groupi_g39885(csa_tree_add_190_195_groupi_n_9104 ,csa_tree_add_190_195_groupi_n_7516 ,csa_tree_add_190_195_groupi_n_8664);
  nor csa_tree_add_190_195_groupi_g39886(csa_tree_add_190_195_groupi_n_9103 ,csa_tree_add_190_195_groupi_n_8820 ,csa_tree_add_190_195_groupi_n_8639);
  or csa_tree_add_190_195_groupi_g39887(csa_tree_add_190_195_groupi_n_9102 ,csa_tree_add_190_195_groupi_n_8744 ,csa_tree_add_190_195_groupi_n_8715);
  or csa_tree_add_190_195_groupi_g39888(csa_tree_add_190_195_groupi_n_9101 ,csa_tree_add_190_195_groupi_n_8543 ,csa_tree_add_190_195_groupi_n_8724);
  nor csa_tree_add_190_195_groupi_g39889(csa_tree_add_190_195_groupi_n_9100 ,csa_tree_add_190_195_groupi_n_8700 ,csa_tree_add_190_195_groupi_n_8741);
  or csa_tree_add_190_195_groupi_g39890(csa_tree_add_190_195_groupi_n_9099 ,csa_tree_add_190_195_groupi_n_7832 ,csa_tree_add_190_195_groupi_n_8616);
  nor csa_tree_add_190_195_groupi_g39891(csa_tree_add_190_195_groupi_n_9098 ,csa_tree_add_190_195_groupi_n_7833 ,csa_tree_add_190_195_groupi_n_8615);
  and csa_tree_add_190_195_groupi_g39892(csa_tree_add_190_195_groupi_n_9097 ,csa_tree_add_190_195_groupi_n_8040 ,csa_tree_add_190_195_groupi_n_8809);
  or csa_tree_add_190_195_groupi_g39893(csa_tree_add_190_195_groupi_n_9096 ,csa_tree_add_190_195_groupi_n_7618 ,csa_tree_add_190_195_groupi_n_8682);
  nor csa_tree_add_190_195_groupi_g39894(csa_tree_add_190_195_groupi_n_9095 ,csa_tree_add_190_195_groupi_n_7619 ,csa_tree_add_190_195_groupi_n_8683);
  and csa_tree_add_190_195_groupi_g39895(csa_tree_add_190_195_groupi_n_9094 ,csa_tree_add_190_195_groupi_n_8734 ,csa_tree_add_190_195_groupi_n_8861);
  or csa_tree_add_190_195_groupi_g39896(csa_tree_add_190_195_groupi_n_9093 ,csa_tree_add_190_195_groupi_n_8510 ,csa_tree_add_190_195_groupi_n_8731);
  and csa_tree_add_190_195_groupi_g39897(csa_tree_add_190_195_groupi_n_9092 ,csa_tree_add_190_195_groupi_n_8359 ,csa_tree_add_190_195_groupi_n_8698);
  and csa_tree_add_190_195_groupi_g39898(csa_tree_add_190_195_groupi_n_9091 ,csa_tree_add_190_195_groupi_n_7702 ,csa_tree_add_190_195_groupi_n_8720);
  or csa_tree_add_190_195_groupi_g39899(csa_tree_add_190_195_groupi_n_9090 ,csa_tree_add_190_195_groupi_n_7507 ,csa_tree_add_190_195_groupi_n_8676);
  nor csa_tree_add_190_195_groupi_g39900(csa_tree_add_190_195_groupi_n_9089 ,csa_tree_add_190_195_groupi_n_7508 ,csa_tree_add_190_195_groupi_n_8677);
  or csa_tree_add_190_195_groupi_g39901(csa_tree_add_190_195_groupi_n_9088 ,csa_tree_add_190_195_groupi_n_7598 ,csa_tree_add_190_195_groupi_n_8633);
  and csa_tree_add_190_195_groupi_g39902(csa_tree_add_190_195_groupi_n_9087 ,csa_tree_add_190_195_groupi_n_7951 ,csa_tree_add_190_195_groupi_n_8873);
  or csa_tree_add_190_195_groupi_g39903(csa_tree_add_190_195_groupi_n_9086 ,csa_tree_add_190_195_groupi_n_7991 ,csa_tree_add_190_195_groupi_n_8635);
  or csa_tree_add_190_195_groupi_g39904(csa_tree_add_190_195_groupi_n_9085 ,csa_tree_add_190_195_groupi_n_7745 ,csa_tree_add_190_195_groupi_n_8701);
  and csa_tree_add_190_195_groupi_g39905(csa_tree_add_190_195_groupi_n_9084 ,csa_tree_add_190_195_groupi_n_8663 ,csa_tree_add_190_195_groupi_n_8489);
  or csa_tree_add_190_195_groupi_g39906(csa_tree_add_190_195_groupi_n_9083 ,csa_tree_add_190_195_groupi_n_8663 ,csa_tree_add_190_195_groupi_n_8489);
  and csa_tree_add_190_195_groupi_g39907(csa_tree_add_190_195_groupi_n_9082 ,csa_tree_add_190_195_groupi_n_7991 ,csa_tree_add_190_195_groupi_n_8635);
  or csa_tree_add_190_195_groupi_g39908(csa_tree_add_190_195_groupi_n_9081 ,csa_tree_add_190_195_groupi_n_7398 ,csa_tree_add_190_195_groupi_n_8728);
  or csa_tree_add_190_195_groupi_g39909(csa_tree_add_190_195_groupi_n_9080 ,csa_tree_add_190_195_groupi_n_7516 ,csa_tree_add_190_195_groupi_n_8664);
  or csa_tree_add_190_195_groupi_g39910(csa_tree_add_190_195_groupi_n_9079 ,csa_tree_add_190_195_groupi_n_8223 ,csa_tree_add_190_195_groupi_n_8771);
  and csa_tree_add_190_195_groupi_g39911(csa_tree_add_190_195_groupi_n_9078 ,csa_tree_add_190_195_groupi_n_8057 ,csa_tree_add_190_195_groupi_n_8739);
  nor csa_tree_add_190_195_groupi_g39912(csa_tree_add_190_195_groupi_n_9077 ,csa_tree_add_190_195_groupi_n_8869 ,csa_tree_add_190_195_groupi_n_8179);
  or csa_tree_add_190_195_groupi_g39913(csa_tree_add_190_195_groupi_n_9076 ,csa_tree_add_190_195_groupi_n_7988 ,csa_tree_add_190_195_groupi_n_8662);
  and csa_tree_add_190_195_groupi_g39914(csa_tree_add_190_195_groupi_n_9075 ,csa_tree_add_190_195_groupi_n_8603 ,csa_tree_add_190_195_groupi_n_8383);
  nor csa_tree_add_190_195_groupi_g39915(csa_tree_add_190_195_groupi_n_9074 ,csa_tree_add_190_195_groupi_n_8498 ,csa_tree_add_190_195_groupi_n_8688);
  or csa_tree_add_190_195_groupi_g39916(csa_tree_add_190_195_groupi_n_9073 ,csa_tree_add_190_195_groupi_n_8038 ,csa_tree_add_190_195_groupi_n_8743);
  and csa_tree_add_190_195_groupi_g39917(csa_tree_add_190_195_groupi_n_9072 ,csa_tree_add_190_195_groupi_n_8656 ,csa_tree_add_190_195_groupi_n_8818);
  or csa_tree_add_190_195_groupi_g39918(csa_tree_add_190_195_groupi_n_9071 ,csa_tree_add_190_195_groupi_n_8656 ,csa_tree_add_190_195_groupi_n_8818);
  nor csa_tree_add_190_195_groupi_g39919(csa_tree_add_190_195_groupi_n_9070 ,csa_tree_add_190_195_groupi_n_8864 ,csa_tree_add_190_195_groupi_n_8754);
  or csa_tree_add_190_195_groupi_g39920(csa_tree_add_190_195_groupi_n_9069 ,csa_tree_add_190_195_groupi_n_7972 ,csa_tree_add_190_195_groupi_n_8863);
  or csa_tree_add_190_195_groupi_g39921(csa_tree_add_190_195_groupi_n_9068 ,csa_tree_add_190_195_groupi_n_7504 ,csa_tree_add_190_195_groupi_n_8654);
  nor csa_tree_add_190_195_groupi_g39922(csa_tree_add_190_195_groupi_n_9067 ,csa_tree_add_190_195_groupi_n_7503 ,csa_tree_add_190_195_groupi_n_8655);
  and csa_tree_add_190_195_groupi_g39923(csa_tree_add_190_195_groupi_n_9066 ,csa_tree_add_190_195_groupi_n_8752 ,csa_tree_add_190_195_groupi_n_8722);
  or csa_tree_add_190_195_groupi_g39924(csa_tree_add_190_195_groupi_n_9065 ,csa_tree_add_190_195_groupi_n_7858 ,csa_tree_add_190_195_groupi_n_8759);
  or csa_tree_add_190_195_groupi_g39925(csa_tree_add_190_195_groupi_n_9064 ,csa_tree_add_190_195_groupi_n_8717 ,csa_tree_add_190_195_groupi_n_8456);
  or csa_tree_add_190_195_groupi_g39926(csa_tree_add_190_195_groupi_n_9063 ,csa_tree_add_190_195_groupi_n_7498 ,csa_tree_add_190_195_groupi_n_8610);
  or csa_tree_add_190_195_groupi_g39927(csa_tree_add_190_195_groupi_n_9062 ,csa_tree_add_190_195_groupi_n_8458 ,csa_tree_add_190_195_groupi_n_8703);
  and csa_tree_add_190_195_groupi_g39928(csa_tree_add_190_195_groupi_n_9061 ,csa_tree_add_190_195_groupi_n_7498 ,csa_tree_add_190_195_groupi_n_8610);
  nor csa_tree_add_190_195_groupi_g39929(csa_tree_add_190_195_groupi_n_9060 ,csa_tree_add_190_195_groupi_n_8359 ,csa_tree_add_190_195_groupi_n_8698);
  nor csa_tree_add_190_195_groupi_g39930(csa_tree_add_190_195_groupi_n_9059 ,csa_tree_add_190_195_groupi_n_7582 ,csa_tree_add_190_195_groupi_n_8833);
  or csa_tree_add_190_195_groupi_g39931(csa_tree_add_190_195_groupi_n_9058 ,csa_tree_add_190_195_groupi_n_7581 ,csa_tree_add_190_195_groupi_n_8834);
  and csa_tree_add_190_195_groupi_g39932(csa_tree_add_190_195_groupi_n_9057 ,csa_tree_add_190_195_groupi_n_8793 ,csa_tree_add_190_195_groupi_n_8706);
  or csa_tree_add_190_195_groupi_g39933(csa_tree_add_190_195_groupi_n_9056 ,csa_tree_add_190_195_groupi_n_8516 ,csa_tree_add_190_195_groupi_n_8777);
  and csa_tree_add_190_195_groupi_g39934(csa_tree_add_190_195_groupi_n_9055 ,csa_tree_add_190_195_groupi_n_7824 ,csa_tree_add_190_195_groupi_n_8642);
  or csa_tree_add_190_195_groupi_g39935(csa_tree_add_190_195_groupi_n_9054 ,csa_tree_add_190_195_groupi_n_7824 ,csa_tree_add_190_195_groupi_n_8642);
  or csa_tree_add_190_195_groupi_g39936(csa_tree_add_190_195_groupi_n_9053 ,csa_tree_add_190_195_groupi_n_8387 ,csa_tree_add_190_195_groupi_n_8791);
  and csa_tree_add_190_195_groupi_g39937(csa_tree_add_190_195_groupi_n_9203 ,csa_tree_add_190_195_groupi_n_7740 ,csa_tree_add_190_195_groupi_n_8756);
  and csa_tree_add_190_195_groupi_g39938(csa_tree_add_190_195_groupi_n_9202 ,csa_tree_add_190_195_groupi_n_6412 ,csa_tree_add_190_195_groupi_n_8764);
  and csa_tree_add_190_195_groupi_g39939(csa_tree_add_190_195_groupi_n_9201 ,csa_tree_add_190_195_groupi_n_8448 ,csa_tree_add_190_195_groupi_n_8761);
  or csa_tree_add_190_195_groupi_g39940(csa_tree_add_190_195_groupi_n_9200 ,csa_tree_add_190_195_groupi_n_8445 ,csa_tree_add_190_195_groupi_n_8779);
  and csa_tree_add_190_195_groupi_g39941(csa_tree_add_190_195_groupi_n_9199 ,csa_tree_add_190_195_groupi_n_5773 ,csa_tree_add_190_195_groupi_n_8776);
  and csa_tree_add_190_195_groupi_g39942(csa_tree_add_190_195_groupi_n_9198 ,csa_tree_add_190_195_groupi_n_8430 ,csa_tree_add_190_195_groupi_n_8740);
  and csa_tree_add_190_195_groupi_g39943(csa_tree_add_190_195_groupi_n_9197 ,csa_tree_add_190_195_groupi_n_6102 ,csa_tree_add_190_195_groupi_n_8762);
  and csa_tree_add_190_195_groupi_g39944(csa_tree_add_190_195_groupi_n_9196 ,csa_tree_add_190_195_groupi_n_8412 ,csa_tree_add_190_195_groupi_n_8763);
  or csa_tree_add_190_195_groupi_g39945(csa_tree_add_190_195_groupi_n_9194 ,csa_tree_add_190_195_groupi_n_8459 ,csa_tree_add_190_195_groupi_n_8765);
  or csa_tree_add_190_195_groupi_g39946(csa_tree_add_190_195_groupi_n_9193 ,csa_tree_add_190_195_groupi_n_6095 ,csa_tree_add_190_195_groupi_n_8769);
  or csa_tree_add_190_195_groupi_g39947(csa_tree_add_190_195_groupi_n_9192 ,csa_tree_add_190_195_groupi_n_7249 ,csa_tree_add_190_195_groupi_n_8733);
  or csa_tree_add_190_195_groupi_g39948(csa_tree_add_190_195_groupi_n_9191 ,csa_tree_add_190_195_groupi_n_8476 ,csa_tree_add_190_195_groupi_n_8785);
  and csa_tree_add_190_195_groupi_g39949(csa_tree_add_190_195_groupi_n_9190 ,csa_tree_add_190_195_groupi_n_8400 ,csa_tree_add_190_195_groupi_n_8735);
  and csa_tree_add_190_195_groupi_g39950(csa_tree_add_190_195_groupi_n_9189 ,csa_tree_add_190_195_groupi_n_8468 ,csa_tree_add_190_195_groupi_n_8799);
  and csa_tree_add_190_195_groupi_g39951(csa_tree_add_190_195_groupi_n_9188 ,csa_tree_add_190_195_groupi_n_7975 ,csa_tree_add_190_195_groupi_n_8747);
  and csa_tree_add_190_195_groupi_g39952(csa_tree_add_190_195_groupi_n_9187 ,csa_tree_add_190_195_groupi_n_8299 ,csa_tree_add_190_195_groupi_n_8798);
  or csa_tree_add_190_195_groupi_g39953(csa_tree_add_190_195_groupi_n_9186 ,csa_tree_add_190_195_groupi_n_8114 ,csa_tree_add_190_195_groupi_n_8726);
  or csa_tree_add_190_195_groupi_g39954(csa_tree_add_190_195_groupi_n_9185 ,csa_tree_add_190_195_groupi_n_8418 ,csa_tree_add_190_195_groupi_n_8729);
  or csa_tree_add_190_195_groupi_g39955(csa_tree_add_190_195_groupi_n_9184 ,csa_tree_add_190_195_groupi_n_8291 ,csa_tree_add_190_195_groupi_n_8755);
  and csa_tree_add_190_195_groupi_g39956(csa_tree_add_190_195_groupi_n_9183 ,csa_tree_add_190_195_groupi_n_8078 ,csa_tree_add_190_195_groupi_n_8780);
  or csa_tree_add_190_195_groupi_g39957(csa_tree_add_190_195_groupi_n_9182 ,csa_tree_add_190_195_groupi_n_8308 ,csa_tree_add_190_195_groupi_n_8784);
  and csa_tree_add_190_195_groupi_g39958(csa_tree_add_190_195_groupi_n_9180 ,csa_tree_add_190_195_groupi_n_8473 ,csa_tree_add_190_195_groupi_n_8782);
  or csa_tree_add_190_195_groupi_g39959(csa_tree_add_190_195_groupi_n_9179 ,csa_tree_add_190_195_groupi_n_5728 ,csa_tree_add_190_195_groupi_n_8774);
  and csa_tree_add_190_195_groupi_g39960(csa_tree_add_190_195_groupi_n_9176 ,csa_tree_add_190_195_groupi_n_8467 ,csa_tree_add_190_195_groupi_n_8772);
  or csa_tree_add_190_195_groupi_g39961(csa_tree_add_190_195_groupi_n_9175 ,csa_tree_add_190_195_groupi_n_6212 ,csa_tree_add_190_195_groupi_n_8730);
  or csa_tree_add_190_195_groupi_g39962(csa_tree_add_190_195_groupi_n_9173 ,csa_tree_add_190_195_groupi_n_2937 ,csa_tree_add_190_195_groupi_n_8757);
  and csa_tree_add_190_195_groupi_g39963(csa_tree_add_190_195_groupi_n_9170 ,csa_tree_add_190_195_groupi_n_8064 ,csa_tree_add_190_195_groupi_n_8789);
  and csa_tree_add_190_195_groupi_g39964(csa_tree_add_190_195_groupi_n_9169 ,csa_tree_add_190_195_groupi_n_6321 ,csa_tree_add_190_195_groupi_n_8767);
  or csa_tree_add_190_195_groupi_g39965(csa_tree_add_190_195_groupi_n_9168 ,csa_tree_add_190_195_groupi_n_8296 ,csa_tree_add_190_195_groupi_n_8768);
  or csa_tree_add_190_195_groupi_g39966(csa_tree_add_190_195_groupi_n_9166 ,csa_tree_add_190_195_groupi_n_6874 ,csa_tree_add_190_195_groupi_n_8783);
  or csa_tree_add_190_195_groupi_g39967(csa_tree_add_190_195_groupi_n_9163 ,csa_tree_add_190_195_groupi_n_7297 ,csa_tree_add_190_195_groupi_n_8800);
  or csa_tree_add_190_195_groupi_g39968(csa_tree_add_190_195_groupi_n_9162 ,csa_tree_add_190_195_groupi_n_8474 ,csa_tree_add_190_195_groupi_n_8805);
  or csa_tree_add_190_195_groupi_g39969(csa_tree_add_190_195_groupi_n_9159 ,csa_tree_add_190_195_groupi_n_8177 ,csa_tree_add_190_195_groupi_n_8806);
  and csa_tree_add_190_195_groupi_g39970(csa_tree_add_190_195_groupi_n_9158 ,csa_tree_add_190_195_groupi_n_8305 ,csa_tree_add_190_195_groupi_n_8808);
  not csa_tree_add_190_195_groupi_g39972(csa_tree_add_190_195_groupi_n_9050 ,csa_tree_add_190_195_groupi_n_9049);
  not csa_tree_add_190_195_groupi_g39973(csa_tree_add_190_195_groupi_n_9047 ,csa_tree_add_190_195_groupi_n_25);
  not csa_tree_add_190_195_groupi_g39975(csa_tree_add_190_195_groupi_n_9041 ,csa_tree_add_190_195_groupi_n_9040);
  not csa_tree_add_190_195_groupi_g39976(csa_tree_add_190_195_groupi_n_9034 ,csa_tree_add_190_195_groupi_n_9033);
  not csa_tree_add_190_195_groupi_g39977(csa_tree_add_190_195_groupi_n_9032 ,csa_tree_add_190_195_groupi_n_9031);
  not csa_tree_add_190_195_groupi_g39978(csa_tree_add_190_195_groupi_n_9029 ,csa_tree_add_190_195_groupi_n_9028);
  not csa_tree_add_190_195_groupi_g39979(csa_tree_add_190_195_groupi_n_9027 ,csa_tree_add_190_195_groupi_n_9026);
  not csa_tree_add_190_195_groupi_g39980(csa_tree_add_190_195_groupi_n_9025 ,csa_tree_add_190_195_groupi_n_9024);
  not csa_tree_add_190_195_groupi_g39981(csa_tree_add_190_195_groupi_n_9023 ,csa_tree_add_190_195_groupi_n_9022);
  not csa_tree_add_190_195_groupi_g39982(csa_tree_add_190_195_groupi_n_9021 ,csa_tree_add_190_195_groupi_n_9020);
  not csa_tree_add_190_195_groupi_g39983(csa_tree_add_190_195_groupi_n_9019 ,csa_tree_add_190_195_groupi_n_9018);
  not csa_tree_add_190_195_groupi_g39984(csa_tree_add_190_195_groupi_n_9016 ,csa_tree_add_190_195_groupi_n_9017);
  not csa_tree_add_190_195_groupi_g39985(csa_tree_add_190_195_groupi_n_9015 ,csa_tree_add_190_195_groupi_n_9014);
  not csa_tree_add_190_195_groupi_g39986(csa_tree_add_190_195_groupi_n_9011 ,csa_tree_add_190_195_groupi_n_9010);
  not csa_tree_add_190_195_groupi_g39987(csa_tree_add_190_195_groupi_n_9008 ,csa_tree_add_190_195_groupi_n_9009);
  not csa_tree_add_190_195_groupi_g39988(csa_tree_add_190_195_groupi_n_9007 ,csa_tree_add_190_195_groupi_n_9006);
  not csa_tree_add_190_195_groupi_g39989(csa_tree_add_190_195_groupi_n_9004 ,csa_tree_add_190_195_groupi_n_9005);
  not csa_tree_add_190_195_groupi_g39990(csa_tree_add_190_195_groupi_n_9003 ,csa_tree_add_190_195_groupi_n_9002);
  not csa_tree_add_190_195_groupi_g39991(csa_tree_add_190_195_groupi_n_9001 ,csa_tree_add_190_195_groupi_n_9000);
  not csa_tree_add_190_195_groupi_g39992(csa_tree_add_190_195_groupi_n_8999 ,csa_tree_add_190_195_groupi_n_8998);
  not csa_tree_add_190_195_groupi_g39993(csa_tree_add_190_195_groupi_n_8997 ,csa_tree_add_190_195_groupi_n_8996);
  not csa_tree_add_190_195_groupi_g39994(csa_tree_add_190_195_groupi_n_8995 ,csa_tree_add_190_195_groupi_n_105);
  not csa_tree_add_190_195_groupi_g39995(csa_tree_add_190_195_groupi_n_8993 ,csa_tree_add_190_195_groupi_n_8994);
  not csa_tree_add_190_195_groupi_g39996(csa_tree_add_190_195_groupi_n_8991 ,csa_tree_add_190_195_groupi_n_8992);
  not csa_tree_add_190_195_groupi_g39997(csa_tree_add_190_195_groupi_n_8990 ,csa_tree_add_190_195_groupi_n_8989);
  not csa_tree_add_190_195_groupi_g39998(csa_tree_add_190_195_groupi_n_8988 ,csa_tree_add_190_195_groupi_n_103);
  not csa_tree_add_190_195_groupi_g39999(csa_tree_add_190_195_groupi_n_8987 ,csa_tree_add_190_195_groupi_n_8986);
  not csa_tree_add_190_195_groupi_g40000(csa_tree_add_190_195_groupi_n_8984 ,csa_tree_add_190_195_groupi_n_8985);
  not csa_tree_add_190_195_groupi_g40001(csa_tree_add_190_195_groupi_n_8983 ,csa_tree_add_190_195_groupi_n_8982);
  not csa_tree_add_190_195_groupi_g40002(csa_tree_add_190_195_groupi_n_8981 ,csa_tree_add_190_195_groupi_n_8980);
  not csa_tree_add_190_195_groupi_g40003(csa_tree_add_190_195_groupi_n_8979 ,csa_tree_add_190_195_groupi_n_8978);
  not csa_tree_add_190_195_groupi_g40004(csa_tree_add_190_195_groupi_n_8977 ,csa_tree_add_190_195_groupi_n_8976);
  not csa_tree_add_190_195_groupi_g40005(csa_tree_add_190_195_groupi_n_8973 ,csa_tree_add_190_195_groupi_n_8972);
  not csa_tree_add_190_195_groupi_g40006(csa_tree_add_190_195_groupi_n_8971 ,csa_tree_add_190_195_groupi_n_8970);
  not csa_tree_add_190_195_groupi_g40007(csa_tree_add_190_195_groupi_n_8968 ,csa_tree_add_190_195_groupi_n_8967);
  not csa_tree_add_190_195_groupi_g40008(csa_tree_add_190_195_groupi_n_8964 ,csa_tree_add_190_195_groupi_n_8963);
  not csa_tree_add_190_195_groupi_g40009(csa_tree_add_190_195_groupi_n_8961 ,csa_tree_add_190_195_groupi_n_8962);
  not csa_tree_add_190_195_groupi_g40010(csa_tree_add_190_195_groupi_n_8958 ,csa_tree_add_190_195_groupi_n_8959);
  not csa_tree_add_190_195_groupi_g40011(csa_tree_add_190_195_groupi_n_8957 ,csa_tree_add_190_195_groupi_n_8956);
  not csa_tree_add_190_195_groupi_g40012(csa_tree_add_190_195_groupi_n_8955 ,csa_tree_add_190_195_groupi_n_8954);
  not csa_tree_add_190_195_groupi_g40013(csa_tree_add_190_195_groupi_n_8952 ,csa_tree_add_190_195_groupi_n_8953);
  not csa_tree_add_190_195_groupi_g40014(csa_tree_add_190_195_groupi_n_8950 ,csa_tree_add_190_195_groupi_n_8951);
  not csa_tree_add_190_195_groupi_g40015(csa_tree_add_190_195_groupi_n_8949 ,csa_tree_add_190_195_groupi_n_8948);
  not csa_tree_add_190_195_groupi_g40016(csa_tree_add_190_195_groupi_n_8946 ,csa_tree_add_190_195_groupi_n_8947);
  nor csa_tree_add_190_195_groupi_g40017(csa_tree_add_190_195_groupi_n_8944 ,csa_tree_add_190_195_groupi_n_8483 ,csa_tree_add_190_195_groupi_n_8694);
  or csa_tree_add_190_195_groupi_g40018(csa_tree_add_190_195_groupi_n_8943 ,csa_tree_add_190_195_groupi_n_8517 ,csa_tree_add_190_195_groupi_n_8807);
  or csa_tree_add_190_195_groupi_g40019(csa_tree_add_190_195_groupi_n_8942 ,csa_tree_add_190_195_groupi_n_6768 ,csa_tree_add_190_195_groupi_n_8647);
  and csa_tree_add_190_195_groupi_g40020(csa_tree_add_190_195_groupi_n_8941 ,csa_tree_add_190_195_groupi_n_6768 ,csa_tree_add_190_195_groupi_n_8647);
  or csa_tree_add_190_195_groupi_g40021(csa_tree_add_190_195_groupi_n_8940 ,csa_tree_add_190_195_groupi_n_6449 ,csa_tree_add_190_195_groupi_n_8711);
  xor csa_tree_add_190_195_groupi_g40022(out1[0] ,csa_tree_add_190_195_groupi_n_5514 ,csa_tree_add_190_195_groupi_n_8268);
  and csa_tree_add_190_195_groupi_g40023(csa_tree_add_190_195_groupi_n_8938 ,csa_tree_add_190_195_groupi_n_8606 ,csa_tree_add_190_195_groupi_n_8852);
  or csa_tree_add_190_195_groupi_g40024(csa_tree_add_190_195_groupi_n_8937 ,csa_tree_add_190_195_groupi_n_7585 ,csa_tree_add_190_195_groupi_n_109);
  nor csa_tree_add_190_195_groupi_g40025(csa_tree_add_190_195_groupi_n_8936 ,csa_tree_add_190_195_groupi_n_7584 ,csa_tree_add_190_195_groupi_n_8634);
  nor csa_tree_add_190_195_groupi_g40026(csa_tree_add_190_195_groupi_n_8935 ,csa_tree_add_190_195_groupi_n_8532 ,csa_tree_add_190_195_groupi_n_8598);
  or csa_tree_add_190_195_groupi_g40027(csa_tree_add_190_195_groupi_n_8934 ,csa_tree_add_190_195_groupi_n_6919 ,csa_tree_add_190_195_groupi_n_8823);
  and csa_tree_add_190_195_groupi_g40028(csa_tree_add_190_195_groupi_n_8933 ,csa_tree_add_190_195_groupi_n_6919 ,csa_tree_add_190_195_groupi_n_8823);
  or csa_tree_add_190_195_groupi_g40029(csa_tree_add_190_195_groupi_n_8932 ,csa_tree_add_190_195_groupi_n_8650 ,csa_tree_add_190_195_groupi_n_8351);
  nor csa_tree_add_190_195_groupi_g40030(csa_tree_add_190_195_groupi_n_8931 ,csa_tree_add_190_195_groupi_n_8651 ,csa_tree_add_190_195_groupi_n_8352);
  or csa_tree_add_190_195_groupi_g40031(csa_tree_add_190_195_groupi_n_8930 ,csa_tree_add_190_195_groupi_n_8500 ,csa_tree_add_190_195_groupi_n_8657);
  or csa_tree_add_190_195_groupi_g40032(csa_tree_add_190_195_groupi_n_8929 ,csa_tree_add_190_195_groupi_n_8646 ,csa_tree_add_190_195_groupi_n_8836);
  nor csa_tree_add_190_195_groupi_g40033(csa_tree_add_190_195_groupi_n_8928 ,csa_tree_add_190_195_groupi_n_8645 ,csa_tree_add_190_195_groupi_n_8837);
  or csa_tree_add_190_195_groupi_g40034(csa_tree_add_190_195_groupi_n_8927 ,csa_tree_add_190_195_groupi_n_8614 ,csa_tree_add_190_195_groupi_n_8826);
  or csa_tree_add_190_195_groupi_g40035(csa_tree_add_190_195_groupi_n_8926 ,csa_tree_add_190_195_groupi_n_8048 ,csa_tree_add_190_195_groupi_n_8781);
  and csa_tree_add_190_195_groupi_g40036(csa_tree_add_190_195_groupi_n_8925 ,csa_tree_add_190_195_groupi_n_8614 ,csa_tree_add_190_195_groupi_n_8826);
  nor csa_tree_add_190_195_groupi_g40037(csa_tree_add_190_195_groupi_n_8924 ,csa_tree_add_190_195_groupi_n_7656 ,csa_tree_add_190_195_groupi_n_8590);
  or csa_tree_add_190_195_groupi_g40038(csa_tree_add_190_195_groupi_n_8923 ,csa_tree_add_190_195_groupi_n_7629 ,csa_tree_add_190_195_groupi_n_8611);
  and csa_tree_add_190_195_groupi_g40039(csa_tree_add_190_195_groupi_n_8922 ,csa_tree_add_190_195_groupi_n_7629 ,csa_tree_add_190_195_groupi_n_8611);
  nor csa_tree_add_190_195_groupi_g40040(csa_tree_add_190_195_groupi_n_8921 ,csa_tree_add_190_195_groupi_n_8501 ,csa_tree_add_190_195_groupi_n_8658);
  or csa_tree_add_190_195_groupi_g40041(csa_tree_add_190_195_groupi_n_8920 ,csa_tree_add_190_195_groupi_n_6304 ,csa_tree_add_190_195_groupi_n_8719);
  or csa_tree_add_190_195_groupi_g40042(csa_tree_add_190_195_groupi_n_8919 ,csa_tree_add_190_195_groupi_n_8341 ,csa_tree_add_190_195_groupi_n_8685);
  nor csa_tree_add_190_195_groupi_g40043(csa_tree_add_190_195_groupi_n_8918 ,csa_tree_add_190_195_groupi_n_8681 ,csa_tree_add_190_195_groupi_n_8679);
  or csa_tree_add_190_195_groupi_g40044(csa_tree_add_190_195_groupi_n_8917 ,csa_tree_add_190_195_groupi_n_8482 ,csa_tree_add_190_195_groupi_n_8695);
  and csa_tree_add_190_195_groupi_g40045(csa_tree_add_190_195_groupi_n_8916 ,csa_tree_add_190_195_groupi_n_6204 ,csa_tree_add_190_195_groupi_n_8721);
  nor csa_tree_add_190_195_groupi_g40046(csa_tree_add_190_195_groupi_n_8915 ,csa_tree_add_190_195_groupi_n_8342 ,csa_tree_add_190_195_groupi_n_8684);
  and csa_tree_add_190_195_groupi_g40047(csa_tree_add_190_195_groupi_n_8914 ,csa_tree_add_190_195_groupi_n_6131 ,csa_tree_add_190_195_groupi_n_72);
  or csa_tree_add_190_195_groupi_g40048(csa_tree_add_190_195_groupi_n_8913 ,csa_tree_add_190_195_groupi_n_8680 ,csa_tree_add_190_195_groupi_n_8678);
  xnor csa_tree_add_190_195_groupi_g40050(csa_tree_add_190_195_groupi_n_8912 ,csa_tree_add_190_195_groupi_n_5451 ,csa_tree_add_190_195_groupi_n_8535);
  xnor csa_tree_add_190_195_groupi_g40051(csa_tree_add_190_195_groupi_n_8911 ,csa_tree_add_190_195_groupi_n_6942 ,csa_tree_add_190_195_groupi_n_8325);
  xnor csa_tree_add_190_195_groupi_g40052(csa_tree_add_190_195_groupi_n_8910 ,csa_tree_add_190_195_groupi_n_7646 ,csa_tree_add_190_195_groupi_n_8386);
  xnor csa_tree_add_190_195_groupi_g40053(csa_tree_add_190_195_groupi_n_8909 ,csa_tree_add_190_195_groupi_n_6918 ,csa_tree_add_190_195_groupi_n_8496);
  xnor csa_tree_add_190_195_groupi_g40054(csa_tree_add_190_195_groupi_n_8908 ,csa_tree_add_190_195_groupi_n_4998 ,csa_tree_add_190_195_groupi_n_8512);
  xnor csa_tree_add_190_195_groupi_g40055(csa_tree_add_190_195_groupi_n_8907 ,csa_tree_add_190_195_groupi_n_8367 ,csa_tree_add_190_195_groupi_n_8223);
  xnor csa_tree_add_190_195_groupi_g40056(csa_tree_add_190_195_groupi_n_8906 ,csa_tree_add_190_195_groupi_n_6762 ,csa_tree_add_190_195_groupi_n_8517);
  xnor csa_tree_add_190_195_groupi_g40057(csa_tree_add_190_195_groupi_n_8905 ,csa_tree_add_190_195_groupi_n_8329 ,csa_tree_add_190_195_groupi_n_7321);
  xnor csa_tree_add_190_195_groupi_g40058(csa_tree_add_190_195_groupi_n_8904 ,csa_tree_add_190_195_groupi_n_5410 ,csa_tree_add_190_195_groupi_n_8538);
  xnor csa_tree_add_190_195_groupi_g40059(csa_tree_add_190_195_groupi_n_8903 ,csa_tree_add_190_195_groupi_n_4675 ,csa_tree_add_190_195_groupi_n_8348);
  xnor csa_tree_add_190_195_groupi_g40060(csa_tree_add_190_195_groupi_n_8902 ,csa_tree_add_190_195_groupi_n_8502 ,csa_tree_add_190_195_groupi_n_7858);
  xor csa_tree_add_190_195_groupi_g40061(csa_tree_add_190_195_groupi_n_8901 ,csa_tree_add_190_195_groupi_n_8320 ,csa_tree_add_190_195_groupi_n_7398);
  xnor csa_tree_add_190_195_groupi_g40062(csa_tree_add_190_195_groupi_n_8900 ,csa_tree_add_190_195_groupi_n_7576 ,csa_tree_add_190_195_groupi_n_8378);
  xnor csa_tree_add_190_195_groupi_g40063(csa_tree_add_190_195_groupi_n_8899 ,csa_tree_add_190_195_groupi_n_7125 ,csa_tree_add_190_195_groupi_n_8545);
  xnor csa_tree_add_190_195_groupi_g40064(csa_tree_add_190_195_groupi_n_8898 ,csa_tree_add_190_195_groupi_n_7093 ,csa_tree_add_190_195_groupi_n_8542);
  xnor csa_tree_add_190_195_groupi_g40066(csa_tree_add_190_195_groupi_n_8897 ,csa_tree_add_190_195_groupi_n_8233 ,csa_tree_add_190_195_groupi_n_8361);
  xnor csa_tree_add_190_195_groupi_g40067(csa_tree_add_190_195_groupi_n_8896 ,csa_tree_add_190_195_groupi_n_7314 ,csa_tree_add_190_195_groupi_n_8486);
  xnor csa_tree_add_190_195_groupi_g40068(csa_tree_add_190_195_groupi_n_8895 ,csa_tree_add_190_195_groupi_n_7303 ,csa_tree_add_190_195_groupi_n_8508);
  xnor csa_tree_add_190_195_groupi_g40069(csa_tree_add_190_195_groupi_n_8894 ,csa_tree_add_190_195_groupi_n_8490 ,csa_tree_add_190_195_groupi_n_8355);
  xnor csa_tree_add_190_195_groupi_g40071(csa_tree_add_190_195_groupi_n_8893 ,csa_tree_add_190_195_groupi_n_7829 ,csa_tree_add_190_195_groupi_n_8516);
  xnor csa_tree_add_190_195_groupi_g40072(csa_tree_add_190_195_groupi_n_8892 ,csa_tree_add_190_195_groupi_n_5536 ,csa_tree_add_190_195_groupi_n_8364);
  xnor csa_tree_add_190_195_groupi_g40073(csa_tree_add_190_195_groupi_n_8891 ,csa_tree_add_190_195_groupi_n_8195 ,csa_tree_add_190_195_groupi_n_8350);
  xnor csa_tree_add_190_195_groupi_g40074(csa_tree_add_190_195_groupi_n_8890 ,csa_tree_add_190_195_groupi_n_8029 ,csa_tree_add_190_195_groupi_n_8531);
  xnor csa_tree_add_190_195_groupi_g40075(csa_tree_add_190_195_groupi_n_8889 ,csa_tree_add_190_195_groupi_n_6962 ,csa_tree_add_190_195_groupi_n_8544);
  xnor csa_tree_add_190_195_groupi_g40076(csa_tree_add_190_195_groupi_n_8888 ,csa_tree_add_190_195_groupi_n_7142 ,csa_tree_add_190_195_groupi_n_8344);
  xnor csa_tree_add_190_195_groupi_g40077(csa_tree_add_190_195_groupi_n_8887 ,csa_tree_add_190_195_groupi_n_50 ,csa_tree_add_190_195_groupi_n_13);
  xnor csa_tree_add_190_195_groupi_g40078(csa_tree_add_190_195_groupi_n_8886 ,csa_tree_add_190_195_groupi_n_7835 ,csa_tree_add_190_195_groupi_n_8480);
  xnor csa_tree_add_190_195_groupi_g40080(csa_tree_add_190_195_groupi_n_8885 ,csa_tree_add_190_195_groupi_n_8002 ,csa_tree_add_190_195_groupi_n_8526);
  xnor csa_tree_add_190_195_groupi_g40081(csa_tree_add_190_195_groupi_n_8884 ,csa_tree_add_190_195_groupi_n_8522 ,csa_tree_add_190_195_groupi_n_7988);
  xnor csa_tree_add_190_195_groupi_g40082(csa_tree_add_190_195_groupi_n_8883 ,csa_tree_add_190_195_groupi_n_7103 ,csa_tree_add_190_195_groupi_n_8392);
  xnor csa_tree_add_190_195_groupi_g40083(csa_tree_add_190_195_groupi_n_8882 ,csa_tree_add_190_195_groupi_n_7538 ,csa_tree_add_190_195_groupi_n_8506);
  xnor csa_tree_add_190_195_groupi_g40084(csa_tree_add_190_195_groupi_n_8881 ,csa_tree_add_190_195_groupi_n_8536 ,csa_tree_add_190_195_groupi_n_7358);
  xnor csa_tree_add_190_195_groupi_g40085(csa_tree_add_190_195_groupi_n_8880 ,csa_tree_add_190_195_groupi_n_7078 ,csa_tree_add_190_195_groupi_n_8499);
  xnor csa_tree_add_190_195_groupi_g40086(csa_tree_add_190_195_groupi_n_8879 ,csa_tree_add_190_195_groupi_n_4699 ,csa_tree_add_190_195_groupi_n_8541);
  xnor csa_tree_add_190_195_groupi_g40087(csa_tree_add_190_195_groupi_n_8878 ,csa_tree_add_190_195_groupi_n_7642 ,csa_tree_add_190_195_groupi_n_8513);
  xnor csa_tree_add_190_195_groupi_g40088(csa_tree_add_190_195_groupi_n_9052 ,csa_tree_add_190_195_groupi_n_7651 ,csa_tree_add_190_195_groupi_n_8269);
  xnor csa_tree_add_190_195_groupi_g40089(csa_tree_add_190_195_groupi_n_9051 ,csa_tree_add_190_195_groupi_n_8394 ,csa_tree_add_190_195_groupi_n_6717);
  xnor csa_tree_add_190_195_groupi_g40090(csa_tree_add_190_195_groupi_n_9049 ,csa_tree_add_190_195_groupi_n_7346 ,csa_tree_add_190_195_groupi_n_8264);
  xnor csa_tree_add_190_195_groupi_g40091(csa_tree_add_190_195_groupi_n_9048 ,csa_tree_add_190_195_groupi_n_7119 ,csa_tree_add_190_195_groupi_n_8285);
  xnor csa_tree_add_190_195_groupi_g40093(csa_tree_add_190_195_groupi_n_9046 ,csa_tree_add_190_195_groupi_n_7862 ,csa_tree_add_190_195_groupi_n_8245);
  xnor csa_tree_add_190_195_groupi_g40094(csa_tree_add_190_195_groupi_n_9045 ,csa_tree_add_190_195_groupi_n_8236 ,csa_tree_add_190_195_groupi_n_1672);
  xnor csa_tree_add_190_195_groupi_g40095(csa_tree_add_190_195_groupi_n_9044 ,csa_tree_add_190_195_groupi_n_5287 ,csa_tree_add_190_195_groupi_n_8272);
  xnor csa_tree_add_190_195_groupi_g40096(csa_tree_add_190_195_groupi_n_9043 ,csa_tree_add_190_195_groupi_n_6953 ,csa_tree_add_190_195_groupi_n_8278);
  xnor csa_tree_add_190_195_groupi_g40097(csa_tree_add_190_195_groupi_n_9042 ,csa_tree_add_190_195_groupi_n_4911 ,csa_tree_add_190_195_groupi_n_8276);
  xnor csa_tree_add_190_195_groupi_g40098(csa_tree_add_190_195_groupi_n_9040 ,csa_tree_add_190_195_groupi_n_4957 ,csa_tree_add_190_195_groupi_n_108);
  xnor csa_tree_add_190_195_groupi_g40099(csa_tree_add_190_195_groupi_n_9039 ,csa_tree_add_190_195_groupi_n_5199 ,csa_tree_add_190_195_groupi_n_8279);
  xnor csa_tree_add_190_195_groupi_g40100(csa_tree_add_190_195_groupi_n_9038 ,csa_tree_add_190_195_groupi_n_8275 ,csa_tree_add_190_195_groupi_n_1002);
  and csa_tree_add_190_195_groupi_g40101(csa_tree_add_190_195_groupi_n_9037 ,csa_tree_add_190_195_groupi_n_6161 ,csa_tree_add_190_195_groupi_n_8589);
  xnor csa_tree_add_190_195_groupi_g40102(csa_tree_add_190_195_groupi_n_9036 ,csa_tree_add_190_195_groupi_n_8280 ,csa_tree_add_190_195_groupi_n_1738);
  or csa_tree_add_190_195_groupi_g40103(csa_tree_add_190_195_groupi_n_9035 ,csa_tree_add_190_195_groupi_n_8397 ,csa_tree_add_190_195_groupi_n_8605);
  xnor csa_tree_add_190_195_groupi_g40104(csa_tree_add_190_195_groupi_n_9033 ,csa_tree_add_190_195_groupi_n_8540 ,csa_tree_add_190_195_groupi_n_7923);
  xnor csa_tree_add_190_195_groupi_g40105(csa_tree_add_190_195_groupi_n_9031 ,csa_tree_add_190_195_groupi_n_5196 ,csa_tree_add_190_195_groupi_n_107);
  xnor csa_tree_add_190_195_groupi_g40106(csa_tree_add_190_195_groupi_n_9030 ,csa_tree_add_190_195_groupi_n_7827 ,csa_tree_add_190_195_groupi_n_8281);
  xnor csa_tree_add_190_195_groupi_g40107(csa_tree_add_190_195_groupi_n_9028 ,csa_tree_add_190_195_groupi_n_7494 ,csa_tree_add_190_195_groupi_n_8237);
  and csa_tree_add_190_195_groupi_g40108(csa_tree_add_190_195_groupi_n_9026 ,csa_tree_add_190_195_groupi_n_8302 ,csa_tree_add_190_195_groupi_n_8594);
  xnor csa_tree_add_190_195_groupi_g40109(csa_tree_add_190_195_groupi_n_9024 ,csa_tree_add_190_195_groupi_n_5452 ,csa_tree_add_190_195_groupi_n_8248);
  xnor csa_tree_add_190_195_groupi_g40110(csa_tree_add_190_195_groupi_n_9022 ,csa_tree_add_190_195_groupi_n_5894 ,csa_tree_add_190_195_groupi_n_8241);
  xnor csa_tree_add_190_195_groupi_g40111(csa_tree_add_190_195_groupi_n_9020 ,csa_tree_add_190_195_groupi_n_8528 ,csa_tree_add_190_195_groupi_n_6683);
  xnor csa_tree_add_190_195_groupi_g40112(csa_tree_add_190_195_groupi_n_9018 ,csa_tree_add_190_195_groupi_n_5049 ,csa_tree_add_190_195_groupi_n_8243);
  xnor csa_tree_add_190_195_groupi_g40113(csa_tree_add_190_195_groupi_n_9017 ,csa_tree_add_190_195_groupi_n_5258 ,csa_tree_add_190_195_groupi_n_8287);
  xnor csa_tree_add_190_195_groupi_g40114(csa_tree_add_190_195_groupi_n_9014 ,csa_tree_add_190_195_groupi_n_8382 ,csa_tree_add_190_195_groupi_n_6665);
  xnor csa_tree_add_190_195_groupi_g40115(csa_tree_add_190_195_groupi_n_9013 ,csa_tree_add_190_195_groupi_n_5508 ,csa_tree_add_190_195_groupi_n_8253);
  xnor csa_tree_add_190_195_groupi_g40116(csa_tree_add_190_195_groupi_n_9012 ,csa_tree_add_190_195_groupi_n_8228 ,csa_tree_add_190_195_groupi_n_8244);
  xnor csa_tree_add_190_195_groupi_g40117(csa_tree_add_190_195_groupi_n_9010 ,csa_tree_add_190_195_groupi_n_4962 ,csa_tree_add_190_195_groupi_n_8284);
  and csa_tree_add_190_195_groupi_g40118(csa_tree_add_190_195_groupi_n_9009 ,csa_tree_add_190_195_groupi_n_7955 ,csa_tree_add_190_195_groupi_n_8604);
  xnor csa_tree_add_190_195_groupi_g40119(csa_tree_add_190_195_groupi_n_9006 ,csa_tree_add_190_195_groupi_n_8530 ,csa_tree_add_190_195_groupi_n_7880);
  xnor csa_tree_add_190_195_groupi_g40120(csa_tree_add_190_195_groupi_n_9005 ,csa_tree_add_190_195_groupi_n_6912 ,csa_tree_add_190_195_groupi_n_8282);
  xnor csa_tree_add_190_195_groupi_g40121(csa_tree_add_190_195_groupi_n_9002 ,csa_tree_add_190_195_groupi_n_7536 ,csa_tree_add_190_195_groupi_n_8246);
  xnor csa_tree_add_190_195_groupi_g40122(csa_tree_add_190_195_groupi_n_9000 ,csa_tree_add_190_195_groupi_n_7110 ,csa_tree_add_190_195_groupi_n_8250);
  xnor csa_tree_add_190_195_groupi_g40123(csa_tree_add_190_195_groupi_n_8998 ,csa_tree_add_190_195_groupi_n_7608 ,csa_tree_add_190_195_groupi_n_8252);
  xnor csa_tree_add_190_195_groupi_g40124(csa_tree_add_190_195_groupi_n_8996 ,csa_tree_add_190_195_groupi_n_4734 ,csa_tree_add_190_195_groupi_n_8257);
  xnor csa_tree_add_190_195_groupi_g40126(csa_tree_add_190_195_groupi_n_8994 ,csa_tree_add_190_195_groupi_n_5935 ,csa_tree_add_190_195_groupi_n_8283);
  xnor csa_tree_add_190_195_groupi_g40127(csa_tree_add_190_195_groupi_n_8992 ,csa_tree_add_190_195_groupi_n_7076 ,csa_tree_add_190_195_groupi_n_8263);
  xnor csa_tree_add_190_195_groupi_g40128(csa_tree_add_190_195_groupi_n_8989 ,csa_tree_add_190_195_groupi_n_7518 ,csa_tree_add_190_195_groupi_n_8259);
  xnor csa_tree_add_190_195_groupi_g40130(csa_tree_add_190_195_groupi_n_8986 ,csa_tree_add_190_195_groupi_n_7823 ,csa_tree_add_190_195_groupi_n_8242);
  xnor csa_tree_add_190_195_groupi_g40131(csa_tree_add_190_195_groupi_n_8985 ,csa_tree_add_190_195_groupi_n_6257 ,csa_tree_add_190_195_groupi_n_8277);
  xnor csa_tree_add_190_195_groupi_g40132(csa_tree_add_190_195_groupi_n_8982 ,csa_tree_add_190_195_groupi_n_7506 ,csa_tree_add_190_195_groupi_n_8260);
  xnor csa_tree_add_190_195_groupi_g40133(csa_tree_add_190_195_groupi_n_8980 ,csa_tree_add_190_195_groupi_n_7594 ,csa_tree_add_190_195_groupi_n_8255);
  xnor csa_tree_add_190_195_groupi_g40134(csa_tree_add_190_195_groupi_n_8978 ,csa_tree_add_190_195_groupi_n_7068 ,csa_tree_add_190_195_groupi_n_8265);
  xnor csa_tree_add_190_195_groupi_g40135(csa_tree_add_190_195_groupi_n_8976 ,csa_tree_add_190_195_groupi_n_4903 ,csa_tree_add_190_195_groupi_n_8261);
  and csa_tree_add_190_195_groupi_g40136(csa_tree_add_190_195_groupi_n_8975 ,csa_tree_add_190_195_groupi_n_7812 ,csa_tree_add_190_195_groupi_n_8602);
  xnor csa_tree_add_190_195_groupi_g40137(csa_tree_add_190_195_groupi_n_8974 ,csa_tree_add_190_195_groupi_n_7547 ,csa_tree_add_190_195_groupi_n_8270);
  xnor csa_tree_add_190_195_groupi_g40138(csa_tree_add_190_195_groupi_n_8972 ,csa_tree_add_190_195_groupi_n_4632 ,csa_tree_add_190_195_groupi_n_8238);
  xnor csa_tree_add_190_195_groupi_g40139(csa_tree_add_190_195_groupi_n_8970 ,csa_tree_add_190_195_groupi_n_4763 ,csa_tree_add_190_195_groupi_n_8256);
  xnor csa_tree_add_190_195_groupi_g40140(csa_tree_add_190_195_groupi_n_8969 ,csa_tree_add_190_195_groupi_n_7571 ,csa_tree_add_190_195_groupi_n_8235);
  and csa_tree_add_190_195_groupi_g40141(csa_tree_add_190_195_groupi_n_8967 ,csa_tree_add_190_195_groupi_n_6470 ,csa_tree_add_190_195_groupi_n_8595);
  and csa_tree_add_190_195_groupi_g40142(csa_tree_add_190_195_groupi_n_8966 ,csa_tree_add_190_195_groupi_n_8464 ,csa_tree_add_190_195_groupi_n_8600);
  xnor csa_tree_add_190_195_groupi_g40143(csa_tree_add_190_195_groupi_n_8965 ,csa_tree_add_190_195_groupi_n_8384 ,csa_tree_add_190_195_groupi_n_34);
  xnor csa_tree_add_190_195_groupi_g40144(csa_tree_add_190_195_groupi_n_8963 ,csa_tree_add_190_195_groupi_n_8514 ,csa_tree_add_190_195_groupi_n_8239);
  xnor csa_tree_add_190_195_groupi_g40145(csa_tree_add_190_195_groupi_n_8962 ,csa_tree_add_190_195_groupi_n_6577 ,csa_tree_add_190_195_groupi_n_8286);
  xnor csa_tree_add_190_195_groupi_g40146(csa_tree_add_190_195_groupi_n_8960 ,csa_tree_add_190_195_groupi_n_8537 ,csa_tree_add_190_195_groupi_n_7022);
  xnor csa_tree_add_190_195_groupi_g40147(csa_tree_add_190_195_groupi_n_8959 ,csa_tree_add_190_195_groupi_n_8529 ,csa_tree_add_190_195_groupi_n_6615);
  xnor csa_tree_add_190_195_groupi_g40148(csa_tree_add_190_195_groupi_n_8956 ,csa_tree_add_190_195_groupi_n_8380 ,csa_tree_add_190_195_groupi_n_6647);
  xnor csa_tree_add_190_195_groupi_g40149(csa_tree_add_190_195_groupi_n_8954 ,csa_tree_add_190_195_groupi_n_5245 ,csa_tree_add_190_195_groupi_n_8254);
  xnor csa_tree_add_190_195_groupi_g40150(csa_tree_add_190_195_groupi_n_8953 ,csa_tree_add_190_195_groupi_n_7660 ,csa_tree_add_190_195_groupi_n_8247);
  xnor csa_tree_add_190_195_groupi_g40151(csa_tree_add_190_195_groupi_n_8951 ,csa_tree_add_190_195_groupi_n_5262 ,csa_tree_add_190_195_groupi_n_8273);
  and csa_tree_add_190_195_groupi_g40152(csa_tree_add_190_195_groupi_n_8948 ,csa_tree_add_190_195_groupi_n_7772 ,csa_tree_add_190_195_groupi_n_8588);
  xnor csa_tree_add_190_195_groupi_g40153(csa_tree_add_190_195_groupi_n_8947 ,csa_tree_add_190_195_groupi_n_8388 ,csa_tree_add_190_195_groupi_n_6643);
  xnor csa_tree_add_190_195_groupi_g40154(csa_tree_add_190_195_groupi_n_8945 ,csa_tree_add_190_195_groupi_n_7843 ,csa_tree_add_190_195_groupi_n_8240);
  not csa_tree_add_190_195_groupi_g40156(csa_tree_add_190_195_groupi_n_8860 ,csa_tree_add_190_195_groupi_n_8859);
  not csa_tree_add_190_195_groupi_g40158(csa_tree_add_190_195_groupi_n_8854 ,csa_tree_add_190_195_groupi_n_8853);
  not csa_tree_add_190_195_groupi_g40159(csa_tree_add_190_195_groupi_n_8849 ,csa_tree_add_190_195_groupi_n_8848);
  not csa_tree_add_190_195_groupi_g40160(csa_tree_add_190_195_groupi_n_8847 ,csa_tree_add_190_195_groupi_n_8846);
  not csa_tree_add_190_195_groupi_g40161(csa_tree_add_190_195_groupi_n_8840 ,csa_tree_add_190_195_groupi_n_8839);
  not csa_tree_add_190_195_groupi_g40162(csa_tree_add_190_195_groupi_n_8836 ,csa_tree_add_190_195_groupi_n_8837);
  not csa_tree_add_190_195_groupi_g40163(csa_tree_add_190_195_groupi_n_8834 ,csa_tree_add_190_195_groupi_n_8833);
  not csa_tree_add_190_195_groupi_g40164(csa_tree_add_190_195_groupi_n_8831 ,csa_tree_add_190_195_groupi_n_8832);
  not csa_tree_add_190_195_groupi_g40165(csa_tree_add_190_195_groupi_n_8830 ,csa_tree_add_190_195_groupi_n_8829);
  not csa_tree_add_190_195_groupi_g40166(csa_tree_add_190_195_groupi_n_8828 ,csa_tree_add_190_195_groupi_n_8827);
  not csa_tree_add_190_195_groupi_g40167(csa_tree_add_190_195_groupi_n_8825 ,csa_tree_add_190_195_groupi_n_8824);
  not csa_tree_add_190_195_groupi_g40168(csa_tree_add_190_195_groupi_n_8821 ,csa_tree_add_190_195_groupi_n_8822);
  not csa_tree_add_190_195_groupi_g40169(csa_tree_add_190_195_groupi_n_8819 ,csa_tree_add_190_195_groupi_n_8820);
  not csa_tree_add_190_195_groupi_g40170(csa_tree_add_190_195_groupi_n_8817 ,csa_tree_add_190_195_groupi_n_8816);
  not csa_tree_add_190_195_groupi_g40171(csa_tree_add_190_195_groupi_n_8815 ,csa_tree_add_190_195_groupi_n_8814);
  not csa_tree_add_190_195_groupi_g40172(csa_tree_add_190_195_groupi_n_8813 ,csa_tree_add_190_195_groupi_n_8812);
  and csa_tree_add_190_195_groupi_g40173(csa_tree_add_190_195_groupi_n_8811 ,csa_tree_add_190_195_groupi_n_8021 ,csa_tree_add_190_195_groupi_n_8481);
  nor csa_tree_add_190_195_groupi_g40174(csa_tree_add_190_195_groupi_n_8810 ,csa_tree_add_190_195_groupi_n_5535 ,csa_tree_add_190_195_groupi_n_8364);
  or csa_tree_add_190_195_groupi_g40175(csa_tree_add_190_195_groupi_n_8809 ,csa_tree_add_190_195_groupi_n_5536 ,csa_tree_add_190_195_groupi_n_8363);
  or csa_tree_add_190_195_groupi_g40176(csa_tree_add_190_195_groupi_n_8808 ,csa_tree_add_190_195_groupi_n_46 ,csa_tree_add_190_195_groupi_n_8304);
  nor csa_tree_add_190_195_groupi_g40177(csa_tree_add_190_195_groupi_n_8807 ,csa_tree_add_190_195_groupi_n_6762 ,csa_tree_add_190_195_groupi_n_8494);
  and csa_tree_add_190_195_groupi_g40178(csa_tree_add_190_195_groupi_n_8806 ,csa_tree_add_190_195_groupi_n_8175 ,csa_tree_add_190_195_groupi_n_8378);
  and csa_tree_add_190_195_groupi_g40179(csa_tree_add_190_195_groupi_n_8805 ,csa_tree_add_190_195_groupi_n_7194 ,csa_tree_add_190_195_groupi_n_8472);
  or csa_tree_add_190_195_groupi_g40180(csa_tree_add_190_195_groupi_n_8804 ,csa_tree_add_190_195_groupi_n_6761 ,csa_tree_add_190_195_groupi_n_8493);
  or csa_tree_add_190_195_groupi_g40181(csa_tree_add_190_195_groupi_n_8803 ,csa_tree_add_190_195_groupi_n_7368 ,csa_tree_add_190_195_groupi_n_8371);
  or csa_tree_add_190_195_groupi_g40182(csa_tree_add_190_195_groupi_n_8802 ,csa_tree_add_190_195_groupi_n_8486 ,csa_tree_add_190_195_groupi_n_7314);
  nor csa_tree_add_190_195_groupi_g40183(csa_tree_add_190_195_groupi_n_8801 ,csa_tree_add_190_195_groupi_n_7367 ,csa_tree_add_190_195_groupi_n_8372);
  and csa_tree_add_190_195_groupi_g40184(csa_tree_add_190_195_groupi_n_8800 ,csa_tree_add_190_195_groupi_n_7295 ,csa_tree_add_190_195_groupi_n_8535);
  or csa_tree_add_190_195_groupi_g40185(csa_tree_add_190_195_groupi_n_8799 ,csa_tree_add_190_195_groupi_n_8466 ,csa_tree_add_190_195_groupi_n_8214);
  or csa_tree_add_190_195_groupi_g40186(csa_tree_add_190_195_groupi_n_8798 ,csa_tree_add_190_195_groupi_n_8395 ,csa_tree_add_190_195_groupi_n_8297);
  and csa_tree_add_190_195_groupi_g40187(csa_tree_add_190_195_groupi_n_8797 ,csa_tree_add_190_195_groupi_n_8486 ,csa_tree_add_190_195_groupi_n_7314);
  nor csa_tree_add_190_195_groupi_g40188(csa_tree_add_190_195_groupi_n_8796 ,csa_tree_add_190_195_groupi_n_6917 ,csa_tree_add_190_195_groupi_n_8496);
  or csa_tree_add_190_195_groupi_g40189(csa_tree_add_190_195_groupi_n_8795 ,csa_tree_add_190_195_groupi_n_6918 ,csa_tree_add_190_195_groupi_n_8495);
  nor csa_tree_add_190_195_groupi_g40190(csa_tree_add_190_195_groupi_n_8794 ,csa_tree_add_190_195_groupi_n_5925 ,csa_tree_add_190_195_groupi_n_8338);
  or csa_tree_add_190_195_groupi_g40191(csa_tree_add_190_195_groupi_n_8793 ,csa_tree_add_190_195_groupi_n_5926 ,csa_tree_add_190_195_groupi_n_8337);
  and csa_tree_add_190_195_groupi_g40192(csa_tree_add_190_195_groupi_n_8792 ,csa_tree_add_190_195_groupi_n_7078 ,csa_tree_add_190_195_groupi_n_8499);
  nor csa_tree_add_190_195_groupi_g40193(csa_tree_add_190_195_groupi_n_8791 ,csa_tree_add_190_195_groupi_n_8195 ,csa_tree_add_190_195_groupi_n_8349);
  or csa_tree_add_190_195_groupi_g40194(csa_tree_add_190_195_groupi_n_8790 ,csa_tree_add_190_195_groupi_n_8194 ,csa_tree_add_190_195_groupi_n_8350);
  or csa_tree_add_190_195_groupi_g40195(csa_tree_add_190_195_groupi_n_8789 ,csa_tree_add_190_195_groupi_n_8137 ,csa_tree_add_190_195_groupi_n_8379);
  or csa_tree_add_190_195_groupi_g40196(csa_tree_add_190_195_groupi_n_8788 ,csa_tree_add_190_195_groupi_n_7078 ,csa_tree_add_190_195_groupi_n_8499);
  nor csa_tree_add_190_195_groupi_g40197(csa_tree_add_190_195_groupi_n_8787 ,csa_tree_add_190_195_groupi_n_7995 ,csa_tree_add_190_195_groupi_n_8361);
  or csa_tree_add_190_195_groupi_g40198(csa_tree_add_190_195_groupi_n_8786 ,csa_tree_add_190_195_groupi_n_7994 ,csa_tree_add_190_195_groupi_n_8360);
  and csa_tree_add_190_195_groupi_g40199(csa_tree_add_190_195_groupi_n_8785 ,csa_tree_add_190_195_groupi_n_8392 ,csa_tree_add_190_195_groupi_n_8288);
  nor csa_tree_add_190_195_groupi_g40200(csa_tree_add_190_195_groupi_n_8784 ,csa_tree_add_190_195_groupi_n_7415 ,csa_tree_add_190_195_groupi_n_8307);
  and csa_tree_add_190_195_groupi_g40201(csa_tree_add_190_195_groupi_n_8783 ,csa_tree_add_190_195_groupi_n_6873 ,csa_tree_add_190_195_groupi_n_8537);
  or csa_tree_add_190_195_groupi_g40202(csa_tree_add_190_195_groupi_n_8782 ,csa_tree_add_190_195_groupi_n_7861 ,csa_tree_add_190_195_groupi_n_8471);
  nor csa_tree_add_190_195_groupi_g40203(csa_tree_add_190_195_groupi_n_8781 ,csa_tree_add_190_195_groupi_n_6942 ,csa_tree_add_190_195_groupi_n_8324);
  or csa_tree_add_190_195_groupi_g40204(csa_tree_add_190_195_groupi_n_8780 ,csa_tree_add_190_195_groupi_n_8386 ,csa_tree_add_190_195_groupi_n_8082);
  nor csa_tree_add_190_195_groupi_g40205(csa_tree_add_190_195_groupi_n_8779 ,csa_tree_add_190_195_groupi_n_8443 ,csa_tree_add_190_195_groupi_n_8508);
  or csa_tree_add_190_195_groupi_g40206(csa_tree_add_190_195_groupi_n_8778 ,csa_tree_add_190_195_groupi_n_5366 ,csa_tree_add_190_195_groupi_n_8362);
  nor csa_tree_add_190_195_groupi_g40207(csa_tree_add_190_195_groupi_n_8777 ,csa_tree_add_190_195_groupi_n_7829 ,csa_tree_add_190_195_groupi_n_8318);
  or csa_tree_add_190_195_groupi_g40208(csa_tree_add_190_195_groupi_n_8776 ,csa_tree_add_190_195_groupi_n_5771 ,csa_tree_add_190_195_groupi_n_8512);
  or csa_tree_add_190_195_groupi_g40209(csa_tree_add_190_195_groupi_n_8775 ,csa_tree_add_190_195_groupi_n_7828 ,csa_tree_add_190_195_groupi_n_8319);
  and csa_tree_add_190_195_groupi_g40210(csa_tree_add_190_195_groupi_n_8774 ,csa_tree_add_190_195_groupi_n_5786 ,csa_tree_add_190_195_groupi_n_8541);
  nor csa_tree_add_190_195_groupi_g40211(csa_tree_add_190_195_groupi_n_8773 ,csa_tree_add_190_195_groupi_n_7996 ,csa_tree_add_190_195_groupi_n_8354);
  or csa_tree_add_190_195_groupi_g40212(csa_tree_add_190_195_groupi_n_8772 ,csa_tree_add_190_195_groupi_n_8393 ,csa_tree_add_190_195_groupi_n_8469);
  and csa_tree_add_190_195_groupi_g40213(csa_tree_add_190_195_groupi_n_8771 ,csa_tree_add_190_195_groupi_n_7096 ,csa_tree_add_190_195_groupi_n_8367);
  or csa_tree_add_190_195_groupi_g40214(csa_tree_add_190_195_groupi_n_8770 ,csa_tree_add_190_195_groupi_n_7096 ,csa_tree_add_190_195_groupi_n_8367);
  nor csa_tree_add_190_195_groupi_g40215(csa_tree_add_190_195_groupi_n_8769 ,csa_tree_add_190_195_groupi_n_6093 ,csa_tree_add_190_195_groupi_n_8529);
  and csa_tree_add_190_195_groupi_g40216(csa_tree_add_190_195_groupi_n_8768 ,csa_tree_add_190_195_groupi_n_7863 ,csa_tree_add_190_195_groupi_n_8295);
  or csa_tree_add_190_195_groupi_g40217(csa_tree_add_190_195_groupi_n_8767 ,csa_tree_add_190_195_groupi_n_6357 ,csa_tree_add_190_195_groupi_n_8394);
  and csa_tree_add_190_195_groupi_g40218(csa_tree_add_190_195_groupi_n_8766 ,csa_tree_add_190_195_groupi_n_8491 ,csa_tree_add_190_195_groupi_n_8355);
  nor csa_tree_add_190_195_groupi_g40219(csa_tree_add_190_195_groupi_n_8765 ,csa_tree_add_190_195_groupi_n_8460 ,csa_tree_add_190_195_groupi_n_7848);
  or csa_tree_add_190_195_groupi_g40220(csa_tree_add_190_195_groupi_n_8764 ,csa_tree_add_190_195_groupi_n_6344 ,csa_tree_add_190_195_groupi_n_8528);
  or csa_tree_add_190_195_groupi_g40221(csa_tree_add_190_195_groupi_n_8763 ,csa_tree_add_190_195_groupi_n_8422 ,csa_tree_add_190_195_groupi_n_8527);
  or csa_tree_add_190_195_groupi_g40222(csa_tree_add_190_195_groupi_n_8762 ,csa_tree_add_190_195_groupi_n_6100 ,csa_tree_add_190_195_groupi_n_8382);
  or csa_tree_add_190_195_groupi_g40223(csa_tree_add_190_195_groupi_n_8761 ,csa_tree_add_190_195_groupi_n_7857 ,csa_tree_add_190_195_groupi_n_8449);
  nor csa_tree_add_190_195_groupi_g40224(csa_tree_add_190_195_groupi_n_8760 ,csa_tree_add_190_195_groupi_n_7539 ,csa_tree_add_190_195_groupi_n_8506);
  and csa_tree_add_190_195_groupi_g40225(csa_tree_add_190_195_groupi_n_8759 ,csa_tree_add_190_195_groupi_n_5200 ,csa_tree_add_190_195_groupi_n_8502);
  or csa_tree_add_190_195_groupi_g40226(csa_tree_add_190_195_groupi_n_8758 ,csa_tree_add_190_195_groupi_n_6941 ,csa_tree_add_190_195_groupi_n_8325);
  nor csa_tree_add_190_195_groupi_g40227(csa_tree_add_190_195_groupi_n_8757 ,csa_tree_add_190_195_groupi_n_3170 ,csa_tree_add_190_195_groupi_n_8384);
  or csa_tree_add_190_195_groupi_g40228(csa_tree_add_190_195_groupi_n_8756 ,csa_tree_add_190_195_groupi_n_8530 ,csa_tree_add_190_195_groupi_n_7736);
  and csa_tree_add_190_195_groupi_g40229(csa_tree_add_190_195_groupi_n_8755 ,csa_tree_add_190_195_groupi_n_8531 ,csa_tree_add_190_195_groupi_n_8294);
  nor csa_tree_add_190_195_groupi_g40230(csa_tree_add_190_195_groupi_n_8754 ,csa_tree_add_190_195_groupi_n_6964 ,csa_tree_add_190_195_groupi_n_8492);
  or csa_tree_add_190_195_groupi_g40231(csa_tree_add_190_195_groupi_n_8753 ,csa_tree_add_190_195_groupi_n_5200 ,csa_tree_add_190_195_groupi_n_8502);
  or csa_tree_add_190_195_groupi_g40232(csa_tree_add_190_195_groupi_n_8752 ,csa_tree_add_190_195_groupi_n_6258 ,csa_tree_add_190_195_groupi_n_8357);
  and csa_tree_add_190_195_groupi_g40233(csa_tree_add_190_195_groupi_n_8751 ,csa_tree_add_190_195_groupi_n_7539 ,csa_tree_add_190_195_groupi_n_8506);
  or csa_tree_add_190_195_groupi_g40234(csa_tree_add_190_195_groupi_n_8750 ,csa_tree_add_190_195_groupi_n_8016 ,csa_tree_add_190_195_groupi_n_8323);
  nor csa_tree_add_190_195_groupi_g40235(csa_tree_add_190_195_groupi_n_8749 ,csa_tree_add_190_195_groupi_n_6259 ,csa_tree_add_190_195_groupi_n_8356);
  nor csa_tree_add_190_195_groupi_g40236(csa_tree_add_190_195_groupi_n_8748 ,csa_tree_add_190_195_groupi_n_8017 ,csa_tree_add_190_195_groupi_n_8322);
  or csa_tree_add_190_195_groupi_g40237(csa_tree_add_190_195_groupi_n_8747 ,csa_tree_add_190_195_groupi_n_7974 ,csa_tree_add_190_195_groupi_n_8546);
  or csa_tree_add_190_195_groupi_g40238(csa_tree_add_190_195_groupi_n_8746 ,csa_tree_add_190_195_groupi_n_4674 ,csa_tree_add_190_195_groupi_n_8348);
  or csa_tree_add_190_195_groupi_g40239(csa_tree_add_190_195_groupi_n_8745 ,csa_tree_add_190_195_groupi_n_7141 ,csa_tree_add_190_195_groupi_n_8344);
  nor csa_tree_add_190_195_groupi_g40240(csa_tree_add_190_195_groupi_n_8744 ,csa_tree_add_190_195_groupi_n_7142 ,csa_tree_add_190_195_groupi_n_8343);
  and csa_tree_add_190_195_groupi_g40241(csa_tree_add_190_195_groupi_n_8743 ,csa_tree_add_190_195_groupi_n_5366 ,csa_tree_add_190_195_groupi_n_8362);
  nor csa_tree_add_190_195_groupi_g40242(csa_tree_add_190_195_groupi_n_8742 ,csa_tree_add_190_195_groupi_n_8491 ,csa_tree_add_190_195_groupi_n_8355);
  nor csa_tree_add_190_195_groupi_g40243(csa_tree_add_190_195_groupi_n_8741 ,csa_tree_add_190_195_groupi_n_8021 ,csa_tree_add_190_195_groupi_n_8481);
  or csa_tree_add_190_195_groupi_g40244(csa_tree_add_190_195_groupi_n_8740 ,csa_tree_add_190_195_groupi_n_8045 ,csa_tree_add_190_195_groupi_n_8453);
  or csa_tree_add_190_195_groupi_g40245(csa_tree_add_190_195_groupi_n_8739 ,csa_tree_add_190_195_groupi_n_7510 ,csa_tree_add_190_195_groupi_n_8345);
  or csa_tree_add_190_195_groupi_g40246(csa_tree_add_190_195_groupi_n_8738 ,csa_tree_add_190_195_groupi_n_7997 ,csa_tree_add_190_195_groupi_n_8353);
  nor csa_tree_add_190_195_groupi_g40247(csa_tree_add_190_195_groupi_n_8737 ,csa_tree_add_190_195_groupi_n_7366 ,csa_tree_add_190_195_groupi_n_8327);
  nor csa_tree_add_190_195_groupi_g40248(csa_tree_add_190_195_groupi_n_8736 ,csa_tree_add_190_195_groupi_n_7509 ,csa_tree_add_190_195_groupi_n_8346);
  or csa_tree_add_190_195_groupi_g40249(csa_tree_add_190_195_groupi_n_8735 ,csa_tree_add_190_195_groupi_n_8208 ,csa_tree_add_190_195_groupi_n_8402);
  or csa_tree_add_190_195_groupi_g40250(csa_tree_add_190_195_groupi_n_8734 ,csa_tree_add_190_195_groupi_n_7365 ,csa_tree_add_190_195_groupi_n_8326);
  and csa_tree_add_190_195_groupi_g40251(csa_tree_add_190_195_groupi_n_8733 ,csa_tree_add_190_195_groupi_n_7245 ,csa_tree_add_190_195_groupi_n_8544);
  or csa_tree_add_190_195_groupi_g40252(csa_tree_add_190_195_groupi_n_8732 ,csa_tree_add_190_195_groupi_n_7835 ,csa_tree_add_190_195_groupi_n_8479);
  nor csa_tree_add_190_195_groupi_g40253(csa_tree_add_190_195_groupi_n_8731 ,csa_tree_add_190_195_groupi_n_7834 ,csa_tree_add_190_195_groupi_n_8480);
  and csa_tree_add_190_195_groupi_g40254(csa_tree_add_190_195_groupi_n_8730 ,csa_tree_add_190_195_groupi_n_6243 ,csa_tree_add_190_195_groupi_n_8388);
  nor csa_tree_add_190_195_groupi_g40255(csa_tree_add_190_195_groupi_n_8729 ,csa_tree_add_190_195_groupi_n_8218 ,csa_tree_add_190_195_groupi_n_8403);
  and csa_tree_add_190_195_groupi_g40256(csa_tree_add_190_195_groupi_n_8728 ,csa_tree_add_190_195_groupi_n_7517 ,csa_tree_add_190_195_groupi_n_8320);
  or csa_tree_add_190_195_groupi_g40257(csa_tree_add_190_195_groupi_n_8727 ,csa_tree_add_190_195_groupi_n_7517 ,csa_tree_add_190_195_groupi_n_8320);
  and csa_tree_add_190_195_groupi_g40258(csa_tree_add_190_195_groupi_n_8726 ,csa_tree_add_190_195_groupi_n_8159 ,csa_tree_add_190_195_groupi_n_8513);
  and csa_tree_add_190_195_groupi_g40259(csa_tree_add_190_195_groupi_n_8725 ,csa_tree_add_190_195_groupi_n_6964 ,csa_tree_add_190_195_groupi_n_8492);
  nor csa_tree_add_190_195_groupi_g40260(csa_tree_add_190_195_groupi_n_8724 ,csa_tree_add_190_195_groupi_n_4675 ,csa_tree_add_190_195_groupi_n_8347);
  and csa_tree_add_190_195_groupi_g40261(csa_tree_add_190_195_groupi_n_8877 ,csa_tree_add_190_195_groupi_n_8111 ,csa_tree_add_190_195_groupi_n_8423);
  and csa_tree_add_190_195_groupi_g40262(csa_tree_add_190_195_groupi_n_8876 ,csa_tree_add_190_195_groupi_n_7815 ,csa_tree_add_190_195_groupi_n_8475);
  or csa_tree_add_190_195_groupi_g40263(csa_tree_add_190_195_groupi_n_8875 ,csa_tree_add_190_195_groupi_n_8173 ,csa_tree_add_190_195_groupi_n_8470);
  and csa_tree_add_190_195_groupi_g40264(csa_tree_add_190_195_groupi_n_8874 ,csa_tree_add_190_195_groupi_n_6208 ,csa_tree_add_190_195_groupi_n_8416);
  or csa_tree_add_190_195_groupi_g40265(csa_tree_add_190_195_groupi_n_8873 ,csa_tree_add_190_195_groupi_n_8139 ,csa_tree_add_190_195_groupi_n_8408);
  and csa_tree_add_190_195_groupi_g40266(csa_tree_add_190_195_groupi_n_8872 ,csa_tree_add_190_195_groupi_n_8160 ,csa_tree_add_190_195_groupi_n_8429);
  and csa_tree_add_190_195_groupi_g40267(csa_tree_add_190_195_groupi_n_8871 ,csa_tree_add_190_195_groupi_n_6516 ,csa_tree_add_190_195_groupi_n_8465);
  and csa_tree_add_190_195_groupi_g40268(csa_tree_add_190_195_groupi_n_8870 ,csa_tree_add_190_195_groupi_n_8068 ,csa_tree_add_190_195_groupi_n_8404);
  and csa_tree_add_190_195_groupi_g40269(csa_tree_add_190_195_groupi_n_8869 ,csa_tree_add_190_195_groupi_n_5673 ,csa_tree_add_190_195_groupi_n_8435);
  and csa_tree_add_190_195_groupi_g40270(csa_tree_add_190_195_groupi_n_8868 ,csa_tree_add_190_195_groupi_n_8158 ,csa_tree_add_190_195_groupi_n_8310);
  and csa_tree_add_190_195_groupi_g40271(csa_tree_add_190_195_groupi_n_8867 ,csa_tree_add_190_195_groupi_n_7796 ,csa_tree_add_190_195_groupi_n_8426);
  and csa_tree_add_190_195_groupi_g40272(csa_tree_add_190_195_groupi_n_8866 ,csa_tree_add_190_195_groupi_n_7724 ,csa_tree_add_190_195_groupi_n_8399);
  and csa_tree_add_190_195_groupi_g40273(csa_tree_add_190_195_groupi_n_8865 ,csa_tree_add_190_195_groupi_n_7254 ,csa_tree_add_190_195_groupi_n_8401);
  and csa_tree_add_190_195_groupi_g40274(csa_tree_add_190_195_groupi_n_8864 ,csa_tree_add_190_195_groupi_n_6138 ,csa_tree_add_190_195_groupi_n_8441);
  and csa_tree_add_190_195_groupi_g40275(csa_tree_add_190_195_groupi_n_8863 ,csa_tree_add_190_195_groupi_n_6136 ,csa_tree_add_190_195_groupi_n_8439);
  and csa_tree_add_190_195_groupi_g40276(csa_tree_add_190_195_groupi_n_8862 ,csa_tree_add_190_195_groupi_n_6129 ,csa_tree_add_190_195_groupi_n_8442);
  or csa_tree_add_190_195_groupi_g40277(csa_tree_add_190_195_groupi_n_8861 ,csa_tree_add_190_195_groupi_n_6124 ,csa_tree_add_190_195_groupi_n_8432);
  or csa_tree_add_190_195_groupi_g40278(csa_tree_add_190_195_groupi_n_8859 ,csa_tree_add_190_195_groupi_n_8087 ,csa_tree_add_190_195_groupi_n_8407);
  and csa_tree_add_190_195_groupi_g40279(csa_tree_add_190_195_groupi_n_8858 ,csa_tree_add_190_195_groupi_n_8089 ,csa_tree_add_190_195_groupi_n_8478);
  and csa_tree_add_190_195_groupi_g40280(csa_tree_add_190_195_groupi_n_8857 ,csa_tree_add_190_195_groupi_n_8075 ,csa_tree_add_190_195_groupi_n_8411);
  or csa_tree_add_190_195_groupi_g40281(csa_tree_add_190_195_groupi_n_8856 ,csa_tree_add_190_195_groupi_n_8091 ,csa_tree_add_190_195_groupi_n_8409);
  and csa_tree_add_190_195_groupi_g40282(csa_tree_add_190_195_groupi_n_8855 ,csa_tree_add_190_195_groupi_n_8149 ,csa_tree_add_190_195_groupi_n_8452);
  or csa_tree_add_190_195_groupi_g40283(csa_tree_add_190_195_groupi_n_8853 ,csa_tree_add_190_195_groupi_n_7945 ,csa_tree_add_190_195_groupi_n_8417);
  or csa_tree_add_190_195_groupi_g40284(csa_tree_add_190_195_groupi_n_8852 ,csa_tree_add_190_195_groupi_n_8106 ,csa_tree_add_190_195_groupi_n_8419);
  or csa_tree_add_190_195_groupi_g40285(csa_tree_add_190_195_groupi_n_8851 ,csa_tree_add_190_195_groupi_n_7978 ,csa_tree_add_190_195_groupi_n_8424);
  and csa_tree_add_190_195_groupi_g40286(csa_tree_add_190_195_groupi_n_8850 ,csa_tree_add_190_195_groupi_n_7789 ,csa_tree_add_190_195_groupi_n_8451);
  or csa_tree_add_190_195_groupi_g40287(csa_tree_add_190_195_groupi_n_8848 ,csa_tree_add_190_195_groupi_n_7966 ,csa_tree_add_190_195_groupi_n_8463);
  or csa_tree_add_190_195_groupi_g40288(csa_tree_add_190_195_groupi_n_8846 ,csa_tree_add_190_195_groupi_n_8079 ,csa_tree_add_190_195_groupi_n_8300);
  and csa_tree_add_190_195_groupi_g40289(csa_tree_add_190_195_groupi_n_8845 ,csa_tree_add_190_195_groupi_n_6394 ,csa_tree_add_190_195_groupi_n_8433);
  and csa_tree_add_190_195_groupi_g40290(csa_tree_add_190_195_groupi_n_8844 ,csa_tree_add_190_195_groupi_n_5755 ,csa_tree_add_190_195_groupi_n_8428);
  and csa_tree_add_190_195_groupi_g40291(csa_tree_add_190_195_groupi_n_8843 ,csa_tree_add_190_195_groupi_n_6465 ,csa_tree_add_190_195_groupi_n_8450);
  and csa_tree_add_190_195_groupi_g40292(csa_tree_add_190_195_groupi_n_8842 ,csa_tree_add_190_195_groupi_n_8128 ,csa_tree_add_190_195_groupi_n_8398);
  and csa_tree_add_190_195_groupi_g40293(csa_tree_add_190_195_groupi_n_8841 ,csa_tree_add_190_195_groupi_n_6434 ,csa_tree_add_190_195_groupi_n_8440);
  or csa_tree_add_190_195_groupi_g40294(csa_tree_add_190_195_groupi_n_8839 ,csa_tree_add_190_195_groupi_n_8135 ,csa_tree_add_190_195_groupi_n_8437);
  or csa_tree_add_190_195_groupi_g40295(csa_tree_add_190_195_groupi_n_8838 ,csa_tree_add_190_195_groupi_n_6448 ,csa_tree_add_190_195_groupi_n_8444);
  or csa_tree_add_190_195_groupi_g40296(csa_tree_add_190_195_groupi_n_8837 ,csa_tree_add_190_195_groupi_n_8134 ,csa_tree_add_190_195_groupi_n_8438);
  and csa_tree_add_190_195_groupi_g40297(csa_tree_add_190_195_groupi_n_8835 ,csa_tree_add_190_195_groupi_n_8125 ,csa_tree_add_190_195_groupi_n_8434);
  and csa_tree_add_190_195_groupi_g40298(csa_tree_add_190_195_groupi_n_8833 ,csa_tree_add_190_195_groupi_n_7766 ,csa_tree_add_190_195_groupi_n_8431);
  or csa_tree_add_190_195_groupi_g40299(csa_tree_add_190_195_groupi_n_8832 ,csa_tree_add_190_195_groupi_n_6191 ,csa_tree_add_190_195_groupi_n_8413);
  and csa_tree_add_190_195_groupi_g40300(csa_tree_add_190_195_groupi_n_8829 ,csa_tree_add_190_195_groupi_n_8144 ,csa_tree_add_190_195_groupi_n_8421);
  and csa_tree_add_190_195_groupi_g40301(csa_tree_add_190_195_groupi_n_8827 ,csa_tree_add_190_195_groupi_n_8157 ,csa_tree_add_190_195_groupi_n_8455);
  and csa_tree_add_190_195_groupi_g40302(csa_tree_add_190_195_groupi_n_8826 ,csa_tree_add_190_195_groupi_n_8099 ,csa_tree_add_190_195_groupi_n_8415);
  or csa_tree_add_190_195_groupi_g40303(csa_tree_add_190_195_groupi_n_8824 ,csa_tree_add_190_195_groupi_n_5715 ,csa_tree_add_190_195_groupi_n_8405);
  and csa_tree_add_190_195_groupi_g40304(csa_tree_add_190_195_groupi_n_8823 ,csa_tree_add_190_195_groupi_n_6880 ,csa_tree_add_190_195_groupi_n_8311);
  or csa_tree_add_190_195_groupi_g40305(csa_tree_add_190_195_groupi_n_8822 ,csa_tree_add_190_195_groupi_n_5735 ,csa_tree_add_190_195_groupi_n_8420);
  or csa_tree_add_190_195_groupi_g40306(csa_tree_add_190_195_groupi_n_8820 ,csa_tree_add_190_195_groupi_n_6312 ,csa_tree_add_190_195_groupi_n_8309);
  or csa_tree_add_190_195_groupi_g40307(csa_tree_add_190_195_groupi_n_8818 ,csa_tree_add_190_195_groupi_n_8180 ,csa_tree_add_190_195_groupi_n_8436);
  and csa_tree_add_190_195_groupi_g40308(csa_tree_add_190_195_groupi_n_8816 ,csa_tree_add_190_195_groupi_n_8153 ,csa_tree_add_190_195_groupi_n_8406);
  and csa_tree_add_190_195_groupi_g40309(csa_tree_add_190_195_groupi_n_8814 ,csa_tree_add_190_195_groupi_n_8122 ,csa_tree_add_190_195_groupi_n_8414);
  and csa_tree_add_190_195_groupi_g40310(csa_tree_add_190_195_groupi_n_8812 ,csa_tree_add_190_195_groupi_n_8098 ,csa_tree_add_190_195_groupi_n_8410);
  not csa_tree_add_190_195_groupi_g40311(csa_tree_add_190_195_groupi_n_8719 ,csa_tree_add_190_195_groupi_n_8718);
  not csa_tree_add_190_195_groupi_g40314(csa_tree_add_190_195_groupi_n_8715 ,csa_tree_add_190_195_groupi_n_8714);
  not csa_tree_add_190_195_groupi_g40315(csa_tree_add_190_195_groupi_n_8711 ,csa_tree_add_190_195_groupi_n_8710);
  not csa_tree_add_190_195_groupi_g40316(csa_tree_add_190_195_groupi_n_8703 ,csa_tree_add_190_195_groupi_n_8702);
  not csa_tree_add_190_195_groupi_g40317(csa_tree_add_190_195_groupi_n_8697 ,csa_tree_add_190_195_groupi_n_8696);
  not csa_tree_add_190_195_groupi_g40318(csa_tree_add_190_195_groupi_n_8695 ,csa_tree_add_190_195_groupi_n_8694);
  not csa_tree_add_190_195_groupi_g40319(csa_tree_add_190_195_groupi_n_8693 ,csa_tree_add_190_195_groupi_n_8692);
  not csa_tree_add_190_195_groupi_g40320(csa_tree_add_190_195_groupi_n_8690 ,csa_tree_add_190_195_groupi_n_8689);
  not csa_tree_add_190_195_groupi_g40321(csa_tree_add_190_195_groupi_n_8686 ,csa_tree_add_190_195_groupi_n_8687);
  not csa_tree_add_190_195_groupi_g40322(csa_tree_add_190_195_groupi_n_8685 ,csa_tree_add_190_195_groupi_n_8684);
  not csa_tree_add_190_195_groupi_g40323(csa_tree_add_190_195_groupi_n_8683 ,csa_tree_add_190_195_groupi_n_8682);
  not csa_tree_add_190_195_groupi_g40324(csa_tree_add_190_195_groupi_n_8681 ,csa_tree_add_190_195_groupi_n_8680);
  not csa_tree_add_190_195_groupi_g40325(csa_tree_add_190_195_groupi_n_8679 ,csa_tree_add_190_195_groupi_n_8678);
  not csa_tree_add_190_195_groupi_g40326(csa_tree_add_190_195_groupi_n_8677 ,csa_tree_add_190_195_groupi_n_8676);
  not csa_tree_add_190_195_groupi_g40327(csa_tree_add_190_195_groupi_n_8675 ,csa_tree_add_190_195_groupi_n_8674);
  not csa_tree_add_190_195_groupi_g40328(csa_tree_add_190_195_groupi_n_8671 ,csa_tree_add_190_195_groupi_n_8672);
  not csa_tree_add_190_195_groupi_g40329(csa_tree_add_190_195_groupi_n_8670 ,csa_tree_add_190_195_groupi_n_8669);
  not csa_tree_add_190_195_groupi_g40330(csa_tree_add_190_195_groupi_n_8668 ,csa_tree_add_190_195_groupi_n_8667);
  not csa_tree_add_190_195_groupi_g40331(csa_tree_add_190_195_groupi_n_8666 ,csa_tree_add_190_195_groupi_n_8665);
  not csa_tree_add_190_195_groupi_g40332(csa_tree_add_190_195_groupi_n_8661 ,csa_tree_add_190_195_groupi_n_112);
  not csa_tree_add_190_195_groupi_g40333(csa_tree_add_190_195_groupi_n_8660 ,csa_tree_add_190_195_groupi_n_8659);
  not csa_tree_add_190_195_groupi_g40334(csa_tree_add_190_195_groupi_n_8658 ,csa_tree_add_190_195_groupi_n_8657);
  not csa_tree_add_190_195_groupi_g40335(csa_tree_add_190_195_groupi_n_8655 ,csa_tree_add_190_195_groupi_n_8654);
  not csa_tree_add_190_195_groupi_g40336(csa_tree_add_190_195_groupi_n_8652 ,csa_tree_add_190_195_groupi_n_8653);
  not csa_tree_add_190_195_groupi_g40337(csa_tree_add_190_195_groupi_n_8651 ,csa_tree_add_190_195_groupi_n_8650);
  not csa_tree_add_190_195_groupi_g40338(csa_tree_add_190_195_groupi_n_8649 ,csa_tree_add_190_195_groupi_n_8648);
  not csa_tree_add_190_195_groupi_g40339(csa_tree_add_190_195_groupi_n_8646 ,csa_tree_add_190_195_groupi_n_8645);
  not csa_tree_add_190_195_groupi_g40340(csa_tree_add_190_195_groupi_n_8643 ,csa_tree_add_190_195_groupi_n_8644);
  not csa_tree_add_190_195_groupi_g40341(csa_tree_add_190_195_groupi_n_8641 ,csa_tree_add_190_195_groupi_n_8640);
  not csa_tree_add_190_195_groupi_g40342(csa_tree_add_190_195_groupi_n_8638 ,csa_tree_add_190_195_groupi_n_8639);
  not csa_tree_add_190_195_groupi_g40343(csa_tree_add_190_195_groupi_n_8637 ,csa_tree_add_190_195_groupi_n_8636);
  not csa_tree_add_190_195_groupi_g40344(csa_tree_add_190_195_groupi_n_8634 ,csa_tree_add_190_195_groupi_n_109);
  not csa_tree_add_190_195_groupi_g40345(csa_tree_add_190_195_groupi_n_8632 ,csa_tree_add_190_195_groupi_n_8631);
  not csa_tree_add_190_195_groupi_g40346(csa_tree_add_190_195_groupi_n_8630 ,csa_tree_add_190_195_groupi_n_8629);
  not csa_tree_add_190_195_groupi_g40347(csa_tree_add_190_195_groupi_n_8628 ,csa_tree_add_190_195_groupi_n_8627);
  not csa_tree_add_190_195_groupi_g40348(csa_tree_add_190_195_groupi_n_8625 ,csa_tree_add_190_195_groupi_n_8626);
  not csa_tree_add_190_195_groupi_g40349(csa_tree_add_190_195_groupi_n_8623 ,csa_tree_add_190_195_groupi_n_8624);
  not csa_tree_add_190_195_groupi_g40350(csa_tree_add_190_195_groupi_n_8622 ,csa_tree_add_190_195_groupi_n_8621);
  not csa_tree_add_190_195_groupi_g40351(csa_tree_add_190_195_groupi_n_8618 ,csa_tree_add_190_195_groupi_n_8619);
  not csa_tree_add_190_195_groupi_g40352(csa_tree_add_190_195_groupi_n_8615 ,csa_tree_add_190_195_groupi_n_8616);
  not csa_tree_add_190_195_groupi_g40353(csa_tree_add_190_195_groupi_n_8613 ,csa_tree_add_190_195_groupi_n_8612);
  not csa_tree_add_190_195_groupi_g40354(csa_tree_add_190_195_groupi_n_8609 ,csa_tree_add_190_195_groupi_n_8608);
  and csa_tree_add_190_195_groupi_g40355(csa_tree_add_190_195_groupi_n_8607 ,csa_tree_add_190_195_groupi_n_7565 ,csa_tree_add_190_195_groupi_n_8315);
  or csa_tree_add_190_195_groupi_g40356(csa_tree_add_190_195_groupi_n_8606 ,csa_tree_add_190_195_groupi_n_7565 ,csa_tree_add_190_195_groupi_n_8315);
  nor csa_tree_add_190_195_groupi_g40357(csa_tree_add_190_195_groupi_n_8605 ,csa_tree_add_190_195_groupi_n_8056 ,csa_tree_add_190_195_groupi_n_8396);
  or csa_tree_add_190_195_groupi_g40358(csa_tree_add_190_195_groupi_n_8604 ,csa_tree_add_190_195_groupi_n_7954 ,csa_tree_add_190_195_groupi_n_8514);
  or csa_tree_add_190_195_groupi_g40359(csa_tree_add_190_195_groupi_n_8603 ,csa_tree_add_190_195_groupi_n_8328 ,csa_tree_add_190_195_groupi_n_7321);
  or csa_tree_add_190_195_groupi_g40360(csa_tree_add_190_195_groupi_n_8602 ,csa_tree_add_190_195_groupi_n_8540 ,csa_tree_add_190_195_groupi_n_7809);
  nor csa_tree_add_190_195_groupi_g40361(csa_tree_add_190_195_groupi_n_8601 ,csa_tree_add_190_195_groupi_n_8329 ,csa_tree_add_190_195_groupi_n_7320);
  or csa_tree_add_190_195_groupi_g40362(csa_tree_add_190_195_groupi_n_8600 ,csa_tree_add_190_195_groupi_n_8534 ,csa_tree_add_190_195_groupi_n_8462);
  nor csa_tree_add_190_195_groupi_g40363(csa_tree_add_190_195_groupi_n_8599 ,csa_tree_add_190_195_groupi_n_8373 ,csa_tree_add_190_195_groupi_n_8375);
  and csa_tree_add_190_195_groupi_g40364(csa_tree_add_190_195_groupi_n_8598 ,csa_tree_add_190_195_groupi_n_8373 ,csa_tree_add_190_195_groupi_n_8375);
  or csa_tree_add_190_195_groupi_g40365(csa_tree_add_190_195_groupi_n_8597 ,csa_tree_add_190_195_groupi_n_7188 ,csa_tree_add_190_195_groupi_n_8376);
  nor csa_tree_add_190_195_groupi_g40366(csa_tree_add_190_195_groupi_n_8596 ,csa_tree_add_190_195_groupi_n_7189 ,csa_tree_add_190_195_groupi_n_8377);
  or csa_tree_add_190_195_groupi_g40367(csa_tree_add_190_195_groupi_n_8595 ,csa_tree_add_190_195_groupi_n_6456 ,csa_tree_add_190_195_groupi_n_8381);
  or csa_tree_add_190_195_groupi_g40368(csa_tree_add_190_195_groupi_n_8594 ,csa_tree_add_190_195_groupi_n_8037 ,csa_tree_add_190_195_groupi_n_8301);
  and csa_tree_add_190_195_groupi_g40369(csa_tree_add_190_195_groupi_n_8593 ,csa_tree_add_190_195_groupi_n_8005 ,csa_tree_add_190_195_groupi_n_8340);
  or csa_tree_add_190_195_groupi_g40370(csa_tree_add_190_195_groupi_n_8592 ,csa_tree_add_190_195_groupi_n_7166 ,csa_tree_add_190_195_groupi_n_8316);
  nor csa_tree_add_190_195_groupi_g40371(csa_tree_add_190_195_groupi_n_8591 ,csa_tree_add_190_195_groupi_n_7165 ,csa_tree_add_190_195_groupi_n_8317);
  nor csa_tree_add_190_195_groupi_g40372(csa_tree_add_190_195_groupi_n_8590 ,csa_tree_add_190_195_groupi_n_8005 ,csa_tree_add_190_195_groupi_n_8340);
  or csa_tree_add_190_195_groupi_g40373(csa_tree_add_190_195_groupi_n_8589 ,csa_tree_add_190_195_groupi_n_6379 ,csa_tree_add_190_195_groupi_n_8539);
  or csa_tree_add_190_195_groupi_g40374(csa_tree_add_190_195_groupi_n_8588 ,csa_tree_add_190_195_groupi_n_7729 ,csa_tree_add_190_195_groupi_n_13);
  xnor csa_tree_add_190_195_groupi_g40375(csa_tree_add_190_195_groupi_n_8587 ,csa_tree_add_190_195_groupi_n_4690 ,csa_tree_add_190_195_groupi_n_101);
  xnor csa_tree_add_190_195_groupi_g40376(csa_tree_add_190_195_groupi_n_8586 ,csa_tree_add_190_195_groupi_n_7535 ,csa_tree_add_190_195_groupi_n_8053);
  xnor csa_tree_add_190_195_groupi_g40377(csa_tree_add_190_195_groupi_n_8585 ,csa_tree_add_190_195_groupi_n_7657 ,csa_tree_add_190_195_groupi_n_7997);
  xnor csa_tree_add_190_195_groupi_g40378(csa_tree_add_190_195_groupi_n_8584 ,csa_tree_add_190_195_groupi_n_8199 ,csa_tree_add_190_195_groupi_n_7522);
  xor csa_tree_add_190_195_groupi_g40379(csa_tree_add_190_195_groupi_n_8583 ,csa_tree_add_190_195_groupi_n_7378 ,csa_tree_add_190_195_groupi_n_8219);
  xnor csa_tree_add_190_195_groupi_g40380(csa_tree_add_190_195_groupi_n_8582 ,csa_tree_add_190_195_groupi_n_4975 ,csa_tree_add_190_195_groupi_n_8227);
  xnor csa_tree_add_190_195_groupi_g40381(csa_tree_add_190_195_groupi_n_8581 ,csa_tree_add_190_195_groupi_n_4771 ,csa_tree_add_190_195_groupi_n_8226);
  xnor csa_tree_add_190_195_groupi_g40382(csa_tree_add_190_195_groupi_n_8580 ,csa_tree_add_190_195_groupi_n_8038 ,csa_tree_add_190_195_groupi_n_5366);
  xnor csa_tree_add_190_195_groupi_g40383(csa_tree_add_190_195_groupi_n_8579 ,csa_tree_add_190_195_groupi_n_8231 ,csa_tree_add_190_195_groupi_n_7534);
  xor csa_tree_add_190_195_groupi_g40384(csa_tree_add_190_195_groupi_n_8578 ,csa_tree_add_190_195_groupi_n_6768 ,csa_tree_add_190_195_groupi_n_8215);
  xnor csa_tree_add_190_195_groupi_g40385(csa_tree_add_190_195_groupi_n_8577 ,csa_tree_add_190_195_groupi_n_7525 ,csa_tree_add_190_195_groupi_n_8055);
  xnor csa_tree_add_190_195_groupi_g40386(csa_tree_add_190_195_groupi_n_8576 ,csa_tree_add_190_195_groupi_n_5039 ,csa_tree_add_190_195_groupi_n_8230);
  xnor csa_tree_add_190_195_groupi_g40387(csa_tree_add_190_195_groupi_n_8575 ,csa_tree_add_190_195_groupi_n_7861 ,csa_tree_add_190_195_groupi_n_8203);
  xnor csa_tree_add_190_195_groupi_g40388(csa_tree_add_190_195_groupi_n_8574 ,csa_tree_add_190_195_groupi_n_4607 ,csa_tree_add_190_195_groupi_n_8035);
  xnor csa_tree_add_190_195_groupi_g40389(csa_tree_add_190_195_groupi_n_8573 ,csa_tree_add_190_195_groupi_n_5384 ,csa_tree_add_190_195_groupi_n_8043);
  xnor csa_tree_add_190_195_groupi_g40390(csa_tree_add_190_195_groupi_n_8572 ,csa_tree_add_190_195_groupi_n_5471 ,csa_tree_add_190_195_groupi_n_7998);
  xnor csa_tree_add_190_195_groupi_g40391(csa_tree_add_190_195_groupi_n_8571 ,csa_tree_add_190_195_groupi_n_6756 ,csa_tree_add_190_195_groupi_n_7990);
  xnor csa_tree_add_190_195_groupi_g40392(csa_tree_add_190_195_groupi_n_8570 ,csa_tree_add_190_195_groupi_n_4649 ,csa_tree_add_190_195_groupi_n_8034);
  xnor csa_tree_add_190_195_groupi_g40393(csa_tree_add_190_195_groupi_n_8569 ,csa_tree_add_190_195_groupi_n_65 ,csa_tree_add_190_195_groupi_n_8193);
  xnor csa_tree_add_190_195_groupi_g40394(csa_tree_add_190_195_groupi_n_8568 ,csa_tree_add_190_195_groupi_n_8046 ,csa_tree_add_190_195_groupi_n_5389);
  xnor csa_tree_add_190_195_groupi_g40395(csa_tree_add_190_195_groupi_n_8567 ,csa_tree_add_190_195_groupi_n_46 ,csa_tree_add_190_195_groupi_n_8009);
  xnor csa_tree_add_190_195_groupi_g40397(csa_tree_add_190_195_groupi_n_8566 ,csa_tree_add_190_195_groupi_n_4712 ,csa_tree_add_190_195_groupi_n_8058);
  xnor csa_tree_add_190_195_groupi_g40398(csa_tree_add_190_195_groupi_n_8565 ,csa_tree_add_190_195_groupi_n_7502 ,csa_tree_add_190_195_groupi_n_8036);
  xnor csa_tree_add_190_195_groupi_g40399(csa_tree_add_190_195_groupi_n_8564 ,csa_tree_add_190_195_groupi_n_20 ,csa_tree_add_190_195_groupi_n_8224);
  xnor csa_tree_add_190_195_groupi_g40400(csa_tree_add_190_195_groupi_n_8563 ,csa_tree_add_190_195_groupi_n_7356 ,csa_tree_add_190_195_groupi_n_8059);
  xnor csa_tree_add_190_195_groupi_g40401(csa_tree_add_190_195_groupi_n_8562 ,csa_tree_add_190_195_groupi_n_5493 ,csa_tree_add_190_195_groupi_n_8221);
  xnor csa_tree_add_190_195_groupi_g40402(csa_tree_add_190_195_groupi_n_8561 ,csa_tree_add_190_195_groupi_n_8220 ,csa_tree_add_190_195_groupi_n_5079);
  xnor csa_tree_add_190_195_groupi_g40403(csa_tree_add_190_195_groupi_n_8560 ,csa_tree_add_190_195_groupi_n_4664 ,csa_tree_add_190_195_groupi_n_8007);
  xnor csa_tree_add_190_195_groupi_g40404(csa_tree_add_190_195_groupi_n_8559 ,csa_tree_add_190_195_groupi_n_5503 ,csa_tree_add_190_195_groupi_n_8052);
  xnor csa_tree_add_190_195_groupi_g40405(csa_tree_add_190_195_groupi_n_8558 ,csa_tree_add_190_195_groupi_n_8005 ,csa_tree_add_190_195_groupi_n_7656);
  xnor csa_tree_add_190_195_groupi_g40406(csa_tree_add_190_195_groupi_n_8557 ,csa_tree_add_190_195_groupi_n_8186 ,csa_tree_add_190_195_groupi_n_7863);
  xnor csa_tree_add_190_195_groupi_g40407(csa_tree_add_190_195_groupi_n_8556 ,csa_tree_add_190_195_groupi_n_5868 ,csa_tree_add_190_195_groupi_n_8013);
  xnor csa_tree_add_190_195_groupi_g40408(csa_tree_add_190_195_groupi_n_8555 ,csa_tree_add_190_195_groupi_n_8218 ,csa_tree_add_190_195_groupi_n_8189);
  xnor csa_tree_add_190_195_groupi_g40409(csa_tree_add_190_195_groupi_n_8554 ,csa_tree_add_190_195_groupi_n_5501 ,csa_tree_add_190_195_groupi_n_8033);
  xnor csa_tree_add_190_195_groupi_g40410(csa_tree_add_190_195_groupi_n_8553 ,csa_tree_add_190_195_groupi_n_5041 ,csa_tree_add_190_195_groupi_n_8205);
  xnor csa_tree_add_190_195_groupi_g40411(csa_tree_add_190_195_groupi_n_8552 ,csa_tree_add_190_195_groupi_n_8041 ,csa_tree_add_190_195_groupi_n_5224);
  xnor csa_tree_add_190_195_groupi_g40412(csa_tree_add_190_195_groupi_n_8551 ,csa_tree_add_190_195_groupi_n_8196 ,csa_tree_add_190_195_groupi_n_7415);
  xnor csa_tree_add_190_195_groupi_g40413(csa_tree_add_190_195_groupi_n_8550 ,csa_tree_add_190_195_groupi_n_5304 ,csa_tree_add_190_195_groupi_n_8232);
  xnor csa_tree_add_190_195_groupi_g40414(csa_tree_add_190_195_groupi_n_8549 ,csa_tree_add_190_195_groupi_n_8210 ,csa_tree_add_190_195_groupi_n_7516);
  xnor csa_tree_add_190_195_groupi_g40415(csa_tree_add_190_195_groupi_n_8548 ,csa_tree_add_190_195_groupi_n_7580 ,csa_tree_add_190_195_groupi_n_7987);
  xnor csa_tree_add_190_195_groupi_g40416(csa_tree_add_190_195_groupi_n_8547 ,csa_tree_add_190_195_groupi_n_7510 ,csa_tree_add_190_195_groupi_n_8057);
  xnor csa_tree_add_190_195_groupi_g40417(csa_tree_add_190_195_groupi_n_8723 ,csa_tree_add_190_195_groupi_n_8042 ,csa_tree_add_190_195_groupi_n_7924);
  xnor csa_tree_add_190_195_groupi_g40418(csa_tree_add_190_195_groupi_n_8722 ,csa_tree_add_190_195_groupi_n_5371 ,csa_tree_add_190_195_groupi_n_7921);
  xnor csa_tree_add_190_195_groupi_g40419(csa_tree_add_190_195_groupi_n_8721 ,csa_tree_add_190_195_groupi_n_7896 ,csa_tree_add_190_195_groupi_n_1228);
  xnor csa_tree_add_190_195_groupi_g40420(csa_tree_add_190_195_groupi_n_8720 ,csa_tree_add_190_195_groupi_n_7894 ,csa_tree_add_190_195_groupi_n_1948);
  xnor csa_tree_add_190_195_groupi_g40421(csa_tree_add_190_195_groupi_n_8718 ,csa_tree_add_190_195_groupi_n_7879 ,csa_tree_add_190_195_groupi_n_574);
  xnor csa_tree_add_190_195_groupi_g40422(csa_tree_add_190_195_groupi_n_8717 ,csa_tree_add_190_195_groupi_n_5922 ,csa_tree_add_190_195_groupi_n_7931);
  and csa_tree_add_190_195_groupi_g40423(csa_tree_add_190_195_groupi_n_8716 ,csa_tree_add_190_195_groupi_n_6324 ,csa_tree_add_190_195_groupi_n_8293);
  xnor csa_tree_add_190_195_groupi_g40424(csa_tree_add_190_195_groupi_n_8714 ,csa_tree_add_190_195_groupi_n_7136 ,csa_tree_add_190_195_groupi_n_7881);
  xnor csa_tree_add_190_195_groupi_g40425(csa_tree_add_190_195_groupi_n_8713 ,csa_tree_add_190_195_groupi_n_5355 ,csa_tree_add_190_195_groupi_n_7889);
  xnor csa_tree_add_190_195_groupi_g40426(csa_tree_add_190_195_groupi_n_8712 ,csa_tree_add_190_195_groupi_n_5037 ,csa_tree_add_190_195_groupi_n_7911);
  xnor csa_tree_add_190_195_groupi_g40427(csa_tree_add_190_195_groupi_n_8710 ,csa_tree_add_190_195_groupi_n_7897 ,csa_tree_add_190_195_groupi_n_2158);
  xnor csa_tree_add_190_195_groupi_g40429(csa_tree_add_190_195_groupi_n_8709 ,csa_tree_add_190_195_groupi_n_104 ,csa_tree_add_190_195_groupi_n_1179);
  xnor csa_tree_add_190_195_groupi_g40430(csa_tree_add_190_195_groupi_n_8708 ,csa_tree_add_190_195_groupi_n_66 ,csa_tree_add_190_195_groupi_n_7925);
  xnor csa_tree_add_190_195_groupi_g40431(csa_tree_add_190_195_groupi_n_8707 ,csa_tree_add_190_195_groupi_n_58 ,csa_tree_add_190_195_groupi_n_7942);
  xnor csa_tree_add_190_195_groupi_g40432(csa_tree_add_190_195_groupi_n_8706 ,csa_tree_add_190_195_groupi_n_7915 ,csa_tree_add_190_195_groupi_n_2041);
  xnor csa_tree_add_190_195_groupi_g40433(csa_tree_add_190_195_groupi_n_8705 ,csa_tree_add_190_195_groupi_n_7936 ,csa_tree_add_190_195_groupi_n_1018);
  xnor csa_tree_add_190_195_groupi_g40434(csa_tree_add_190_195_groupi_n_8704 ,csa_tree_add_190_195_groupi_n_6996 ,csa_tree_add_190_195_groupi_n_7900);
  xnor csa_tree_add_190_195_groupi_g40435(csa_tree_add_190_195_groupi_n_8702 ,csa_tree_add_190_195_groupi_n_7934 ,csa_tree_add_190_195_groupi_n_1827);
  and csa_tree_add_190_195_groupi_g40436(csa_tree_add_190_195_groupi_n_8701 ,csa_tree_add_190_195_groupi_n_6193 ,csa_tree_add_190_195_groupi_n_8290);
  and csa_tree_add_190_195_groupi_g40437(csa_tree_add_190_195_groupi_n_8700 ,csa_tree_add_190_195_groupi_n_8176 ,csa_tree_add_190_195_groupi_n_8292);
  and csa_tree_add_190_195_groupi_g40438(csa_tree_add_190_195_groupi_n_8699 ,csa_tree_add_190_195_groupi_n_5810 ,csa_tree_add_190_195_groupi_n_8303);
  xnor csa_tree_add_190_195_groupi_g40439(csa_tree_add_190_195_groupi_n_8698 ,csa_tree_add_190_195_groupi_n_4891 ,csa_tree_add_190_195_groupi_n_7885);
  xnor csa_tree_add_190_195_groupi_g40440(csa_tree_add_190_195_groupi_n_8696 ,csa_tree_add_190_195_groupi_n_7558 ,csa_tree_add_190_195_groupi_n_7883);
  xnor csa_tree_add_190_195_groupi_g40441(csa_tree_add_190_195_groupi_n_8694 ,csa_tree_add_190_195_groupi_n_5487 ,csa_tree_add_190_195_groupi_n_7882);
  xnor csa_tree_add_190_195_groupi_g40442(csa_tree_add_190_195_groupi_n_8692 ,csa_tree_add_190_195_groupi_n_7232 ,csa_tree_add_190_195_groupi_n_7903);
  or csa_tree_add_190_195_groupi_g40443(csa_tree_add_190_195_groupi_n_8691 ,csa_tree_add_190_195_groupi_n_114 ,csa_tree_add_190_195_groupi_n_1332);
  xnor csa_tree_add_190_195_groupi_g40444(csa_tree_add_190_195_groupi_n_8689 ,csa_tree_add_190_195_groupi_n_6951 ,csa_tree_add_190_195_groupi_n_7928);
  xnor csa_tree_add_190_195_groupi_g40445(csa_tree_add_190_195_groupi_n_8688 ,csa_tree_add_190_195_groupi_n_7106 ,csa_tree_add_190_195_groupi_n_7902);
  xnor csa_tree_add_190_195_groupi_g40446(csa_tree_add_190_195_groupi_n_8687 ,csa_tree_add_190_195_groupi_n_4916 ,csa_tree_add_190_195_groupi_n_7926);
  xnor csa_tree_add_190_195_groupi_g40447(csa_tree_add_190_195_groupi_n_8684 ,csa_tree_add_190_195_groupi_n_5236 ,csa_tree_add_190_195_groupi_n_102);
  xnor csa_tree_add_190_195_groupi_g40448(csa_tree_add_190_195_groupi_n_8682 ,csa_tree_add_190_195_groupi_n_5348 ,csa_tree_add_190_195_groupi_n_7878);
  xnor csa_tree_add_190_195_groupi_g40449(csa_tree_add_190_195_groupi_n_8680 ,csa_tree_add_190_195_groupi_n_5406 ,csa_tree_add_190_195_groupi_n_7888);
  xnor csa_tree_add_190_195_groupi_g40450(csa_tree_add_190_195_groupi_n_8678 ,csa_tree_add_190_195_groupi_n_7850 ,csa_tree_add_190_195_groupi_n_7890);
  xnor csa_tree_add_190_195_groupi_g40451(csa_tree_add_190_195_groupi_n_8676 ,csa_tree_add_190_195_groupi_n_6757 ,csa_tree_add_190_195_groupi_n_7892);
  xnor csa_tree_add_190_195_groupi_g40452(csa_tree_add_190_195_groupi_n_8674 ,csa_tree_add_190_195_groupi_n_22 ,csa_tree_add_190_195_groupi_n_1232);
  xnor csa_tree_add_190_195_groupi_g40453(csa_tree_add_190_195_groupi_n_8673 ,csa_tree_add_190_195_groupi_n_6281 ,csa_tree_add_190_195_groupi_n_7901);
  xnor csa_tree_add_190_195_groupi_g40454(csa_tree_add_190_195_groupi_n_8672 ,csa_tree_add_190_195_groupi_n_5484 ,csa_tree_add_190_195_groupi_n_7935);
  xnor csa_tree_add_190_195_groupi_g40455(csa_tree_add_190_195_groupi_n_8669 ,csa_tree_add_190_195_groupi_n_8216 ,csa_tree_add_190_195_groupi_n_6075);
  xnor csa_tree_add_190_195_groupi_g40456(csa_tree_add_190_195_groupi_n_8667 ,csa_tree_add_190_195_groupi_n_7133 ,csa_tree_add_190_195_groupi_n_7914);
  xnor csa_tree_add_190_195_groupi_g40457(csa_tree_add_190_195_groupi_n_8665 ,csa_tree_add_190_195_groupi_n_7555 ,csa_tree_add_190_195_groupi_n_7899);
  xnor csa_tree_add_190_195_groupi_g40458(csa_tree_add_190_195_groupi_n_8664 ,csa_tree_add_190_195_groupi_n_6969 ,csa_tree_add_190_195_groupi_n_7905);
  xnor csa_tree_add_190_195_groupi_g40459(csa_tree_add_190_195_groupi_n_8663 ,csa_tree_add_190_195_groupi_n_6773 ,csa_tree_add_190_195_groupi_n_7933);
  xnor csa_tree_add_190_195_groupi_g40460(csa_tree_add_190_195_groupi_n_8662 ,csa_tree_add_190_195_groupi_n_7513 ,csa_tree_add_190_195_groupi_n_7907);
  and csa_tree_add_190_195_groupi_g40462(csa_tree_add_190_195_groupi_n_8659 ,csa_tree_add_190_195_groupi_n_7962 ,csa_tree_add_190_195_groupi_n_8306);
  xnor csa_tree_add_190_195_groupi_g40463(csa_tree_add_190_195_groupi_n_8657 ,csa_tree_add_190_195_groupi_n_7390 ,csa_tree_add_190_195_groupi_n_7913);
  xnor csa_tree_add_190_195_groupi_g40464(csa_tree_add_190_195_groupi_n_8656 ,csa_tree_add_190_195_groupi_n_8054 ,csa_tree_add_190_195_groupi_n_6711);
  xnor csa_tree_add_190_195_groupi_g40465(csa_tree_add_190_195_groupi_n_8654 ,csa_tree_add_190_195_groupi_n_7615 ,csa_tree_add_190_195_groupi_n_7929);
  xnor csa_tree_add_190_195_groupi_g40466(csa_tree_add_190_195_groupi_n_8653 ,csa_tree_add_190_195_groupi_n_6280 ,csa_tree_add_190_195_groupi_n_7912);
  xnor csa_tree_add_190_195_groupi_g40467(csa_tree_add_190_195_groupi_n_8650 ,csa_tree_add_190_195_groupi_n_5387 ,csa_tree_add_190_195_groupi_n_106);
  xnor csa_tree_add_190_195_groupi_g40468(csa_tree_add_190_195_groupi_n_8648 ,csa_tree_add_190_195_groupi_n_7500 ,csa_tree_add_190_195_groupi_n_7898);
  or csa_tree_add_190_195_groupi_g40469(csa_tree_add_190_195_groupi_n_8647 ,csa_tree_add_190_195_groupi_n_5802 ,csa_tree_add_190_195_groupi_n_8289);
  xnor csa_tree_add_190_195_groupi_g40470(csa_tree_add_190_195_groupi_n_8645 ,csa_tree_add_190_195_groupi_n_7872 ,csa_tree_add_190_195_groupi_n_7895);
  xnor csa_tree_add_190_195_groupi_g40471(csa_tree_add_190_195_groupi_n_8644 ,csa_tree_add_190_195_groupi_n_7597 ,csa_tree_add_190_195_groupi_n_7937);
  xnor csa_tree_add_190_195_groupi_g40472(csa_tree_add_190_195_groupi_n_8642 ,csa_tree_add_190_195_groupi_n_6925 ,csa_tree_add_190_195_groupi_n_7886);
  xnor csa_tree_add_190_195_groupi_g40473(csa_tree_add_190_195_groupi_n_8640 ,csa_tree_add_190_195_groupi_n_5365 ,csa_tree_add_190_195_groupi_n_7891);
  xnor csa_tree_add_190_195_groupi_g40474(csa_tree_add_190_195_groupi_n_8639 ,csa_tree_add_190_195_groupi_n_8222 ,csa_tree_add_190_195_groupi_n_6668);
  xnor csa_tree_add_190_195_groupi_g40475(csa_tree_add_190_195_groupi_n_8636 ,csa_tree_add_190_195_groupi_n_5352 ,csa_tree_add_190_195_groupi_n_7908);
  xnor csa_tree_add_190_195_groupi_g40476(csa_tree_add_190_195_groupi_n_8635 ,csa_tree_add_190_195_groupi_n_7405 ,csa_tree_add_190_195_groupi_n_7938);
  xnor csa_tree_add_190_195_groupi_g40478(csa_tree_add_190_195_groupi_n_8633 ,csa_tree_add_190_195_groupi_n_8050 ,csa_tree_add_190_195_groupi_n_6680);
  xnor csa_tree_add_190_195_groupi_g40479(csa_tree_add_190_195_groupi_n_8631 ,csa_tree_add_190_195_groupi_n_8047 ,csa_tree_add_190_195_groupi_n_6619);
  xnor csa_tree_add_190_195_groupi_g40480(csa_tree_add_190_195_groupi_n_8629 ,csa_tree_add_190_195_groupi_n_7426 ,csa_tree_add_190_195_groupi_n_7906);
  xnor csa_tree_add_190_195_groupi_g40481(csa_tree_add_190_195_groupi_n_8627 ,csa_tree_add_190_195_groupi_n_7411 ,csa_tree_add_190_195_groupi_n_7940);
  xnor csa_tree_add_190_195_groupi_g40482(csa_tree_add_190_195_groupi_n_8626 ,csa_tree_add_190_195_groupi_n_7075 ,csa_tree_add_190_195_groupi_n_7927);
  xnor csa_tree_add_190_195_groupi_g40483(csa_tree_add_190_195_groupi_n_8624 ,csa_tree_add_190_195_groupi_n_8049 ,csa_tree_add_190_195_groupi_n_6693);
  xnor csa_tree_add_190_195_groupi_g40484(csa_tree_add_190_195_groupi_n_8621 ,csa_tree_add_190_195_groupi_n_7196 ,csa_tree_add_190_195_groupi_n_7939);
  xnor csa_tree_add_190_195_groupi_g40485(csa_tree_add_190_195_groupi_n_8620 ,csa_tree_add_190_195_groupi_n_4655 ,csa_tree_add_190_195_groupi_n_7922);
  xnor csa_tree_add_190_195_groupi_g40486(csa_tree_add_190_195_groupi_n_8619 ,csa_tree_add_190_195_groupi_n_4977 ,csa_tree_add_190_195_groupi_n_7920);
  xnor csa_tree_add_190_195_groupi_g40487(csa_tree_add_190_195_groupi_n_8617 ,csa_tree_add_190_195_groupi_n_7864 ,csa_tree_add_190_195_groupi_n_7909);
  xnor csa_tree_add_190_195_groupi_g40488(csa_tree_add_190_195_groupi_n_8616 ,csa_tree_add_190_195_groupi_n_5223 ,csa_tree_add_190_195_groupi_n_7943);
  xnor csa_tree_add_190_195_groupi_g40489(csa_tree_add_190_195_groupi_n_8614 ,csa_tree_add_190_195_groupi_n_5358 ,csa_tree_add_190_195_groupi_n_7930);
  xnor csa_tree_add_190_195_groupi_g40490(csa_tree_add_190_195_groupi_n_8612 ,csa_tree_add_190_195_groupi_n_7178 ,csa_tree_add_190_195_groupi_n_7904);
  xnor csa_tree_add_190_195_groupi_g40491(csa_tree_add_190_195_groupi_n_8611 ,csa_tree_add_190_195_groupi_n_7174 ,csa_tree_add_190_195_groupi_n_7884);
  xnor csa_tree_add_190_195_groupi_g40492(csa_tree_add_190_195_groupi_n_8610 ,csa_tree_add_190_195_groupi_n_4898 ,csa_tree_add_190_195_groupi_n_7944);
  xnor csa_tree_add_190_195_groupi_g40493(csa_tree_add_190_195_groupi_n_8608 ,csa_tree_add_190_195_groupi_n_7342 ,csa_tree_add_190_195_groupi_n_7932);
  not csa_tree_add_190_195_groupi_g40494(csa_tree_add_190_195_groupi_n_8546 ,csa_tree_add_190_195_groupi_n_8545);
  not csa_tree_add_190_195_groupi_g40495(csa_tree_add_190_195_groupi_n_8539 ,csa_tree_add_190_195_groupi_n_8538);
  not csa_tree_add_190_195_groupi_g40498(csa_tree_add_190_195_groupi_n_8527 ,csa_tree_add_190_195_groupi_n_8526);
  not csa_tree_add_190_195_groupi_g40499(csa_tree_add_190_195_groupi_n_8520 ,csa_tree_add_190_195_groupi_n_8519);
  not csa_tree_add_190_195_groupi_g40501(csa_tree_add_190_195_groupi_n_8503 ,csa_tree_add_190_195_groupi_n_8504);
  not csa_tree_add_190_195_groupi_g40502(csa_tree_add_190_195_groupi_n_8501 ,csa_tree_add_190_195_groupi_n_8500);
  not csa_tree_add_190_195_groupi_g40503(csa_tree_add_190_195_groupi_n_8498 ,csa_tree_add_190_195_groupi_n_8497);
  not csa_tree_add_190_195_groupi_g40504(csa_tree_add_190_195_groupi_n_8495 ,csa_tree_add_190_195_groupi_n_8496);
  not csa_tree_add_190_195_groupi_g40505(csa_tree_add_190_195_groupi_n_8494 ,csa_tree_add_190_195_groupi_n_8493);
  not csa_tree_add_190_195_groupi_g40506(csa_tree_add_190_195_groupi_n_8491 ,csa_tree_add_190_195_groupi_n_8490);
  not csa_tree_add_190_195_groupi_g40507(csa_tree_add_190_195_groupi_n_8487 ,csa_tree_add_190_195_groupi_n_8488);
  not csa_tree_add_190_195_groupi_g40508(csa_tree_add_190_195_groupi_n_8485 ,csa_tree_add_190_195_groupi_n_8484);
  not csa_tree_add_190_195_groupi_g40509(csa_tree_add_190_195_groupi_n_8482 ,csa_tree_add_190_195_groupi_n_8483);
  not csa_tree_add_190_195_groupi_g40510(csa_tree_add_190_195_groupi_n_8480 ,csa_tree_add_190_195_groupi_n_8479);
  or csa_tree_add_190_195_groupi_g40511(csa_tree_add_190_195_groupi_n_8478 ,csa_tree_add_190_195_groupi_n_7655 ,csa_tree_add_190_195_groupi_n_8088);
  or csa_tree_add_190_195_groupi_g40512(csa_tree_add_190_195_groupi_n_8477 ,csa_tree_add_190_195_groupi_n_7495 ,csa_tree_add_190_195_groupi_n_8025);
  nor csa_tree_add_190_195_groupi_g40513(csa_tree_add_190_195_groupi_n_8476 ,csa_tree_add_190_195_groupi_n_7103 ,csa_tree_add_190_195_groupi_n_8019);
  or csa_tree_add_190_195_groupi_g40514(csa_tree_add_190_195_groupi_n_8475 ,csa_tree_add_190_195_groupi_n_7814 ,csa_tree_add_190_195_groupi_n_8209);
  nor csa_tree_add_190_195_groupi_g40515(csa_tree_add_190_195_groupi_n_8474 ,csa_tree_add_190_195_groupi_n_5867 ,csa_tree_add_190_195_groupi_n_8013);
  or csa_tree_add_190_195_groupi_g40516(csa_tree_add_190_195_groupi_n_8473 ,csa_tree_add_190_195_groupi_n_7333 ,csa_tree_add_190_195_groupi_n_8202);
  or csa_tree_add_190_195_groupi_g40517(csa_tree_add_190_195_groupi_n_8472 ,csa_tree_add_190_195_groupi_n_5868 ,csa_tree_add_190_195_groupi_n_8012);
  nor csa_tree_add_190_195_groupi_g40518(csa_tree_add_190_195_groupi_n_8471 ,csa_tree_add_190_195_groupi_n_7334 ,csa_tree_add_190_195_groupi_n_8203);
  and csa_tree_add_190_195_groupi_g40519(csa_tree_add_190_195_groupi_n_8470 ,csa_tree_add_190_195_groupi_n_6791 ,csa_tree_add_190_195_groupi_n_8171);
  nor csa_tree_add_190_195_groupi_g40520(csa_tree_add_190_195_groupi_n_8469 ,csa_tree_add_190_195_groupi_n_7992 ,csa_tree_add_190_195_groupi_n_7612);
  or csa_tree_add_190_195_groupi_g40521(csa_tree_add_190_195_groupi_n_8468 ,csa_tree_add_190_195_groupi_n_65 ,csa_tree_add_190_195_groupi_n_8192);
  or csa_tree_add_190_195_groupi_g40522(csa_tree_add_190_195_groupi_n_8467 ,csa_tree_add_190_195_groupi_n_7993 ,csa_tree_add_190_195_groupi_n_7611);
  nor csa_tree_add_190_195_groupi_g40523(csa_tree_add_190_195_groupi_n_8466 ,csa_tree_add_190_195_groupi_n_5954 ,csa_tree_add_190_195_groupi_n_8193);
  or csa_tree_add_190_195_groupi_g40524(csa_tree_add_190_195_groupi_n_8465 ,csa_tree_add_190_195_groupi_n_6515 ,csa_tree_add_190_195_groupi_n_8046);
  or csa_tree_add_190_195_groupi_g40525(csa_tree_add_190_195_groupi_n_8464 ,csa_tree_add_190_195_groupi_n_8199 ,csa_tree_add_190_195_groupi_n_7521);
  nor csa_tree_add_190_195_groupi_g40526(csa_tree_add_190_195_groupi_n_8463 ,csa_tree_add_190_195_groupi_n_7877 ,csa_tree_add_190_195_groupi_n_7965);
  nor csa_tree_add_190_195_groupi_g40527(csa_tree_add_190_195_groupi_n_8462 ,csa_tree_add_190_195_groupi_n_8198 ,csa_tree_add_190_195_groupi_n_7522);
  nor csa_tree_add_190_195_groupi_g40528(csa_tree_add_190_195_groupi_n_8461 ,csa_tree_add_190_195_groupi_n_7496 ,csa_tree_add_190_195_groupi_n_8024);
  nor csa_tree_add_190_195_groupi_g40529(csa_tree_add_190_195_groupi_n_8460 ,csa_tree_add_190_195_groupi_n_5471 ,csa_tree_add_190_195_groupi_n_7998);
  and csa_tree_add_190_195_groupi_g40530(csa_tree_add_190_195_groupi_n_8459 ,csa_tree_add_190_195_groupi_n_5471 ,csa_tree_add_190_195_groupi_n_7998);
  nor csa_tree_add_190_195_groupi_g40531(csa_tree_add_190_195_groupi_n_8458 ,csa_tree_add_190_195_groupi_n_4611 ,csa_tree_add_190_195_groupi_n_8000);
  or csa_tree_add_190_195_groupi_g40532(csa_tree_add_190_195_groupi_n_8457 ,csa_tree_add_190_195_groupi_n_4610 ,csa_tree_add_190_195_groupi_n_7999);
  and csa_tree_add_190_195_groupi_g40533(csa_tree_add_190_195_groupi_n_8456 ,csa_tree_add_190_195_groupi_n_8030 ,csa_tree_add_190_195_groupi_n_7981);
  or csa_tree_add_190_195_groupi_g40534(csa_tree_add_190_195_groupi_n_8455 ,csa_tree_add_190_195_groupi_n_7388 ,csa_tree_add_190_195_groupi_n_8154);
  or csa_tree_add_190_195_groupi_g40535(csa_tree_add_190_195_groupi_n_8454 ,csa_tree_add_190_195_groupi_n_8030 ,csa_tree_add_190_195_groupi_n_7981);
  nor csa_tree_add_190_195_groupi_g40536(csa_tree_add_190_195_groupi_n_8453 ,csa_tree_add_190_195_groupi_n_4664 ,csa_tree_add_190_195_groupi_n_8006);
  or csa_tree_add_190_195_groupi_g40537(csa_tree_add_190_195_groupi_n_8452 ,csa_tree_add_190_195_groupi_n_7660 ,csa_tree_add_190_195_groupi_n_8147);
  or csa_tree_add_190_195_groupi_g40538(csa_tree_add_190_195_groupi_n_8451 ,csa_tree_add_190_195_groupi_n_7788 ,csa_tree_add_190_195_groupi_n_8221);
  or csa_tree_add_190_195_groupi_g40539(csa_tree_add_190_195_groupi_n_8450 ,csa_tree_add_190_195_groupi_n_6463 ,csa_tree_add_190_195_groupi_n_8222);
  nor csa_tree_add_190_195_groupi_g40540(csa_tree_add_190_195_groupi_n_8449 ,csa_tree_add_190_195_groupi_n_6756 ,csa_tree_add_190_195_groupi_n_7989);
  or csa_tree_add_190_195_groupi_g40541(csa_tree_add_190_195_groupi_n_8448 ,csa_tree_add_190_195_groupi_n_6755 ,csa_tree_add_190_195_groupi_n_7990);
  nor csa_tree_add_190_195_groupi_g40542(csa_tree_add_190_195_groupi_n_8447 ,csa_tree_add_190_195_groupi_n_8031 ,csa_tree_add_190_195_groupi_n_8004);
  or csa_tree_add_190_195_groupi_g40543(csa_tree_add_190_195_groupi_n_8446 ,csa_tree_add_190_195_groupi_n_8032 ,csa_tree_add_190_195_groupi_n_8003);
  and csa_tree_add_190_195_groupi_g40544(csa_tree_add_190_195_groupi_n_8445 ,csa_tree_add_190_195_groupi_n_7303 ,csa_tree_add_190_195_groupi_n_7979);
  and csa_tree_add_190_195_groupi_g40545(csa_tree_add_190_195_groupi_n_8444 ,csa_tree_add_190_195_groupi_n_6441 ,csa_tree_add_190_195_groupi_n_8049);
  nor csa_tree_add_190_195_groupi_g40546(csa_tree_add_190_195_groupi_n_8443 ,csa_tree_add_190_195_groupi_n_7303 ,csa_tree_add_190_195_groupi_n_7979);
  or csa_tree_add_190_195_groupi_g40547(csa_tree_add_190_195_groupi_n_8442 ,csa_tree_add_190_195_groupi_n_6128 ,csa_tree_add_190_195_groupi_n_8034);
  or csa_tree_add_190_195_groupi_g40548(csa_tree_add_190_195_groupi_n_8441 ,csa_tree_add_190_195_groupi_n_6132 ,csa_tree_add_190_195_groupi_n_8033);
  or csa_tree_add_190_195_groupi_g40549(csa_tree_add_190_195_groupi_n_8440 ,csa_tree_add_190_195_groupi_n_6424 ,csa_tree_add_190_195_groupi_n_8051);
  or csa_tree_add_190_195_groupi_g40550(csa_tree_add_190_195_groupi_n_8439 ,csa_tree_add_190_195_groupi_n_6134 ,csa_tree_add_190_195_groupi_n_8052);
  and csa_tree_add_190_195_groupi_g40551(csa_tree_add_190_195_groupi_n_8438 ,csa_tree_add_190_195_groupi_n_7212 ,csa_tree_add_190_195_groupi_n_8132);
  and csa_tree_add_190_195_groupi_g40552(csa_tree_add_190_195_groupi_n_8437 ,csa_tree_add_190_195_groupi_n_7210 ,csa_tree_add_190_195_groupi_n_8130);
  nor csa_tree_add_190_195_groupi_g40553(csa_tree_add_190_195_groupi_n_8436 ,csa_tree_add_190_195_groupi_n_7868 ,csa_tree_add_190_195_groupi_n_7977);
  or csa_tree_add_190_195_groupi_g40554(csa_tree_add_190_195_groupi_n_8435 ,csa_tree_add_190_195_groupi_n_5688 ,csa_tree_add_190_195_groupi_n_101);
  or csa_tree_add_190_195_groupi_g40555(csa_tree_add_190_195_groupi_n_8434 ,csa_tree_add_190_195_groupi_n_7844 ,csa_tree_add_190_195_groupi_n_8124);
  or csa_tree_add_190_195_groupi_g40556(csa_tree_add_190_195_groupi_n_8433 ,csa_tree_add_190_195_groupi_n_6530 ,csa_tree_add_190_195_groupi_n_8224);
  nor csa_tree_add_190_195_groupi_g40557(csa_tree_add_190_195_groupi_n_8432 ,csa_tree_add_190_195_groupi_n_6221 ,csa_tree_add_190_195_groupi_n_8047);
  or csa_tree_add_190_195_groupi_g40558(csa_tree_add_190_195_groupi_n_8431 ,csa_tree_add_190_195_groupi_n_8225 ,csa_tree_add_190_195_groupi_n_7763);
  or csa_tree_add_190_195_groupi_g40559(csa_tree_add_190_195_groupi_n_8430 ,csa_tree_add_190_195_groupi_n_4663 ,csa_tree_add_190_195_groupi_n_8007);
  or csa_tree_add_190_195_groupi_g40560(csa_tree_add_190_195_groupi_n_8429 ,csa_tree_add_190_195_groupi_n_7407 ,csa_tree_add_190_195_groupi_n_8165);
  or csa_tree_add_190_195_groupi_g40561(csa_tree_add_190_195_groupi_n_8428 ,csa_tree_add_190_195_groupi_n_5796 ,csa_tree_add_190_195_groupi_n_8226);
  nor csa_tree_add_190_195_groupi_g40562(csa_tree_add_190_195_groupi_n_8427 ,csa_tree_add_190_195_groupi_n_5963 ,csa_tree_add_190_195_groupi_n_8201);
  or csa_tree_add_190_195_groupi_g40563(csa_tree_add_190_195_groupi_n_8426 ,csa_tree_add_190_195_groupi_n_7751 ,csa_tree_add_190_195_groupi_n_8059);
  or csa_tree_add_190_195_groupi_g40564(csa_tree_add_190_195_groupi_n_8425 ,csa_tree_add_190_195_groupi_n_5964 ,csa_tree_add_190_195_groupi_n_8200);
  nor csa_tree_add_190_195_groupi_g40565(csa_tree_add_190_195_groupi_n_8424 ,csa_tree_add_190_195_groupi_n_7414 ,csa_tree_add_190_195_groupi_n_8109);
  or csa_tree_add_190_195_groupi_g40566(csa_tree_add_190_195_groupi_n_8423 ,csa_tree_add_190_195_groupi_n_7663 ,csa_tree_add_190_195_groupi_n_8104);
  nor csa_tree_add_190_195_groupi_g40567(csa_tree_add_190_195_groupi_n_8422 ,csa_tree_add_190_195_groupi_n_5439 ,csa_tree_add_190_195_groupi_n_8002);
  or csa_tree_add_190_195_groupi_g40568(csa_tree_add_190_195_groupi_n_8421 ,csa_tree_add_190_195_groupi_n_7417 ,csa_tree_add_190_195_groupi_n_8152);
  and csa_tree_add_190_195_groupi_g40569(csa_tree_add_190_195_groupi_n_8420 ,csa_tree_add_190_195_groupi_n_5817 ,csa_tree_add_190_195_groupi_n_8227);
  and csa_tree_add_190_195_groupi_g40570(csa_tree_add_190_195_groupi_n_8419 ,csa_tree_add_190_195_groupi_n_7862 ,csa_tree_add_190_195_groupi_n_8103);
  nor csa_tree_add_190_195_groupi_g40571(csa_tree_add_190_195_groupi_n_8418 ,csa_tree_add_190_195_groupi_n_5073 ,csa_tree_add_190_195_groupi_n_8189);
  and csa_tree_add_190_195_groupi_g40572(csa_tree_add_190_195_groupi_n_8417 ,csa_tree_add_190_195_groupi_n_6993 ,csa_tree_add_190_195_groupi_n_8100);
  or csa_tree_add_190_195_groupi_g40573(csa_tree_add_190_195_groupi_n_8416 ,csa_tree_add_190_195_groupi_n_6171 ,csa_tree_add_190_195_groupi_n_8041);
  or csa_tree_add_190_195_groupi_g40574(csa_tree_add_190_195_groupi_n_8415 ,csa_tree_add_190_195_groupi_n_8229 ,csa_tree_add_190_195_groupi_n_8096);
  or csa_tree_add_190_195_groupi_g40575(csa_tree_add_190_195_groupi_n_8414 ,csa_tree_add_190_195_groupi_n_7397 ,csa_tree_add_190_195_groupi_n_8123);
  and csa_tree_add_190_195_groupi_g40576(csa_tree_add_190_195_groupi_n_8413 ,csa_tree_add_190_195_groupi_n_6330 ,csa_tree_add_190_195_groupi_n_8054);
  or csa_tree_add_190_195_groupi_g40577(csa_tree_add_190_195_groupi_n_8412 ,csa_tree_add_190_195_groupi_n_64 ,csa_tree_add_190_195_groupi_n_8001);
  or csa_tree_add_190_195_groupi_g40578(csa_tree_add_190_195_groupi_n_8411 ,csa_tree_add_190_195_groupi_n_6979 ,csa_tree_add_190_195_groupi_n_8146);
  or csa_tree_add_190_195_groupi_g40579(csa_tree_add_190_195_groupi_n_8410 ,csa_tree_add_190_195_groupi_n_7855 ,csa_tree_add_190_195_groupi_n_8113);
  and csa_tree_add_190_195_groupi_g40580(csa_tree_add_190_195_groupi_n_8409 ,csa_tree_add_190_195_groupi_n_8090 ,csa_tree_add_190_195_groupi_n_8053);
  nor csa_tree_add_190_195_groupi_g40581(csa_tree_add_190_195_groupi_n_8408 ,csa_tree_add_190_195_groupi_n_7213 ,csa_tree_add_190_195_groupi_n_8105);
  nor csa_tree_add_190_195_groupi_g40582(csa_tree_add_190_195_groupi_n_8407 ,csa_tree_add_190_195_groupi_n_7222 ,csa_tree_add_190_195_groupi_n_8081);
  or csa_tree_add_190_195_groupi_g40583(csa_tree_add_190_195_groupi_n_8406 ,csa_tree_add_190_195_groupi_n_7403 ,csa_tree_add_190_195_groupi_n_8074);
  nor csa_tree_add_190_195_groupi_g40584(csa_tree_add_190_195_groupi_n_8405 ,csa_tree_add_190_195_groupi_n_5685 ,csa_tree_add_190_195_groupi_n_8230);
  or csa_tree_add_190_195_groupi_g40585(csa_tree_add_190_195_groupi_n_8404 ,csa_tree_add_190_195_groupi_n_7404 ,csa_tree_add_190_195_groupi_n_8069);
  and csa_tree_add_190_195_groupi_g40586(csa_tree_add_190_195_groupi_n_8403 ,csa_tree_add_190_195_groupi_n_5073 ,csa_tree_add_190_195_groupi_n_8189);
  nor csa_tree_add_190_195_groupi_g40587(csa_tree_add_190_195_groupi_n_8402 ,csa_tree_add_190_195_groupi_n_5041 ,csa_tree_add_190_195_groupi_n_8204);
  or csa_tree_add_190_195_groupi_g40588(csa_tree_add_190_195_groupi_n_8401 ,csa_tree_add_190_195_groupi_n_7253 ,csa_tree_add_190_195_groupi_n_8232);
  or csa_tree_add_190_195_groupi_g40589(csa_tree_add_190_195_groupi_n_8400 ,csa_tree_add_190_195_groupi_n_5040 ,csa_tree_add_190_195_groupi_n_8205);
  or csa_tree_add_190_195_groupi_g40590(csa_tree_add_190_195_groupi_n_8399 ,csa_tree_add_190_195_groupi_n_7722 ,csa_tree_add_190_195_groupi_n_8042);
  or csa_tree_add_190_195_groupi_g40591(csa_tree_add_190_195_groupi_n_8398 ,csa_tree_add_190_195_groupi_n_7651 ,csa_tree_add_190_195_groupi_n_8102);
  nor csa_tree_add_190_195_groupi_g40592(csa_tree_add_190_195_groupi_n_8397 ,csa_tree_add_190_195_groupi_n_8188 ,csa_tree_add_190_195_groupi_n_7525);
  and csa_tree_add_190_195_groupi_g40593(csa_tree_add_190_195_groupi_n_8396 ,csa_tree_add_190_195_groupi_n_8188 ,csa_tree_add_190_195_groupi_n_7525);
  or csa_tree_add_190_195_groupi_g40594(csa_tree_add_190_195_groupi_n_8545 ,csa_tree_add_190_195_groupi_n_7690 ,csa_tree_add_190_195_groupi_n_7973);
  or csa_tree_add_190_195_groupi_g40595(csa_tree_add_190_195_groupi_n_8544 ,csa_tree_add_190_195_groupi_n_6222 ,csa_tree_add_190_195_groupi_n_8063);
  and csa_tree_add_190_195_groupi_g40596(csa_tree_add_190_195_groupi_n_8543 ,csa_tree_add_190_195_groupi_n_3349 ,csa_tree_add_190_195_groupi_n_8086);
  and csa_tree_add_190_195_groupi_g40597(csa_tree_add_190_195_groupi_n_8542 ,csa_tree_add_190_195_groupi_n_6545 ,csa_tree_add_190_195_groupi_n_8178);
  or csa_tree_add_190_195_groupi_g40598(csa_tree_add_190_195_groupi_n_8541 ,csa_tree_add_190_195_groupi_n_3452 ,csa_tree_add_190_195_groupi_n_8065);
  and csa_tree_add_190_195_groupi_g40599(csa_tree_add_190_195_groupi_n_8540 ,csa_tree_add_190_195_groupi_n_5829 ,csa_tree_add_190_195_groupi_n_8174);
  or csa_tree_add_190_195_groupi_g40600(csa_tree_add_190_195_groupi_n_8538 ,csa_tree_add_190_195_groupi_n_5689 ,csa_tree_add_190_195_groupi_n_8115);
  or csa_tree_add_190_195_groupi_g40601(csa_tree_add_190_195_groupi_n_8537 ,csa_tree_add_190_195_groupi_n_7783 ,csa_tree_add_190_195_groupi_n_7969);
  and csa_tree_add_190_195_groupi_g40602(csa_tree_add_190_195_groupi_n_8536 ,csa_tree_add_190_195_groupi_n_7768 ,csa_tree_add_190_195_groupi_n_8083);
  or csa_tree_add_190_195_groupi_g40603(csa_tree_add_190_195_groupi_n_8535 ,csa_tree_add_190_195_groupi_n_3403 ,csa_tree_add_190_195_groupi_n_8169);
  and csa_tree_add_190_195_groupi_g40604(csa_tree_add_190_195_groupi_n_8534 ,csa_tree_add_190_195_groupi_n_7804 ,csa_tree_add_190_195_groupi_n_8164);
  or csa_tree_add_190_195_groupi_g40605(csa_tree_add_190_195_groupi_n_8533 ,csa_tree_add_190_195_groupi_n_7711 ,csa_tree_add_190_195_groupi_n_8118);
  and csa_tree_add_190_195_groupi_g40606(csa_tree_add_190_195_groupi_n_8532 ,csa_tree_add_190_195_groupi_n_7801 ,csa_tree_add_190_195_groupi_n_8163);
  or csa_tree_add_190_195_groupi_g40607(csa_tree_add_190_195_groupi_n_8531 ,csa_tree_add_190_195_groupi_n_7739 ,csa_tree_add_190_195_groupi_n_8092);
  and csa_tree_add_190_195_groupi_g40608(csa_tree_add_190_195_groupi_n_8530 ,csa_tree_add_190_195_groupi_n_6830 ,csa_tree_add_190_195_groupi_n_8093);
  and csa_tree_add_190_195_groupi_g40609(csa_tree_add_190_195_groupi_n_8529 ,csa_tree_add_190_195_groupi_n_7491 ,csa_tree_add_190_195_groupi_n_8182);
  and csa_tree_add_190_195_groupi_g40610(csa_tree_add_190_195_groupi_n_8528 ,csa_tree_add_190_195_groupi_n_7744 ,csa_tree_add_190_195_groupi_n_8085);
  or csa_tree_add_190_195_groupi_g40611(csa_tree_add_190_195_groupi_n_8526 ,csa_tree_add_190_195_groupi_n_6843 ,csa_tree_add_190_195_groupi_n_8107);
  and csa_tree_add_190_195_groupi_g40612(csa_tree_add_190_195_groupi_n_8525 ,csa_tree_add_190_195_groupi_n_3618 ,csa_tree_add_190_195_groupi_n_8161);
  or csa_tree_add_190_195_groupi_g40613(csa_tree_add_190_195_groupi_n_8524 ,csa_tree_add_190_195_groupi_n_7758 ,csa_tree_add_190_195_groupi_n_8116);
  or csa_tree_add_190_195_groupi_g40614(csa_tree_add_190_195_groupi_n_8523 ,csa_tree_add_190_195_groupi_n_2891 ,csa_tree_add_190_195_groupi_n_8155);
  and csa_tree_add_190_195_groupi_g40615(csa_tree_add_190_195_groupi_n_8522 ,csa_tree_add_190_195_groupi_n_7695 ,csa_tree_add_190_195_groupi_n_8181);
  or csa_tree_add_190_195_groupi_g40616(csa_tree_add_190_195_groupi_n_8521 ,csa_tree_add_190_195_groupi_n_7761 ,csa_tree_add_190_195_groupi_n_8119);
  or csa_tree_add_190_195_groupi_g40617(csa_tree_add_190_195_groupi_n_8519 ,csa_tree_add_190_195_groupi_n_6103 ,csa_tree_add_190_195_groupi_n_7970);
  and csa_tree_add_190_195_groupi_g40618(csa_tree_add_190_195_groupi_n_8518 ,csa_tree_add_190_195_groupi_n_5747 ,csa_tree_add_190_195_groupi_n_8120);
  and csa_tree_add_190_195_groupi_g40619(csa_tree_add_190_195_groupi_n_8517 ,csa_tree_add_190_195_groupi_n_7697 ,csa_tree_add_190_195_groupi_n_8166);
  and csa_tree_add_190_195_groupi_g40620(csa_tree_add_190_195_groupi_n_8516 ,csa_tree_add_190_195_groupi_n_6397 ,csa_tree_add_190_195_groupi_n_8127);
  and csa_tree_add_190_195_groupi_g40621(csa_tree_add_190_195_groupi_n_8515 ,csa_tree_add_190_195_groupi_n_7777 ,csa_tree_add_190_195_groupi_n_8066);
  and csa_tree_add_190_195_groupi_g40622(csa_tree_add_190_195_groupi_n_8514 ,csa_tree_add_190_195_groupi_n_7049 ,csa_tree_add_190_195_groupi_n_8129);
  or csa_tree_add_190_195_groupi_g40623(csa_tree_add_190_195_groupi_n_8513 ,csa_tree_add_190_195_groupi_n_6736 ,csa_tree_add_190_195_groupi_n_8117);
  and csa_tree_add_190_195_groupi_g40624(csa_tree_add_190_195_groupi_n_8512 ,csa_tree_add_190_195_groupi_n_3627 ,csa_tree_add_190_195_groupi_n_8136);
  and csa_tree_add_190_195_groupi_g40625(csa_tree_add_190_195_groupi_n_8511 ,csa_tree_add_190_195_groupi_n_6475 ,csa_tree_add_190_195_groupi_n_8148);
  and csa_tree_add_190_195_groupi_g40626(csa_tree_add_190_195_groupi_n_8510 ,csa_tree_add_190_195_groupi_n_7708 ,csa_tree_add_190_195_groupi_n_8061);
  and csa_tree_add_190_195_groupi_g40627(csa_tree_add_190_195_groupi_n_8509 ,csa_tree_add_190_195_groupi_n_7725 ,csa_tree_add_190_195_groupi_n_8071);
  and csa_tree_add_190_195_groupi_g40628(csa_tree_add_190_195_groupi_n_8508 ,csa_tree_add_190_195_groupi_n_7781 ,csa_tree_add_190_195_groupi_n_8138);
  and csa_tree_add_190_195_groupi_g40629(csa_tree_add_190_195_groupi_n_8507 ,csa_tree_add_190_195_groupi_n_7284 ,csa_tree_add_190_195_groupi_n_8140);
  and csa_tree_add_190_195_groupi_g40630(csa_tree_add_190_195_groupi_n_8506 ,csa_tree_add_190_195_groupi_n_7743 ,csa_tree_add_190_195_groupi_n_8095);
  and csa_tree_add_190_195_groupi_g40631(csa_tree_add_190_195_groupi_n_8505 ,csa_tree_add_190_195_groupi_n_7785 ,csa_tree_add_190_195_groupi_n_8150);
  and csa_tree_add_190_195_groupi_g40632(csa_tree_add_190_195_groupi_n_8504 ,csa_tree_add_190_195_groupi_n_7792 ,csa_tree_add_190_195_groupi_n_8151);
  and csa_tree_add_190_195_groupi_g40633(csa_tree_add_190_195_groupi_n_8502 ,csa_tree_add_190_195_groupi_n_7057 ,csa_tree_add_190_195_groupi_n_7971);
  or csa_tree_add_190_195_groupi_g40634(csa_tree_add_190_195_groupi_n_8500 ,csa_tree_add_190_195_groupi_n_6239 ,csa_tree_add_190_195_groupi_n_8170);
  or csa_tree_add_190_195_groupi_g40635(csa_tree_add_190_195_groupi_n_8499 ,csa_tree_add_190_195_groupi_n_7794 ,csa_tree_add_190_195_groupi_n_8156);
  or csa_tree_add_190_195_groupi_g40636(csa_tree_add_190_195_groupi_n_8497 ,csa_tree_add_190_195_groupi_n_7694 ,csa_tree_add_190_195_groupi_n_8183);
  and csa_tree_add_190_195_groupi_g40637(csa_tree_add_190_195_groupi_n_8496 ,csa_tree_add_190_195_groupi_n_6382 ,csa_tree_add_190_195_groupi_n_8162);
  and csa_tree_add_190_195_groupi_g40638(csa_tree_add_190_195_groupi_n_8493 ,csa_tree_add_190_195_groupi_n_7238 ,csa_tree_add_190_195_groupi_n_8101);
  or csa_tree_add_190_195_groupi_g40639(csa_tree_add_190_195_groupi_n_8492 ,csa_tree_add_190_195_groupi_n_6170 ,csa_tree_add_190_195_groupi_n_8184);
  or csa_tree_add_190_195_groupi_g40640(csa_tree_add_190_195_groupi_n_8490 ,csa_tree_add_190_195_groupi_n_7800 ,csa_tree_add_190_195_groupi_n_8070);
  or csa_tree_add_190_195_groupi_g40641(csa_tree_add_190_195_groupi_n_8489 ,csa_tree_add_190_195_groupi_n_7481 ,csa_tree_add_190_195_groupi_n_8121);
  or csa_tree_add_190_195_groupi_g40642(csa_tree_add_190_195_groupi_n_8488 ,csa_tree_add_190_195_groupi_n_7719 ,csa_tree_add_190_195_groupi_n_8084);
  and csa_tree_add_190_195_groupi_g40643(csa_tree_add_190_195_groupi_n_8486 ,csa_tree_add_190_195_groupi_n_5816 ,csa_tree_add_190_195_groupi_n_8167);
  or csa_tree_add_190_195_groupi_g40644(csa_tree_add_190_195_groupi_n_8484 ,csa_tree_add_190_195_groupi_n_7298 ,csa_tree_add_190_195_groupi_n_8172);
  or csa_tree_add_190_195_groupi_g40645(csa_tree_add_190_195_groupi_n_8483 ,csa_tree_add_190_195_groupi_n_7718 ,csa_tree_add_190_195_groupi_n_8080);
  or csa_tree_add_190_195_groupi_g40646(csa_tree_add_190_195_groupi_n_8481 ,csa_tree_add_190_195_groupi_n_7728 ,csa_tree_add_190_195_groupi_n_8073);
  and csa_tree_add_190_195_groupi_g40647(csa_tree_add_190_195_groupi_n_8479 ,csa_tree_add_190_195_groupi_n_7710 ,csa_tree_add_190_195_groupi_n_8062);
  not csa_tree_add_190_195_groupi_g40649(csa_tree_add_190_195_groupi_n_8381 ,csa_tree_add_190_195_groupi_n_8380);
  not csa_tree_add_190_195_groupi_g40651(csa_tree_add_190_195_groupi_n_8377 ,csa_tree_add_190_195_groupi_n_8376);
  not csa_tree_add_190_195_groupi_g40652(csa_tree_add_190_195_groupi_n_8375 ,csa_tree_add_190_195_groupi_n_8374);
  not csa_tree_add_190_195_groupi_g40653(csa_tree_add_190_195_groupi_n_8372 ,csa_tree_add_190_195_groupi_n_8371);
  not csa_tree_add_190_195_groupi_g40654(csa_tree_add_190_195_groupi_n_8369 ,csa_tree_add_190_195_groupi_n_8368);
  not csa_tree_add_190_195_groupi_g40655(csa_tree_add_190_195_groupi_n_8366 ,csa_tree_add_190_195_groupi_n_8365);
  not csa_tree_add_190_195_groupi_g40656(csa_tree_add_190_195_groupi_n_8364 ,csa_tree_add_190_195_groupi_n_8363);
  not csa_tree_add_190_195_groupi_g40657(csa_tree_add_190_195_groupi_n_8360 ,csa_tree_add_190_195_groupi_n_8361);
  not csa_tree_add_190_195_groupi_g40658(csa_tree_add_190_195_groupi_n_8359 ,csa_tree_add_190_195_groupi_n_8358);
  not csa_tree_add_190_195_groupi_g40659(csa_tree_add_190_195_groupi_n_8357 ,csa_tree_add_190_195_groupi_n_8356);
  not csa_tree_add_190_195_groupi_g40660(csa_tree_add_190_195_groupi_n_8354 ,csa_tree_add_190_195_groupi_n_8353);
  not csa_tree_add_190_195_groupi_g40661(csa_tree_add_190_195_groupi_n_8352 ,csa_tree_add_190_195_groupi_n_8351);
  not csa_tree_add_190_195_groupi_g40662(csa_tree_add_190_195_groupi_n_8349 ,csa_tree_add_190_195_groupi_n_8350);
  not csa_tree_add_190_195_groupi_g40663(csa_tree_add_190_195_groupi_n_8348 ,csa_tree_add_190_195_groupi_n_8347);
  not csa_tree_add_190_195_groupi_g40664(csa_tree_add_190_195_groupi_n_8345 ,csa_tree_add_190_195_groupi_n_8346);
  not csa_tree_add_190_195_groupi_g40665(csa_tree_add_190_195_groupi_n_8344 ,csa_tree_add_190_195_groupi_n_8343);
  not csa_tree_add_190_195_groupi_g40666(csa_tree_add_190_195_groupi_n_8342 ,csa_tree_add_190_195_groupi_n_8341);
  not csa_tree_add_190_195_groupi_g40667(csa_tree_add_190_195_groupi_n_8337 ,csa_tree_add_190_195_groupi_n_8338);
  not csa_tree_add_190_195_groupi_g40668(csa_tree_add_190_195_groupi_n_8335 ,csa_tree_add_190_195_groupi_n_8336);
  not csa_tree_add_190_195_groupi_g40669(csa_tree_add_190_195_groupi_n_8333 ,csa_tree_add_190_195_groupi_n_8334);
  not csa_tree_add_190_195_groupi_g40670(csa_tree_add_190_195_groupi_n_8332 ,csa_tree_add_190_195_groupi_n_8331);
  not csa_tree_add_190_195_groupi_g40671(csa_tree_add_190_195_groupi_n_8329 ,csa_tree_add_190_195_groupi_n_8328);
  not csa_tree_add_190_195_groupi_g40672(csa_tree_add_190_195_groupi_n_8327 ,csa_tree_add_190_195_groupi_n_8326);
  not csa_tree_add_190_195_groupi_g40673(csa_tree_add_190_195_groupi_n_8324 ,csa_tree_add_190_195_groupi_n_8325);
  not csa_tree_add_190_195_groupi_g40674(csa_tree_add_190_195_groupi_n_8322 ,csa_tree_add_190_195_groupi_n_8323);
  not csa_tree_add_190_195_groupi_g40675(csa_tree_add_190_195_groupi_n_8319 ,csa_tree_add_190_195_groupi_n_8318);
  not csa_tree_add_190_195_groupi_g40676(csa_tree_add_190_195_groupi_n_8317 ,csa_tree_add_190_195_groupi_n_8316);
  not csa_tree_add_190_195_groupi_g40677(csa_tree_add_190_195_groupi_n_8313 ,csa_tree_add_190_195_groupi_n_8314);
  or csa_tree_add_190_195_groupi_g40678(csa_tree_add_190_195_groupi_n_8312 ,csa_tree_add_190_195_groupi_n_8020 ,csa_tree_add_190_195_groupi_n_8197);
  or csa_tree_add_190_195_groupi_g40679(csa_tree_add_190_195_groupi_n_8311 ,csa_tree_add_190_195_groupi_n_6877 ,csa_tree_add_190_195_groupi_n_8220);
  or csa_tree_add_190_195_groupi_g40680(csa_tree_add_190_195_groupi_n_8310 ,csa_tree_add_190_195_groupi_n_7387 ,csa_tree_add_190_195_groupi_n_8168);
  and csa_tree_add_190_195_groupi_g40681(csa_tree_add_190_195_groupi_n_8309 ,csa_tree_add_190_195_groupi_n_6310 ,csa_tree_add_190_195_groupi_n_8043);
  nor csa_tree_add_190_195_groupi_g40682(csa_tree_add_190_195_groupi_n_8308 ,csa_tree_add_190_195_groupi_n_7599 ,csa_tree_add_190_195_groupi_n_8196);
  and csa_tree_add_190_195_groupi_g40683(csa_tree_add_190_195_groupi_n_8307 ,csa_tree_add_190_195_groupi_n_7599 ,csa_tree_add_190_195_groupi_n_8196);
  or csa_tree_add_190_195_groupi_g40684(csa_tree_add_190_195_groupi_n_8306 ,csa_tree_add_190_195_groupi_n_7670 ,csa_tree_add_190_195_groupi_n_7960);
  or csa_tree_add_190_195_groupi_g40685(csa_tree_add_190_195_groupi_n_8305 ,csa_tree_add_190_195_groupi_n_7578 ,csa_tree_add_190_195_groupi_n_8008);
  nor csa_tree_add_190_195_groupi_g40686(csa_tree_add_190_195_groupi_n_8304 ,csa_tree_add_190_195_groupi_n_7577 ,csa_tree_add_190_195_groupi_n_8009);
  or csa_tree_add_190_195_groupi_g40688(csa_tree_add_190_195_groupi_n_8303 ,csa_tree_add_190_195_groupi_n_5808 ,csa_tree_add_190_195_groupi_n_8217);
  or csa_tree_add_190_195_groupi_g40689(csa_tree_add_190_195_groupi_n_8302 ,csa_tree_add_190_195_groupi_n_7502 ,csa_tree_add_190_195_groupi_n_8014);
  nor csa_tree_add_190_195_groupi_g40690(csa_tree_add_190_195_groupi_n_8301 ,csa_tree_add_190_195_groupi_n_7501 ,csa_tree_add_190_195_groupi_n_8015);
  and csa_tree_add_190_195_groupi_g40691(csa_tree_add_190_195_groupi_n_8300 ,csa_tree_add_190_195_groupi_n_8231 ,csa_tree_add_190_195_groupi_n_8108);
  or csa_tree_add_190_195_groupi_g40692(csa_tree_add_190_195_groupi_n_8299 ,csa_tree_add_190_195_groupi_n_7580 ,csa_tree_add_190_195_groupi_n_7986);
  and csa_tree_add_190_195_groupi_g40693(csa_tree_add_190_195_groupi_n_8298 ,csa_tree_add_190_195_groupi_n_8020 ,csa_tree_add_190_195_groupi_n_8197);
  nor csa_tree_add_190_195_groupi_g40694(csa_tree_add_190_195_groupi_n_8297 ,csa_tree_add_190_195_groupi_n_7579 ,csa_tree_add_190_195_groupi_n_7987);
  nor csa_tree_add_190_195_groupi_g40695(csa_tree_add_190_195_groupi_n_8296 ,csa_tree_add_190_195_groupi_n_8186 ,csa_tree_add_190_195_groupi_n_8190);
  or csa_tree_add_190_195_groupi_g40696(csa_tree_add_190_195_groupi_n_8295 ,csa_tree_add_190_195_groupi_n_8185 ,csa_tree_add_190_195_groupi_n_8191);
  or csa_tree_add_190_195_groupi_g40697(csa_tree_add_190_195_groupi_n_8294 ,csa_tree_add_190_195_groupi_n_8023 ,csa_tree_add_190_195_groupi_n_8028);
  or csa_tree_add_190_195_groupi_g40698(csa_tree_add_190_195_groupi_n_8293 ,csa_tree_add_190_195_groupi_n_93 ,csa_tree_add_190_195_groupi_n_8039);
  or csa_tree_add_190_195_groupi_g40699(csa_tree_add_190_195_groupi_n_8292 ,csa_tree_add_190_195_groupi_n_7422 ,csa_tree_add_190_195_groupi_n_8072);
  nor csa_tree_add_190_195_groupi_g40700(csa_tree_add_190_195_groupi_n_8291 ,csa_tree_add_190_195_groupi_n_8022 ,csa_tree_add_190_195_groupi_n_8029);
  or csa_tree_add_190_195_groupi_g40701(csa_tree_add_190_195_groupi_n_8290 ,csa_tree_add_190_195_groupi_n_6188 ,csa_tree_add_190_195_groupi_n_8058);
  and csa_tree_add_190_195_groupi_g40702(csa_tree_add_190_195_groupi_n_8289 ,csa_tree_add_190_195_groupi_n_5815 ,csa_tree_add_190_195_groupi_n_8035);
  or csa_tree_add_190_195_groupi_g40703(csa_tree_add_190_195_groupi_n_8288 ,csa_tree_add_190_195_groupi_n_7102 ,csa_tree_add_190_195_groupi_n_8018);
  xnor csa_tree_add_190_195_groupi_g40704(csa_tree_add_190_195_groupi_n_8287 ,csa_tree_add_190_195_groupi_n_4676 ,csa_tree_add_190_195_groupi_n_7870);
  xnor csa_tree_add_190_195_groupi_g40705(csa_tree_add_190_195_groupi_n_8286 ,csa_tree_add_190_195_groupi_n_5474 ,csa_tree_add_190_195_groupi_n_7661);
  xnor csa_tree_add_190_195_groupi_g40706(csa_tree_add_190_195_groupi_n_8285 ,csa_tree_add_190_195_groupi_n_7666 ,csa_tree_add_190_195_groupi_n_1676);
  xnor csa_tree_add_190_195_groupi_g40707(csa_tree_add_190_195_groupi_n_8284 ,csa_tree_add_190_195_groupi_n_4603 ,csa_tree_add_190_195_groupi_n_7859);
  xnor csa_tree_add_190_195_groupi_g40708(csa_tree_add_190_195_groupi_n_8283 ,csa_tree_add_190_195_groupi_n_7869 ,csa_tree_add_190_195_groupi_n_5335);
  xnor csa_tree_add_190_195_groupi_g40709(csa_tree_add_190_195_groupi_n_8282 ,csa_tree_add_190_195_groupi_n_7672 ,csa_tree_add_190_195_groupi_n_753);
  xor csa_tree_add_190_195_groupi_g40710(csa_tree_add_190_195_groupi_n_8281 ,csa_tree_add_190_195_groupi_n_7868 ,csa_tree_add_190_195_groupi_n_7836);
  xnor csa_tree_add_190_195_groupi_g40711(csa_tree_add_190_195_groupi_n_8280 ,csa_tree_add_190_195_groupi_n_7653 ,csa_tree_add_190_195_groupi_n_1789);
  xnor csa_tree_add_190_195_groupi_g40712(csa_tree_add_190_195_groupi_n_8279 ,csa_tree_add_190_195_groupi_n_7649 ,csa_tree_add_190_195_groupi_n_6763);
  xnor csa_tree_add_190_195_groupi_g40713(csa_tree_add_190_195_groupi_n_8278 ,csa_tree_add_190_195_groupi_n_5331 ,csa_tree_add_190_195_groupi_n_7652);
  xnor csa_tree_add_190_195_groupi_g40714(csa_tree_add_190_195_groupi_n_8277 ,csa_tree_add_190_195_groupi_n_7564 ,csa_tree_add_190_195_groupi_n_7844);
  xnor csa_tree_add_190_195_groupi_g40715(csa_tree_add_190_195_groupi_n_8276 ,csa_tree_add_190_195_groupi_n_4599 ,csa_tree_add_190_195_groupi_n_7676);
  xnor csa_tree_add_190_195_groupi_g40716(csa_tree_add_190_195_groupi_n_8275 ,csa_tree_add_190_195_groupi_n_7671 ,csa_tree_add_190_195_groupi_n_1804);
  xnor csa_tree_add_190_195_groupi_g40717(csa_tree_add_190_195_groupi_n_8274 ,csa_tree_add_190_195_groupi_n_4 ,csa_tree_add_190_195_groupi_n_1859);
  xnor csa_tree_add_190_195_groupi_g40718(csa_tree_add_190_195_groupi_n_8273 ,csa_tree_add_190_195_groupi_n_5915 ,csa_tree_add_190_195_groupi_n_43);
  xnor csa_tree_add_190_195_groupi_g40719(csa_tree_add_190_195_groupi_n_8272 ,csa_tree_add_190_195_groupi_n_4706 ,csa_tree_add_190_195_groupi_n_7849);
  xnor csa_tree_add_190_195_groupi_g40720(csa_tree_add_190_195_groupi_n_8271 ,csa_tree_add_190_195_groupi_n_7146 ,csa_tree_add_190_195_groupi_n_7531);
  xnor csa_tree_add_190_195_groupi_g40721(csa_tree_add_190_195_groupi_n_8270 ,csa_tree_add_190_195_groupi_n_7663 ,csa_tree_add_190_195_groupi_n_4931);
  xnor csa_tree_add_190_195_groupi_g40722(csa_tree_add_190_195_groupi_n_8269 ,csa_tree_add_190_195_groupi_n_7628 ,csa_tree_add_190_195_groupi_n_7567);
  xnor csa_tree_add_190_195_groupi_g40723(csa_tree_add_190_195_groupi_n_8268 ,csa_tree_add_190_195_groupi_n_4570 ,csa_tree_add_190_195_groupi_n_7650);
  xnor csa_tree_add_190_195_groupi_g40724(csa_tree_add_190_195_groupi_n_8267 ,csa_tree_add_190_195_groupi_n_7158 ,csa_tree_add_190_195_groupi_n_7527);
  xnor csa_tree_add_190_195_groupi_g40725(csa_tree_add_190_195_groupi_n_8266 ,csa_tree_add_190_195_groupi_n_7310 ,csa_tree_add_190_195_groupi_n_7621);
  xnor csa_tree_add_190_195_groupi_g40726(csa_tree_add_190_195_groupi_n_8265 ,csa_tree_add_190_195_groupi_n_7609 ,csa_tree_add_190_195_groupi_n_7407);
  xnor csa_tree_add_190_195_groupi_g40727(csa_tree_add_190_195_groupi_n_8264 ,csa_tree_add_190_195_groupi_n_7403 ,csa_tree_add_190_195_groupi_n_7587);
  xnor csa_tree_add_190_195_groupi_g40728(csa_tree_add_190_195_groupi_n_8263 ,csa_tree_add_190_195_groupi_n_7364 ,csa_tree_add_190_195_groupi_n_7667);
  xnor csa_tree_add_190_195_groupi_g40729(csa_tree_add_190_195_groupi_n_8262 ,csa_tree_add_190_195_groupi_n_7170 ,csa_tree_add_190_195_groupi_n_7524);
  xnor csa_tree_add_190_195_groupi_g40730(csa_tree_add_190_195_groupi_n_8261 ,csa_tree_add_190_195_groupi_n_4780 ,csa_tree_add_190_195_groupi_n_7873);
  xnor csa_tree_add_190_195_groupi_g40731(csa_tree_add_190_195_groupi_n_8260 ,csa_tree_add_190_195_groupi_n_7397 ,csa_tree_add_190_195_groupi_n_7635);
  xnor csa_tree_add_190_195_groupi_g40733(csa_tree_add_190_195_groupi_n_8259 ,csa_tree_add_190_195_groupi_n_7855 ,csa_tree_add_190_195_groupi_n_7183);
  xnor csa_tree_add_190_195_groupi_g40734(csa_tree_add_190_195_groupi_n_8258 ,csa_tree_add_190_195_groupi_n_7319 ,csa_tree_add_190_195_groupi_n_7831);
  xnor csa_tree_add_190_195_groupi_g40735(csa_tree_add_190_195_groupi_n_8257 ,csa_tree_add_190_195_groupi_n_6571 ,csa_tree_add_190_195_groupi_n_7847);
  xnor csa_tree_add_190_195_groupi_g40736(csa_tree_add_190_195_groupi_n_8256 ,csa_tree_add_190_195_groupi_n_7325 ,csa_tree_add_190_195_groupi_n_7875);
  xnor csa_tree_add_190_195_groupi_g40737(csa_tree_add_190_195_groupi_n_8255 ,csa_tree_add_190_195_groupi_n_7610 ,csa_tree_add_190_195_groupi_n_7877);
  xnor csa_tree_add_190_195_groupi_g40738(csa_tree_add_190_195_groupi_n_8254 ,csa_tree_add_190_195_groupi_n_7647 ,csa_tree_add_190_195_groupi_n_4752);
  xnor csa_tree_add_190_195_groupi_g40739(csa_tree_add_190_195_groupi_n_8253 ,csa_tree_add_190_195_groupi_n_7846 ,csa_tree_add_190_195_groupi_n_74);
  xnor csa_tree_add_190_195_groupi_g40741(csa_tree_add_190_195_groupi_n_8252 ,csa_tree_add_190_195_groupi_n_6993 ,csa_tree_add_190_195_groupi_n_7541);
  xnor csa_tree_add_190_195_groupi_g40742(csa_tree_add_190_195_groupi_n_8251 ,csa_tree_add_190_195_groupi_n_7532 ,csa_tree_add_190_195_groupi_n_7147);
  xnor csa_tree_add_190_195_groupi_g40743(csa_tree_add_190_195_groupi_n_8250 ,csa_tree_add_190_195_groupi_n_7529 ,csa_tree_add_190_195_groupi_n_7655);
  xnor csa_tree_add_190_195_groupi_g40744(csa_tree_add_190_195_groupi_n_8249 ,csa_tree_add_190_195_groupi_n_6923 ,csa_tree_add_190_195_groupi_n_7604);
  xnor csa_tree_add_190_195_groupi_g40745(csa_tree_add_190_195_groupi_n_8248 ,csa_tree_add_190_195_groupi_n_4759 ,csa_tree_add_190_195_groupi_n_7866);
  xnor csa_tree_add_190_195_groupi_g40746(csa_tree_add_190_195_groupi_n_8247 ,csa_tree_add_190_195_groupi_n_53 ,csa_tree_add_190_195_groupi_n_7606);
  xnor csa_tree_add_190_195_groupi_g40747(csa_tree_add_190_195_groupi_n_8246 ,csa_tree_add_190_195_groupi_n_7537 ,csa_tree_add_190_195_groupi_n_6979);
  xnor csa_tree_add_190_195_groupi_g40748(csa_tree_add_190_195_groupi_n_8245 ,csa_tree_add_190_195_groupi_n_7087 ,csa_tree_add_190_195_groupi_n_7544);
  xnor csa_tree_add_190_195_groupi_g40749(csa_tree_add_190_195_groupi_n_8244 ,csa_tree_add_190_195_groupi_n_7633 ,csa_tree_add_190_195_groupi_n_7540);
  xnor csa_tree_add_190_195_groupi_g40750(csa_tree_add_190_195_groupi_n_8243 ,csa_tree_add_190_195_groupi_n_4946 ,csa_tree_add_190_195_groupi_n_7871);
  xnor csa_tree_add_190_195_groupi_g40751(csa_tree_add_190_195_groupi_n_8242 ,csa_tree_add_190_195_groupi_n_7388 ,csa_tree_add_190_195_groupi_n_7821);
  xnor csa_tree_add_190_195_groupi_g40752(csa_tree_add_190_195_groupi_n_8241 ,csa_tree_add_190_195_groupi_n_4906 ,csa_tree_add_190_195_groupi_n_7674);
  xnor csa_tree_add_190_195_groupi_g40753(csa_tree_add_190_195_groupi_n_8240 ,csa_tree_add_190_195_groupi_n_6911 ,csa_tree_add_190_195_groupi_n_7669);
  xnor csa_tree_add_190_195_groupi_g40754(csa_tree_add_190_195_groupi_n_8239 ,csa_tree_add_190_195_groupi_n_7344 ,csa_tree_add_190_195_groupi_n_7644);
  xnor csa_tree_add_190_195_groupi_g40755(csa_tree_add_190_195_groupi_n_8238 ,csa_tree_add_190_195_groupi_n_4724 ,csa_tree_add_190_195_groupi_n_7851);
  xnor csa_tree_add_190_195_groupi_g40756(csa_tree_add_190_195_groupi_n_8237 ,csa_tree_add_190_195_groupi_n_7212 ,csa_tree_add_190_195_groupi_n_7557);
  xnor csa_tree_add_190_195_groupi_g40757(csa_tree_add_190_195_groupi_n_8236 ,csa_tree_add_190_195_groupi_n_7648 ,csa_tree_add_190_195_groupi_n_1226);
  xor csa_tree_add_190_195_groupi_g40758(csa_tree_add_190_195_groupi_n_8235 ,csa_tree_add_190_195_groupi_n_7573 ,csa_tree_add_190_195_groupi_n_6791);
  and csa_tree_add_190_195_groupi_g40759(csa_tree_add_190_195_groupi_n_8395 ,csa_tree_add_190_195_groupi_n_7479 ,csa_tree_add_190_195_groupi_n_7964);
  xnor csa_tree_add_190_195_groupi_g40760(csa_tree_add_190_195_groupi_n_8394 ,csa_tree_add_190_195_groupi_n_5005 ,csa_tree_add_190_195_groupi_n_7454);
  xnor csa_tree_add_190_195_groupi_g40761(csa_tree_add_190_195_groupi_n_8393 ,csa_tree_add_190_195_groupi_n_4657 ,csa_tree_add_190_195_groupi_n_7433);
  xnor csa_tree_add_190_195_groupi_g40762(csa_tree_add_190_195_groupi_n_8392 ,csa_tree_add_190_195_groupi_n_5043 ,csa_tree_add_190_195_groupi_n_7455);
  or csa_tree_add_190_195_groupi_g40763(csa_tree_add_190_195_groupi_n_8391 ,csa_tree_add_190_195_groupi_n_6160 ,csa_tree_add_190_195_groupi_n_7963);
  and csa_tree_add_190_195_groupi_g40764(csa_tree_add_190_195_groupi_n_8390 ,csa_tree_add_190_195_groupi_n_7753 ,csa_tree_add_190_195_groupi_n_7953);
  and csa_tree_add_190_195_groupi_g40765(csa_tree_add_190_195_groupi_n_8389 ,csa_tree_add_190_195_groupi_n_5699 ,csa_tree_add_190_195_groupi_n_7950);
  xnor csa_tree_add_190_195_groupi_g40766(csa_tree_add_190_195_groupi_n_8388 ,csa_tree_add_190_195_groupi_n_4671 ,csa_tree_add_190_195_groupi_n_7435);
  xnor csa_tree_add_190_195_groupi_g40767(csa_tree_add_190_195_groupi_n_8387 ,csa_tree_add_190_195_groupi_n_5482 ,csa_tree_add_190_195_groupi_n_7473);
  xnor csa_tree_add_190_195_groupi_g40768(csa_tree_add_190_195_groupi_n_8386 ,csa_tree_add_190_195_groupi_n_5227 ,csa_tree_add_190_195_groupi_n_7472);
  xnor csa_tree_add_190_195_groupi_g40769(csa_tree_add_190_195_groupi_n_8385 ,csa_tree_add_190_195_groupi_n_7406 ,csa_tree_add_190_195_groupi_n_7459);
  xnor csa_tree_add_190_195_groupi_g40770(csa_tree_add_190_195_groupi_n_8384 ,csa_tree_add_190_195_groupi_n_7443 ,csa_tree_add_190_195_groupi_n_1093);
  xnor csa_tree_add_190_195_groupi_g40772(csa_tree_add_190_195_groupi_n_8383 ,csa_tree_add_190_195_groupi_n_7662 ,csa_tree_add_190_195_groupi_n_3956);
  xnor csa_tree_add_190_195_groupi_g40773(csa_tree_add_190_195_groupi_n_8382 ,csa_tree_add_190_195_groupi_n_5034 ,csa_tree_add_190_195_groupi_n_7445);
  xnor csa_tree_add_190_195_groupi_g40774(csa_tree_add_190_195_groupi_n_8380 ,csa_tree_add_190_195_groupi_n_7463 ,csa_tree_add_190_195_groupi_n_1033);
  xnor csa_tree_add_190_195_groupi_g40775(csa_tree_add_190_195_groupi_n_8379 ,csa_tree_add_190_195_groupi_n_7449 ,csa_tree_add_190_195_groupi_n_900);
  xnor csa_tree_add_190_195_groupi_g40776(csa_tree_add_190_195_groupi_n_8378 ,csa_tree_add_190_195_groupi_n_7675 ,csa_tree_add_190_195_groupi_n_7019);
  xnor csa_tree_add_190_195_groupi_g40777(csa_tree_add_190_195_groupi_n_8376 ,csa_tree_add_190_195_groupi_n_4627 ,csa_tree_add_190_195_groupi_n_7440);
  xnor csa_tree_add_190_195_groupi_g40778(csa_tree_add_190_195_groupi_n_8374 ,csa_tree_add_190_195_groupi_n_4612 ,csa_tree_add_190_195_groupi_n_7465);
  xnor csa_tree_add_190_195_groupi_g40779(csa_tree_add_190_195_groupi_n_8373 ,csa_tree_add_190_195_groupi_n_5216 ,csa_tree_add_190_195_groupi_n_7466);
  xnor csa_tree_add_190_195_groupi_g40780(csa_tree_add_190_195_groupi_n_8371 ,csa_tree_add_190_195_groupi_n_7216 ,csa_tree_add_190_195_groupi_n_7468);
  xnor csa_tree_add_190_195_groupi_g40781(csa_tree_add_190_195_groupi_n_8370 ,csa_tree_add_190_195_groupi_n_5458 ,csa_tree_add_190_195_groupi_n_7438);
  xnor csa_tree_add_190_195_groupi_g40782(csa_tree_add_190_195_groupi_n_8368 ,csa_tree_add_190_195_groupi_n_7845 ,csa_tree_add_190_195_groupi_n_6070);
  xnor csa_tree_add_190_195_groupi_g40783(csa_tree_add_190_195_groupi_n_8367 ,csa_tree_add_190_195_groupi_n_4992 ,csa_tree_add_190_195_groupi_n_7446);
  xnor csa_tree_add_190_195_groupi_g40784(csa_tree_add_190_195_groupi_n_8365 ,csa_tree_add_190_195_groupi_n_4718 ,csa_tree_add_190_195_groupi_n_7469);
  xnor csa_tree_add_190_195_groupi_g40785(csa_tree_add_190_195_groupi_n_8363 ,csa_tree_add_190_195_groupi_n_7470 ,csa_tree_add_190_195_groupi_n_1775);
  xnor csa_tree_add_190_195_groupi_g40786(csa_tree_add_190_195_groupi_n_8362 ,csa_tree_add_190_195_groupi_n_100 ,csa_tree_add_190_195_groupi_n_1116);
  xnor csa_tree_add_190_195_groupi_g40787(csa_tree_add_190_195_groupi_n_8361 ,csa_tree_add_190_195_groupi_n_5323 ,csa_tree_add_190_195_groupi_n_7471);
  xnor csa_tree_add_190_195_groupi_g40788(csa_tree_add_190_195_groupi_n_8358 ,csa_tree_add_190_195_groupi_n_5485 ,csa_tree_add_190_195_groupi_n_7441);
  xnor csa_tree_add_190_195_groupi_g40789(csa_tree_add_190_195_groupi_n_8356 ,csa_tree_add_190_195_groupi_n_6963 ,csa_tree_add_190_195_groupi_n_7448);
  xnor csa_tree_add_190_195_groupi_g40790(csa_tree_add_190_195_groupi_n_8355 ,csa_tree_add_190_195_groupi_n_7395 ,csa_tree_add_190_195_groupi_n_7434);
  xnor csa_tree_add_190_195_groupi_g40791(csa_tree_add_190_195_groupi_n_8353 ,csa_tree_add_190_195_groupi_n_5094 ,csa_tree_add_190_195_groupi_n_7447);
  xnor csa_tree_add_190_195_groupi_g40792(csa_tree_add_190_195_groupi_n_8351 ,csa_tree_add_190_195_groupi_n_78 ,csa_tree_add_190_195_groupi_n_7439);
  xnor csa_tree_add_190_195_groupi_g40793(csa_tree_add_190_195_groupi_n_8350 ,csa_tree_add_190_195_groupi_n_7658 ,csa_tree_add_190_195_groupi_n_7444);
  xnor csa_tree_add_190_195_groupi_g40794(csa_tree_add_190_195_groupi_n_8347 ,csa_tree_add_190_195_groupi_n_7450 ,csa_tree_add_190_195_groupi_n_1746);
  xnor csa_tree_add_190_195_groupi_g40795(csa_tree_add_190_195_groupi_n_8346 ,csa_tree_add_190_195_groupi_n_5441 ,csa_tree_add_190_195_groupi_n_7442);
  xnor csa_tree_add_190_195_groupi_g40796(csa_tree_add_190_195_groupi_n_8343 ,csa_tree_add_190_195_groupi_n_6947 ,csa_tree_add_190_195_groupi_n_7451);
  xnor csa_tree_add_190_195_groupi_g40797(csa_tree_add_190_195_groupi_n_8341 ,csa_tree_add_190_195_groupi_n_7228 ,csa_tree_add_190_195_groupi_n_7464);
  xnor csa_tree_add_190_195_groupi_g40798(csa_tree_add_190_195_groupi_n_8340 ,csa_tree_add_190_195_groupi_n_6938 ,csa_tree_add_190_195_groupi_n_7456);
  xnor csa_tree_add_190_195_groupi_g40799(csa_tree_add_190_195_groupi_n_8339 ,csa_tree_add_190_195_groupi_n_7673 ,csa_tree_add_190_195_groupi_n_6696);
  xnor csa_tree_add_190_195_groupi_g40800(csa_tree_add_190_195_groupi_n_8338 ,csa_tree_add_190_195_groupi_n_7474 ,csa_tree_add_190_195_groupi_n_2002);
  xnor csa_tree_add_190_195_groupi_g40801(csa_tree_add_190_195_groupi_n_8336 ,csa_tree_add_190_195_groupi_n_7664 ,csa_tree_add_190_195_groupi_n_6609);
  xnor csa_tree_add_190_195_groupi_g40802(csa_tree_add_190_195_groupi_n_8334 ,csa_tree_add_190_195_groupi_n_7654 ,csa_tree_add_190_195_groupi_n_4010);
  and csa_tree_add_190_195_groupi_g40803(csa_tree_add_190_195_groupi_n_8331 ,csa_tree_add_190_195_groupi_n_7684 ,csa_tree_add_190_195_groupi_n_7946);
  xnor csa_tree_add_190_195_groupi_g40804(csa_tree_add_190_195_groupi_n_8330 ,csa_tree_add_190_195_groupi_n_5311 ,csa_tree_add_190_195_groupi_n_7462);
  or csa_tree_add_190_195_groupi_g40805(csa_tree_add_190_195_groupi_n_8328 ,csa_tree_add_190_195_groupi_n_5736 ,csa_tree_add_190_195_groupi_n_7961);
  or csa_tree_add_190_195_groupi_g40806(csa_tree_add_190_195_groupi_n_8326 ,csa_tree_add_190_195_groupi_n_6315 ,csa_tree_add_190_195_groupi_n_7948);
  xnor csa_tree_add_190_195_groupi_g40807(csa_tree_add_190_195_groupi_n_8325 ,csa_tree_add_190_195_groupi_n_5414 ,csa_tree_add_190_195_groupi_n_7437);
  xnor csa_tree_add_190_195_groupi_g40808(csa_tree_add_190_195_groupi_n_8323 ,csa_tree_add_190_195_groupi_n_5183 ,csa_tree_add_190_195_groupi_n_7436);
  xnor csa_tree_add_190_195_groupi_g40809(csa_tree_add_190_195_groupi_n_8321 ,csa_tree_add_190_195_groupi_n_4907 ,csa_tree_add_190_195_groupi_n_7458);
  xnor csa_tree_add_190_195_groupi_g40810(csa_tree_add_190_195_groupi_n_8320 ,csa_tree_add_190_195_groupi_n_5885 ,csa_tree_add_190_195_groupi_n_7432);
  xnor csa_tree_add_190_195_groupi_g40811(csa_tree_add_190_195_groupi_n_8318 ,csa_tree_add_190_195_groupi_n_5051 ,csa_tree_add_190_195_groupi_n_7457);
  xnor csa_tree_add_190_195_groupi_g40812(csa_tree_add_190_195_groupi_n_8316 ,csa_tree_add_190_195_groupi_n_7659 ,csa_tree_add_190_195_groupi_n_7452);
  xnor csa_tree_add_190_195_groupi_g40813(csa_tree_add_190_195_groupi_n_8315 ,csa_tree_add_190_195_groupi_n_4971 ,csa_tree_add_190_195_groupi_n_7453);
  or csa_tree_add_190_195_groupi_g40814(csa_tree_add_190_195_groupi_n_8314 ,csa_tree_add_190_195_groupi_n_5983 ,csa_tree_add_190_195_groupi_n_8234);
  not csa_tree_add_190_195_groupi_g40816(csa_tree_add_190_195_groupi_n_8229 ,csa_tree_add_190_195_groupi_n_8228);
  not csa_tree_add_190_195_groupi_g40818(csa_tree_add_190_195_groupi_n_8217 ,csa_tree_add_190_195_groupi_n_8216);
  not csa_tree_add_190_195_groupi_g40819(csa_tree_add_190_195_groupi_n_8214 ,csa_tree_add_190_195_groupi_n_8213);
  not csa_tree_add_190_195_groupi_g40820(csa_tree_add_190_195_groupi_n_8212 ,csa_tree_add_190_195_groupi_n_8211);
  not csa_tree_add_190_195_groupi_g40823(csa_tree_add_190_195_groupi_n_8206 ,csa_tree_add_190_195_groupi_n_8207);
  not csa_tree_add_190_195_groupi_g40824(csa_tree_add_190_195_groupi_n_8205 ,csa_tree_add_190_195_groupi_n_8204);
  not csa_tree_add_190_195_groupi_g40825(csa_tree_add_190_195_groupi_n_8203 ,csa_tree_add_190_195_groupi_n_8202);
  not csa_tree_add_190_195_groupi_g40826(csa_tree_add_190_195_groupi_n_8200 ,csa_tree_add_190_195_groupi_n_8201);
  not csa_tree_add_190_195_groupi_g40827(csa_tree_add_190_195_groupi_n_8198 ,csa_tree_add_190_195_groupi_n_8199);
  not csa_tree_add_190_195_groupi_g40828(csa_tree_add_190_195_groupi_n_8195 ,csa_tree_add_190_195_groupi_n_8194);
  not csa_tree_add_190_195_groupi_g40829(csa_tree_add_190_195_groupi_n_8193 ,csa_tree_add_190_195_groupi_n_8192);
  not csa_tree_add_190_195_groupi_g40830(csa_tree_add_190_195_groupi_n_8191 ,csa_tree_add_190_195_groupi_n_8190);
  not csa_tree_add_190_195_groupi_g40831(csa_tree_add_190_195_groupi_n_8188 ,csa_tree_add_190_195_groupi_n_8187);
  not csa_tree_add_190_195_groupi_g40832(csa_tree_add_190_195_groupi_n_8185 ,csa_tree_add_190_195_groupi_n_8186);
  and csa_tree_add_190_195_groupi_g40833(csa_tree_add_190_195_groupi_n_8184 ,csa_tree_add_190_195_groupi_n_6148 ,csa_tree_add_190_195_groupi_n_7870);
  and csa_tree_add_190_195_groupi_g40834(csa_tree_add_190_195_groupi_n_8183 ,csa_tree_add_190_195_groupi_n_7411 ,csa_tree_add_190_195_groupi_n_7806);
  or csa_tree_add_190_195_groupi_g40835(csa_tree_add_190_195_groupi_n_8182 ,csa_tree_add_190_195_groupi_n_7413 ,csa_tree_add_190_195_groupi_n_7490);
  or csa_tree_add_190_195_groupi_g40836(csa_tree_add_190_195_groupi_n_8181 ,csa_tree_add_190_195_groupi_n_7390 ,csa_tree_add_190_195_groupi_n_7791);
  nor csa_tree_add_190_195_groupi_g40837(csa_tree_add_190_195_groupi_n_8180 ,csa_tree_add_190_195_groupi_n_7827 ,csa_tree_add_190_195_groupi_n_7837);
  nor csa_tree_add_190_195_groupi_g40838(csa_tree_add_190_195_groupi_n_8179 ,csa_tree_add_190_195_groupi_n_7607 ,csa_tree_add_190_195_groupi_n_7638);
  or csa_tree_add_190_195_groupi_g40839(csa_tree_add_190_195_groupi_n_8178 ,csa_tree_add_190_195_groupi_n_6543 ,csa_tree_add_190_195_groupi_n_7867);
  nor csa_tree_add_190_195_groupi_g40840(csa_tree_add_190_195_groupi_n_8177 ,csa_tree_add_190_195_groupi_n_7362 ,csa_tree_add_190_195_groupi_n_7575);
  or csa_tree_add_190_195_groupi_g40841(csa_tree_add_190_195_groupi_n_8176 ,csa_tree_add_190_195_groupi_n_7145 ,csa_tree_add_190_195_groupi_n_7531);
  or csa_tree_add_190_195_groupi_g40842(csa_tree_add_190_195_groupi_n_8175 ,csa_tree_add_190_195_groupi_n_7361 ,csa_tree_add_190_195_groupi_n_7576);
  or csa_tree_add_190_195_groupi_g40843(csa_tree_add_190_195_groupi_n_8174 ,csa_tree_add_190_195_groupi_n_5827 ,csa_tree_add_190_195_groupi_n_7871);
  nor csa_tree_add_190_195_groupi_g40844(csa_tree_add_190_195_groupi_n_8173 ,csa_tree_add_190_195_groupi_n_7573 ,csa_tree_add_190_195_groupi_n_7571);
  and csa_tree_add_190_195_groupi_g40845(csa_tree_add_190_195_groupi_n_8172 ,csa_tree_add_190_195_groupi_n_7296 ,csa_tree_add_190_195_groupi_n_7672);
  or csa_tree_add_190_195_groupi_g40846(csa_tree_add_190_195_groupi_n_8171 ,csa_tree_add_190_195_groupi_n_7572 ,csa_tree_add_190_195_groupi_n_7570);
  nor csa_tree_add_190_195_groupi_g40847(csa_tree_add_190_195_groupi_n_8170 ,csa_tree_add_190_195_groupi_n_6444 ,csa_tree_add_190_195_groupi_n_7650);
  and csa_tree_add_190_195_groupi_g40848(csa_tree_add_190_195_groupi_n_8169 ,csa_tree_add_190_195_groupi_n_3424 ,csa_tree_add_190_195_groupi_n_7671);
  nor csa_tree_add_190_195_groupi_g40849(csa_tree_add_190_195_groupi_n_8168 ,csa_tree_add_190_195_groupi_n_7158 ,csa_tree_add_190_195_groupi_n_7526);
  or csa_tree_add_190_195_groupi_g40850(csa_tree_add_190_195_groupi_n_8167 ,csa_tree_add_190_195_groupi_n_5760 ,csa_tree_add_190_195_groupi_n_7852);
  or csa_tree_add_190_195_groupi_g40851(csa_tree_add_190_195_groupi_n_8166 ,csa_tree_add_190_195_groupi_n_7778 ,csa_tree_add_190_195_groupi_n_7876);
  and csa_tree_add_190_195_groupi_g40852(csa_tree_add_190_195_groupi_n_8165 ,csa_tree_add_190_195_groupi_n_7068 ,csa_tree_add_190_195_groupi_n_7609);
  or csa_tree_add_190_195_groupi_g40853(csa_tree_add_190_195_groupi_n_8164 ,csa_tree_add_190_195_groupi_n_7196 ,csa_tree_add_190_195_groupi_n_7802);
  or csa_tree_add_190_195_groupi_g40854(csa_tree_add_190_195_groupi_n_8163 ,csa_tree_add_190_195_groupi_n_7872 ,csa_tree_add_190_195_groupi_n_7799);
  or csa_tree_add_190_195_groupi_g40855(csa_tree_add_190_195_groupi_n_8162 ,csa_tree_add_190_195_groupi_n_6500 ,csa_tree_add_190_195_groupi_n_7869);
  or csa_tree_add_190_195_groupi_g40856(csa_tree_add_190_195_groupi_n_8161 ,csa_tree_add_190_195_groupi_n_3616 ,csa_tree_add_190_195_groupi_n_7648);
  or csa_tree_add_190_195_groupi_g40857(csa_tree_add_190_195_groupi_n_8160 ,csa_tree_add_190_195_groupi_n_7068 ,csa_tree_add_190_195_groupi_n_7609);
  or csa_tree_add_190_195_groupi_g40858(csa_tree_add_190_195_groupi_n_8159 ,csa_tree_add_190_195_groupi_n_7335 ,csa_tree_add_190_195_groupi_n_7642);
  or csa_tree_add_190_195_groupi_g40859(csa_tree_add_190_195_groupi_n_8158 ,csa_tree_add_190_195_groupi_n_7157 ,csa_tree_add_190_195_groupi_n_7527);
  or csa_tree_add_190_195_groupi_g40860(csa_tree_add_190_195_groupi_n_8157 ,csa_tree_add_190_195_groupi_n_7821 ,csa_tree_add_190_195_groupi_n_7822);
  and csa_tree_add_190_195_groupi_g40861(csa_tree_add_190_195_groupi_n_8156 ,csa_tree_add_190_195_groupi_n_7793 ,csa_tree_add_190_195_groupi_n_7666);
  and csa_tree_add_190_195_groupi_g40862(csa_tree_add_190_195_groupi_n_8155 ,csa_tree_add_190_195_groupi_n_3171 ,csa_tree_add_190_195_groupi_n_4);
  nor csa_tree_add_190_195_groupi_g40863(csa_tree_add_190_195_groupi_n_8154 ,csa_tree_add_190_195_groupi_n_7820 ,csa_tree_add_190_195_groupi_n_7823);
  or csa_tree_add_190_195_groupi_g40864(csa_tree_add_190_195_groupi_n_8153 ,csa_tree_add_190_195_groupi_n_7346 ,csa_tree_add_190_195_groupi_n_7586);
  and csa_tree_add_190_195_groupi_g40865(csa_tree_add_190_195_groupi_n_8152 ,csa_tree_add_190_195_groupi_n_7190 ,csa_tree_add_190_195_groupi_n_7513);
  or csa_tree_add_190_195_groupi_g40866(csa_tree_add_190_195_groupi_n_8151 ,csa_tree_add_190_195_groupi_n_7865 ,csa_tree_add_190_195_groupi_n_7786);
  or csa_tree_add_190_195_groupi_g40867(csa_tree_add_190_195_groupi_n_8150 ,csa_tree_add_190_195_groupi_n_7427 ,csa_tree_add_190_195_groupi_n_7774);
  or csa_tree_add_190_195_groupi_g40868(csa_tree_add_190_195_groupi_n_8149 ,csa_tree_add_190_195_groupi_n_5913 ,csa_tree_add_190_195_groupi_n_7605);
  or csa_tree_add_190_195_groupi_g40869(csa_tree_add_190_195_groupi_n_8148 ,csa_tree_add_190_195_groupi_n_6474 ,csa_tree_add_190_195_groupi_n_43);
  nor csa_tree_add_190_195_groupi_g40870(csa_tree_add_190_195_groupi_n_8147 ,csa_tree_add_190_195_groupi_n_53 ,csa_tree_add_190_195_groupi_n_7606);
  and csa_tree_add_190_195_groupi_g40871(csa_tree_add_190_195_groupi_n_8146 ,csa_tree_add_190_195_groupi_n_7537 ,csa_tree_add_190_195_groupi_n_7536);
  and csa_tree_add_190_195_groupi_g40872(csa_tree_add_190_195_groupi_n_8145 ,csa_tree_add_190_195_groupi_n_7607 ,csa_tree_add_190_195_groupi_n_7638);
  or csa_tree_add_190_195_groupi_g40873(csa_tree_add_190_195_groupi_n_8144 ,csa_tree_add_190_195_groupi_n_7190 ,csa_tree_add_190_195_groupi_n_7513);
  or csa_tree_add_190_195_groupi_g40874(csa_tree_add_190_195_groupi_n_8143 ,csa_tree_add_190_195_groupi_n_7338 ,csa_tree_add_190_195_groupi_n_7625);
  nor csa_tree_add_190_195_groupi_g40875(csa_tree_add_190_195_groupi_n_8142 ,csa_tree_add_190_195_groupi_n_7560 ,csa_tree_add_190_195_groupi_n_7595);
  or csa_tree_add_190_195_groupi_g40876(csa_tree_add_190_195_groupi_n_8141 ,csa_tree_add_190_195_groupi_n_7559 ,csa_tree_add_190_195_groupi_n_7596);
  or csa_tree_add_190_195_groupi_g40877(csa_tree_add_190_195_groupi_n_8140 ,csa_tree_add_190_195_groupi_n_7283 ,csa_tree_add_190_195_groupi_n_7659);
  nor csa_tree_add_190_195_groupi_g40878(csa_tree_add_190_195_groupi_n_8139 ,csa_tree_add_190_195_groupi_n_6265 ,csa_tree_add_190_195_groupi_n_7615);
  or csa_tree_add_190_195_groupi_g40879(csa_tree_add_190_195_groupi_n_8138 ,csa_tree_add_190_195_groupi_n_7780 ,csa_tree_add_190_195_groupi_n_7209);
  nor csa_tree_add_190_195_groupi_g40880(csa_tree_add_190_195_groupi_n_8137 ,csa_tree_add_190_195_groupi_n_4788 ,csa_tree_add_190_195_groupi_n_7841);
  or csa_tree_add_190_195_groupi_g40881(csa_tree_add_190_195_groupi_n_8136 ,csa_tree_add_190_195_groupi_n_3659 ,csa_tree_add_190_195_groupi_n_7662);
  nor csa_tree_add_190_195_groupi_g40882(csa_tree_add_190_195_groupi_n_8135 ,csa_tree_add_190_195_groupi_n_7359 ,csa_tree_add_190_195_groupi_n_7555);
  nor csa_tree_add_190_195_groupi_g40883(csa_tree_add_190_195_groupi_n_8134 ,csa_tree_add_190_195_groupi_n_7493 ,csa_tree_add_190_195_groupi_n_7557);
  nor csa_tree_add_190_195_groupi_g40884(csa_tree_add_190_195_groupi_n_8133 ,csa_tree_add_190_195_groupi_n_7337 ,csa_tree_add_190_195_groupi_n_7626);
  or csa_tree_add_190_195_groupi_g40885(csa_tree_add_190_195_groupi_n_8132 ,csa_tree_add_190_195_groupi_n_7494 ,csa_tree_add_190_195_groupi_n_7556);
  or csa_tree_add_190_195_groupi_g40886(csa_tree_add_190_195_groupi_n_8131 ,csa_tree_add_190_195_groupi_n_7349 ,csa_tree_add_190_195_groupi_n_7553);
  or csa_tree_add_190_195_groupi_g40887(csa_tree_add_190_195_groupi_n_8130 ,csa_tree_add_190_195_groupi_n_7360 ,csa_tree_add_190_195_groupi_n_7554);
  or csa_tree_add_190_195_groupi_g40888(csa_tree_add_190_195_groupi_n_8129 ,csa_tree_add_190_195_groupi_n_7050 ,csa_tree_add_190_195_groupi_n_7658);
  or csa_tree_add_190_195_groupi_g40889(csa_tree_add_190_195_groupi_n_8128 ,csa_tree_add_190_195_groupi_n_7627 ,csa_tree_add_190_195_groupi_n_7567);
  or csa_tree_add_190_195_groupi_g40890(csa_tree_add_190_195_groupi_n_8127 ,csa_tree_add_190_195_groupi_n_6240 ,csa_tree_add_190_195_groupi_n_7665);
  nor csa_tree_add_190_195_groupi_g40891(csa_tree_add_190_195_groupi_n_8126 ,csa_tree_add_190_195_groupi_n_7350 ,csa_tree_add_190_195_groupi_n_7552);
  or csa_tree_add_190_195_groupi_g40892(csa_tree_add_190_195_groupi_n_8125 ,csa_tree_add_190_195_groupi_n_6257 ,csa_tree_add_190_195_groupi_n_7563);
  nor csa_tree_add_190_195_groupi_g40893(csa_tree_add_190_195_groupi_n_8124 ,csa_tree_add_190_195_groupi_n_6256 ,csa_tree_add_190_195_groupi_n_7564);
  nor csa_tree_add_190_195_groupi_g40894(csa_tree_add_190_195_groupi_n_8123 ,csa_tree_add_190_195_groupi_n_7506 ,csa_tree_add_190_195_groupi_n_7635);
  or csa_tree_add_190_195_groupi_g40895(csa_tree_add_190_195_groupi_n_8122 ,csa_tree_add_190_195_groupi_n_7505 ,csa_tree_add_190_195_groupi_n_7634);
  and csa_tree_add_190_195_groupi_g40896(csa_tree_add_190_195_groupi_n_8121 ,csa_tree_add_190_195_groupi_n_6969 ,csa_tree_add_190_195_groupi_n_7480);
  or csa_tree_add_190_195_groupi_g40897(csa_tree_add_190_195_groupi_n_8120 ,csa_tree_add_190_195_groupi_n_5821 ,csa_tree_add_190_195_groupi_n_7874);
  nor csa_tree_add_190_195_groupi_g40898(csa_tree_add_190_195_groupi_n_8119 ,csa_tree_add_190_195_groupi_n_6976 ,csa_tree_add_190_195_groupi_n_7760);
  and csa_tree_add_190_195_groupi_g40899(csa_tree_add_190_195_groupi_n_8118 ,csa_tree_add_190_195_groupi_n_7425 ,csa_tree_add_190_195_groupi_n_7692);
  and csa_tree_add_190_195_groupi_g40900(csa_tree_add_190_195_groupi_n_8117 ,csa_tree_add_190_195_groupi_n_6735 ,csa_tree_add_190_195_groupi_n_7675);
  and csa_tree_add_190_195_groupi_g40901(csa_tree_add_190_195_groupi_n_8116 ,csa_tree_add_190_195_groupi_n_7757 ,csa_tree_add_190_195_groupi_n_7423);
  and csa_tree_add_190_195_groupi_g40902(csa_tree_add_190_195_groupi_n_8115 ,csa_tree_add_190_195_groupi_n_5717 ,csa_tree_add_190_195_groupi_n_7676);
  nor csa_tree_add_190_195_groupi_g40903(csa_tree_add_190_195_groupi_n_8114 ,csa_tree_add_190_195_groupi_n_7336 ,csa_tree_add_190_195_groupi_n_7641);
  and csa_tree_add_190_195_groupi_g40904(csa_tree_add_190_195_groupi_n_8113 ,csa_tree_add_190_195_groupi_n_7183 ,csa_tree_add_190_195_groupi_n_7518);
  and csa_tree_add_190_195_groupi_g40905(csa_tree_add_190_195_groupi_n_8112 ,csa_tree_add_190_195_groupi_n_7825 ,csa_tree_add_190_195_groupi_n_7826);
  or csa_tree_add_190_195_groupi_g40906(csa_tree_add_190_195_groupi_n_8111 ,csa_tree_add_190_195_groupi_n_4931 ,csa_tree_add_190_195_groupi_n_7547);
  or csa_tree_add_190_195_groupi_g40907(csa_tree_add_190_195_groupi_n_8110 ,csa_tree_add_190_195_groupi_n_7825 ,csa_tree_add_190_195_groupi_n_7826);
  nor csa_tree_add_190_195_groupi_g40908(csa_tree_add_190_195_groupi_n_8109 ,csa_tree_add_190_195_groupi_n_4888 ,csa_tree_add_190_195_groupi_n_7558);
  or csa_tree_add_190_195_groupi_g40909(csa_tree_add_190_195_groupi_n_8108 ,csa_tree_add_190_195_groupi_n_7332 ,csa_tree_add_190_195_groupi_n_7533);
  and csa_tree_add_190_195_groupi_g40910(csa_tree_add_190_195_groupi_n_8107 ,csa_tree_add_190_195_groupi_n_6807 ,csa_tree_add_190_195_groupi_n_7661);
  nor csa_tree_add_190_195_groupi_g40911(csa_tree_add_190_195_groupi_n_8106 ,csa_tree_add_190_195_groupi_n_7086 ,csa_tree_add_190_195_groupi_n_7544);
  and csa_tree_add_190_195_groupi_g40912(csa_tree_add_190_195_groupi_n_8105 ,csa_tree_add_190_195_groupi_n_6265 ,csa_tree_add_190_195_groupi_n_7615);
  and csa_tree_add_190_195_groupi_g40913(csa_tree_add_190_195_groupi_n_8104 ,csa_tree_add_190_195_groupi_n_4931 ,csa_tree_add_190_195_groupi_n_7547);
  or csa_tree_add_190_195_groupi_g40914(csa_tree_add_190_195_groupi_n_8103 ,csa_tree_add_190_195_groupi_n_7087 ,csa_tree_add_190_195_groupi_n_7543);
  nor csa_tree_add_190_195_groupi_g40915(csa_tree_add_190_195_groupi_n_8102 ,csa_tree_add_190_195_groupi_n_7628 ,csa_tree_add_190_195_groupi_n_7566);
  or csa_tree_add_190_195_groupi_g40916(csa_tree_add_190_195_groupi_n_8101 ,csa_tree_add_190_195_groupi_n_7056 ,csa_tree_add_190_195_groupi_n_7652);
  or csa_tree_add_190_195_groupi_g40917(csa_tree_add_190_195_groupi_n_8100 ,csa_tree_add_190_195_groupi_n_7608 ,csa_tree_add_190_195_groupi_n_7542);
  or csa_tree_add_190_195_groupi_g40918(csa_tree_add_190_195_groupi_n_8099 ,csa_tree_add_190_195_groupi_n_7540 ,csa_tree_add_190_195_groupi_n_7633);
  or csa_tree_add_190_195_groupi_g40919(csa_tree_add_190_195_groupi_n_8098 ,csa_tree_add_190_195_groupi_n_7183 ,csa_tree_add_190_195_groupi_n_7518);
  or csa_tree_add_190_195_groupi_g40920(csa_tree_add_190_195_groupi_n_8097 ,csa_tree_add_190_195_groupi_n_7354 ,csa_tree_add_190_195_groupi_n_7632);
  and csa_tree_add_190_195_groupi_g40921(csa_tree_add_190_195_groupi_n_8096 ,csa_tree_add_190_195_groupi_n_7540 ,csa_tree_add_190_195_groupi_n_7633);
  or csa_tree_add_190_195_groupi_g40922(csa_tree_add_190_195_groupi_n_8095 ,csa_tree_add_190_195_groupi_n_7232 ,csa_tree_add_190_195_groupi_n_7741);
  and csa_tree_add_190_195_groupi_g40923(csa_tree_add_190_195_groupi_n_8094 ,csa_tree_add_190_195_groupi_n_7354 ,csa_tree_add_190_195_groupi_n_7632);
  or csa_tree_add_190_195_groupi_g40924(csa_tree_add_190_195_groupi_n_8093 ,csa_tree_add_190_195_groupi_n_6829 ,csa_tree_add_190_195_groupi_n_7847);
  nor csa_tree_add_190_195_groupi_g40925(csa_tree_add_190_195_groupi_n_8092 ,csa_tree_add_190_195_groupi_n_6590 ,csa_tree_add_190_195_groupi_n_7737);
  and csa_tree_add_190_195_groupi_g40926(csa_tree_add_190_195_groupi_n_8091 ,csa_tree_add_190_195_groupi_n_4700 ,csa_tree_add_190_195_groupi_n_7535);
  or csa_tree_add_190_195_groupi_g40927(csa_tree_add_190_195_groupi_n_8090 ,csa_tree_add_190_195_groupi_n_4700 ,csa_tree_add_190_195_groupi_n_7535);
  or csa_tree_add_190_195_groupi_g40928(csa_tree_add_190_195_groupi_n_8089 ,csa_tree_add_190_195_groupi_n_7109 ,csa_tree_add_190_195_groupi_n_7528);
  nor csa_tree_add_190_195_groupi_g40929(csa_tree_add_190_195_groupi_n_8088 ,csa_tree_add_190_195_groupi_n_7110 ,csa_tree_add_190_195_groupi_n_7529);
  and csa_tree_add_190_195_groupi_g40930(csa_tree_add_190_195_groupi_n_8087 ,csa_tree_add_190_195_groupi_n_7152 ,csa_tree_add_190_195_groupi_n_7597);
  or csa_tree_add_190_195_groupi_g40931(csa_tree_add_190_195_groupi_n_8086 ,csa_tree_add_190_195_groupi_n_3359 ,csa_tree_add_190_195_groupi_n_7654);
  or csa_tree_add_190_195_groupi_g40932(csa_tree_add_190_195_groupi_n_8085 ,csa_tree_add_190_195_groupi_n_7854 ,csa_tree_add_190_195_groupi_n_7701);
  and csa_tree_add_190_195_groupi_g40933(csa_tree_add_190_195_groupi_n_8084 ,csa_tree_add_190_195_groupi_n_7221 ,csa_tree_add_190_195_groupi_n_7735);
  or csa_tree_add_190_195_groupi_g40934(csa_tree_add_190_195_groupi_n_8083 ,csa_tree_add_190_195_groupi_n_7226 ,csa_tree_add_190_195_groupi_n_7734);
  nor csa_tree_add_190_195_groupi_g40935(csa_tree_add_190_195_groupi_n_8082 ,csa_tree_add_190_195_groupi_n_7519 ,csa_tree_add_190_195_groupi_n_7646);
  nor csa_tree_add_190_195_groupi_g40936(csa_tree_add_190_195_groupi_n_8081 ,csa_tree_add_190_195_groupi_n_7152 ,csa_tree_add_190_195_groupi_n_7597);
  and csa_tree_add_190_195_groupi_g40937(csa_tree_add_190_195_groupi_n_8080 ,csa_tree_add_190_195_groupi_n_7850 ,csa_tree_add_190_195_groupi_n_7731);
  nor csa_tree_add_190_195_groupi_g40938(csa_tree_add_190_195_groupi_n_8079 ,csa_tree_add_190_195_groupi_n_7331 ,csa_tree_add_190_195_groupi_n_7534);
  or csa_tree_add_190_195_groupi_g40939(csa_tree_add_190_195_groupi_n_8078 ,csa_tree_add_190_195_groupi_n_7520 ,csa_tree_add_190_195_groupi_n_7645);
  or csa_tree_add_190_195_groupi_g40940(csa_tree_add_190_195_groupi_n_8077 ,csa_tree_add_190_195_groupi_n_7147 ,csa_tree_add_190_195_groupi_n_7532);
  and csa_tree_add_190_195_groupi_g40941(csa_tree_add_190_195_groupi_n_8076 ,csa_tree_add_190_195_groupi_n_7147 ,csa_tree_add_190_195_groupi_n_7532);
  or csa_tree_add_190_195_groupi_g40942(csa_tree_add_190_195_groupi_n_8075 ,csa_tree_add_190_195_groupi_n_7537 ,csa_tree_add_190_195_groupi_n_7536);
  nor csa_tree_add_190_195_groupi_g40943(csa_tree_add_190_195_groupi_n_8074 ,csa_tree_add_190_195_groupi_n_7345 ,csa_tree_add_190_195_groupi_n_7587);
  nor csa_tree_add_190_195_groupi_g40944(csa_tree_add_190_195_groupi_n_8073 ,csa_tree_add_190_195_groupi_n_7424 ,csa_tree_add_190_195_groupi_n_7797);
  nor csa_tree_add_190_195_groupi_g40945(csa_tree_add_190_195_groupi_n_8072 ,csa_tree_add_190_195_groupi_n_7146 ,csa_tree_add_190_195_groupi_n_7530);
  or csa_tree_add_190_195_groupi_g40946(csa_tree_add_190_195_groupi_n_8071 ,csa_tree_add_190_195_groupi_n_6996 ,csa_tree_add_190_195_groupi_n_7723);
  nor csa_tree_add_190_195_groupi_g40947(csa_tree_add_190_195_groupi_n_8070 ,csa_tree_add_190_195_groupi_n_7412 ,csa_tree_add_190_195_groupi_n_7776);
  nor csa_tree_add_190_195_groupi_g40948(csa_tree_add_190_195_groupi_n_8069 ,csa_tree_add_190_195_groupi_n_7181 ,csa_tree_add_190_195_groupi_n_7500);
  or csa_tree_add_190_195_groupi_g40949(csa_tree_add_190_195_groupi_n_8068 ,csa_tree_add_190_195_groupi_n_7180 ,csa_tree_add_190_195_groupi_n_7499);
  nor csa_tree_add_190_195_groupi_g40950(csa_tree_add_190_195_groupi_n_8067 ,csa_tree_add_190_195_groupi_n_7170 ,csa_tree_add_190_195_groupi_n_7523);
  or csa_tree_add_190_195_groupi_g40951(csa_tree_add_190_195_groupi_n_8066 ,csa_tree_add_190_195_groupi_n_7668 ,csa_tree_add_190_195_groupi_n_7716);
  and csa_tree_add_190_195_groupi_g40952(csa_tree_add_190_195_groupi_n_8065 ,csa_tree_add_190_195_groupi_n_3416 ,csa_tree_add_190_195_groupi_n_7653);
  or csa_tree_add_190_195_groupi_g40953(csa_tree_add_190_195_groupi_n_8064 ,csa_tree_add_190_195_groupi_n_4789 ,csa_tree_add_190_195_groupi_n_7840);
  and csa_tree_add_190_195_groupi_g40954(csa_tree_add_190_195_groupi_n_8063 ,csa_tree_add_190_195_groupi_n_6216 ,csa_tree_add_190_195_groupi_n_7674);
  or csa_tree_add_190_195_groupi_g40955(csa_tree_add_190_195_groupi_n_8062 ,csa_tree_add_190_195_groupi_n_7405 ,csa_tree_add_190_195_groupi_n_7709);
  or csa_tree_add_190_195_groupi_g40956(csa_tree_add_190_195_groupi_n_8061 ,csa_tree_add_190_195_groupi_n_6774 ,csa_tree_add_190_195_groupi_n_7707);
  or csa_tree_add_190_195_groupi_g40957(csa_tree_add_190_195_groupi_n_8060 ,csa_tree_add_190_195_groupi_n_7169 ,csa_tree_add_190_195_groupi_n_7524);
  or csa_tree_add_190_195_groupi_g40958(csa_tree_add_190_195_groupi_n_8234 ,csa_tree_add_190_195_groupi_n_7280 ,csa_tree_add_190_195_groupi_n_7811);
  and csa_tree_add_190_195_groupi_g40959(csa_tree_add_190_195_groupi_n_8233 ,csa_tree_add_190_195_groupi_n_6809 ,csa_tree_add_190_195_groupi_n_7720);
  and csa_tree_add_190_195_groupi_g40960(csa_tree_add_190_195_groupi_n_8232 ,csa_tree_add_190_195_groupi_n_3161 ,csa_tree_add_190_195_groupi_n_7727);
  or csa_tree_add_190_195_groupi_g40961(csa_tree_add_190_195_groupi_n_8231 ,csa_tree_add_190_195_groupi_n_7256 ,csa_tree_add_190_195_groupi_n_7730);
  and csa_tree_add_190_195_groupi_g40962(csa_tree_add_190_195_groupi_n_8230 ,csa_tree_add_190_195_groupi_n_2735 ,csa_tree_add_190_195_groupi_n_7733);
  or csa_tree_add_190_195_groupi_g40963(csa_tree_add_190_195_groupi_n_8228 ,csa_tree_add_190_195_groupi_n_6342 ,csa_tree_add_190_195_groupi_n_7742);
  or csa_tree_add_190_195_groupi_g40964(csa_tree_add_190_195_groupi_n_8227 ,csa_tree_add_190_195_groupi_n_2819 ,csa_tree_add_190_195_groupi_n_7712);
  and csa_tree_add_190_195_groupi_g40965(csa_tree_add_190_195_groupi_n_8226 ,csa_tree_add_190_195_groupi_n_3282 ,csa_tree_add_190_195_groupi_n_7756);
  and csa_tree_add_190_195_groupi_g40966(csa_tree_add_190_195_groupi_n_8225 ,csa_tree_add_190_195_groupi_n_5750 ,csa_tree_add_190_195_groupi_n_7764);
  and csa_tree_add_190_195_groupi_g40967(csa_tree_add_190_195_groupi_n_8224 ,csa_tree_add_190_195_groupi_n_7277 ,csa_tree_add_190_195_groupi_n_7765);
  and csa_tree_add_190_195_groupi_g40968(csa_tree_add_190_195_groupi_n_8223 ,csa_tree_add_190_195_groupi_n_6169 ,csa_tree_add_190_195_groupi_n_7698);
  and csa_tree_add_190_195_groupi_g40969(csa_tree_add_190_195_groupi_n_8222 ,csa_tree_add_190_195_groupi_n_2770 ,csa_tree_add_190_195_groupi_n_7784);
  and csa_tree_add_190_195_groupi_g40970(csa_tree_add_190_195_groupi_n_8221 ,csa_tree_add_190_195_groupi_n_7286 ,csa_tree_add_190_195_groupi_n_7787);
  and csa_tree_add_190_195_groupi_g40971(csa_tree_add_190_195_groupi_n_8220 ,csa_tree_add_190_195_groupi_n_2756 ,csa_tree_add_190_195_groupi_n_7790);
  or csa_tree_add_190_195_groupi_g40972(csa_tree_add_190_195_groupi_n_8219 ,csa_tree_add_190_195_groupi_n_6496 ,csa_tree_add_190_195_groupi_n_7798);
  and csa_tree_add_190_195_groupi_g40973(csa_tree_add_190_195_groupi_n_8218 ,csa_tree_add_190_195_groupi_n_3680 ,csa_tree_add_190_195_groupi_n_7696);
  or csa_tree_add_190_195_groupi_g40974(csa_tree_add_190_195_groupi_n_8216 ,csa_tree_add_190_195_groupi_n_2894 ,csa_tree_add_190_195_groupi_n_7803);
  or csa_tree_add_190_195_groupi_g40975(csa_tree_add_190_195_groupi_n_8215 ,csa_tree_add_190_195_groupi_n_5844 ,csa_tree_add_190_195_groupi_n_7816);
  or csa_tree_add_190_195_groupi_g40976(csa_tree_add_190_195_groupi_n_8213 ,csa_tree_add_190_195_groupi_n_7294 ,csa_tree_add_190_195_groupi_n_7807);
  or csa_tree_add_190_195_groupi_g40977(csa_tree_add_190_195_groupi_n_8211 ,csa_tree_add_190_195_groupi_n_7250 ,csa_tree_add_190_195_groupi_n_7732);
  or csa_tree_add_190_195_groupi_g40978(csa_tree_add_190_195_groupi_n_8210 ,csa_tree_add_190_195_groupi_n_6151 ,csa_tree_add_190_195_groupi_n_7706);
  and csa_tree_add_190_195_groupi_g40979(csa_tree_add_190_195_groupi_n_8209 ,csa_tree_add_190_195_groupi_n_7233 ,csa_tree_add_190_195_groupi_n_7813);
  and csa_tree_add_190_195_groupi_g40980(csa_tree_add_190_195_groupi_n_8208 ,csa_tree_add_190_195_groupi_n_7247 ,csa_tree_add_190_195_groupi_n_7715);
  or csa_tree_add_190_195_groupi_g40981(csa_tree_add_190_195_groupi_n_8207 ,csa_tree_add_190_195_groupi_n_6428 ,csa_tree_add_190_195_groupi_n_7773);
  or csa_tree_add_190_195_groupi_g40982(csa_tree_add_190_195_groupi_n_8204 ,csa_tree_add_190_195_groupi_n_6319 ,csa_tree_add_190_195_groupi_n_7746);
  and csa_tree_add_190_195_groupi_g40983(csa_tree_add_190_195_groupi_n_8202 ,csa_tree_add_190_195_groupi_n_6178 ,csa_tree_add_190_195_groupi_n_7700);
  and csa_tree_add_190_195_groupi_g40984(csa_tree_add_190_195_groupi_n_8201 ,csa_tree_add_190_195_groupi_n_6366 ,csa_tree_add_190_195_groupi_n_7749);
  and csa_tree_add_190_195_groupi_g40985(csa_tree_add_190_195_groupi_n_8199 ,csa_tree_add_190_195_groupi_n_6509 ,csa_tree_add_190_195_groupi_n_7805);
  and csa_tree_add_190_195_groupi_g40986(csa_tree_add_190_195_groupi_n_8197 ,csa_tree_add_190_195_groupi_n_6422 ,csa_tree_add_190_195_groupi_n_7770);
  and csa_tree_add_190_195_groupi_g40987(csa_tree_add_190_195_groupi_n_8196 ,csa_tree_add_190_195_groupi_n_7246 ,csa_tree_add_190_195_groupi_n_7713);
  and csa_tree_add_190_195_groupi_g40988(csa_tree_add_190_195_groupi_n_8194 ,csa_tree_add_190_195_groupi_n_6871 ,csa_tree_add_190_195_groupi_n_7754);
  and csa_tree_add_190_195_groupi_g40989(csa_tree_add_190_195_groupi_n_8192 ,csa_tree_add_190_195_groupi_n_6526 ,csa_tree_add_190_195_groupi_n_7808);
  and csa_tree_add_190_195_groupi_g40990(csa_tree_add_190_195_groupi_n_8190 ,csa_tree_add_190_195_groupi_n_5798 ,csa_tree_add_190_195_groupi_n_7755);
  and csa_tree_add_190_195_groupi_g40991(csa_tree_add_190_195_groupi_n_8189 ,csa_tree_add_190_195_groupi_n_3074 ,csa_tree_add_190_195_groupi_n_7699);
  or csa_tree_add_190_195_groupi_g40992(csa_tree_add_190_195_groupi_n_8187 ,csa_tree_add_190_195_groupi_n_6237 ,csa_tree_add_190_195_groupi_n_7717);
  and csa_tree_add_190_195_groupi_g40993(csa_tree_add_190_195_groupi_n_8186 ,csa_tree_add_190_195_groupi_n_6376 ,csa_tree_add_190_195_groupi_n_7759);
  not csa_tree_add_190_195_groupi_g40994(csa_tree_add_190_195_groupi_n_8056 ,csa_tree_add_190_195_groupi_n_8055);
  not csa_tree_add_190_195_groupi_g40995(csa_tree_add_190_195_groupi_n_8051 ,csa_tree_add_190_195_groupi_n_8050);
  not csa_tree_add_190_195_groupi_g40997(csa_tree_add_190_195_groupi_n_8045 ,csa_tree_add_190_195_groupi_n_8044);
  not csa_tree_add_190_195_groupi_g40999(csa_tree_add_190_195_groupi_n_8037 ,csa_tree_add_190_195_groupi_n_8036);
  not csa_tree_add_190_195_groupi_g41000(csa_tree_add_190_195_groupi_n_8032 ,csa_tree_add_190_195_groupi_n_8031);
  not csa_tree_add_190_195_groupi_g41001(csa_tree_add_190_195_groupi_n_8029 ,csa_tree_add_190_195_groupi_n_8028);
  not csa_tree_add_190_195_groupi_g41002(csa_tree_add_190_195_groupi_n_8027 ,csa_tree_add_190_195_groupi_n_8026);
  not csa_tree_add_190_195_groupi_g41003(csa_tree_add_190_195_groupi_n_8025 ,csa_tree_add_190_195_groupi_n_8024);
  not csa_tree_add_190_195_groupi_g41004(csa_tree_add_190_195_groupi_n_8023 ,csa_tree_add_190_195_groupi_n_8022);
  not csa_tree_add_190_195_groupi_g41005(csa_tree_add_190_195_groupi_n_8018 ,csa_tree_add_190_195_groupi_n_8019);
  not csa_tree_add_190_195_groupi_g41006(csa_tree_add_190_195_groupi_n_8017 ,csa_tree_add_190_195_groupi_n_8016);
  not csa_tree_add_190_195_groupi_g41007(csa_tree_add_190_195_groupi_n_8014 ,csa_tree_add_190_195_groupi_n_8015);
  not csa_tree_add_190_195_groupi_g41008(csa_tree_add_190_195_groupi_n_8013 ,csa_tree_add_190_195_groupi_n_8012);
  not csa_tree_add_190_195_groupi_g41009(csa_tree_add_190_195_groupi_n_8010 ,csa_tree_add_190_195_groupi_n_8011);
  not csa_tree_add_190_195_groupi_g41010(csa_tree_add_190_195_groupi_n_8009 ,csa_tree_add_190_195_groupi_n_8008);
  not csa_tree_add_190_195_groupi_g41011(csa_tree_add_190_195_groupi_n_8006 ,csa_tree_add_190_195_groupi_n_8007);
  not csa_tree_add_190_195_groupi_g41012(csa_tree_add_190_195_groupi_n_8003 ,csa_tree_add_190_195_groupi_n_8004);
  not csa_tree_add_190_195_groupi_g41013(csa_tree_add_190_195_groupi_n_8002 ,csa_tree_add_190_195_groupi_n_8001);
  not csa_tree_add_190_195_groupi_g41014(csa_tree_add_190_195_groupi_n_7999 ,csa_tree_add_190_195_groupi_n_8000);
  not csa_tree_add_190_195_groupi_g41015(csa_tree_add_190_195_groupi_n_7996 ,csa_tree_add_190_195_groupi_n_7997);
  not csa_tree_add_190_195_groupi_g41016(csa_tree_add_190_195_groupi_n_7995 ,csa_tree_add_190_195_groupi_n_7994);
  not csa_tree_add_190_195_groupi_g41017(csa_tree_add_190_195_groupi_n_7993 ,csa_tree_add_190_195_groupi_n_7992);
  not csa_tree_add_190_195_groupi_g41018(csa_tree_add_190_195_groupi_n_7990 ,csa_tree_add_190_195_groupi_n_7989);
  not csa_tree_add_190_195_groupi_g41019(csa_tree_add_190_195_groupi_n_7987 ,csa_tree_add_190_195_groupi_n_7986);
  not csa_tree_add_190_195_groupi_g41020(csa_tree_add_190_195_groupi_n_7985 ,csa_tree_add_190_195_groupi_n_7984);
  not csa_tree_add_190_195_groupi_g41021(csa_tree_add_190_195_groupi_n_7983 ,csa_tree_add_190_195_groupi_n_7982);
  and csa_tree_add_190_195_groupi_g41022(csa_tree_add_190_195_groupi_n_7978 ,csa_tree_add_190_195_groupi_n_4888 ,csa_tree_add_190_195_groupi_n_7558);
  and csa_tree_add_190_195_groupi_g41023(csa_tree_add_190_195_groupi_n_7977 ,csa_tree_add_190_195_groupi_n_7827 ,csa_tree_add_190_195_groupi_n_7837);
  or csa_tree_add_190_195_groupi_g41024(csa_tree_add_190_195_groupi_n_7976 ,csa_tree_add_190_195_groupi_n_6922 ,csa_tree_add_190_195_groupi_n_7604);
  or csa_tree_add_190_195_groupi_g41025(csa_tree_add_190_195_groupi_n_7975 ,csa_tree_add_190_195_groupi_n_7124 ,csa_tree_add_190_195_groupi_n_7838);
  nor csa_tree_add_190_195_groupi_g41026(csa_tree_add_190_195_groupi_n_7974 ,csa_tree_add_190_195_groupi_n_7125 ,csa_tree_add_190_195_groupi_n_7839);
  and csa_tree_add_190_195_groupi_g41027(csa_tree_add_190_195_groupi_n_7973 ,csa_tree_add_190_195_groupi_n_7382 ,csa_tree_add_190_195_groupi_n_7689);
  nor csa_tree_add_190_195_groupi_g41028(csa_tree_add_190_195_groupi_n_7972 ,csa_tree_add_190_195_groupi_n_6923 ,csa_tree_add_190_195_groupi_n_89);
  or csa_tree_add_190_195_groupi_g41029(csa_tree_add_190_195_groupi_n_7971 ,csa_tree_add_190_195_groupi_n_7037 ,csa_tree_add_190_195_groupi_n_7649);
  and csa_tree_add_190_195_groupi_g41030(csa_tree_add_190_195_groupi_n_7970 ,csa_tree_add_190_195_groupi_n_6101 ,csa_tree_add_190_195_groupi_n_7673);
  nor csa_tree_add_190_195_groupi_g41031(csa_tree_add_190_195_groupi_n_7969 ,csa_tree_add_190_195_groupi_n_6999 ,csa_tree_add_190_195_groupi_n_7782);
  or csa_tree_add_190_195_groupi_g41032(csa_tree_add_190_195_groupi_n_7968 ,csa_tree_add_190_195_groupi_n_7179 ,csa_tree_add_190_195_groupi_n_7583);
  and csa_tree_add_190_195_groupi_g41033(csa_tree_add_190_195_groupi_n_7967 ,csa_tree_add_190_195_groupi_n_7179 ,csa_tree_add_190_195_groupi_n_7583);
  nor csa_tree_add_190_195_groupi_g41034(csa_tree_add_190_195_groupi_n_7966 ,csa_tree_add_190_195_groupi_n_7610 ,csa_tree_add_190_195_groupi_n_7594);
  and csa_tree_add_190_195_groupi_g41035(csa_tree_add_190_195_groupi_n_7965 ,csa_tree_add_190_195_groupi_n_7610 ,csa_tree_add_190_195_groupi_n_7594);
  or csa_tree_add_190_195_groupi_g41036(csa_tree_add_190_195_groupi_n_7964 ,csa_tree_add_190_195_groupi_n_7391 ,csa_tree_add_190_195_groupi_n_7485);
  and csa_tree_add_190_195_groupi_g41037(csa_tree_add_190_195_groupi_n_7963 ,csa_tree_add_190_195_groupi_n_6299 ,csa_tree_add_190_195_groupi_n_7849);
  or csa_tree_add_190_195_groupi_g41038(csa_tree_add_190_195_groupi_n_7962 ,csa_tree_add_190_195_groupi_n_6911 ,csa_tree_add_190_195_groupi_n_7842);
  and csa_tree_add_190_195_groupi_g41039(csa_tree_add_190_195_groupi_n_7961 ,csa_tree_add_190_195_groupi_n_5669 ,csa_tree_add_190_195_groupi_n_7845);
  nor csa_tree_add_190_195_groupi_g41040(csa_tree_add_190_195_groupi_n_7960 ,csa_tree_add_190_195_groupi_n_6910 ,csa_tree_add_190_195_groupi_n_7843);
  or csa_tree_add_190_195_groupi_g41041(csa_tree_add_190_195_groupi_n_7959 ,csa_tree_add_190_195_groupi_n_7310 ,csa_tree_add_190_195_groupi_n_7620);
  or csa_tree_add_190_195_groupi_g41042(csa_tree_add_190_195_groupi_n_7958 ,csa_tree_add_190_195_groupi_n_7318 ,csa_tree_add_190_195_groupi_n_7830);
  or csa_tree_add_190_195_groupi_g41043(csa_tree_add_190_195_groupi_n_7957 ,csa_tree_add_190_195_groupi_n_7569 ,csa_tree_add_190_195_groupi_n_7511);
  nor csa_tree_add_190_195_groupi_g41044(csa_tree_add_190_195_groupi_n_7956 ,csa_tree_add_190_195_groupi_n_7568 ,csa_tree_add_190_195_groupi_n_7512);
  or csa_tree_add_190_195_groupi_g41045(csa_tree_add_190_195_groupi_n_7955 ,csa_tree_add_190_195_groupi_n_7344 ,csa_tree_add_190_195_groupi_n_7643);
  nor csa_tree_add_190_195_groupi_g41046(csa_tree_add_190_195_groupi_n_7954 ,csa_tree_add_190_195_groupi_n_7343 ,csa_tree_add_190_195_groupi_n_7644);
  or csa_tree_add_190_195_groupi_g41047(csa_tree_add_190_195_groupi_n_7953 ,csa_tree_add_190_195_groupi_n_7752 ,csa_tree_add_190_195_groupi_n_7846);
  nor csa_tree_add_190_195_groupi_g41048(csa_tree_add_190_195_groupi_n_7952 ,csa_tree_add_190_195_groupi_n_7309 ,csa_tree_add_190_195_groupi_n_7621);
  or csa_tree_add_190_195_groupi_g41049(csa_tree_add_190_195_groupi_n_7951 ,csa_tree_add_190_195_groupi_n_7347 ,csa_tree_add_190_195_groupi_n_7617);
  or csa_tree_add_190_195_groupi_g41050(csa_tree_add_190_195_groupi_n_7950 ,csa_tree_add_190_195_groupi_n_5739 ,csa_tree_add_190_195_groupi_n_7860);
  nor csa_tree_add_190_195_groupi_g41051(csa_tree_add_190_195_groupi_n_7949 ,csa_tree_add_190_195_groupi_n_7319 ,csa_tree_add_190_195_groupi_n_7831);
  nor csa_tree_add_190_195_groupi_g41052(csa_tree_add_190_195_groupi_n_7948 ,csa_tree_add_190_195_groupi_n_6227 ,csa_tree_add_190_195_groupi_n_7647);
  nor csa_tree_add_190_195_groupi_g41053(csa_tree_add_190_195_groupi_n_7947 ,csa_tree_add_190_195_groupi_n_7348 ,csa_tree_add_190_195_groupi_n_7616);
  or csa_tree_add_190_195_groupi_g41054(csa_tree_add_190_195_groupi_n_7946 ,csa_tree_add_190_195_groupi_n_7853 ,csa_tree_add_190_195_groupi_n_7682);
  and csa_tree_add_190_195_groupi_g41055(csa_tree_add_190_195_groupi_n_7945 ,csa_tree_add_190_195_groupi_n_7608 ,csa_tree_add_190_195_groupi_n_7542);
  xnor csa_tree_add_190_195_groupi_g41056(csa_tree_add_190_195_groupi_n_7944 ,csa_tree_add_190_195_groupi_n_7227 ,csa_tree_add_190_195_groupi_n_5429);
  xnor csa_tree_add_190_195_groupi_g41057(csa_tree_add_190_195_groupi_n_7943 ,csa_tree_add_190_195_groupi_n_5438 ,csa_tree_add_190_195_groupi_n_7399);
  xnor csa_tree_add_190_195_groupi_g41058(csa_tree_add_190_195_groupi_n_7942 ,csa_tree_add_190_195_groupi_n_5931 ,csa_tree_add_190_195_groupi_n_7410);
  xnor csa_tree_add_190_195_groupi_g41059(csa_tree_add_190_195_groupi_n_7941 ,csa_tree_add_190_195_groupi_n_7094 ,csa_tree_add_190_195_groupi_n_7317);
  xnor csa_tree_add_190_195_groupi_g41060(csa_tree_add_190_195_groupi_n_7940 ,csa_tree_add_190_195_groupi_n_6943 ,csa_tree_add_190_195_groupi_n_7154);
  xnor csa_tree_add_190_195_groupi_g41061(csa_tree_add_190_195_groupi_n_7939 ,csa_tree_add_190_195_groupi_n_5940 ,csa_tree_add_190_195_groupi_n_7108);
  xnor csa_tree_add_190_195_groupi_g41062(csa_tree_add_190_195_groupi_n_7938 ,csa_tree_add_190_195_groupi_n_5209 ,csa_tree_add_190_195_groupi_n_7176);
  xor csa_tree_add_190_195_groupi_g41063(csa_tree_add_190_195_groupi_n_7937 ,csa_tree_add_190_195_groupi_n_7222 ,csa_tree_add_190_195_groupi_n_7152);
  xnor csa_tree_add_190_195_groupi_g41064(csa_tree_add_190_195_groupi_n_7936 ,csa_tree_add_190_195_groupi_n_7428 ,csa_tree_add_190_195_groupi_n_1951);
  xnor csa_tree_add_190_195_groupi_g41065(csa_tree_add_190_195_groupi_n_7935 ,csa_tree_add_190_195_groupi_n_7198 ,csa_tree_add_190_195_groupi_n_5189);
  xnor csa_tree_add_190_195_groupi_g41066(csa_tree_add_190_195_groupi_n_7934 ,csa_tree_add_190_195_groupi_n_7392 ,csa_tree_add_190_195_groupi_n_2041);
  xnor csa_tree_add_190_195_groupi_g41067(csa_tree_add_190_195_groupi_n_7933 ,csa_tree_add_190_195_groupi_n_7073 ,csa_tree_add_190_195_groupi_n_52);
  xnor csa_tree_add_190_195_groupi_g41068(csa_tree_add_190_195_groupi_n_7932 ,csa_tree_add_190_195_groupi_n_7226 ,csa_tree_add_190_195_groupi_n_7);
  xnor csa_tree_add_190_195_groupi_g41069(csa_tree_add_190_195_groupi_n_7931 ,csa_tree_add_190_195_groupi_n_4922 ,csa_tree_add_190_195_groupi_n_7383);
  xnor csa_tree_add_190_195_groupi_g41070(csa_tree_add_190_195_groupi_n_7930 ,csa_tree_add_190_195_groupi_n_5883 ,csa_tree_add_190_195_groupi_n_7215);
  xnor csa_tree_add_190_195_groupi_g41071(csa_tree_add_190_195_groupi_n_7929 ,csa_tree_add_190_195_groupi_n_7213 ,csa_tree_add_190_195_groupi_n_6265);
  xnor csa_tree_add_190_195_groupi_g41072(csa_tree_add_190_195_groupi_n_7928 ,csa_tree_add_190_195_groupi_n_5531 ,csa_tree_add_190_195_groupi_n_7386);
  xnor csa_tree_add_190_195_groupi_g41073(csa_tree_add_190_195_groupi_n_7927 ,csa_tree_add_190_195_groupi_n_7140 ,csa_tree_add_190_195_groupi_n_7221);
  xnor csa_tree_add_190_195_groupi_g41074(csa_tree_add_190_195_groupi_n_7926 ,csa_tree_add_190_195_groupi_n_4897 ,csa_tree_add_190_195_groupi_n_7409);
  xnor csa_tree_add_190_195_groupi_g41075(csa_tree_add_190_195_groupi_n_7925 ,csa_tree_add_190_195_groupi_n_5526 ,csa_tree_add_190_195_groupi_n_7218);
  xnor csa_tree_add_190_195_groupi_g41076(csa_tree_add_190_195_groupi_n_7924 ,csa_tree_add_190_195_groupi_n_5928 ,csa_tree_add_190_195_groupi_n_7380);
  xnor csa_tree_add_190_195_groupi_g41077(csa_tree_add_190_195_groupi_n_7923 ,csa_tree_add_190_195_groupi_n_5404 ,csa_tree_add_190_195_groupi_n_7105);
  xnor csa_tree_add_190_195_groupi_g41078(csa_tree_add_190_195_groupi_n_7922 ,csa_tree_add_190_195_groupi_n_7382 ,csa_tree_add_190_195_groupi_n_7065);
  xnor csa_tree_add_190_195_groupi_g41079(csa_tree_add_190_195_groupi_n_7921 ,csa_tree_add_190_195_groupi_n_7400 ,csa_tree_add_190_195_groupi_n_2152);
  xnor csa_tree_add_190_195_groupi_g41080(csa_tree_add_190_195_groupi_n_7920 ,csa_tree_add_190_195_groupi_n_5953 ,csa_tree_add_190_195_groupi_n_84);
  xnor csa_tree_add_190_195_groupi_g41081(csa_tree_add_190_195_groupi_n_7919 ,csa_tree_add_190_195_groupi_n_5241 ,csa_tree_add_190_195_groupi_n_7224);
  xnor csa_tree_add_190_195_groupi_g41082(csa_tree_add_190_195_groupi_n_7918 ,csa_tree_add_190_195_groupi_n_7351 ,csa_tree_add_190_195_groupi_n_7135);
  xnor csa_tree_add_190_195_groupi_g41083(csa_tree_add_190_195_groupi_n_7917 ,csa_tree_add_190_195_groupi_n_7370 ,csa_tree_add_190_195_groupi_n_7085);
  xnor csa_tree_add_190_195_groupi_g41084(csa_tree_add_190_195_groupi_n_7916 ,csa_tree_add_190_195_groupi_n_7307 ,csa_tree_add_190_195_groupi_n_7080);
  xnor csa_tree_add_190_195_groupi_g41085(csa_tree_add_190_195_groupi_n_7915 ,csa_tree_add_190_195_groupi_n_6269 ,csa_tree_add_190_195_groupi_n_7389);
  xnor csa_tree_add_190_195_groupi_g41086(csa_tree_add_190_195_groupi_n_7914 ,csa_tree_add_190_195_groupi_n_7425 ,csa_tree_add_190_195_groupi_n_7101);
  xnor csa_tree_add_190_195_groupi_g41087(csa_tree_add_190_195_groupi_n_7913 ,csa_tree_add_190_195_groupi_n_6272 ,csa_tree_add_190_195_groupi_n_7192);
  xnor csa_tree_add_190_195_groupi_g41088(csa_tree_add_190_195_groupi_n_7912 ,csa_tree_add_190_195_groupi_n_5326 ,csa_tree_add_190_195_groupi_n_7205);
  xnor csa_tree_add_190_195_groupi_g41089(csa_tree_add_190_195_groupi_n_7911 ,csa_tree_add_190_195_groupi_n_6998 ,csa_tree_add_190_195_groupi_n_7088);
  xnor csa_tree_add_190_195_groupi_g41090(csa_tree_add_190_195_groupi_n_7910 ,csa_tree_add_190_195_groupi_n_7373 ,csa_tree_add_190_195_groupi_n_5400);
  xnor csa_tree_add_190_195_groupi_g41091(csa_tree_add_190_195_groupi_n_7909 ,csa_tree_add_190_195_groupi_n_7127 ,csa_tree_add_190_195_groupi_n_7312);
  xnor csa_tree_add_190_195_groupi_g41092(csa_tree_add_190_195_groupi_n_7908 ,csa_tree_add_190_195_groupi_n_7204 ,csa_tree_add_190_195_groupi_n_5353);
  xnor csa_tree_add_190_195_groupi_g41093(csa_tree_add_190_195_groupi_n_7907 ,csa_tree_add_190_195_groupi_n_7190 ,csa_tree_add_190_195_groupi_n_7417);
  xnor csa_tree_add_190_195_groupi_g41094(csa_tree_add_190_195_groupi_n_7906 ,csa_tree_add_190_195_groupi_n_7187 ,csa_tree_add_190_195_groupi_n_7149);
  xnor csa_tree_add_190_195_groupi_g41095(csa_tree_add_190_195_groupi_n_7905 ,csa_tree_add_190_195_groupi_n_7091 ,csa_tree_add_190_195_groupi_n_7134);
  xnor csa_tree_add_190_195_groupi_g41096(csa_tree_add_190_195_groupi_n_7904 ,csa_tree_add_190_195_groupi_n_6968 ,csa_tree_add_190_195_groupi_n_7413);
  xnor csa_tree_add_190_195_groupi_g41097(csa_tree_add_190_195_groupi_n_7903 ,csa_tree_add_190_195_groupi_n_6940 ,csa_tree_add_190_195_groupi_n_7160);
  xnor csa_tree_add_190_195_groupi_g41100(csa_tree_add_190_195_groupi_n_7902 ,csa_tree_add_190_195_groupi_n_7412 ,csa_tree_add_190_195_groupi_n_7363);
  xnor csa_tree_add_190_195_groupi_g41101(csa_tree_add_190_195_groupi_n_7901 ,csa_tree_add_190_195_groupi_n_4633 ,csa_tree_add_190_195_groupi_n_7231);
  xnor csa_tree_add_190_195_groupi_g41103(csa_tree_add_190_195_groupi_n_7900 ,csa_tree_add_190_195_groupi_n_7077 ,csa_tree_add_190_195_groupi_n_5281);
  xnor csa_tree_add_190_195_groupi_g41104(csa_tree_add_190_195_groupi_n_7899 ,csa_tree_add_190_195_groupi_n_7360 ,csa_tree_add_190_195_groupi_n_7210);
  xnor csa_tree_add_190_195_groupi_g41105(csa_tree_add_190_195_groupi_n_7898 ,csa_tree_add_190_195_groupi_n_7404 ,csa_tree_add_190_195_groupi_n_7181);
  xnor csa_tree_add_190_195_groupi_g41106(csa_tree_add_190_195_groupi_n_7897 ,csa_tree_add_190_195_groupi_n_7229 ,csa_tree_add_190_195_groupi_n_2040);
  xnor csa_tree_add_190_195_groupi_g41107(csa_tree_add_190_195_groupi_n_7896 ,csa_tree_add_190_195_groupi_n_7385 ,csa_tree_add_190_195_groupi_n_470);
  xnor csa_tree_add_190_195_groupi_g41108(csa_tree_add_190_195_groupi_n_7895 ,csa_tree_add_190_195_groupi_n_6754 ,csa_tree_add_190_195_groupi_n_7185);
  xnor csa_tree_add_190_195_groupi_g41109(csa_tree_add_190_195_groupi_n_7894 ,csa_tree_add_190_195_groupi_n_73 ,csa_tree_add_190_195_groupi_n_2042);
  xnor csa_tree_add_190_195_groupi_g41110(csa_tree_add_190_195_groupi_n_7893 ,csa_tree_add_190_195_groupi_n_7341 ,csa_tree_add_190_195_groupi_n_7164);
  xnor csa_tree_add_190_195_groupi_g41111(csa_tree_add_190_195_groupi_n_7892 ,csa_tree_add_190_195_groupi_n_7424 ,csa_tree_add_190_195_groupi_n_7315);
  xnor csa_tree_add_190_195_groupi_g41112(csa_tree_add_190_195_groupi_n_7891 ,csa_tree_add_190_195_groupi_n_7209 ,csa_tree_add_190_195_groupi_n_7182);
  xnor csa_tree_add_190_195_groupi_g41113(csa_tree_add_190_195_groupi_n_7890 ,csa_tree_add_190_195_groupi_n_7339 ,csa_tree_add_190_195_groupi_n_7150);
  xnor csa_tree_add_190_195_groupi_g41114(csa_tree_add_190_195_groupi_n_7889 ,csa_tree_add_190_195_groupi_n_6929 ,csa_tree_add_190_195_groupi_n_7200);
  xnor csa_tree_add_190_195_groupi_g41115(csa_tree_add_190_195_groupi_n_7888 ,csa_tree_add_190_195_groupi_n_7394 ,csa_tree_add_190_195_groupi_n_5412);
  xnor csa_tree_add_190_195_groupi_g41117(csa_tree_add_190_195_groupi_n_7887 ,csa_tree_add_190_195_groupi_n_7114 ,csa_tree_add_190_195_groupi_n_7305);
  xnor csa_tree_add_190_195_groupi_g41118(csa_tree_add_190_195_groupi_n_7886 ,csa_tree_add_190_195_groupi_n_7429 ,csa_tree_add_190_195_groupi_n_5058);
  xnor csa_tree_add_190_195_groupi_g41119(csa_tree_add_190_195_groupi_n_7885 ,csa_tree_add_190_195_groupi_n_6976 ,csa_tree_add_190_195_groupi_n_30);
  xnor csa_tree_add_190_195_groupi_g41120(csa_tree_add_190_195_groupi_n_7884 ,csa_tree_add_190_195_groupi_n_6931 ,csa_tree_add_190_195_groupi_n_7391);
  xnor csa_tree_add_190_195_groupi_g41121(csa_tree_add_190_195_groupi_n_7883 ,csa_tree_add_190_195_groupi_n_4888 ,csa_tree_add_190_195_groupi_n_7414);
  xnor csa_tree_add_190_195_groupi_g41122(csa_tree_add_190_195_groupi_n_7882 ,csa_tree_add_190_195_groupi_n_7082 ,csa_tree_add_190_195_groupi_n_7423);
  xnor csa_tree_add_190_195_groupi_g41123(csa_tree_add_190_195_groupi_n_7881 ,csa_tree_add_190_195_groupi_n_7153 ,csa_tree_add_190_195_groupi_n_6590);
  xnor csa_tree_add_190_195_groupi_g41124(csa_tree_add_190_195_groupi_n_7880 ,csa_tree_add_190_195_groupi_n_7156 ,csa_tree_add_190_195_groupi_n_7121);
  xnor csa_tree_add_190_195_groupi_g41125(csa_tree_add_190_195_groupi_n_7879 ,csa_tree_add_190_195_groupi_n_7199 ,csa_tree_add_190_195_groupi_n_1745);
  xnor csa_tree_add_190_195_groupi_g41126(csa_tree_add_190_195_groupi_n_7878 ,csa_tree_add_190_195_groupi_n_7396 ,csa_tree_add_190_195_groupi_n_5350);
  xnor csa_tree_add_190_195_groupi_g41128(csa_tree_add_190_195_groupi_n_8059 ,csa_tree_add_190_195_groupi_n_4944 ,csa_tree_add_190_195_groupi_n_7020);
  xnor csa_tree_add_190_195_groupi_g41129(csa_tree_add_190_195_groupi_n_8058 ,csa_tree_add_190_195_groupi_n_7419 ,csa_tree_add_190_195_groupi_n_3780);
  xnor csa_tree_add_190_195_groupi_g41130(csa_tree_add_190_195_groupi_n_8057 ,csa_tree_add_190_195_groupi_n_7408 ,csa_tree_add_190_195_groupi_n_6720);
  xnor csa_tree_add_190_195_groupi_g41131(csa_tree_add_190_195_groupi_n_8055 ,csa_tree_add_190_195_groupi_n_4783 ,csa_tree_add_190_195_groupi_n_7032);
  xnor csa_tree_add_190_195_groupi_g41133(csa_tree_add_190_195_groupi_n_8054 ,csa_tree_add_190_195_groupi_n_7418 ,csa_tree_add_190_195_groupi_n_4077);
  xnor csa_tree_add_190_195_groupi_g41134(csa_tree_add_190_195_groupi_n_8053 ,csa_tree_add_190_195_groupi_n_36 ,csa_tree_add_190_195_groupi_n_1961);
  xnor csa_tree_add_190_195_groupi_g41135(csa_tree_add_190_195_groupi_n_8052 ,csa_tree_add_190_195_groupi_n_7225 ,csa_tree_add_190_195_groupi_n_3758);
  xnor csa_tree_add_190_195_groupi_g41136(csa_tree_add_190_195_groupi_n_8050 ,csa_tree_add_190_195_groupi_n_7211 ,csa_tree_add_190_195_groupi_n_47);
  xnor csa_tree_add_190_195_groupi_g41137(csa_tree_add_190_195_groupi_n_8049 ,csa_tree_add_190_195_groupi_n_7402 ,csa_tree_add_190_195_groupi_n_3793);
  and csa_tree_add_190_195_groupi_g41138(csa_tree_add_190_195_groupi_n_8048 ,csa_tree_add_190_195_groupi_n_7263 ,csa_tree_add_190_195_groupi_n_7484);
  xnor csa_tree_add_190_195_groupi_g41139(csa_tree_add_190_195_groupi_n_8047 ,csa_tree_add_190_195_groupi_n_7381 ,csa_tree_add_190_195_groupi_n_3773);
  and csa_tree_add_190_195_groupi_g41140(csa_tree_add_190_195_groupi_n_8046 ,csa_tree_add_190_195_groupi_n_6163 ,csa_tree_add_190_195_groupi_n_7488);
  or csa_tree_add_190_195_groupi_g41141(csa_tree_add_190_195_groupi_n_8044 ,csa_tree_add_190_195_groupi_n_3265 ,csa_tree_add_190_195_groupi_n_7492);
  or csa_tree_add_190_195_groupi_g41142(csa_tree_add_190_195_groupi_n_8043 ,csa_tree_add_190_195_groupi_n_7041 ,csa_tree_add_190_195_groupi_n_7810);
  and csa_tree_add_190_195_groupi_g41143(csa_tree_add_190_195_groupi_n_8042 ,csa_tree_add_190_195_groupi_n_3318 ,csa_tree_add_190_195_groupi_n_7795);
  and csa_tree_add_190_195_groupi_g41144(csa_tree_add_190_195_groupi_n_8041 ,csa_tree_add_190_195_groupi_n_6565 ,csa_tree_add_190_195_groupi_n_7762);
  or csa_tree_add_190_195_groupi_g41145(csa_tree_add_190_195_groupi_n_8040 ,csa_tree_add_190_195_groupi_n_3430 ,csa_tree_add_190_195_groupi_n_7726);
  and csa_tree_add_190_195_groupi_g41146(csa_tree_add_190_195_groupi_n_8039 ,csa_tree_add_190_195_groupi_n_3633 ,csa_tree_add_190_195_groupi_n_7691);
  and csa_tree_add_190_195_groupi_g41147(csa_tree_add_190_195_groupi_n_8038 ,csa_tree_add_190_195_groupi_n_6849 ,csa_tree_add_190_195_groupi_n_7677);
  or csa_tree_add_190_195_groupi_g41148(csa_tree_add_190_195_groupi_n_8036 ,csa_tree_add_190_195_groupi_n_7282 ,csa_tree_add_190_195_groupi_n_7679);
  or csa_tree_add_190_195_groupi_g41149(csa_tree_add_190_195_groupi_n_8035 ,csa_tree_add_190_195_groupi_n_3147 ,csa_tree_add_190_195_groupi_n_7680);
  and csa_tree_add_190_195_groupi_g41150(csa_tree_add_190_195_groupi_n_8034 ,csa_tree_add_190_195_groupi_n_2853 ,csa_tree_add_190_195_groupi_n_7686);
  and csa_tree_add_190_195_groupi_g41151(csa_tree_add_190_195_groupi_n_8033 ,csa_tree_add_190_195_groupi_n_2878 ,csa_tree_add_190_195_groupi_n_7687);
  xnor csa_tree_add_190_195_groupi_g41152(csa_tree_add_190_195_groupi_n_8031 ,csa_tree_add_190_195_groupi_n_7009 ,csa_tree_add_190_195_groupi_n_7018);
  xnor csa_tree_add_190_195_groupi_g41153(csa_tree_add_190_195_groupi_n_8030 ,csa_tree_add_190_195_groupi_n_7430 ,csa_tree_add_190_195_groupi_n_5996);
  or csa_tree_add_190_195_groupi_g41154(csa_tree_add_190_195_groupi_n_8028 ,csa_tree_add_190_195_groupi_n_6326 ,csa_tree_add_190_195_groupi_n_7482);
  xnor csa_tree_add_190_195_groupi_g41155(csa_tree_add_190_195_groupi_n_8026 ,csa_tree_add_190_195_groupi_n_7207 ,csa_tree_add_190_195_groupi_n_6659);
  xnor csa_tree_add_190_195_groupi_g41156(csa_tree_add_190_195_groupi_n_8024 ,csa_tree_add_190_195_groupi_n_7420 ,csa_tree_add_190_195_groupi_n_6002);
  and csa_tree_add_190_195_groupi_g41157(csa_tree_add_190_195_groupi_n_8022 ,csa_tree_add_190_195_groupi_n_6420 ,csa_tree_add_190_195_groupi_n_7483);
  xnor csa_tree_add_190_195_groupi_g41158(csa_tree_add_190_195_groupi_n_8021 ,csa_tree_add_190_195_groupi_n_7214 ,csa_tree_add_190_195_groupi_n_6666);
  and csa_tree_add_190_195_groupi_g41159(csa_tree_add_190_195_groupi_n_8020 ,csa_tree_add_190_195_groupi_n_6398 ,csa_tree_add_190_195_groupi_n_7486);
  xnor csa_tree_add_190_195_groupi_g41160(csa_tree_add_190_195_groupi_n_8019 ,csa_tree_add_190_195_groupi_n_5082 ,csa_tree_add_190_195_groupi_n_7021);
  xnor csa_tree_add_190_195_groupi_g41161(csa_tree_add_190_195_groupi_n_8016 ,csa_tree_add_190_195_groupi_n_6994 ,csa_tree_add_190_195_groupi_n_7024);
  or csa_tree_add_190_195_groupi_g41162(csa_tree_add_190_195_groupi_n_8015 ,csa_tree_add_190_195_groupi_n_6436 ,csa_tree_add_190_195_groupi_n_7487);
  xnor csa_tree_add_190_195_groupi_g41163(csa_tree_add_190_195_groupi_n_8012 ,csa_tree_add_190_195_groupi_n_6775 ,csa_tree_add_190_195_groupi_n_7033);
  xnor csa_tree_add_190_195_groupi_g41164(csa_tree_add_190_195_groupi_n_8011 ,csa_tree_add_190_195_groupi_n_7195 ,csa_tree_add_190_195_groupi_n_6617);
  xnor csa_tree_add_190_195_groupi_g41165(csa_tree_add_190_195_groupi_n_8008 ,csa_tree_add_190_195_groupi_n_97 ,csa_tree_add_190_195_groupi_n_1944);
  and csa_tree_add_190_195_groupi_g41166(csa_tree_add_190_195_groupi_n_8007 ,csa_tree_add_190_195_groupi_n_3227 ,csa_tree_add_190_195_groupi_n_7475);
  xnor csa_tree_add_190_195_groupi_g41167(csa_tree_add_190_195_groupi_n_8005 ,csa_tree_add_190_195_groupi_n_4893 ,csa_tree_add_190_195_groupi_n_7023);
  xnor csa_tree_add_190_195_groupi_g41168(csa_tree_add_190_195_groupi_n_8004 ,csa_tree_add_190_195_groupi_n_14 ,csa_tree_add_190_195_groupi_n_7028);
  xnor csa_tree_add_190_195_groupi_g41169(csa_tree_add_190_195_groupi_n_8001 ,csa_tree_add_190_195_groupi_n_7193 ,csa_tree_add_190_195_groupi_n_4123);
  xnor csa_tree_add_190_195_groupi_g41170(csa_tree_add_190_195_groupi_n_8000 ,csa_tree_add_190_195_groupi_n_7202 ,csa_tree_add_190_195_groupi_n_3799);
  xnor csa_tree_add_190_195_groupi_g41171(csa_tree_add_190_195_groupi_n_7998 ,csa_tree_add_190_195_groupi_n_7030 ,csa_tree_add_190_195_groupi_n_2015);
  xnor csa_tree_add_190_195_groupi_g41172(csa_tree_add_190_195_groupi_n_7997 ,csa_tree_add_190_195_groupi_n_4582 ,csa_tree_add_190_195_groupi_n_7027);
  xnor csa_tree_add_190_195_groupi_g41173(csa_tree_add_190_195_groupi_n_7994 ,csa_tree_add_190_195_groupi_n_4755 ,csa_tree_add_190_195_groupi_n_7026);
  xnor csa_tree_add_190_195_groupi_g41174(csa_tree_add_190_195_groupi_n_7992 ,csa_tree_add_190_195_groupi_n_4933 ,csa_tree_add_190_195_groupi_n_7025);
  xnor csa_tree_add_190_195_groupi_g41175(csa_tree_add_190_195_groupi_n_7991 ,csa_tree_add_190_195_groupi_n_7401 ,csa_tree_add_190_195_groupi_n_6658);
  or csa_tree_add_190_195_groupi_g41176(csa_tree_add_190_195_groupi_n_7989 ,csa_tree_add_190_195_groupi_n_6743 ,csa_tree_add_190_195_groupi_n_7678);
  xnor csa_tree_add_190_195_groupi_g41177(csa_tree_add_190_195_groupi_n_7988 ,csa_tree_add_190_195_groupi_n_5230 ,csa_tree_add_190_195_groupi_n_7034);
  xnor csa_tree_add_190_195_groupi_g41178(csa_tree_add_190_195_groupi_n_7986 ,csa_tree_add_190_195_groupi_n_5456 ,csa_tree_add_190_195_groupi_n_7017);
  xnor csa_tree_add_190_195_groupi_g41179(csa_tree_add_190_195_groupi_n_7984 ,csa_tree_add_190_195_groupi_n_7197 ,csa_tree_add_190_195_groupi_n_6681);
  and csa_tree_add_190_195_groupi_g41180(csa_tree_add_190_195_groupi_n_7982 ,csa_tree_add_190_195_groupi_n_7054 ,csa_tree_add_190_195_groupi_n_7681);
  and csa_tree_add_190_195_groupi_g41181(csa_tree_add_190_195_groupi_n_7981 ,csa_tree_add_190_195_groupi_n_6109 ,csa_tree_add_190_195_groupi_n_7683);
  xnor csa_tree_add_190_195_groupi_g41182(csa_tree_add_190_195_groupi_n_7980 ,csa_tree_add_190_195_groupi_n_4761 ,csa_tree_add_190_195_groupi_n_7029);
  xnor csa_tree_add_190_195_groupi_g41183(csa_tree_add_190_195_groupi_n_7979 ,csa_tree_add_190_195_groupi_n_98 ,csa_tree_add_190_195_groupi_n_1945);
  not csa_tree_add_190_195_groupi_g41184(csa_tree_add_190_195_groupi_n_7876 ,csa_tree_add_190_195_groupi_n_7875);
  not csa_tree_add_190_195_groupi_g41185(csa_tree_add_190_195_groupi_n_7874 ,csa_tree_add_190_195_groupi_n_7873);
  not csa_tree_add_190_195_groupi_g41186(csa_tree_add_190_195_groupi_n_7867 ,csa_tree_add_190_195_groupi_n_7866);
  not csa_tree_add_190_195_groupi_g41187(csa_tree_add_190_195_groupi_n_7865 ,csa_tree_add_190_195_groupi_n_7864);
  not csa_tree_add_190_195_groupi_g41188(csa_tree_add_190_195_groupi_n_7860 ,csa_tree_add_190_195_groupi_n_7859);
  not csa_tree_add_190_195_groupi_g41189(csa_tree_add_190_195_groupi_n_7857 ,csa_tree_add_190_195_groupi_n_7856);
  not csa_tree_add_190_195_groupi_g41192(csa_tree_add_190_195_groupi_n_7852 ,csa_tree_add_190_195_groupi_n_7851);
  not csa_tree_add_190_195_groupi_g41193(csa_tree_add_190_195_groupi_n_7842 ,csa_tree_add_190_195_groupi_n_7843);
  not csa_tree_add_190_195_groupi_g41194(csa_tree_add_190_195_groupi_n_7840 ,csa_tree_add_190_195_groupi_n_7841);
  not csa_tree_add_190_195_groupi_g41195(csa_tree_add_190_195_groupi_n_7838 ,csa_tree_add_190_195_groupi_n_7839);
  not csa_tree_add_190_195_groupi_g41196(csa_tree_add_190_195_groupi_n_7837 ,csa_tree_add_190_195_groupi_n_7836);
  not csa_tree_add_190_195_groupi_g41197(csa_tree_add_190_195_groupi_n_7834 ,csa_tree_add_190_195_groupi_n_7835);
  not csa_tree_add_190_195_groupi_g41198(csa_tree_add_190_195_groupi_n_7832 ,csa_tree_add_190_195_groupi_n_7833);
  not csa_tree_add_190_195_groupi_g41199(csa_tree_add_190_195_groupi_n_7830 ,csa_tree_add_190_195_groupi_n_7831);
  not csa_tree_add_190_195_groupi_g41200(csa_tree_add_190_195_groupi_n_7828 ,csa_tree_add_190_195_groupi_n_7829);
  not csa_tree_add_190_195_groupi_g41201(csa_tree_add_190_195_groupi_n_7822 ,csa_tree_add_190_195_groupi_n_7823);
  not csa_tree_add_190_195_groupi_g41202(csa_tree_add_190_195_groupi_n_7821 ,csa_tree_add_190_195_groupi_n_7820);
  not csa_tree_add_190_195_groupi_g41203(csa_tree_add_190_195_groupi_n_7818 ,csa_tree_add_190_195_groupi_n_7819);
  and csa_tree_add_190_195_groupi_g41204(csa_tree_add_190_195_groupi_n_7817 ,csa_tree_add_190_195_groupi_n_5400 ,csa_tree_add_190_195_groupi_n_7373);
  and csa_tree_add_190_195_groupi_g41205(csa_tree_add_190_195_groupi_n_7816 ,csa_tree_add_190_195_groupi_n_5834 ,csa_tree_add_190_195_groupi_n_7409);
  or csa_tree_add_190_195_groupi_g41206(csa_tree_add_190_195_groupi_n_7815 ,csa_tree_add_190_195_groupi_n_7317 ,csa_tree_add_190_195_groupi_n_7094);
  and csa_tree_add_190_195_groupi_g41207(csa_tree_add_190_195_groupi_n_7814 ,csa_tree_add_190_195_groupi_n_7317 ,csa_tree_add_190_195_groupi_n_7094);
  or csa_tree_add_190_195_groupi_g41208(csa_tree_add_190_195_groupi_n_7813 ,csa_tree_add_190_195_groupi_n_7300 ,csa_tree_add_190_195_groupi_n_78);
  or csa_tree_add_190_195_groupi_g41209(csa_tree_add_190_195_groupi_n_7812 ,csa_tree_add_190_195_groupi_n_5404 ,csa_tree_add_190_195_groupi_n_7104);
  nor csa_tree_add_190_195_groupi_g41210(csa_tree_add_190_195_groupi_n_7811 ,csa_tree_add_190_195_groupi_n_7272 ,csa_tree_add_190_195_groupi_n_7395);
  nor csa_tree_add_190_195_groupi_g41211(csa_tree_add_190_195_groupi_n_7810 ,csa_tree_add_190_195_groupi_n_6972 ,csa_tree_add_190_195_groupi_n_7040);
  nor csa_tree_add_190_195_groupi_g41212(csa_tree_add_190_195_groupi_n_7809 ,csa_tree_add_190_195_groupi_n_5403 ,csa_tree_add_190_195_groupi_n_7105);
  or csa_tree_add_190_195_groupi_g41213(csa_tree_add_190_195_groupi_n_7808 ,csa_tree_add_190_195_groupi_n_6525 ,csa_tree_add_190_195_groupi_n_84);
  and csa_tree_add_190_195_groupi_g41214(csa_tree_add_190_195_groupi_n_7807 ,csa_tree_add_190_195_groupi_n_7293 ,csa_tree_add_190_195_groupi_n_7406);
  or csa_tree_add_190_195_groupi_g41215(csa_tree_add_190_195_groupi_n_7806 ,csa_tree_add_190_195_groupi_n_6943 ,csa_tree_add_190_195_groupi_n_7154);
  or csa_tree_add_190_195_groupi_g41216(csa_tree_add_190_195_groupi_n_7805 ,csa_tree_add_190_195_groupi_n_6508 ,csa_tree_add_190_195_groupi_n_7197);
  or csa_tree_add_190_195_groupi_g41217(csa_tree_add_190_195_groupi_n_7804 ,csa_tree_add_190_195_groupi_n_5939 ,csa_tree_add_190_195_groupi_n_7107);
  nor csa_tree_add_190_195_groupi_g41218(csa_tree_add_190_195_groupi_n_7803 ,csa_tree_add_190_195_groupi_n_3049 ,csa_tree_add_190_195_groupi_n_7419);
  nor csa_tree_add_190_195_groupi_g41219(csa_tree_add_190_195_groupi_n_7802 ,csa_tree_add_190_195_groupi_n_5940 ,csa_tree_add_190_195_groupi_n_7108);
  or csa_tree_add_190_195_groupi_g41220(csa_tree_add_190_195_groupi_n_7801 ,csa_tree_add_190_195_groupi_n_6754 ,csa_tree_add_190_195_groupi_n_7184);
  and csa_tree_add_190_195_groupi_g41221(csa_tree_add_190_195_groupi_n_7800 ,csa_tree_add_190_195_groupi_n_7106 ,csa_tree_add_190_195_groupi_n_7363);
  nor csa_tree_add_190_195_groupi_g41222(csa_tree_add_190_195_groupi_n_7799 ,csa_tree_add_190_195_groupi_n_6753 ,csa_tree_add_190_195_groupi_n_7185);
  and csa_tree_add_190_195_groupi_g41223(csa_tree_add_190_195_groupi_n_7798 ,csa_tree_add_190_195_groupi_n_6495 ,csa_tree_add_190_195_groupi_n_7410);
  nor csa_tree_add_190_195_groupi_g41224(csa_tree_add_190_195_groupi_n_7797 ,csa_tree_add_190_195_groupi_n_7315 ,csa_tree_add_190_195_groupi_n_6757);
  or csa_tree_add_190_195_groupi_g41225(csa_tree_add_190_195_groupi_n_7796 ,csa_tree_add_190_195_groupi_n_7355 ,csa_tree_add_190_195_groupi_n_7374);
  or csa_tree_add_190_195_groupi_g41226(csa_tree_add_190_195_groupi_n_7795 ,csa_tree_add_190_195_groupi_n_3364 ,csa_tree_add_190_195_groupi_n_7418);
  and csa_tree_add_190_195_groupi_g41227(csa_tree_add_190_195_groupi_n_7794 ,csa_tree_add_190_195_groupi_n_1676 ,csa_tree_add_190_195_groupi_n_7119);
  or csa_tree_add_190_195_groupi_g41228(csa_tree_add_190_195_groupi_n_7793 ,csa_tree_add_190_195_groupi_n_1676 ,csa_tree_add_190_195_groupi_n_7119);
  or csa_tree_add_190_195_groupi_g41229(csa_tree_add_190_195_groupi_n_7792 ,csa_tree_add_190_195_groupi_n_7127 ,csa_tree_add_190_195_groupi_n_7311);
  nor csa_tree_add_190_195_groupi_g41230(csa_tree_add_190_195_groupi_n_7791 ,csa_tree_add_190_195_groupi_n_6272 ,csa_tree_add_190_195_groupi_n_7191);
  or csa_tree_add_190_195_groupi_g41231(csa_tree_add_190_195_groupi_n_7790 ,csa_tree_add_190_195_groupi_n_2939 ,csa_tree_add_190_195_groupi_n_7193);
  or csa_tree_add_190_195_groupi_g41232(csa_tree_add_190_195_groupi_n_7789 ,csa_tree_add_190_195_groupi_n_5492 ,csa_tree_add_190_195_groupi_n_7328);
  nor csa_tree_add_190_195_groupi_g41233(csa_tree_add_190_195_groupi_n_7788 ,csa_tree_add_190_195_groupi_n_5493 ,csa_tree_add_190_195_groupi_n_7329);
  or csa_tree_add_190_195_groupi_g41234(csa_tree_add_190_195_groupi_n_7787 ,csa_tree_add_190_195_groupi_n_7285 ,csa_tree_add_190_195_groupi_n_7429);
  nor csa_tree_add_190_195_groupi_g41235(csa_tree_add_190_195_groupi_n_7786 ,csa_tree_add_190_195_groupi_n_7126 ,csa_tree_add_190_195_groupi_n_7312);
  or csa_tree_add_190_195_groupi_g41236(csa_tree_add_190_195_groupi_n_7785 ,csa_tree_add_190_195_groupi_n_7187 ,csa_tree_add_190_195_groupi_n_7148);
  or csa_tree_add_190_195_groupi_g41237(csa_tree_add_190_195_groupi_n_7784 ,csa_tree_add_190_195_groupi_n_3132 ,csa_tree_add_190_195_groupi_n_7428);
  nor csa_tree_add_190_195_groupi_g41238(csa_tree_add_190_195_groupi_n_7783 ,csa_tree_add_190_195_groupi_n_5038 ,csa_tree_add_190_195_groupi_n_7088);
  and csa_tree_add_190_195_groupi_g41239(csa_tree_add_190_195_groupi_n_7782 ,csa_tree_add_190_195_groupi_n_5038 ,csa_tree_add_190_195_groupi_n_7088);
  or csa_tree_add_190_195_groupi_g41240(csa_tree_add_190_195_groupi_n_7781 ,csa_tree_add_190_195_groupi_n_5365 ,csa_tree_add_190_195_groupi_n_7182);
  and csa_tree_add_190_195_groupi_g41241(csa_tree_add_190_195_groupi_n_7780 ,csa_tree_add_190_195_groupi_n_5365 ,csa_tree_add_190_195_groupi_n_7182);
  nor csa_tree_add_190_195_groupi_g41242(csa_tree_add_190_195_groupi_n_7779 ,csa_tree_add_190_195_groupi_n_7097 ,csa_tree_add_190_195_groupi_n_7377);
  nor csa_tree_add_190_195_groupi_g41243(csa_tree_add_190_195_groupi_n_7778 ,csa_tree_add_190_195_groupi_n_4763 ,csa_tree_add_190_195_groupi_n_7324);
  or csa_tree_add_190_195_groupi_g41244(csa_tree_add_190_195_groupi_n_7777 ,csa_tree_add_190_195_groupi_n_7076 ,csa_tree_add_190_195_groupi_n_7364);
  nor csa_tree_add_190_195_groupi_g41245(csa_tree_add_190_195_groupi_n_7776 ,csa_tree_add_190_195_groupi_n_7106 ,csa_tree_add_190_195_groupi_n_7363);
  nor csa_tree_add_190_195_groupi_g41246(csa_tree_add_190_195_groupi_n_7775 ,csa_tree_add_190_195_groupi_n_7370 ,csa_tree_add_190_195_groupi_n_7084);
  nor csa_tree_add_190_195_groupi_g41247(csa_tree_add_190_195_groupi_n_7774 ,csa_tree_add_190_195_groupi_n_7186 ,csa_tree_add_190_195_groupi_n_7149);
  nor csa_tree_add_190_195_groupi_g41248(csa_tree_add_190_195_groupi_n_7773 ,csa_tree_add_190_195_groupi_n_6426 ,csa_tree_add_190_195_groupi_n_7204);
  or csa_tree_add_190_195_groupi_g41249(csa_tree_add_190_195_groupi_n_7772 ,csa_tree_add_190_195_groupi_n_5955 ,csa_tree_add_190_195_groupi_n_7090);
  and csa_tree_add_190_195_groupi_g41250(csa_tree_add_190_195_groupi_n_7771 ,csa_tree_add_190_195_groupi_n_7097 ,csa_tree_add_190_195_groupi_n_7377);
  or csa_tree_add_190_195_groupi_g41251(csa_tree_add_190_195_groupi_n_7770 ,csa_tree_add_190_195_groupi_n_6418 ,csa_tree_add_190_195_groupi_n_7396);
  and csa_tree_add_190_195_groupi_g41252(csa_tree_add_190_195_groupi_n_7769 ,csa_tree_add_190_195_groupi_n_7352 ,csa_tree_add_190_195_groupi_n_7083);
  or csa_tree_add_190_195_groupi_g41253(csa_tree_add_190_195_groupi_n_7768 ,csa_tree_add_190_195_groupi_n_7 ,csa_tree_add_190_195_groupi_n_7342);
  nor csa_tree_add_190_195_groupi_g41254(csa_tree_add_190_195_groupi_n_7767 ,csa_tree_add_190_195_groupi_n_7352 ,csa_tree_add_190_195_groupi_n_7083);
  or csa_tree_add_190_195_groupi_g41255(csa_tree_add_190_195_groupi_n_7766 ,csa_tree_add_190_195_groupi_n_5382 ,csa_tree_add_190_195_groupi_n_7330);
  or csa_tree_add_190_195_groupi_g41256(csa_tree_add_190_195_groupi_n_7765 ,csa_tree_add_190_195_groupi_n_6987 ,csa_tree_add_190_195_groupi_n_7276);
  or csa_tree_add_190_195_groupi_g41257(csa_tree_add_190_195_groupi_n_7764 ,csa_tree_add_190_195_groupi_n_5746 ,csa_tree_add_190_195_groupi_n_7430);
  and csa_tree_add_190_195_groupi_g41258(csa_tree_add_190_195_groupi_n_7763 ,csa_tree_add_190_195_groupi_n_5382 ,csa_tree_add_190_195_groupi_n_7330);
  or csa_tree_add_190_195_groupi_g41259(csa_tree_add_190_195_groupi_n_7762 ,csa_tree_add_190_195_groupi_n_6562 ,csa_tree_add_190_195_groupi_n_7400);
  and csa_tree_add_190_195_groupi_g41260(csa_tree_add_190_195_groupi_n_7761 ,csa_tree_add_190_195_groupi_n_4891 ,csa_tree_add_190_195_groupi_n_30);
  nor csa_tree_add_190_195_groupi_g41261(csa_tree_add_190_195_groupi_n_7760 ,csa_tree_add_190_195_groupi_n_4891 ,csa_tree_add_190_195_groupi_n_30);
  or csa_tree_add_190_195_groupi_g41262(csa_tree_add_190_195_groupi_n_7759 ,csa_tree_add_190_195_groupi_n_7384 ,csa_tree_add_190_195_groupi_n_6372);
  nor csa_tree_add_190_195_groupi_g41263(csa_tree_add_190_195_groupi_n_7758 ,csa_tree_add_190_195_groupi_n_5487 ,csa_tree_add_190_195_groupi_n_7082);
  or csa_tree_add_190_195_groupi_g41264(csa_tree_add_190_195_groupi_n_7757 ,csa_tree_add_190_195_groupi_n_5486 ,csa_tree_add_190_195_groupi_n_7081);
  or csa_tree_add_190_195_groupi_g41265(csa_tree_add_190_195_groupi_n_7756 ,csa_tree_add_190_195_groupi_n_3279 ,csa_tree_add_190_195_groupi_n_7211);
  or csa_tree_add_190_195_groupi_g41266(csa_tree_add_190_195_groupi_n_7755 ,csa_tree_add_190_195_groupi_n_5653 ,csa_tree_add_190_195_groupi_n_7421);
  or csa_tree_add_190_195_groupi_g41267(csa_tree_add_190_195_groupi_n_7754 ,csa_tree_add_190_195_groupi_n_6848 ,csa_tree_add_190_195_groupi_n_7206);
  or csa_tree_add_190_195_groupi_g41268(csa_tree_add_190_195_groupi_n_7753 ,csa_tree_add_190_195_groupi_n_5507 ,csa_tree_add_190_195_groupi_n_74);
  nor csa_tree_add_190_195_groupi_g41269(csa_tree_add_190_195_groupi_n_7752 ,csa_tree_add_190_195_groupi_n_5508 ,csa_tree_add_190_195_groupi_n_7095);
  nor csa_tree_add_190_195_groupi_g41270(csa_tree_add_190_195_groupi_n_7751 ,csa_tree_add_190_195_groupi_n_7356 ,csa_tree_add_190_195_groupi_n_7375);
  nor csa_tree_add_190_195_groupi_g41271(csa_tree_add_190_195_groupi_n_7750 ,csa_tree_add_190_195_groupi_n_5400 ,csa_tree_add_190_195_groupi_n_7373);
  or csa_tree_add_190_195_groupi_g41272(csa_tree_add_190_195_groupi_n_7749 ,csa_tree_add_190_195_groupi_n_6196 ,csa_tree_add_190_195_groupi_n_7227);
  and csa_tree_add_190_195_groupi_g41273(csa_tree_add_190_195_groupi_n_7748 ,csa_tree_add_190_195_groupi_n_7067 ,csa_tree_add_190_195_groupi_n_7308);
  or csa_tree_add_190_195_groupi_g41274(csa_tree_add_190_195_groupi_n_7747 ,csa_tree_add_190_195_groupi_n_7369 ,csa_tree_add_190_195_groupi_n_7085);
  and csa_tree_add_190_195_groupi_g41275(csa_tree_add_190_195_groupi_n_7746 ,csa_tree_add_190_195_groupi_n_6229 ,csa_tree_add_190_195_groupi_n_7224);
  nor csa_tree_add_190_195_groupi_g41276(csa_tree_add_190_195_groupi_n_7745 ,csa_tree_add_190_195_groupi_n_7340 ,csa_tree_add_190_195_groupi_n_7164);
  or csa_tree_add_190_195_groupi_g41277(csa_tree_add_190_195_groupi_n_7744 ,csa_tree_add_190_195_groupi_n_4956 ,csa_tree_add_190_195_groupi_n_21);
  or csa_tree_add_190_195_groupi_g41278(csa_tree_add_190_195_groupi_n_7743 ,csa_tree_add_190_195_groupi_n_6939 ,csa_tree_add_190_195_groupi_n_7160);
  and csa_tree_add_190_195_groupi_g41279(csa_tree_add_190_195_groupi_n_7742 ,csa_tree_add_190_195_groupi_n_6340 ,csa_tree_add_190_195_groupi_n_7399);
  nor csa_tree_add_190_195_groupi_g41280(csa_tree_add_190_195_groupi_n_7741 ,csa_tree_add_190_195_groupi_n_6940 ,csa_tree_add_190_195_groupi_n_7159);
  or csa_tree_add_190_195_groupi_g41281(csa_tree_add_190_195_groupi_n_7740 ,csa_tree_add_190_195_groupi_n_7156 ,csa_tree_add_190_195_groupi_n_7120);
  nor csa_tree_add_190_195_groupi_g41282(csa_tree_add_190_195_groupi_n_7739 ,csa_tree_add_190_195_groupi_n_7153 ,csa_tree_add_190_195_groupi_n_7137);
  nor csa_tree_add_190_195_groupi_g41283(csa_tree_add_190_195_groupi_n_7738 ,csa_tree_add_190_195_groupi_n_7067 ,csa_tree_add_190_195_groupi_n_7308);
  and csa_tree_add_190_195_groupi_g41284(csa_tree_add_190_195_groupi_n_7737 ,csa_tree_add_190_195_groupi_n_7153 ,csa_tree_add_190_195_groupi_n_7137);
  nor csa_tree_add_190_195_groupi_g41285(csa_tree_add_190_195_groupi_n_7736 ,csa_tree_add_190_195_groupi_n_7155 ,csa_tree_add_190_195_groupi_n_7121);
  or csa_tree_add_190_195_groupi_g41286(csa_tree_add_190_195_groupi_n_7735 ,csa_tree_add_190_195_groupi_n_7074 ,csa_tree_add_190_195_groupi_n_7140);
  and csa_tree_add_190_195_groupi_g41287(csa_tree_add_190_195_groupi_n_7734 ,csa_tree_add_190_195_groupi_n_7 ,csa_tree_add_190_195_groupi_n_7342);
  or csa_tree_add_190_195_groupi_g41288(csa_tree_add_190_195_groupi_n_7733 ,csa_tree_add_190_195_groupi_n_2787 ,csa_tree_add_190_195_groupi_n_7225);
  and csa_tree_add_190_195_groupi_g41289(csa_tree_add_190_195_groupi_n_7732 ,csa_tree_add_190_195_groupi_n_7386 ,csa_tree_add_190_195_groupi_n_7258);
  or csa_tree_add_190_195_groupi_g41290(csa_tree_add_190_195_groupi_n_7731 ,csa_tree_add_190_195_groupi_n_7339 ,csa_tree_add_190_195_groupi_n_7150);
  and csa_tree_add_190_195_groupi_g41291(csa_tree_add_190_195_groupi_n_7730 ,csa_tree_add_190_195_groupi_n_7228 ,csa_tree_add_190_195_groupi_n_7255);
  nor csa_tree_add_190_195_groupi_g41292(csa_tree_add_190_195_groupi_n_7729 ,csa_tree_add_190_195_groupi_n_50 ,csa_tree_add_190_195_groupi_n_7089);
  and csa_tree_add_190_195_groupi_g41293(csa_tree_add_190_195_groupi_n_7728 ,csa_tree_add_190_195_groupi_n_7315 ,csa_tree_add_190_195_groupi_n_6757);
  or csa_tree_add_190_195_groupi_g41294(csa_tree_add_190_195_groupi_n_7727 ,csa_tree_add_190_195_groupi_n_3186 ,csa_tree_add_190_195_groupi_n_7220);
  nor csa_tree_add_190_195_groupi_g41295(csa_tree_add_190_195_groupi_n_7726 ,csa_tree_add_190_195_groupi_n_3437 ,csa_tree_add_190_195_groupi_n_7199);
  or csa_tree_add_190_195_groupi_g41296(csa_tree_add_190_195_groupi_n_7725 ,csa_tree_add_190_195_groupi_n_5281 ,csa_tree_add_190_195_groupi_n_7077);
  or csa_tree_add_190_195_groupi_g41297(csa_tree_add_190_195_groupi_n_7724 ,csa_tree_add_190_195_groupi_n_5927 ,csa_tree_add_190_195_groupi_n_7379);
  and csa_tree_add_190_195_groupi_g41298(csa_tree_add_190_195_groupi_n_7723 ,csa_tree_add_190_195_groupi_n_5281 ,csa_tree_add_190_195_groupi_n_7077);
  nor csa_tree_add_190_195_groupi_g41299(csa_tree_add_190_195_groupi_n_7722 ,csa_tree_add_190_195_groupi_n_5928 ,csa_tree_add_190_195_groupi_n_7380);
  or csa_tree_add_190_195_groupi_g41300(csa_tree_add_190_195_groupi_n_7721 ,csa_tree_add_190_195_groupi_n_7143 ,csa_tree_add_190_195_groupi_n_7371);
  or csa_tree_add_190_195_groupi_g41301(csa_tree_add_190_195_groupi_n_7720 ,csa_tree_add_190_195_groupi_n_6887 ,csa_tree_add_190_195_groupi_n_7223);
  nor csa_tree_add_190_195_groupi_g41302(csa_tree_add_190_195_groupi_n_7719 ,csa_tree_add_190_195_groupi_n_7075 ,csa_tree_add_190_195_groupi_n_7139);
  and csa_tree_add_190_195_groupi_g41303(csa_tree_add_190_195_groupi_n_7718 ,csa_tree_add_190_195_groupi_n_7339 ,csa_tree_add_190_195_groupi_n_7150);
  and csa_tree_add_190_195_groupi_g41304(csa_tree_add_190_195_groupi_n_7717 ,csa_tree_add_190_195_groupi_n_6201 ,csa_tree_add_190_195_groupi_n_7401);
  and csa_tree_add_190_195_groupi_g41305(csa_tree_add_190_195_groupi_n_7716 ,csa_tree_add_190_195_groupi_n_7076 ,csa_tree_add_190_195_groupi_n_7364);
  or csa_tree_add_190_195_groupi_g41306(csa_tree_add_190_195_groupi_n_7715 ,csa_tree_add_190_195_groupi_n_7002 ,csa_tree_add_190_195_groupi_n_7244);
  nor csa_tree_add_190_195_groupi_g41307(csa_tree_add_190_195_groupi_n_7714 ,csa_tree_add_190_195_groupi_n_7144 ,csa_tree_add_190_195_groupi_n_7372);
  or csa_tree_add_190_195_groupi_g41308(csa_tree_add_190_195_groupi_n_7713 ,csa_tree_add_190_195_groupi_n_6776 ,csa_tree_add_190_195_groupi_n_7269);
  and csa_tree_add_190_195_groupi_g41309(csa_tree_add_190_195_groupi_n_7712 ,csa_tree_add_190_195_groupi_n_3181 ,csa_tree_add_190_195_groupi_n_7402);
  nor csa_tree_add_190_195_groupi_g41310(csa_tree_add_190_195_groupi_n_7711 ,csa_tree_add_190_195_groupi_n_7133 ,csa_tree_add_190_195_groupi_n_7101);
  or csa_tree_add_190_195_groupi_g41311(csa_tree_add_190_195_groupi_n_7710 ,csa_tree_add_190_195_groupi_n_5208 ,csa_tree_add_190_195_groupi_n_7175);
  nor csa_tree_add_190_195_groupi_g41312(csa_tree_add_190_195_groupi_n_7709 ,csa_tree_add_190_195_groupi_n_5209 ,csa_tree_add_190_195_groupi_n_7176);
  or csa_tree_add_190_195_groupi_g41313(csa_tree_add_190_195_groupi_n_7708 ,csa_tree_add_190_195_groupi_n_52 ,csa_tree_add_190_195_groupi_n_7073);
  and csa_tree_add_190_195_groupi_g41314(csa_tree_add_190_195_groupi_n_7707 ,csa_tree_add_190_195_groupi_n_52 ,csa_tree_add_190_195_groupi_n_7073);
  and csa_tree_add_190_195_groupi_g41315(csa_tree_add_190_195_groupi_n_7706 ,csa_tree_add_190_195_groupi_n_6323 ,csa_tree_add_190_195_groupi_n_7408);
  and csa_tree_add_190_195_groupi_g41316(csa_tree_add_190_195_groupi_n_7705 ,csa_tree_add_190_195_groupi_n_7351 ,csa_tree_add_190_195_groupi_n_7135);
  or csa_tree_add_190_195_groupi_g41317(csa_tree_add_190_195_groupi_n_7704 ,csa_tree_add_190_195_groupi_n_7341 ,csa_tree_add_190_195_groupi_n_7163);
  or csa_tree_add_190_195_groupi_g41318(csa_tree_add_190_195_groupi_n_7703 ,csa_tree_add_190_195_groupi_n_5417 ,csa_tree_add_190_195_groupi_n_7316);
  or csa_tree_add_190_195_groupi_g41319(csa_tree_add_190_195_groupi_n_7702 ,csa_tree_add_190_195_groupi_n_7351 ,csa_tree_add_190_195_groupi_n_7135);
  nor csa_tree_add_190_195_groupi_g41320(csa_tree_add_190_195_groupi_n_7701 ,csa_tree_add_190_195_groupi_n_4957 ,csa_tree_add_190_195_groupi_n_7151);
  or csa_tree_add_190_195_groupi_g41321(csa_tree_add_190_195_groupi_n_7700 ,csa_tree_add_190_195_groupi_n_6175 ,csa_tree_add_190_195_groupi_n_7195);
  or csa_tree_add_190_195_groupi_g41322(csa_tree_add_190_195_groupi_n_7699 ,csa_tree_add_190_195_groupi_n_3037 ,csa_tree_add_190_195_groupi_n_7203);
  or csa_tree_add_190_195_groupi_g41323(csa_tree_add_190_195_groupi_n_7698 ,csa_tree_add_190_195_groupi_n_6197 ,csa_tree_add_190_195_groupi_n_7219);
  or csa_tree_add_190_195_groupi_g41324(csa_tree_add_190_195_groupi_n_7697 ,csa_tree_add_190_195_groupi_n_4762 ,csa_tree_add_190_195_groupi_n_7325);
  or csa_tree_add_190_195_groupi_g41325(csa_tree_add_190_195_groupi_n_7696 ,csa_tree_add_190_195_groupi_n_2817 ,csa_tree_add_190_195_groupi_n_7393);
  or csa_tree_add_190_195_groupi_g41326(csa_tree_add_190_195_groupi_n_7695 ,csa_tree_add_190_195_groupi_n_6271 ,csa_tree_add_190_195_groupi_n_7192);
  and csa_tree_add_190_195_groupi_g41327(csa_tree_add_190_195_groupi_n_7694 ,csa_tree_add_190_195_groupi_n_6943 ,csa_tree_add_190_195_groupi_n_7154);
  and csa_tree_add_190_195_groupi_g41328(csa_tree_add_190_195_groupi_n_7693 ,csa_tree_add_190_195_groupi_n_5417 ,csa_tree_add_190_195_groupi_n_7316);
  or csa_tree_add_190_195_groupi_g41329(csa_tree_add_190_195_groupi_n_7692 ,csa_tree_add_190_195_groupi_n_7132 ,csa_tree_add_190_195_groupi_n_7100);
  or csa_tree_add_190_195_groupi_g41330(csa_tree_add_190_195_groupi_n_7691 ,csa_tree_add_190_195_groupi_n_3645 ,csa_tree_add_190_195_groupi_n_7416);
  nor csa_tree_add_190_195_groupi_g41331(csa_tree_add_190_195_groupi_n_7690 ,csa_tree_add_190_195_groupi_n_4654 ,csa_tree_add_190_195_groupi_n_7065);
  or csa_tree_add_190_195_groupi_g41332(csa_tree_add_190_195_groupi_n_7689 ,csa_tree_add_190_195_groupi_n_4655 ,csa_tree_add_190_195_groupi_n_7064);
  nor csa_tree_add_190_195_groupi_g41333(csa_tree_add_190_195_groupi_n_7688 ,csa_tree_add_190_195_groupi_n_7305 ,csa_tree_add_190_195_groupi_n_7114);
  or csa_tree_add_190_195_groupi_g41334(csa_tree_add_190_195_groupi_n_7687 ,csa_tree_add_190_195_groupi_n_2844 ,csa_tree_add_190_195_groupi_n_7381);
  or csa_tree_add_190_195_groupi_g41335(csa_tree_add_190_195_groupi_n_7686 ,csa_tree_add_190_195_groupi_n_3024 ,csa_tree_add_190_195_groupi_n_7230);
  or csa_tree_add_190_195_groupi_g41336(csa_tree_add_190_195_groupi_n_7685 ,csa_tree_add_190_195_groupi_n_7304 ,csa_tree_add_190_195_groupi_n_7113);
  or csa_tree_add_190_195_groupi_g41337(csa_tree_add_190_195_groupi_n_7684 ,csa_tree_add_190_195_groupi_n_5196 ,csa_tree_add_190_195_groupi_n_7062);
  or csa_tree_add_190_195_groupi_g41338(csa_tree_add_190_195_groupi_n_7683 ,csa_tree_add_190_195_groupi_n_6108 ,csa_tree_add_190_195_groupi_n_7198);
  nor csa_tree_add_190_195_groupi_g41339(csa_tree_add_190_195_groupi_n_7682 ,csa_tree_add_190_195_groupi_n_5195 ,csa_tree_add_190_195_groupi_n_7063);
  or csa_tree_add_190_195_groupi_g41340(csa_tree_add_190_195_groupi_n_7681 ,csa_tree_add_190_195_groupi_n_7217 ,csa_tree_add_190_195_groupi_n_7053);
  and csa_tree_add_190_195_groupi_g41341(csa_tree_add_190_195_groupi_n_7680 ,csa_tree_add_190_195_groupi_n_2781 ,csa_tree_add_190_195_groupi_n_7201);
  and csa_tree_add_190_195_groupi_g41342(csa_tree_add_190_195_groupi_n_7679 ,csa_tree_add_190_195_groupi_n_7281 ,csa_tree_add_190_195_groupi_n_7200);
  nor csa_tree_add_190_195_groupi_g41343(csa_tree_add_190_195_groupi_n_7678 ,csa_tree_add_190_195_groupi_n_6742 ,csa_tree_add_190_195_groupi_n_7231);
  or csa_tree_add_190_195_groupi_g41344(csa_tree_add_190_195_groupi_n_7677 ,csa_tree_add_190_195_groupi_n_6840 ,csa_tree_add_190_195_groupi_n_7389);
  and csa_tree_add_190_195_groupi_g41345(csa_tree_add_190_195_groupi_n_7877 ,csa_tree_add_190_195_groupi_n_6177 ,csa_tree_add_190_195_groupi_n_7042);
  or csa_tree_add_190_195_groupi_g41346(csa_tree_add_190_195_groupi_n_7875 ,csa_tree_add_190_195_groupi_n_6839 ,csa_tree_add_190_195_groupi_n_7237);
  or csa_tree_add_190_195_groupi_g41347(csa_tree_add_190_195_groupi_n_7873 ,csa_tree_add_190_195_groupi_n_6567 ,csa_tree_add_190_195_groupi_n_7045);
  and csa_tree_add_190_195_groupi_g41348(csa_tree_add_190_195_groupi_n_7872 ,csa_tree_add_190_195_groupi_n_6503 ,csa_tree_add_190_195_groupi_n_7291);
  and csa_tree_add_190_195_groupi_g41349(csa_tree_add_190_195_groupi_n_7871 ,csa_tree_add_190_195_groupi_n_3343 ,csa_tree_add_190_195_groupi_n_7043);
  or csa_tree_add_190_195_groupi_g41350(csa_tree_add_190_195_groupi_n_7870 ,csa_tree_add_190_195_groupi_n_5661 ,csa_tree_add_190_195_groupi_n_7234);
  and csa_tree_add_190_195_groupi_g41351(csa_tree_add_190_195_groupi_n_7869 ,csa_tree_add_190_195_groupi_n_5784 ,csa_tree_add_190_195_groupi_n_7290);
  and csa_tree_add_190_195_groupi_g41352(csa_tree_add_190_195_groupi_n_7868 ,csa_tree_add_190_195_groupi_n_6865 ,csa_tree_add_190_195_groupi_n_7235);
  or csa_tree_add_190_195_groupi_g41353(csa_tree_add_190_195_groupi_n_7866 ,csa_tree_add_190_195_groupi_n_3667 ,csa_tree_add_190_195_groupi_n_7301);
  or csa_tree_add_190_195_groupi_g41354(csa_tree_add_190_195_groupi_n_7864 ,csa_tree_add_190_195_groupi_n_6228 ,csa_tree_add_190_195_groupi_n_7287);
  or csa_tree_add_190_195_groupi_g41355(csa_tree_add_190_195_groupi_n_7863 ,csa_tree_add_190_195_groupi_n_6370 ,csa_tree_add_190_195_groupi_n_7271);
  or csa_tree_add_190_195_groupi_g41356(csa_tree_add_190_195_groupi_n_7862 ,csa_tree_add_190_195_groupi_n_6210 ,csa_tree_add_190_195_groupi_n_7265);
  and csa_tree_add_190_195_groupi_g41357(csa_tree_add_190_195_groupi_n_7861 ,csa_tree_add_190_195_groupi_n_5684 ,csa_tree_add_190_195_groupi_n_7240);
  or csa_tree_add_190_195_groupi_g41358(csa_tree_add_190_195_groupi_n_7859 ,csa_tree_add_190_195_groupi_n_2778 ,csa_tree_add_190_195_groupi_n_7260);
  and csa_tree_add_190_195_groupi_g41359(csa_tree_add_190_195_groupi_n_7858 ,csa_tree_add_190_195_groupi_n_6905 ,csa_tree_add_190_195_groupi_n_7059);
  or csa_tree_add_190_195_groupi_g41360(csa_tree_add_190_195_groupi_n_7856 ,csa_tree_add_190_195_groupi_n_5646 ,csa_tree_add_190_195_groupi_n_7058);
  and csa_tree_add_190_195_groupi_g41361(csa_tree_add_190_195_groupi_n_7855 ,csa_tree_add_190_195_groupi_n_6446 ,csa_tree_add_190_195_groupi_n_7242);
  and csa_tree_add_190_195_groupi_g41362(csa_tree_add_190_195_groupi_n_7854 ,csa_tree_add_190_195_groupi_n_6185 ,csa_tree_add_190_195_groupi_n_7248);
  and csa_tree_add_190_195_groupi_g41363(csa_tree_add_190_195_groupi_n_7853 ,csa_tree_add_190_195_groupi_n_5706 ,csa_tree_add_190_195_groupi_n_7055);
  or csa_tree_add_190_195_groupi_g41364(csa_tree_add_190_195_groupi_n_7851 ,csa_tree_add_190_195_groupi_n_5814 ,csa_tree_add_190_195_groupi_n_7292);
  or csa_tree_add_190_195_groupi_g41365(csa_tree_add_190_195_groupi_n_7850 ,csa_tree_add_190_195_groupi_n_6300 ,csa_tree_add_190_195_groupi_n_7259);
  or csa_tree_add_190_195_groupi_g41366(csa_tree_add_190_195_groupi_n_7849 ,csa_tree_add_190_195_groupi_n_5710 ,csa_tree_add_190_195_groupi_n_7257);
  and csa_tree_add_190_195_groupi_g41367(csa_tree_add_190_195_groupi_n_7848 ,csa_tree_add_190_195_groupi_n_6747 ,csa_tree_add_190_195_groupi_n_7052);
  and csa_tree_add_190_195_groupi_g41368(csa_tree_add_190_195_groupi_n_7847 ,csa_tree_add_190_195_groupi_n_5721 ,csa_tree_add_190_195_groupi_n_7261);
  and csa_tree_add_190_195_groupi_g41369(csa_tree_add_190_195_groupi_n_7846 ,csa_tree_add_190_195_groupi_n_6232 ,csa_tree_add_190_195_groupi_n_7270);
  or csa_tree_add_190_195_groupi_g41370(csa_tree_add_190_195_groupi_n_7845 ,csa_tree_add_190_195_groupi_n_3061 ,csa_tree_add_190_195_groupi_n_7051);
  and csa_tree_add_190_195_groupi_g41371(csa_tree_add_190_195_groupi_n_7844 ,csa_tree_add_190_195_groupi_n_6381 ,csa_tree_add_190_195_groupi_n_7278);
  or csa_tree_add_190_195_groupi_g41372(csa_tree_add_190_195_groupi_n_7843 ,csa_tree_add_190_195_groupi_n_5741 ,csa_tree_add_190_195_groupi_n_7266);
  or csa_tree_add_190_195_groupi_g41373(csa_tree_add_190_195_groupi_n_7841 ,csa_tree_add_190_195_groupi_n_4878 ,csa_tree_add_190_195_groupi_n_7046);
  or csa_tree_add_190_195_groupi_g41374(csa_tree_add_190_195_groupi_n_7839 ,csa_tree_add_190_195_groupi_n_6141 ,csa_tree_add_190_195_groupi_n_7302);
  or csa_tree_add_190_195_groupi_g41375(csa_tree_add_190_195_groupi_n_7836 ,csa_tree_add_190_195_groupi_n_6858 ,csa_tree_add_190_195_groupi_n_7236);
  and csa_tree_add_190_195_groupi_g41376(csa_tree_add_190_195_groupi_n_7835 ,csa_tree_add_190_195_groupi_n_6492 ,csa_tree_add_190_195_groupi_n_7243);
  or csa_tree_add_190_195_groupi_g41377(csa_tree_add_190_195_groupi_n_7833 ,csa_tree_add_190_195_groupi_n_6487 ,csa_tree_add_190_195_groupi_n_7251);
  or csa_tree_add_190_195_groupi_g41378(csa_tree_add_190_195_groupi_n_7831 ,csa_tree_add_190_195_groupi_n_5702 ,csa_tree_add_190_195_groupi_n_7252);
  or csa_tree_add_190_195_groupi_g41379(csa_tree_add_190_195_groupi_n_7829 ,csa_tree_add_190_195_groupi_n_6401 ,csa_tree_add_190_195_groupi_n_7048);
  and csa_tree_add_190_195_groupi_g41380(csa_tree_add_190_195_groupi_n_7827 ,csa_tree_add_190_195_groupi_n_6154 ,csa_tree_add_190_195_groupi_n_7044);
  or csa_tree_add_190_195_groupi_g41381(csa_tree_add_190_195_groupi_n_7826 ,csa_tree_add_190_195_groupi_n_6361 ,csa_tree_add_190_195_groupi_n_7267);
  or csa_tree_add_190_195_groupi_g41382(csa_tree_add_190_195_groupi_n_7825 ,csa_tree_add_190_195_groupi_n_6329 ,csa_tree_add_190_195_groupi_n_7268);
  or csa_tree_add_190_195_groupi_g41383(csa_tree_add_190_195_groupi_n_7824 ,csa_tree_add_190_195_groupi_n_6731 ,csa_tree_add_190_195_groupi_n_7273);
  or csa_tree_add_190_195_groupi_g41384(csa_tree_add_190_195_groupi_n_7823 ,csa_tree_add_190_195_groupi_n_5770 ,csa_tree_add_190_195_groupi_n_7288);
  or csa_tree_add_190_195_groupi_g41385(csa_tree_add_190_195_groupi_n_7820 ,csa_tree_add_190_195_groupi_n_5794 ,csa_tree_add_190_195_groupi_n_7289);
  or csa_tree_add_190_195_groupi_g41386(csa_tree_add_190_195_groupi_n_7819 ,csa_tree_add_190_195_groupi_n_5624 ,csa_tree_add_190_195_groupi_n_7299);
  not csa_tree_add_190_195_groupi_g41387(csa_tree_add_190_195_groupi_n_7670 ,csa_tree_add_190_195_groupi_n_7669);
  not csa_tree_add_190_195_groupi_g41388(csa_tree_add_190_195_groupi_n_7668 ,csa_tree_add_190_195_groupi_n_7667);
  not csa_tree_add_190_195_groupi_g41389(csa_tree_add_190_195_groupi_n_7665 ,csa_tree_add_190_195_groupi_n_7664);
  not csa_tree_add_190_195_groupi_g41390(csa_tree_add_190_195_groupi_n_7645 ,csa_tree_add_190_195_groupi_n_7646);
  not csa_tree_add_190_195_groupi_g41391(csa_tree_add_190_195_groupi_n_7644 ,csa_tree_add_190_195_groupi_n_7643);
  not csa_tree_add_190_195_groupi_g41392(csa_tree_add_190_195_groupi_n_7641 ,csa_tree_add_190_195_groupi_n_7642);
  not csa_tree_add_190_195_groupi_g41393(csa_tree_add_190_195_groupi_n_7639 ,csa_tree_add_190_195_groupi_n_7640);
  not csa_tree_add_190_195_groupi_g41394(csa_tree_add_190_195_groupi_n_7636 ,csa_tree_add_190_195_groupi_n_7637);
  not csa_tree_add_190_195_groupi_g41395(csa_tree_add_190_195_groupi_n_7634 ,csa_tree_add_190_195_groupi_n_7635);
  not csa_tree_add_190_195_groupi_g41396(csa_tree_add_190_195_groupi_n_7630 ,csa_tree_add_190_195_groupi_n_7631);
  not csa_tree_add_190_195_groupi_g41397(csa_tree_add_190_195_groupi_n_7627 ,csa_tree_add_190_195_groupi_n_7628);
  not csa_tree_add_190_195_groupi_g41398(csa_tree_add_190_195_groupi_n_7626 ,csa_tree_add_190_195_groupi_n_7625);
  not csa_tree_add_190_195_groupi_g41399(csa_tree_add_190_195_groupi_n_7623 ,csa_tree_add_190_195_groupi_n_7624);
  not csa_tree_add_190_195_groupi_g41400(csa_tree_add_190_195_groupi_n_7621 ,csa_tree_add_190_195_groupi_n_7620);
  not csa_tree_add_190_195_groupi_g41401(csa_tree_add_190_195_groupi_n_7618 ,csa_tree_add_190_195_groupi_n_7619);
  not csa_tree_add_190_195_groupi_g41402(csa_tree_add_190_195_groupi_n_7617 ,csa_tree_add_190_195_groupi_n_7616);
  not csa_tree_add_190_195_groupi_g41403(csa_tree_add_190_195_groupi_n_7614 ,csa_tree_add_190_195_groupi_n_7613);
  not csa_tree_add_190_195_groupi_g41404(csa_tree_add_190_195_groupi_n_7611 ,csa_tree_add_190_195_groupi_n_7612);
  not csa_tree_add_190_195_groupi_g41405(csa_tree_add_190_195_groupi_n_7605 ,csa_tree_add_190_195_groupi_n_7606);
  not csa_tree_add_190_195_groupi_g41406(csa_tree_add_190_195_groupi_n_7604 ,csa_tree_add_190_195_groupi_n_89);
  not csa_tree_add_190_195_groupi_g41407(csa_tree_add_190_195_groupi_n_7602 ,csa_tree_add_190_195_groupi_n_7603);
  not csa_tree_add_190_195_groupi_g41408(csa_tree_add_190_195_groupi_n_7600 ,csa_tree_add_190_195_groupi_n_7601);
  not csa_tree_add_190_195_groupi_g41409(csa_tree_add_190_195_groupi_n_7595 ,csa_tree_add_190_195_groupi_n_7596);
  not csa_tree_add_190_195_groupi_g41410(csa_tree_add_190_195_groupi_n_7592 ,csa_tree_add_190_195_groupi_n_7593);
  not csa_tree_add_190_195_groupi_g41411(csa_tree_add_190_195_groupi_n_7590 ,csa_tree_add_190_195_groupi_n_7591);
  not csa_tree_add_190_195_groupi_g41412(csa_tree_add_190_195_groupi_n_7588 ,csa_tree_add_190_195_groupi_n_7589);
  not csa_tree_add_190_195_groupi_g41413(csa_tree_add_190_195_groupi_n_7587 ,csa_tree_add_190_195_groupi_n_7586);
  not csa_tree_add_190_195_groupi_g41414(csa_tree_add_190_195_groupi_n_7585 ,csa_tree_add_190_195_groupi_n_7584);
  not csa_tree_add_190_195_groupi_g41415(csa_tree_add_190_195_groupi_n_7581 ,csa_tree_add_190_195_groupi_n_7582);
  not csa_tree_add_190_195_groupi_g41416(csa_tree_add_190_195_groupi_n_7580 ,csa_tree_add_190_195_groupi_n_7579);
  not csa_tree_add_190_195_groupi_g41417(csa_tree_add_190_195_groupi_n_7578 ,csa_tree_add_190_195_groupi_n_7577);
  not csa_tree_add_190_195_groupi_g41418(csa_tree_add_190_195_groupi_n_7576 ,csa_tree_add_190_195_groupi_n_7575);
  not csa_tree_add_190_195_groupi_g41419(csa_tree_add_190_195_groupi_n_7572 ,csa_tree_add_190_195_groupi_n_7573);
  not csa_tree_add_190_195_groupi_g41420(csa_tree_add_190_195_groupi_n_7570 ,csa_tree_add_190_195_groupi_n_7571);
  not csa_tree_add_190_195_groupi_g41421(csa_tree_add_190_195_groupi_n_7569 ,csa_tree_add_190_195_groupi_n_7568);
  not csa_tree_add_190_195_groupi_g41422(csa_tree_add_190_195_groupi_n_7566 ,csa_tree_add_190_195_groupi_n_7567);
  not csa_tree_add_190_195_groupi_g41423(csa_tree_add_190_195_groupi_n_7563 ,csa_tree_add_190_195_groupi_n_7564);
  not csa_tree_add_190_195_groupi_g41424(csa_tree_add_190_195_groupi_n_7561 ,csa_tree_add_190_195_groupi_n_7562);
  not csa_tree_add_190_195_groupi_g41425(csa_tree_add_190_195_groupi_n_7559 ,csa_tree_add_190_195_groupi_n_7560);
  not csa_tree_add_190_195_groupi_g41426(csa_tree_add_190_195_groupi_n_7556 ,csa_tree_add_190_195_groupi_n_7557);
  not csa_tree_add_190_195_groupi_g41427(csa_tree_add_190_195_groupi_n_7554 ,csa_tree_add_190_195_groupi_n_7555);
  not csa_tree_add_190_195_groupi_g41428(csa_tree_add_190_195_groupi_n_7552 ,csa_tree_add_190_195_groupi_n_7553);
  not csa_tree_add_190_195_groupi_g41429(csa_tree_add_190_195_groupi_n_7550 ,csa_tree_add_190_195_groupi_n_7551);
  not csa_tree_add_190_195_groupi_g41430(csa_tree_add_190_195_groupi_n_7548 ,csa_tree_add_190_195_groupi_n_7549);
  not csa_tree_add_190_195_groupi_g41431(csa_tree_add_190_195_groupi_n_7546 ,csa_tree_add_190_195_groupi_n_7545);
  not csa_tree_add_190_195_groupi_g41432(csa_tree_add_190_195_groupi_n_7543 ,csa_tree_add_190_195_groupi_n_7544);
  not csa_tree_add_190_195_groupi_g41433(csa_tree_add_190_195_groupi_n_7542 ,csa_tree_add_190_195_groupi_n_7541);
  not csa_tree_add_190_195_groupi_g41434(csa_tree_add_190_195_groupi_n_7539 ,csa_tree_add_190_195_groupi_n_7538);
  not csa_tree_add_190_195_groupi_g41435(csa_tree_add_190_195_groupi_n_7533 ,csa_tree_add_190_195_groupi_n_7534);
  not csa_tree_add_190_195_groupi_g41436(csa_tree_add_190_195_groupi_n_7530 ,csa_tree_add_190_195_groupi_n_7531);
  not csa_tree_add_190_195_groupi_g41437(csa_tree_add_190_195_groupi_n_7528 ,csa_tree_add_190_195_groupi_n_7529);
  not csa_tree_add_190_195_groupi_g41438(csa_tree_add_190_195_groupi_n_7526 ,csa_tree_add_190_195_groupi_n_7527);
  not csa_tree_add_190_195_groupi_g41439(csa_tree_add_190_195_groupi_n_7523 ,csa_tree_add_190_195_groupi_n_7524);
  not csa_tree_add_190_195_groupi_g41440(csa_tree_add_190_195_groupi_n_7521 ,csa_tree_add_190_195_groupi_n_7522);
  not csa_tree_add_190_195_groupi_g41441(csa_tree_add_190_195_groupi_n_7519 ,csa_tree_add_190_195_groupi_n_7520);
  not csa_tree_add_190_195_groupi_g41442(csa_tree_add_190_195_groupi_n_7514 ,csa_tree_add_190_195_groupi_n_7515);
  not csa_tree_add_190_195_groupi_g41443(csa_tree_add_190_195_groupi_n_7512 ,csa_tree_add_190_195_groupi_n_7511);
  not csa_tree_add_190_195_groupi_g41444(csa_tree_add_190_195_groupi_n_7510 ,csa_tree_add_190_195_groupi_n_7509);
  not csa_tree_add_190_195_groupi_g41445(csa_tree_add_190_195_groupi_n_7507 ,csa_tree_add_190_195_groupi_n_7508);
  not csa_tree_add_190_195_groupi_g41446(csa_tree_add_190_195_groupi_n_7506 ,csa_tree_add_190_195_groupi_n_7505);
  not csa_tree_add_190_195_groupi_g41447(csa_tree_add_190_195_groupi_n_7503 ,csa_tree_add_190_195_groupi_n_7504);
  not csa_tree_add_190_195_groupi_g41448(csa_tree_add_190_195_groupi_n_7502 ,csa_tree_add_190_195_groupi_n_7501);
  not csa_tree_add_190_195_groupi_g41449(csa_tree_add_190_195_groupi_n_7499 ,csa_tree_add_190_195_groupi_n_7500);
  not csa_tree_add_190_195_groupi_g41450(csa_tree_add_190_195_groupi_n_7495 ,csa_tree_add_190_195_groupi_n_7496);
  not csa_tree_add_190_195_groupi_g41451(csa_tree_add_190_195_groupi_n_7494 ,csa_tree_add_190_195_groupi_n_7493);
  nor csa_tree_add_190_195_groupi_g41452(csa_tree_add_190_195_groupi_n_7492 ,csa_tree_add_190_195_groupi_n_3266 ,csa_tree_add_190_195_groupi_n_7385);
  or csa_tree_add_190_195_groupi_g41453(csa_tree_add_190_195_groupi_n_7491 ,csa_tree_add_190_195_groupi_n_6967 ,csa_tree_add_190_195_groupi_n_7178);
  nor csa_tree_add_190_195_groupi_g41454(csa_tree_add_190_195_groupi_n_7490 ,csa_tree_add_190_195_groupi_n_6968 ,csa_tree_add_190_195_groupi_n_7177);
  nor csa_tree_add_190_195_groupi_g41455(csa_tree_add_190_195_groupi_n_7489 ,csa_tree_add_190_195_groupi_n_7307 ,csa_tree_add_190_195_groupi_n_7080);
  or csa_tree_add_190_195_groupi_g41456(csa_tree_add_190_195_groupi_n_7488 ,csa_tree_add_190_195_groupi_n_6513 ,csa_tree_add_190_195_groupi_n_7431);
  and csa_tree_add_190_195_groupi_g41457(csa_tree_add_190_195_groupi_n_7487 ,csa_tree_add_190_195_groupi_n_6435 ,csa_tree_add_190_195_groupi_n_7215);
  or csa_tree_add_190_195_groupi_g41458(csa_tree_add_190_195_groupi_n_7486 ,csa_tree_add_190_195_groupi_n_6195 ,csa_tree_add_190_195_groupi_n_7208);
  nor csa_tree_add_190_195_groupi_g41459(csa_tree_add_190_195_groupi_n_7485 ,csa_tree_add_190_195_groupi_n_6931 ,csa_tree_add_190_195_groupi_n_7174);
  or csa_tree_add_190_195_groupi_g41460(csa_tree_add_190_195_groupi_n_7484 ,csa_tree_add_190_195_groupi_n_6985 ,csa_tree_add_190_195_groupi_n_7279);
  or csa_tree_add_190_195_groupi_g41461(csa_tree_add_190_195_groupi_n_7483 ,csa_tree_add_190_195_groupi_n_6328 ,csa_tree_add_190_195_groupi_n_7394);
  nor csa_tree_add_190_195_groupi_g41462(csa_tree_add_190_195_groupi_n_7482 ,csa_tree_add_190_195_groupi_n_6457 ,csa_tree_add_190_195_groupi_n_7214);
  and csa_tree_add_190_195_groupi_g41463(csa_tree_add_190_195_groupi_n_7481 ,csa_tree_add_190_195_groupi_n_7091 ,csa_tree_add_190_195_groupi_n_7134);
  or csa_tree_add_190_195_groupi_g41464(csa_tree_add_190_195_groupi_n_7480 ,csa_tree_add_190_195_groupi_n_7091 ,csa_tree_add_190_195_groupi_n_7134);
  or csa_tree_add_190_195_groupi_g41465(csa_tree_add_190_195_groupi_n_7479 ,csa_tree_add_190_195_groupi_n_6930 ,csa_tree_add_190_195_groupi_n_7173);
  nor csa_tree_add_190_195_groupi_g41466(csa_tree_add_190_195_groupi_n_7478 ,csa_tree_add_190_195_groupi_n_7117 ,csa_tree_add_190_195_groupi_n_7116);
  or csa_tree_add_190_195_groupi_g41467(csa_tree_add_190_195_groupi_n_7477 ,csa_tree_add_190_195_groupi_n_7118 ,csa_tree_add_190_195_groupi_n_7115);
  or csa_tree_add_190_195_groupi_g41468(csa_tree_add_190_195_groupi_n_7476 ,csa_tree_add_190_195_groupi_n_7306 ,csa_tree_add_190_195_groupi_n_7079);
  or csa_tree_add_190_195_groupi_g41469(csa_tree_add_190_195_groupi_n_7475 ,csa_tree_add_190_195_groupi_n_3228 ,csa_tree_add_190_195_groupi_n_86);
  xnor csa_tree_add_190_195_groupi_g41470(csa_tree_add_190_195_groupi_n_7474 ,csa_tree_add_190_195_groupi_n_7008 ,csa_tree_add_190_195_groupi_n_2156);
  xnor csa_tree_add_190_195_groupi_g41471(csa_tree_add_190_195_groupi_n_7473 ,csa_tree_add_190_195_groupi_n_5340 ,csa_tree_add_190_195_groupi_n_6992);
  xnor csa_tree_add_190_195_groupi_g41472(csa_tree_add_190_195_groupi_n_7472 ,csa_tree_add_190_195_groupi_n_6776 ,csa_tree_add_190_195_groupi_n_6770);
  xnor csa_tree_add_190_195_groupi_g41473(csa_tree_add_190_195_groupi_n_7471 ,csa_tree_add_190_195_groupi_n_4628 ,csa_tree_add_190_195_groupi_n_7014);
  xnor csa_tree_add_190_195_groupi_g41474(csa_tree_add_190_195_groupi_n_7470 ,csa_tree_add_190_195_groupi_n_7016 ,csa_tree_add_190_195_groupi_n_5278);
  xnor csa_tree_add_190_195_groupi_g41475(csa_tree_add_190_195_groupi_n_7469 ,csa_tree_add_190_195_groupi_n_4983 ,csa_tree_add_190_195_groupi_n_6982);
  xnor csa_tree_add_190_195_groupi_g41476(csa_tree_add_190_195_groupi_n_7468 ,csa_tree_add_190_195_groupi_n_4609 ,csa_tree_add_190_195_groupi_n_6772);
  xnor csa_tree_add_190_195_groupi_g41477(csa_tree_add_190_195_groupi_n_7467 ,csa_tree_add_190_195_groupi_n_6983 ,csa_tree_add_190_195_groupi_n_1960);
  xnor csa_tree_add_190_195_groupi_g41478(csa_tree_add_190_195_groupi_n_7466 ,csa_tree_add_190_195_groupi_n_4966 ,csa_tree_add_190_195_groupi_n_6989);
  xnor csa_tree_add_190_195_groupi_g41479(csa_tree_add_190_195_groupi_n_7465 ,csa_tree_add_190_195_groupi_n_6260 ,csa_tree_add_190_195_groupi_n_6784);
  xnor csa_tree_add_190_195_groupi_g41480(csa_tree_add_190_195_groupi_n_7464 ,csa_tree_add_190_195_groupi_n_5250 ,csa_tree_add_190_195_groupi_n_6958);
  xnor csa_tree_add_190_195_groupi_g41481(csa_tree_add_190_195_groupi_n_7463 ,csa_tree_add_190_195_groupi_n_6988 ,csa_tree_add_190_195_groupi_n_1143);
  xnor csa_tree_add_190_195_groupi_g41482(csa_tree_add_190_195_groupi_n_7462 ,csa_tree_add_190_195_groupi_n_6997 ,csa_tree_add_190_195_groupi_n_5266);
  xnor csa_tree_add_190_195_groupi_g41483(csa_tree_add_190_195_groupi_n_7461 ,csa_tree_add_190_195_groupi_n_6921 ,csa_tree_add_190_195_groupi_n_6966);
  xnor csa_tree_add_190_195_groupi_g41484(csa_tree_add_190_195_groupi_n_7460 ,csa_tree_add_190_195_groupi_n_56 ,csa_tree_add_190_195_groupi_n_6949);
  xnor csa_tree_add_190_195_groupi_g41485(csa_tree_add_190_195_groupi_n_7459 ,csa_tree_add_190_195_groupi_n_6914 ,csa_tree_add_190_195_groupi_n_6916);
  xnor csa_tree_add_190_195_groupi_g41486(csa_tree_add_190_195_groupi_n_7458 ,csa_tree_add_190_195_groupi_n_4988 ,csa_tree_add_190_195_groupi_n_6991);
  xnor csa_tree_add_190_195_groupi_g41487(csa_tree_add_190_195_groupi_n_7457 ,csa_tree_add_190_195_groupi_n_4952 ,csa_tree_add_190_195_groupi_n_6974);
  xnor csa_tree_add_190_195_groupi_g41488(csa_tree_add_190_195_groupi_n_7456 ,csa_tree_add_190_195_groupi_n_4915 ,csa_tree_add_190_195_groupi_n_6987);
  xnor csa_tree_add_190_195_groupi_g41489(csa_tree_add_190_195_groupi_n_7455 ,csa_tree_add_190_195_groupi_n_5077 ,csa_tree_add_190_195_groupi_n_6981);
  xnor csa_tree_add_190_195_groupi_g41490(csa_tree_add_190_195_groupi_n_7454 ,csa_tree_add_190_195_groupi_n_6777 ,csa_tree_add_190_195_groupi_n_865);
  xnor csa_tree_add_190_195_groupi_g41491(csa_tree_add_190_195_groupi_n_7453 ,csa_tree_add_190_195_groupi_n_4973 ,csa_tree_add_190_195_groupi_n_6995);
  xnor csa_tree_add_190_195_groupi_g41492(csa_tree_add_190_195_groupi_n_7452 ,csa_tree_add_190_195_groupi_n_5891 ,csa_tree_add_190_195_groupi_n_6765);
  xnor csa_tree_add_190_195_groupi_g41493(csa_tree_add_190_195_groupi_n_7451 ,csa_tree_add_190_195_groupi_n_6985 ,csa_tree_add_190_195_groupi_n_6945);
  xnor csa_tree_add_190_195_groupi_g41494(csa_tree_add_190_195_groupi_n_7450 ,csa_tree_add_190_195_groupi_n_6973 ,csa_tree_add_190_195_groupi_n_459);
  xnor csa_tree_add_190_195_groupi_g41495(csa_tree_add_190_195_groupi_n_7449 ,csa_tree_add_190_195_groupi_n_6778 ,csa_tree_add_190_195_groupi_n_5283);
  xnor csa_tree_add_190_195_groupi_g41497(csa_tree_add_190_195_groupi_n_7448 ,csa_tree_add_190_195_groupi_n_7002 ,csa_tree_add_190_195_groupi_n_4782);
  xnor csa_tree_add_190_195_groupi_g41498(csa_tree_add_190_195_groupi_n_7447 ,csa_tree_add_190_195_groupi_n_5957 ,csa_tree_add_190_195_groupi_n_7012);
  xnor csa_tree_add_190_195_groupi_g41499(csa_tree_add_190_195_groupi_n_7446 ,csa_tree_add_190_195_groupi_n_6950 ,csa_tree_add_190_195_groupi_n_6972);
  xnor csa_tree_add_190_195_groupi_g41500(csa_tree_add_190_195_groupi_n_7445 ,csa_tree_add_190_195_groupi_n_5016 ,csa_tree_add_190_195_groupi_n_7007);
  xnor csa_tree_add_190_195_groupi_g41501(csa_tree_add_190_195_groupi_n_7444 ,csa_tree_add_190_195_groupi_n_6575 ,csa_tree_add_190_195_groupi_n_6934);
  xnor csa_tree_add_190_195_groupi_g41502(csa_tree_add_190_195_groupi_n_7443 ,csa_tree_add_190_195_groupi_n_4136 ,csa_tree_add_190_195_groupi_n_6975);
  xnor csa_tree_add_190_195_groupi_g41503(csa_tree_add_190_195_groupi_n_7442 ,csa_tree_add_190_195_groupi_n_5538 ,csa_tree_add_190_195_groupi_n_7005);
  xnor csa_tree_add_190_195_groupi_g41504(csa_tree_add_190_195_groupi_n_7441 ,csa_tree_add_190_195_groupi_n_4892 ,csa_tree_add_190_195_groupi_n_7013);
  xnor csa_tree_add_190_195_groupi_g41505(csa_tree_add_190_195_groupi_n_7440 ,csa_tree_add_190_195_groupi_n_4623 ,csa_tree_add_190_195_groupi_n_6790);
  xnor csa_tree_add_190_195_groupi_g41506(csa_tree_add_190_195_groupi_n_7439 ,csa_tree_add_190_195_groupi_n_6278 ,csa_tree_add_190_195_groupi_n_35);
  xnor csa_tree_add_190_195_groupi_g41507(csa_tree_add_190_195_groupi_n_7438 ,csa_tree_add_190_195_groupi_n_4659 ,csa_tree_add_190_195_groupi_n_6786);
  xnor csa_tree_add_190_195_groupi_g41508(csa_tree_add_190_195_groupi_n_7437 ,csa_tree_add_190_195_groupi_n_6789 ,csa_tree_add_190_195_groupi_n_5442);
  xnor csa_tree_add_190_195_groupi_g41509(csa_tree_add_190_195_groupi_n_7436 ,csa_tree_add_190_195_groupi_n_4920 ,csa_tree_add_190_195_groupi_n_6781);
  xnor csa_tree_add_190_195_groupi_g41510(csa_tree_add_190_195_groupi_n_7435 ,csa_tree_add_190_195_groupi_n_4669 ,csa_tree_add_190_195_groupi_n_6978);
  xnor csa_tree_add_190_195_groupi_g41511(csa_tree_add_190_195_groupi_n_7434 ,csa_tree_add_190_195_groupi_n_6276 ,csa_tree_add_190_195_groupi_n_6932);
  xnor csa_tree_add_190_195_groupi_g41512(csa_tree_add_190_195_groupi_n_7433 ,csa_tree_add_190_195_groupi_n_4791 ,csa_tree_add_190_195_groupi_n_7004);
  xnor csa_tree_add_190_195_groupi_g41513(csa_tree_add_190_195_groupi_n_7432 ,csa_tree_add_190_195_groupi_n_5879 ,csa_tree_add_190_195_groupi_n_6971);
  xnor csa_tree_add_190_195_groupi_g41514(csa_tree_add_190_195_groupi_n_7676 ,csa_tree_add_190_195_groupi_n_6596 ,csa_tree_add_190_195_groupi_n_1170);
  xnor csa_tree_add_190_195_groupi_g41515(csa_tree_add_190_195_groupi_n_7675 ,csa_tree_add_190_195_groupi_n_6716 ,csa_tree_add_190_195_groupi_n_1750);
  or csa_tree_add_190_195_groupi_g41516(csa_tree_add_190_195_groupi_n_7674 ,csa_tree_add_190_195_groupi_n_3358 ,csa_tree_add_190_195_groupi_n_7039);
  xnor csa_tree_add_190_195_groupi_g41517(csa_tree_add_190_195_groupi_n_7673 ,csa_tree_add_190_195_groupi_n_5504 ,csa_tree_add_190_195_groupi_n_6721);
  xnor csa_tree_add_190_195_groupi_g41518(csa_tree_add_190_195_groupi_n_7672 ,csa_tree_add_190_195_groupi_n_4135 ,csa_tree_add_190_195_groupi_n_6698);
  xnor csa_tree_add_190_195_groupi_g41519(csa_tree_add_190_195_groupi_n_7671 ,csa_tree_add_190_195_groupi_n_5263 ,csa_tree_add_190_195_groupi_n_6697);
  or csa_tree_add_190_195_groupi_g41520(csa_tree_add_190_195_groupi_n_7669 ,csa_tree_add_190_195_groupi_n_5842 ,csa_tree_add_190_195_groupi_n_7036);
  xnor csa_tree_add_190_195_groupi_g41521(csa_tree_add_190_195_groupi_n_7667 ,csa_tree_add_190_195_groupi_n_4978 ,csa_tree_add_190_195_groupi_n_6637);
  xnor csa_tree_add_190_195_groupi_g41522(csa_tree_add_190_195_groupi_n_7666 ,csa_tree_add_190_195_groupi_n_5553 ,csa_tree_add_190_195_groupi_n_6691);
  xnor csa_tree_add_190_195_groupi_g41524(csa_tree_add_190_195_groupi_n_7664 ,csa_tree_add_190_195_groupi_n_6656 ,csa_tree_add_190_195_groupi_n_2059);
  and csa_tree_add_190_195_groupi_g41525(csa_tree_add_190_195_groupi_n_7663 ,csa_tree_add_190_195_groupi_n_3408 ,csa_tree_add_190_195_groupi_n_7038);
  xnor csa_tree_add_190_195_groupi_g41527(csa_tree_add_190_195_groupi_n_7662 ,csa_tree_add_190_195_groupi_n_4127 ,csa_tree_add_190_195_groupi_n_6605);
  xnor csa_tree_add_190_195_groupi_g41528(csa_tree_add_190_195_groupi_n_7661 ,csa_tree_add_190_195_groupi_n_5579 ,csa_tree_add_190_195_groupi_n_6704);
  xnor csa_tree_add_190_195_groupi_g41529(csa_tree_add_190_195_groupi_n_7660 ,csa_tree_add_190_195_groupi_n_6669 ,csa_tree_add_190_195_groupi_n_2117);
  xnor csa_tree_add_190_195_groupi_g41530(csa_tree_add_190_195_groupi_n_7659 ,csa_tree_add_190_195_groupi_n_5944 ,csa_tree_add_190_195_groupi_n_6682);
  xnor csa_tree_add_190_195_groupi_g41531(csa_tree_add_190_195_groupi_n_7658 ,csa_tree_add_190_195_groupi_n_57 ,csa_tree_add_190_195_groupi_n_1749);
  xnor csa_tree_add_190_195_groupi_g41532(csa_tree_add_190_195_groupi_n_7657 ,csa_tree_add_190_195_groupi_n_5541 ,csa_tree_add_190_195_groupi_n_6661);
  xnor csa_tree_add_190_195_groupi_g41533(csa_tree_add_190_195_groupi_n_7656 ,csa_tree_add_190_195_groupi_n_7011 ,csa_tree_add_190_195_groupi_n_6673);
  xnor csa_tree_add_190_195_groupi_g41534(csa_tree_add_190_195_groupi_n_7655 ,csa_tree_add_190_195_groupi_n_5151 ,csa_tree_add_190_195_groupi_n_6623);
  xnor csa_tree_add_190_195_groupi_g41535(csa_tree_add_190_195_groupi_n_7654 ,csa_tree_add_190_195_groupi_n_4565 ,csa_tree_add_190_195_groupi_n_6648);
  xnor csa_tree_add_190_195_groupi_g41536(csa_tree_add_190_195_groupi_n_7653 ,csa_tree_add_190_195_groupi_n_5419 ,csa_tree_add_190_195_groupi_n_6677);
  xnor csa_tree_add_190_195_groupi_g41537(csa_tree_add_190_195_groupi_n_7652 ,csa_tree_add_190_195_groupi_n_6662 ,csa_tree_add_190_195_groupi_n_1691);
  xnor csa_tree_add_190_195_groupi_g41538(csa_tree_add_190_195_groupi_n_7651 ,csa_tree_add_190_195_groupi_n_5557 ,csa_tree_add_190_195_groupi_n_6707);
  xnor csa_tree_add_190_195_groupi_g41539(csa_tree_add_190_195_groupi_n_7650 ,csa_tree_add_190_195_groupi_n_18 ,csa_tree_add_190_195_groupi_n_6650);
  xnor csa_tree_add_190_195_groupi_g41540(csa_tree_add_190_195_groupi_n_7649 ,csa_tree_add_190_195_groupi_n_6645 ,csa_tree_add_190_195_groupi_n_1928);
  xnor csa_tree_add_190_195_groupi_g41541(csa_tree_add_190_195_groupi_n_7648 ,csa_tree_add_190_195_groupi_n_5379 ,csa_tree_add_190_195_groupi_n_6634);
  xnor csa_tree_add_190_195_groupi_g41542(csa_tree_add_190_195_groupi_n_7647 ,csa_tree_add_190_195_groupi_n_6977 ,csa_tree_add_190_195_groupi_n_4087);
  xnor csa_tree_add_190_195_groupi_g41543(csa_tree_add_190_195_groupi_n_7646 ,csa_tree_add_190_195_groupi_n_6980 ,csa_tree_add_190_195_groupi_n_6722);
  and csa_tree_add_190_195_groupi_g41544(csa_tree_add_190_195_groupi_n_7643 ,csa_tree_add_190_195_groupi_n_5662 ,csa_tree_add_190_195_groupi_n_7047);
  xnor csa_tree_add_190_195_groupi_g41545(csa_tree_add_190_195_groupi_n_7642 ,csa_tree_add_190_195_groupi_n_5117 ,csa_tree_add_190_195_groupi_n_79);
  xnor csa_tree_add_190_195_groupi_g41546(csa_tree_add_190_195_groupi_n_7640 ,csa_tree_add_190_195_groupi_n_5872 ,csa_tree_add_190_195_groupi_n_6705);
  xnor csa_tree_add_190_195_groupi_g41547(csa_tree_add_190_195_groupi_n_7638 ,csa_tree_add_190_195_groupi_n_5968 ,csa_tree_add_190_195_groupi_n_6713);
  xnor csa_tree_add_190_195_groupi_g41548(csa_tree_add_190_195_groupi_n_7637 ,csa_tree_add_190_195_groupi_n_5932 ,csa_tree_add_190_195_groupi_n_6593);
  xnor csa_tree_add_190_195_groupi_g41549(csa_tree_add_190_195_groupi_n_7635 ,csa_tree_add_190_195_groupi_n_5252 ,csa_tree_add_190_195_groupi_n_6644);
  xnor csa_tree_add_190_195_groupi_g41550(csa_tree_add_190_195_groupi_n_7633 ,csa_tree_add_190_195_groupi_n_6626 ,csa_tree_add_190_195_groupi_n_943);
  xnor csa_tree_add_190_195_groupi_g41551(csa_tree_add_190_195_groupi_n_7632 ,csa_tree_add_190_195_groupi_n_6970 ,csa_tree_add_190_195_groupi_n_6026);
  xnor csa_tree_add_190_195_groupi_g41552(csa_tree_add_190_195_groupi_n_7631 ,csa_tree_add_190_195_groupi_n_5491 ,csa_tree_add_190_195_groupi_n_6709);
  xnor csa_tree_add_190_195_groupi_g41553(csa_tree_add_190_195_groupi_n_7629 ,csa_tree_add_190_195_groupi_n_5349 ,csa_tree_add_190_195_groupi_n_6629);
  xnor csa_tree_add_190_195_groupi_g41554(csa_tree_add_190_195_groupi_n_7628 ,csa_tree_add_190_195_groupi_n_5185 ,csa_tree_add_190_195_groupi_n_6694);
  xnor csa_tree_add_190_195_groupi_g41555(csa_tree_add_190_195_groupi_n_7625 ,csa_tree_add_190_195_groupi_n_5127 ,csa_tree_add_190_195_groupi_n_6632);
  xnor csa_tree_add_190_195_groupi_g41556(csa_tree_add_190_195_groupi_n_7624 ,csa_tree_add_190_195_groupi_n_32 ,csa_tree_add_190_195_groupi_n_6701);
  xor csa_tree_add_190_195_groupi_g41557(csa_tree_add_190_195_groupi_n_7622 ,csa_tree_add_190_195_groupi_n_5969 ,csa_tree_add_190_195_groupi_n_6718);
  xnor csa_tree_add_190_195_groupi_g41558(csa_tree_add_190_195_groupi_n_7620 ,csa_tree_add_190_195_groupi_n_5593 ,csa_tree_add_190_195_groupi_n_6678);
  xnor csa_tree_add_190_195_groupi_g41559(csa_tree_add_190_195_groupi_n_7619 ,csa_tree_add_190_195_groupi_n_5269 ,csa_tree_add_190_195_groupi_n_6690);
  xnor csa_tree_add_190_195_groupi_g41560(csa_tree_add_190_195_groupi_n_7616 ,csa_tree_add_190_195_groupi_n_4705 ,csa_tree_add_190_195_groupi_n_87);
  xnor csa_tree_add_190_195_groupi_g41561(csa_tree_add_190_195_groupi_n_7615 ,csa_tree_add_190_195_groupi_n_7000 ,csa_tree_add_190_195_groupi_n_6084);
  xnor csa_tree_add_190_195_groupi_g41562(csa_tree_add_190_195_groupi_n_7613 ,csa_tree_add_190_195_groupi_n_4820 ,csa_tree_add_190_195_groupi_n_6630);
  xnor csa_tree_add_190_195_groupi_g41563(csa_tree_add_190_195_groupi_n_7612 ,csa_tree_add_190_195_groupi_n_7001 ,csa_tree_add_190_195_groupi_n_5993);
  xnor csa_tree_add_190_195_groupi_g41564(csa_tree_add_190_195_groupi_n_7610 ,csa_tree_add_190_195_groupi_n_5157 ,csa_tree_add_190_195_groupi_n_6627);
  xnor csa_tree_add_190_195_groupi_g41565(csa_tree_add_190_195_groupi_n_7609 ,csa_tree_add_190_195_groupi_n_4872 ,csa_tree_add_190_195_groupi_n_6653);
  xnor csa_tree_add_190_195_groupi_g41566(csa_tree_add_190_195_groupi_n_7608 ,csa_tree_add_190_195_groupi_n_6779 ,csa_tree_add_190_195_groupi_n_6028);
  xnor csa_tree_add_190_195_groupi_g41567(csa_tree_add_190_195_groupi_n_7607 ,csa_tree_add_190_195_groupi_n_5129 ,csa_tree_add_190_195_groupi_n_6652);
  xnor csa_tree_add_190_195_groupi_g41568(csa_tree_add_190_195_groupi_n_7606 ,csa_tree_add_190_195_groupi_n_5895 ,csa_tree_add_190_195_groupi_n_19);
  xnor csa_tree_add_190_195_groupi_g41570(csa_tree_add_190_195_groupi_n_7603 ,csa_tree_add_190_195_groupi_n_5411 ,csa_tree_add_190_195_groupi_n_6676);
  xnor csa_tree_add_190_195_groupi_g41571(csa_tree_add_190_195_groupi_n_7601 ,csa_tree_add_190_195_groupi_n_6787 ,csa_tree_add_190_195_groupi_n_6687);
  xnor csa_tree_add_190_195_groupi_g41572(csa_tree_add_190_195_groupi_n_7599 ,csa_tree_add_190_195_groupi_n_4621 ,csa_tree_add_190_195_groupi_n_6636);
  xnor csa_tree_add_190_195_groupi_g41573(csa_tree_add_190_195_groupi_n_7598 ,csa_tree_add_190_195_groupi_n_5896 ,csa_tree_add_190_195_groupi_n_6624);
  xnor csa_tree_add_190_195_groupi_g41574(csa_tree_add_190_195_groupi_n_7597 ,csa_tree_add_190_195_groupi_n_26 ,csa_tree_add_190_195_groupi_n_6639);
  xnor csa_tree_add_190_195_groupi_g41575(csa_tree_add_190_195_groupi_n_7596 ,csa_tree_add_190_195_groupi_n_5556 ,csa_tree_add_190_195_groupi_n_6688);
  xnor csa_tree_add_190_195_groupi_g41576(csa_tree_add_190_195_groupi_n_7594 ,csa_tree_add_190_195_groupi_n_5607 ,csa_tree_add_190_195_groupi_n_6638);
  xnor csa_tree_add_190_195_groupi_g41577(csa_tree_add_190_195_groupi_n_7593 ,csa_tree_add_190_195_groupi_n_5877 ,csa_tree_add_190_195_groupi_n_6602);
  xnor csa_tree_add_190_195_groupi_g41578(csa_tree_add_190_195_groupi_n_7591 ,csa_tree_add_190_195_groupi_n_4640 ,csa_tree_add_190_195_groupi_n_6598);
  xnor csa_tree_add_190_195_groupi_g41579(csa_tree_add_190_195_groupi_n_7589 ,csa_tree_add_190_195_groupi_n_5962 ,csa_tree_add_190_195_groupi_n_6719);
  xnor csa_tree_add_190_195_groupi_g41580(csa_tree_add_190_195_groupi_n_7586 ,csa_tree_add_190_195_groupi_n_4566 ,csa_tree_add_190_195_groupi_n_6625);
  xnor csa_tree_add_190_195_groupi_g41581(csa_tree_add_190_195_groupi_n_7584 ,csa_tree_add_190_195_groupi_n_5156 ,csa_tree_add_190_195_groupi_n_6640);
  xnor csa_tree_add_190_195_groupi_g41582(csa_tree_add_190_195_groupi_n_7583 ,csa_tree_add_190_195_groupi_n_4618 ,csa_tree_add_190_195_groupi_n_6649);
  xnor csa_tree_add_190_195_groupi_g41583(csa_tree_add_190_195_groupi_n_7582 ,csa_tree_add_190_195_groupi_n_5103 ,csa_tree_add_190_195_groupi_n_6685);
  or csa_tree_add_190_195_groupi_g41584(csa_tree_add_190_195_groupi_n_7579 ,csa_tree_add_190_195_groupi_n_6419 ,csa_tree_add_190_195_groupi_n_7035);
  xnor csa_tree_add_190_195_groupi_g41585(csa_tree_add_190_195_groupi_n_7577 ,csa_tree_add_190_195_groupi_n_4605 ,csa_tree_add_190_195_groupi_n_6702);
  xnor csa_tree_add_190_195_groupi_g41586(csa_tree_add_190_195_groupi_n_7575 ,csa_tree_add_190_195_groupi_n_4746 ,csa_tree_add_190_195_groupi_n_6700);
  xnor csa_tree_add_190_195_groupi_g41587(csa_tree_add_190_195_groupi_n_7574 ,csa_tree_add_190_195_groupi_n_5552 ,csa_tree_add_190_195_groupi_n_6597);
  xnor csa_tree_add_190_195_groupi_g41588(csa_tree_add_190_195_groupi_n_7573 ,csa_tree_add_190_195_groupi_n_6699 ,csa_tree_add_190_195_groupi_n_1847);
  xnor csa_tree_add_190_195_groupi_g41589(csa_tree_add_190_195_groupi_n_7571 ,csa_tree_add_190_195_groupi_n_6594 ,csa_tree_add_190_195_groupi_n_1099);
  xnor csa_tree_add_190_195_groupi_g41590(csa_tree_add_190_195_groupi_n_7568 ,csa_tree_add_190_195_groupi_n_4853 ,csa_tree_add_190_195_groupi_n_6631);
  xnor csa_tree_add_190_195_groupi_g41591(csa_tree_add_190_195_groupi_n_7567 ,csa_tree_add_190_195_groupi_n_5528 ,csa_tree_add_190_195_groupi_n_6651);
  or csa_tree_add_190_195_groupi_g41592(csa_tree_add_190_195_groupi_n_7565 ,csa_tree_add_190_195_groupi_n_6353 ,csa_tree_add_190_195_groupi_n_7060);
  xnor csa_tree_add_190_195_groupi_g41593(csa_tree_add_190_195_groupi_n_7564 ,csa_tree_add_190_195_groupi_n_6599 ,csa_tree_add_190_195_groupi_n_1077);
  xnor csa_tree_add_190_195_groupi_g41594(csa_tree_add_190_195_groupi_n_7562 ,csa_tree_add_190_195_groupi_n_5583 ,csa_tree_add_190_195_groupi_n_6610);
  xnor csa_tree_add_190_195_groupi_g41595(csa_tree_add_190_195_groupi_n_7560 ,csa_tree_add_190_195_groupi_n_4825 ,csa_tree_add_190_195_groupi_n_6608);
  xnor csa_tree_add_190_195_groupi_g41596(csa_tree_add_190_195_groupi_n_7558 ,csa_tree_add_190_195_groupi_n_4134 ,csa_tree_add_190_195_groupi_n_6655);
  xnor csa_tree_add_190_195_groupi_g41597(csa_tree_add_190_195_groupi_n_7557 ,csa_tree_add_190_195_groupi_n_24 ,csa_tree_add_190_195_groupi_n_6603);
  xnor csa_tree_add_190_195_groupi_g41598(csa_tree_add_190_195_groupi_n_7555 ,csa_tree_add_190_195_groupi_n_5385 ,csa_tree_add_190_195_groupi_n_6601);
  xnor csa_tree_add_190_195_groupi_g41599(csa_tree_add_190_195_groupi_n_7553 ,csa_tree_add_190_195_groupi_n_16 ,csa_tree_add_190_195_groupi_n_6672);
  xnor csa_tree_add_190_195_groupi_g41600(csa_tree_add_190_195_groupi_n_7551 ,csa_tree_add_190_195_groupi_n_5961 ,csa_tree_add_190_195_groupi_n_6607);
  xnor csa_tree_add_190_195_groupi_g41601(csa_tree_add_190_195_groupi_n_7549 ,csa_tree_add_190_195_groupi_n_6580 ,csa_tree_add_190_195_groupi_n_6595);
  xnor csa_tree_add_190_195_groupi_g41602(csa_tree_add_190_195_groupi_n_7547 ,csa_tree_add_190_195_groupi_n_6679 ,csa_tree_add_190_195_groupi_n_2057);
  xnor csa_tree_add_190_195_groupi_g41603(csa_tree_add_190_195_groupi_n_7545 ,csa_tree_add_190_195_groupi_n_5559 ,csa_tree_add_190_195_groupi_n_6695);
  xnor csa_tree_add_190_195_groupi_g41604(csa_tree_add_190_195_groupi_n_7544 ,csa_tree_add_190_195_groupi_n_6663 ,csa_tree_add_190_195_groupi_n_1868);
  xnor csa_tree_add_190_195_groupi_g41605(csa_tree_add_190_195_groupi_n_7541 ,csa_tree_add_190_195_groupi_n_49 ,csa_tree_add_190_195_groupi_n_6675);
  xnor csa_tree_add_190_195_groupi_g41606(csa_tree_add_190_195_groupi_n_7540 ,csa_tree_add_190_195_groupi_n_6712 ,csa_tree_add_190_195_groupi_n_1816);
  xnor csa_tree_add_190_195_groupi_g41607(csa_tree_add_190_195_groupi_n_7538 ,csa_tree_add_190_195_groupi_n_5918 ,csa_tree_add_190_195_groupi_n_6600);
  xnor csa_tree_add_190_195_groupi_g41608(csa_tree_add_190_195_groupi_n_7537 ,csa_tree_add_190_195_groupi_n_6671 ,csa_tree_add_190_195_groupi_n_589);
  xnor csa_tree_add_190_195_groupi_g41609(csa_tree_add_190_195_groupi_n_7536 ,csa_tree_add_190_195_groupi_n_6670 ,csa_tree_add_190_195_groupi_n_1751);
  xnor csa_tree_add_190_195_groupi_g41610(csa_tree_add_190_195_groupi_n_7535 ,csa_tree_add_190_195_groupi_n_23 ,csa_tree_add_190_195_groupi_n_1962);
  xnor csa_tree_add_190_195_groupi_g41611(csa_tree_add_190_195_groupi_n_7534 ,csa_tree_add_190_195_groupi_n_6782 ,csa_tree_add_190_195_groupi_n_6667);
  xnor csa_tree_add_190_195_groupi_g41612(csa_tree_add_190_195_groupi_n_7532 ,csa_tree_add_190_195_groupi_n_5408 ,csa_tree_add_190_195_groupi_n_6635);
  xnor csa_tree_add_190_195_groupi_g41613(csa_tree_add_190_195_groupi_n_7531 ,csa_tree_add_190_195_groupi_n_5609 ,csa_tree_add_190_195_groupi_n_6664);
  xnor csa_tree_add_190_195_groupi_g41614(csa_tree_add_190_195_groupi_n_7529 ,csa_tree_add_190_195_groupi_n_5170 ,csa_tree_add_190_195_groupi_n_6622);
  xnor csa_tree_add_190_195_groupi_g41615(csa_tree_add_190_195_groupi_n_7527 ,csa_tree_add_190_195_groupi_n_4686 ,csa_tree_add_190_195_groupi_n_6660);
  xnor csa_tree_add_190_195_groupi_g41616(csa_tree_add_190_195_groupi_n_7525 ,csa_tree_add_190_195_groupi_n_5378 ,csa_tree_add_190_195_groupi_n_6674);
  xnor csa_tree_add_190_195_groupi_g41617(csa_tree_add_190_195_groupi_n_7524 ,csa_tree_add_190_195_groupi_n_4817 ,csa_tree_add_190_195_groupi_n_6606);
  xnor csa_tree_add_190_195_groupi_g41618(csa_tree_add_190_195_groupi_n_7522 ,csa_tree_add_190_195_groupi_n_6274 ,csa_tree_add_190_195_groupi_n_6614);
  xnor csa_tree_add_190_195_groupi_g41619(csa_tree_add_190_195_groupi_n_7520 ,csa_tree_add_190_195_groupi_n_5259 ,csa_tree_add_190_195_groupi_n_6612);
  xnor csa_tree_add_190_195_groupi_g41620(csa_tree_add_190_195_groupi_n_7518 ,csa_tree_add_190_195_groupi_n_4991 ,csa_tree_add_190_195_groupi_n_6686);
  xnor csa_tree_add_190_195_groupi_g41621(csa_tree_add_190_195_groupi_n_7517 ,csa_tree_add_190_195_groupi_n_5243 ,csa_tree_add_190_195_groupi_n_6618);
  xor csa_tree_add_190_195_groupi_g41622(csa_tree_add_190_195_groupi_n_7516 ,csa_tree_add_190_195_groupi_n_5586 ,csa_tree_add_190_195_groupi_n_6654);
  xnor csa_tree_add_190_195_groupi_g41623(csa_tree_add_190_195_groupi_n_7515 ,csa_tree_add_190_195_groupi_n_5887 ,csa_tree_add_190_195_groupi_n_6692);
  xnor csa_tree_add_190_195_groupi_g41624(csa_tree_add_190_195_groupi_n_7513 ,csa_tree_add_190_195_groupi_n_5546 ,csa_tree_add_190_195_groupi_n_6657);
  xnor csa_tree_add_190_195_groupi_g41625(csa_tree_add_190_195_groupi_n_7511 ,csa_tree_add_190_195_groupi_n_6783 ,csa_tree_add_190_195_groupi_n_6033);
  xnor csa_tree_add_190_195_groupi_g41626(csa_tree_add_190_195_groupi_n_7509 ,csa_tree_add_190_195_groupi_n_5558 ,csa_tree_add_190_195_groupi_n_6714);
  xnor csa_tree_add_190_195_groupi_g41627(csa_tree_add_190_195_groupi_n_7508 ,csa_tree_add_190_195_groupi_n_6788 ,csa_tree_add_190_195_groupi_n_6715);
  xnor csa_tree_add_190_195_groupi_g41628(csa_tree_add_190_195_groupi_n_7505 ,csa_tree_add_190_195_groupi_n_4870 ,csa_tree_add_190_195_groupi_n_6628);
  xnor csa_tree_add_190_195_groupi_g41629(csa_tree_add_190_195_groupi_n_7504 ,csa_tree_add_190_195_groupi_n_5549 ,csa_tree_add_190_195_groupi_n_6646);
  xnor csa_tree_add_190_195_groupi_g41630(csa_tree_add_190_195_groupi_n_7501 ,csa_tree_add_190_195_groupi_n_4863 ,csa_tree_add_190_195_groupi_n_6633);
  xnor csa_tree_add_190_195_groupi_g41631(csa_tree_add_190_195_groupi_n_7500 ,csa_tree_add_190_195_groupi_n_5110 ,csa_tree_add_190_195_groupi_n_6620);
  xnor csa_tree_add_190_195_groupi_g41632(csa_tree_add_190_195_groupi_n_7498 ,csa_tree_add_190_195_groupi_n_6780 ,csa_tree_add_190_195_groupi_n_6684);
  xnor csa_tree_add_190_195_groupi_g41633(csa_tree_add_190_195_groupi_n_7497 ,csa_tree_add_190_195_groupi_n_5225 ,csa_tree_add_190_195_groupi_n_6710);
  xnor csa_tree_add_190_195_groupi_g41634(csa_tree_add_190_195_groupi_n_7496 ,csa_tree_add_190_195_groupi_n_5588 ,csa_tree_add_190_195_groupi_n_6706);
  xnor csa_tree_add_190_195_groupi_g41635(csa_tree_add_190_195_groupi_n_7493 ,csa_tree_add_190_195_groupi_n_6986 ,csa_tree_add_190_195_groupi_n_6604);
  not csa_tree_add_190_195_groupi_g41637(csa_tree_add_190_195_groupi_n_7427 ,csa_tree_add_190_195_groupi_n_7426);
  not csa_tree_add_190_195_groupi_g41639(csa_tree_add_190_195_groupi_n_7421 ,csa_tree_add_190_195_groupi_n_7420);
  not csa_tree_add_190_195_groupi_g41641(csa_tree_add_190_195_groupi_n_7393 ,csa_tree_add_190_195_groupi_n_7392);
  not csa_tree_add_190_195_groupi_g41643(csa_tree_add_190_195_groupi_n_7384 ,csa_tree_add_190_195_groupi_n_7383);
  not csa_tree_add_190_195_groupi_g41644(csa_tree_add_190_195_groupi_n_7379 ,csa_tree_add_190_195_groupi_n_7380);
  not csa_tree_add_190_195_groupi_g41645(csa_tree_add_190_195_groupi_n_7377 ,csa_tree_add_190_195_groupi_n_7376);
  not csa_tree_add_190_195_groupi_g41646(csa_tree_add_190_195_groupi_n_7374 ,csa_tree_add_190_195_groupi_n_7375);
  not csa_tree_add_190_195_groupi_g41647(csa_tree_add_190_195_groupi_n_7371 ,csa_tree_add_190_195_groupi_n_7372);
  not csa_tree_add_190_195_groupi_g41648(csa_tree_add_190_195_groupi_n_7369 ,csa_tree_add_190_195_groupi_n_7370);
  not csa_tree_add_190_195_groupi_g41649(csa_tree_add_190_195_groupi_n_7367 ,csa_tree_add_190_195_groupi_n_7368);
  not csa_tree_add_190_195_groupi_g41650(csa_tree_add_190_195_groupi_n_7365 ,csa_tree_add_190_195_groupi_n_7366);
  not csa_tree_add_190_195_groupi_g41651(csa_tree_add_190_195_groupi_n_7361 ,csa_tree_add_190_195_groupi_n_7362);
  not csa_tree_add_190_195_groupi_g41652(csa_tree_add_190_195_groupi_n_7360 ,csa_tree_add_190_195_groupi_n_7359);
  not csa_tree_add_190_195_groupi_g41653(csa_tree_add_190_195_groupi_n_7357 ,csa_tree_add_190_195_groupi_n_7358);
  not csa_tree_add_190_195_groupi_g41654(csa_tree_add_190_195_groupi_n_7355 ,csa_tree_add_190_195_groupi_n_7356);
  not csa_tree_add_190_195_groupi_g41655(csa_tree_add_190_195_groupi_n_7349 ,csa_tree_add_190_195_groupi_n_7350);
  not csa_tree_add_190_195_groupi_g41656(csa_tree_add_190_195_groupi_n_7348 ,csa_tree_add_190_195_groupi_n_7347);
  not csa_tree_add_190_195_groupi_g41657(csa_tree_add_190_195_groupi_n_7345 ,csa_tree_add_190_195_groupi_n_7346);
  not csa_tree_add_190_195_groupi_g41658(csa_tree_add_190_195_groupi_n_7344 ,csa_tree_add_190_195_groupi_n_7343);
  not csa_tree_add_190_195_groupi_g41659(csa_tree_add_190_195_groupi_n_7340 ,csa_tree_add_190_195_groupi_n_7341);
  not csa_tree_add_190_195_groupi_g41660(csa_tree_add_190_195_groupi_n_7337 ,csa_tree_add_190_195_groupi_n_7338);
  not csa_tree_add_190_195_groupi_g41661(csa_tree_add_190_195_groupi_n_7335 ,csa_tree_add_190_195_groupi_n_7336);
  not csa_tree_add_190_195_groupi_g41662(csa_tree_add_190_195_groupi_n_7333 ,csa_tree_add_190_195_groupi_n_7334);
  not csa_tree_add_190_195_groupi_g41663(csa_tree_add_190_195_groupi_n_7331 ,csa_tree_add_190_195_groupi_n_7332);
  not csa_tree_add_190_195_groupi_g41664(csa_tree_add_190_195_groupi_n_7329 ,csa_tree_add_190_195_groupi_n_7328);
  not csa_tree_add_190_195_groupi_g41665(csa_tree_add_190_195_groupi_n_7326 ,csa_tree_add_190_195_groupi_n_7327);
  not csa_tree_add_190_195_groupi_g41666(csa_tree_add_190_195_groupi_n_7324 ,csa_tree_add_190_195_groupi_n_7325);
  not csa_tree_add_190_195_groupi_g41667(csa_tree_add_190_195_groupi_n_7322 ,csa_tree_add_190_195_groupi_n_7323);
  not csa_tree_add_190_195_groupi_g41668(csa_tree_add_190_195_groupi_n_7321 ,csa_tree_add_190_195_groupi_n_7320);
  not csa_tree_add_190_195_groupi_g41669(csa_tree_add_190_195_groupi_n_7319 ,csa_tree_add_190_195_groupi_n_7318);
  not csa_tree_add_190_195_groupi_g41670(csa_tree_add_190_195_groupi_n_7311 ,csa_tree_add_190_195_groupi_n_7312);
  not csa_tree_add_190_195_groupi_g41671(csa_tree_add_190_195_groupi_n_7310 ,csa_tree_add_190_195_groupi_n_7309);
  not csa_tree_add_190_195_groupi_g41672(csa_tree_add_190_195_groupi_n_7307 ,csa_tree_add_190_195_groupi_n_7306);
  not csa_tree_add_190_195_groupi_g41673(csa_tree_add_190_195_groupi_n_7304 ,csa_tree_add_190_195_groupi_n_7305);
  and csa_tree_add_190_195_groupi_g41674(csa_tree_add_190_195_groupi_n_7302 ,csa_tree_add_190_195_groupi_n_6139 ,csa_tree_add_190_195_groupi_n_6786);
  and csa_tree_add_190_195_groupi_g41675(csa_tree_add_190_195_groupi_n_7301 ,csa_tree_add_190_195_groupi_n_3647 ,csa_tree_add_190_195_groupi_n_7008);
  nor csa_tree_add_190_195_groupi_g41676(csa_tree_add_190_195_groupi_n_7300 ,csa_tree_add_190_195_groupi_n_6278 ,csa_tree_add_190_195_groupi_n_35);
  and csa_tree_add_190_195_groupi_g41677(csa_tree_add_190_195_groupi_n_7299 ,csa_tree_add_190_195_groupi_n_5623 ,csa_tree_add_190_195_groupi_n_6974);
  and csa_tree_add_190_195_groupi_g41678(csa_tree_add_190_195_groupi_n_7298 ,csa_tree_add_190_195_groupi_n_753 ,csa_tree_add_190_195_groupi_n_6912);
  nor csa_tree_add_190_195_groupi_g41679(csa_tree_add_190_195_groupi_n_7297 ,csa_tree_add_190_195_groupi_n_5451 ,csa_tree_add_190_195_groupi_n_6767);
  or csa_tree_add_190_195_groupi_g41680(csa_tree_add_190_195_groupi_n_7296 ,csa_tree_add_190_195_groupi_n_855 ,csa_tree_add_190_195_groupi_n_6912);
  or csa_tree_add_190_195_groupi_g41681(csa_tree_add_190_195_groupi_n_7295 ,csa_tree_add_190_195_groupi_n_5450 ,csa_tree_add_190_195_groupi_n_6766);
  nor csa_tree_add_190_195_groupi_g41682(csa_tree_add_190_195_groupi_n_7294 ,csa_tree_add_190_195_groupi_n_6914 ,csa_tree_add_190_195_groupi_n_6915);
  or csa_tree_add_190_195_groupi_g41683(csa_tree_add_190_195_groupi_n_7293 ,csa_tree_add_190_195_groupi_n_6913 ,csa_tree_add_190_195_groupi_n_6916);
  nor csa_tree_add_190_195_groupi_g41684(csa_tree_add_190_195_groupi_n_7292 ,csa_tree_add_190_195_groupi_n_5812 ,csa_tree_add_190_195_groupi_n_6777);
  or csa_tree_add_190_195_groupi_g41685(csa_tree_add_190_195_groupi_n_7291 ,csa_tree_add_190_195_groupi_n_6502 ,csa_tree_add_190_195_groupi_n_6986);
  or csa_tree_add_190_195_groupi_g41686(csa_tree_add_190_195_groupi_n_7290 ,csa_tree_add_190_195_groupi_n_5803 ,csa_tree_add_190_195_groupi_n_6981);
  and csa_tree_add_190_195_groupi_g41687(csa_tree_add_190_195_groupi_n_7289 ,csa_tree_add_190_195_groupi_n_5729 ,csa_tree_add_190_195_groupi_n_7004);
  and csa_tree_add_190_195_groupi_g41688(csa_tree_add_190_195_groupi_n_7288 ,csa_tree_add_190_195_groupi_n_5793 ,csa_tree_add_190_195_groupi_n_7001);
  nor csa_tree_add_190_195_groupi_g41689(csa_tree_add_190_195_groupi_n_7287 ,csa_tree_add_190_195_groupi_n_6997 ,csa_tree_add_190_195_groupi_n_6466);
  or csa_tree_add_190_195_groupi_g41690(csa_tree_add_190_195_groupi_n_7286 ,csa_tree_add_190_195_groupi_n_5058 ,csa_tree_add_190_195_groupi_n_6924);
  nor csa_tree_add_190_195_groupi_g41691(csa_tree_add_190_195_groupi_n_7285 ,csa_tree_add_190_195_groupi_n_5057 ,csa_tree_add_190_195_groupi_n_6925);
  or csa_tree_add_190_195_groupi_g41692(csa_tree_add_190_195_groupi_n_7284 ,csa_tree_add_190_195_groupi_n_5890 ,csa_tree_add_190_195_groupi_n_6764);
  nor csa_tree_add_190_195_groupi_g41693(csa_tree_add_190_195_groupi_n_7283 ,csa_tree_add_190_195_groupi_n_5891 ,csa_tree_add_190_195_groupi_n_6765);
  nor csa_tree_add_190_195_groupi_g41694(csa_tree_add_190_195_groupi_n_7282 ,csa_tree_add_190_195_groupi_n_5355 ,csa_tree_add_190_195_groupi_n_6928);
  or csa_tree_add_190_195_groupi_g41695(csa_tree_add_190_195_groupi_n_7281 ,csa_tree_add_190_195_groupi_n_5354 ,csa_tree_add_190_195_groupi_n_6929);
  and csa_tree_add_190_195_groupi_g41696(csa_tree_add_190_195_groupi_n_7280 ,csa_tree_add_190_195_groupi_n_6276 ,csa_tree_add_190_195_groupi_n_6932);
  nor csa_tree_add_190_195_groupi_g41697(csa_tree_add_190_195_groupi_n_7279 ,csa_tree_add_190_195_groupi_n_6944 ,csa_tree_add_190_195_groupi_n_6947);
  or csa_tree_add_190_195_groupi_g41698(csa_tree_add_190_195_groupi_n_7278 ,csa_tree_add_190_195_groupi_n_6439 ,csa_tree_add_190_195_groupi_n_6789);
  or csa_tree_add_190_195_groupi_g41699(csa_tree_add_190_195_groupi_n_7277 ,csa_tree_add_190_195_groupi_n_4914 ,csa_tree_add_190_195_groupi_n_6938);
  nor csa_tree_add_190_195_groupi_g41700(csa_tree_add_190_195_groupi_n_7276 ,csa_tree_add_190_195_groupi_n_4915 ,csa_tree_add_190_195_groupi_n_6937);
  nor csa_tree_add_190_195_groupi_g41701(csa_tree_add_190_195_groupi_n_7275 ,csa_tree_add_190_195_groupi_n_5193 ,csa_tree_add_190_195_groupi_n_6759);
  or csa_tree_add_190_195_groupi_g41702(csa_tree_add_190_195_groupi_n_7274 ,csa_tree_add_190_195_groupi_n_5192 ,csa_tree_add_190_195_groupi_n_6760);
  and csa_tree_add_190_195_groupi_g41703(csa_tree_add_190_195_groupi_n_7273 ,csa_tree_add_190_195_groupi_n_6994 ,csa_tree_add_190_195_groupi_n_6732);
  nor csa_tree_add_190_195_groupi_g41704(csa_tree_add_190_195_groupi_n_7272 ,csa_tree_add_190_195_groupi_n_6276 ,csa_tree_add_190_195_groupi_n_6932);
  and csa_tree_add_190_195_groupi_g41705(csa_tree_add_190_195_groupi_n_7271 ,csa_tree_add_190_195_groupi_n_6369 ,csa_tree_add_190_195_groupi_n_6780);
  or csa_tree_add_190_195_groupi_g41706(csa_tree_add_190_195_groupi_n_7270 ,csa_tree_add_190_195_groupi_n_6368 ,csa_tree_add_190_195_groupi_n_7015);
  nor csa_tree_add_190_195_groupi_g41707(csa_tree_add_190_195_groupi_n_7269 ,csa_tree_add_190_195_groupi_n_5227 ,csa_tree_add_190_195_groupi_n_6770);
  and csa_tree_add_190_195_groupi_g41708(csa_tree_add_190_195_groupi_n_7268 ,csa_tree_add_190_195_groupi_n_6364 ,csa_tree_add_190_195_groupi_n_7013);
  and csa_tree_add_190_195_groupi_g41709(csa_tree_add_190_195_groupi_n_7267 ,csa_tree_add_190_195_groupi_n_6122 ,csa_tree_add_190_195_groupi_n_6781);
  nor csa_tree_add_190_195_groupi_g41710(csa_tree_add_190_195_groupi_n_7266 ,csa_tree_add_190_195_groupi_n_5845 ,csa_tree_add_190_195_groupi_n_6970);
  and csa_tree_add_190_195_groupi_g41711(csa_tree_add_190_195_groupi_n_7265 ,csa_tree_add_190_195_groupi_n_6348 ,csa_tree_add_190_195_groupi_n_6782);
  nor csa_tree_add_190_195_groupi_g41712(csa_tree_add_190_195_groupi_n_7264 ,csa_tree_add_190_195_groupi_n_5251 ,csa_tree_add_190_195_groupi_n_6949);
  or csa_tree_add_190_195_groupi_g41713(csa_tree_add_190_195_groupi_n_7263 ,csa_tree_add_190_195_groupi_n_6945 ,csa_tree_add_190_195_groupi_n_6946);
  or csa_tree_add_190_195_groupi_g41714(csa_tree_add_190_195_groupi_n_7262 ,csa_tree_add_190_195_groupi_n_56 ,csa_tree_add_190_195_groupi_n_6948);
  or csa_tree_add_190_195_groupi_g41715(csa_tree_add_190_195_groupi_n_7261 ,csa_tree_add_190_195_groupi_n_5787 ,csa_tree_add_190_195_groupi_n_7000);
  and csa_tree_add_190_195_groupi_g41716(csa_tree_add_190_195_groupi_n_7260 ,csa_tree_add_190_195_groupi_n_2753 ,csa_tree_add_190_195_groupi_n_6973);
  and csa_tree_add_190_195_groupi_g41717(csa_tree_add_190_195_groupi_n_7259 ,csa_tree_add_190_195_groupi_n_6116 ,csa_tree_add_190_195_groupi_n_7012);
  or csa_tree_add_190_195_groupi_g41718(csa_tree_add_190_195_groupi_n_7258 ,csa_tree_add_190_195_groupi_n_5531 ,csa_tree_add_190_195_groupi_n_6951);
  and csa_tree_add_190_195_groupi_g41719(csa_tree_add_190_195_groupi_n_7257 ,csa_tree_add_190_195_groupi_n_5704 ,csa_tree_add_190_195_groupi_n_7007);
  nor csa_tree_add_190_195_groupi_g41720(csa_tree_add_190_195_groupi_n_7256 ,csa_tree_add_190_195_groupi_n_5249 ,csa_tree_add_190_195_groupi_n_6958);
  or csa_tree_add_190_195_groupi_g41721(csa_tree_add_190_195_groupi_n_7255 ,csa_tree_add_190_195_groupi_n_5250 ,csa_tree_add_190_195_groupi_n_6957);
  or csa_tree_add_190_195_groupi_g41722(csa_tree_add_190_195_groupi_n_7254 ,csa_tree_add_190_195_groupi_n_5303 ,csa_tree_add_190_195_groupi_n_6927);
  nor csa_tree_add_190_195_groupi_g41723(csa_tree_add_190_195_groupi_n_7253 ,csa_tree_add_190_195_groupi_n_5304 ,csa_tree_add_190_195_groupi_n_6926);
  and csa_tree_add_190_195_groupi_g41724(csa_tree_add_190_195_groupi_n_7252 ,csa_tree_add_190_195_groupi_n_5647 ,csa_tree_add_190_195_groupi_n_6783);
  and csa_tree_add_190_195_groupi_g41725(csa_tree_add_190_195_groupi_n_7251 ,csa_tree_add_190_195_groupi_n_6535 ,csa_tree_add_190_195_groupi_n_6788);
  and csa_tree_add_190_195_groupi_g41726(csa_tree_add_190_195_groupi_n_7250 ,csa_tree_add_190_195_groupi_n_5531 ,csa_tree_add_190_195_groupi_n_6951);
  nor csa_tree_add_190_195_groupi_g41727(csa_tree_add_190_195_groupi_n_7249 ,csa_tree_add_190_195_groupi_n_6936 ,csa_tree_add_190_195_groupi_n_6961);
  or csa_tree_add_190_195_groupi_g41728(csa_tree_add_190_195_groupi_n_7248 ,csa_tree_add_190_195_groupi_n_6236 ,csa_tree_add_190_195_groupi_n_6778);
  or csa_tree_add_190_195_groupi_g41729(csa_tree_add_190_195_groupi_n_7247 ,csa_tree_add_190_195_groupi_n_4782 ,csa_tree_add_190_195_groupi_n_6963);
  or csa_tree_add_190_195_groupi_g41730(csa_tree_add_190_195_groupi_n_7246 ,csa_tree_add_190_195_groupi_n_5226 ,csa_tree_add_190_195_groupi_n_6769);
  or csa_tree_add_190_195_groupi_g41731(csa_tree_add_190_195_groupi_n_7245 ,csa_tree_add_190_195_groupi_n_6935 ,csa_tree_add_190_195_groupi_n_6962);
  and csa_tree_add_190_195_groupi_g41732(csa_tree_add_190_195_groupi_n_7244 ,csa_tree_add_190_195_groupi_n_4782 ,csa_tree_add_190_195_groupi_n_6963);
  or csa_tree_add_190_195_groupi_g41733(csa_tree_add_190_195_groupi_n_7243 ,csa_tree_add_190_195_groupi_n_6980 ,csa_tree_add_190_195_groupi_n_6218);
  or csa_tree_add_190_195_groupi_g41734(csa_tree_add_190_195_groupi_n_7242 ,csa_tree_add_190_195_groupi_n_6111 ,csa_tree_add_190_195_groupi_n_6971);
  nor csa_tree_add_190_195_groupi_g41735(csa_tree_add_190_195_groupi_n_7241 ,csa_tree_add_190_195_groupi_n_6966 ,csa_tree_add_190_195_groupi_n_6921);
  or csa_tree_add_190_195_groupi_g41736(csa_tree_add_190_195_groupi_n_7240 ,csa_tree_add_190_195_groupi_n_5759 ,csa_tree_add_190_195_groupi_n_6982);
  or csa_tree_add_190_195_groupi_g41737(csa_tree_add_190_195_groupi_n_7239 ,csa_tree_add_190_195_groupi_n_6965 ,csa_tree_add_190_195_groupi_n_6920);
  or csa_tree_add_190_195_groupi_g41738(csa_tree_add_190_195_groupi_n_7238 ,csa_tree_add_190_195_groupi_n_5330 ,csa_tree_add_190_195_groupi_n_6952);
  and csa_tree_add_190_195_groupi_g41739(csa_tree_add_190_195_groupi_n_7237 ,csa_tree_add_190_195_groupi_n_6852 ,csa_tree_add_190_195_groupi_n_6775);
  and csa_tree_add_190_195_groupi_g41740(csa_tree_add_190_195_groupi_n_7236 ,csa_tree_add_190_195_groupi_n_27 ,csa_tree_add_190_195_groupi_n_6862);
  or csa_tree_add_190_195_groupi_g41741(csa_tree_add_190_195_groupi_n_7235 ,csa_tree_add_190_195_groupi_n_6868 ,csa_tree_add_190_195_groupi_n_7010);
  and csa_tree_add_190_195_groupi_g41742(csa_tree_add_190_195_groupi_n_7234 ,csa_tree_add_190_195_groupi_n_5658 ,csa_tree_add_190_195_groupi_n_6978);
  or csa_tree_add_190_195_groupi_g41743(csa_tree_add_190_195_groupi_n_7233 ,csa_tree_add_190_195_groupi_n_6277 ,csa_tree_add_190_195_groupi_n_6758);
  and csa_tree_add_190_195_groupi_g41744(csa_tree_add_190_195_groupi_n_7431 ,csa_tree_add_190_195_groupi_n_6512 ,csa_tree_add_190_195_groupi_n_6889);
  and csa_tree_add_190_195_groupi_g41745(csa_tree_add_190_195_groupi_n_7430 ,csa_tree_add_190_195_groupi_n_5865 ,csa_tree_add_190_195_groupi_n_6851);
  and csa_tree_add_190_195_groupi_g41746(csa_tree_add_190_195_groupi_n_7429 ,csa_tree_add_190_195_groupi_n_6458 ,csa_tree_add_190_195_groupi_n_6875);
  and csa_tree_add_190_195_groupi_g41747(csa_tree_add_190_195_groupi_n_7428 ,csa_tree_add_190_195_groupi_n_6462 ,csa_tree_add_190_195_groupi_n_6745);
  or csa_tree_add_190_195_groupi_g41748(csa_tree_add_190_195_groupi_n_7426 ,csa_tree_add_190_195_groupi_n_6303 ,csa_tree_add_190_195_groupi_n_6867);
  or csa_tree_add_190_195_groupi_g41749(csa_tree_add_190_195_groupi_n_7425 ,csa_tree_add_190_195_groupi_n_96 ,csa_tree_add_190_195_groupi_n_6792);
  and csa_tree_add_190_195_groupi_g41750(csa_tree_add_190_195_groupi_n_7424 ,csa_tree_add_190_195_groupi_n_6407 ,csa_tree_add_190_195_groupi_n_6814);
  or csa_tree_add_190_195_groupi_g41751(csa_tree_add_190_195_groupi_n_7423 ,csa_tree_add_190_195_groupi_n_6373 ,csa_tree_add_190_195_groupi_n_6907);
  and csa_tree_add_190_195_groupi_g41752(csa_tree_add_190_195_groupi_n_7422 ,csa_tree_add_190_195_groupi_n_6471 ,csa_tree_add_190_195_groupi_n_6813);
  or csa_tree_add_190_195_groupi_g41753(csa_tree_add_190_195_groupi_n_7420 ,csa_tree_add_190_195_groupi_n_6356 ,csa_tree_add_190_195_groupi_n_6749);
  and csa_tree_add_190_195_groupi_g41754(csa_tree_add_190_195_groupi_n_7419 ,csa_tree_add_190_195_groupi_n_6504 ,csa_tree_add_190_195_groupi_n_6884);
  and csa_tree_add_190_195_groupi_g41755(csa_tree_add_190_195_groupi_n_7418 ,csa_tree_add_190_195_groupi_n_6564 ,csa_tree_add_190_195_groupi_n_6810);
  and csa_tree_add_190_195_groupi_g41756(csa_tree_add_190_195_groupi_n_7417 ,csa_tree_add_190_195_groupi_n_6211 ,csa_tree_add_190_195_groupi_n_6821);
  and csa_tree_add_190_195_groupi_g41757(csa_tree_add_190_195_groupi_n_7416 ,csa_tree_add_190_195_groupi_n_6317 ,csa_tree_add_190_195_groupi_n_6900);
  and csa_tree_add_190_195_groupi_g41758(csa_tree_add_190_195_groupi_n_7415 ,csa_tree_add_190_195_groupi_n_6380 ,csa_tree_add_190_195_groupi_n_6799);
  and csa_tree_add_190_195_groupi_g41759(csa_tree_add_190_195_groupi_n_7414 ,csa_tree_add_190_195_groupi_n_6360 ,csa_tree_add_190_195_groupi_n_6846);
  and csa_tree_add_190_195_groupi_g41760(csa_tree_add_190_195_groupi_n_7413 ,csa_tree_add_190_195_groupi_n_6557 ,csa_tree_add_190_195_groupi_n_6904);
  and csa_tree_add_190_195_groupi_g41761(csa_tree_add_190_195_groupi_n_7412 ,csa_tree_add_190_195_groupi_n_2936 ,csa_tree_add_190_195_groupi_n_6820);
  or csa_tree_add_190_195_groupi_g41762(csa_tree_add_190_195_groupi_n_7411 ,csa_tree_add_190_195_groupi_n_6548 ,csa_tree_add_190_195_groupi_n_6893);
  or csa_tree_add_190_195_groupi_g41763(csa_tree_add_190_195_groupi_n_7410 ,csa_tree_add_190_195_groupi_n_6494 ,csa_tree_add_190_195_groupi_n_6885);
  or csa_tree_add_190_195_groupi_g41764(csa_tree_add_190_195_groupi_n_7409 ,csa_tree_add_190_195_groupi_n_3153 ,csa_tree_add_190_195_groupi_n_6902);
  or csa_tree_add_190_195_groupi_g41765(csa_tree_add_190_195_groupi_n_7408 ,csa_tree_add_190_195_groupi_n_6305 ,csa_tree_add_190_195_groupi_n_6841);
  and csa_tree_add_190_195_groupi_g41766(csa_tree_add_190_195_groupi_n_7407 ,csa_tree_add_190_195_groupi_n_6167 ,csa_tree_add_190_195_groupi_n_6823);
  or csa_tree_add_190_195_groupi_g41767(csa_tree_add_190_195_groupi_n_7406 ,csa_tree_add_190_195_groupi_n_6322 ,csa_tree_add_190_195_groupi_n_6890);
  and csa_tree_add_190_195_groupi_g41768(csa_tree_add_190_195_groupi_n_7405 ,csa_tree_add_190_195_groupi_n_6217 ,csa_tree_add_190_195_groupi_n_6798);
  and csa_tree_add_190_195_groupi_g41769(csa_tree_add_190_195_groupi_n_7404 ,csa_tree_add_190_195_groupi_n_6207 ,csa_tree_add_190_195_groupi_n_6824);
  and csa_tree_add_190_195_groupi_g41770(csa_tree_add_190_195_groupi_n_7403 ,csa_tree_add_190_195_groupi_n_6386 ,csa_tree_add_190_195_groupi_n_6793);
  or csa_tree_add_190_195_groupi_g41771(csa_tree_add_190_195_groupi_n_7402 ,csa_tree_add_190_195_groupi_n_6345 ,csa_tree_add_190_195_groupi_n_6838);
  or csa_tree_add_190_195_groupi_g41772(csa_tree_add_190_195_groupi_n_7401 ,csa_tree_add_190_195_groupi_n_6235 ,csa_tree_add_190_195_groupi_n_6805);
  and csa_tree_add_190_195_groupi_g41773(csa_tree_add_190_195_groupi_n_7400 ,csa_tree_add_190_195_groupi_n_6384 ,csa_tree_add_190_195_groupi_n_6903);
  or csa_tree_add_190_195_groupi_g41774(csa_tree_add_190_195_groupi_n_7399 ,csa_tree_add_190_195_groupi_n_6339 ,csa_tree_add_190_195_groupi_n_6837);
  and csa_tree_add_190_195_groupi_g41775(csa_tree_add_190_195_groupi_n_7398 ,csa_tree_add_190_195_groupi_n_6387 ,csa_tree_add_190_195_groupi_n_6804);
  and csa_tree_add_190_195_groupi_g41776(csa_tree_add_190_195_groupi_n_7397 ,csa_tree_add_190_195_groupi_n_6180 ,csa_tree_add_190_195_groupi_n_6817);
  and csa_tree_add_190_195_groupi_g41777(csa_tree_add_190_195_groupi_n_7396 ,csa_tree_add_190_195_groupi_n_6417 ,csa_tree_add_190_195_groupi_n_6863);
  and csa_tree_add_190_195_groupi_g41778(csa_tree_add_190_195_groupi_n_7395 ,csa_tree_add_190_195_groupi_n_6365 ,csa_tree_add_190_195_groupi_n_6797);
  and csa_tree_add_190_195_groupi_g41779(csa_tree_add_190_195_groupi_n_7394 ,csa_tree_add_190_195_groupi_n_6106 ,csa_tree_add_190_195_groupi_n_6831);
  or csa_tree_add_190_195_groupi_g41780(csa_tree_add_190_195_groupi_n_7392 ,csa_tree_add_190_195_groupi_n_6551 ,csa_tree_add_190_195_groupi_n_6833);
  and csa_tree_add_190_195_groupi_g41781(csa_tree_add_190_195_groupi_n_7391 ,csa_tree_add_190_195_groupi_n_6202 ,csa_tree_add_190_195_groupi_n_6861);
  and csa_tree_add_190_195_groupi_g41782(csa_tree_add_190_195_groupi_n_7390 ,csa_tree_add_190_195_groupi_n_6199 ,csa_tree_add_190_195_groupi_n_6878);
  and csa_tree_add_190_195_groupi_g41783(csa_tree_add_190_195_groupi_n_7389 ,csa_tree_add_190_195_groupi_n_6561 ,csa_tree_add_190_195_groupi_n_6857);
  and csa_tree_add_190_195_groupi_g41784(csa_tree_add_190_195_groupi_n_7388 ,csa_tree_add_190_195_groupi_n_6238 ,csa_tree_add_190_195_groupi_n_6882);
  and csa_tree_add_190_195_groupi_g41785(csa_tree_add_190_195_groupi_n_7387 ,csa_tree_add_190_195_groupi_n_6549 ,csa_tree_add_190_195_groupi_n_6806);
  or csa_tree_add_190_195_groupi_g41786(csa_tree_add_190_195_groupi_n_7386 ,csa_tree_add_190_195_groupi_n_6298 ,csa_tree_add_190_195_groupi_n_6819);
  and csa_tree_add_190_195_groupi_g41787(csa_tree_add_190_195_groupi_n_7385 ,csa_tree_add_190_195_groupi_n_6143 ,csa_tree_add_190_195_groupi_n_6891);
  or csa_tree_add_190_195_groupi_g41788(csa_tree_add_190_195_groupi_n_7383 ,csa_tree_add_190_195_groupi_n_3517 ,csa_tree_add_190_195_groupi_n_6850);
  or csa_tree_add_190_195_groupi_g41789(csa_tree_add_190_195_groupi_n_7382 ,csa_tree_add_190_195_groupi_n_6137 ,csa_tree_add_190_195_groupi_n_6881);
  and csa_tree_add_190_195_groupi_g41790(csa_tree_add_190_195_groupi_n_7381 ,csa_tree_add_190_195_groupi_n_6130 ,csa_tree_add_190_195_groupi_n_6896);
  or csa_tree_add_190_195_groupi_g41791(csa_tree_add_190_195_groupi_n_7380 ,csa_tree_add_190_195_groupi_n_3259 ,csa_tree_add_190_195_groupi_n_6811);
  or csa_tree_add_190_195_groupi_g41792(csa_tree_add_190_195_groupi_n_7378 ,csa_tree_add_190_195_groupi_n_6499 ,csa_tree_add_190_195_groupi_n_6886);
  or csa_tree_add_190_195_groupi_g41793(csa_tree_add_190_195_groupi_n_7376 ,csa_tree_add_190_195_groupi_n_6443 ,csa_tree_add_190_195_groupi_n_6866);
  or csa_tree_add_190_195_groupi_g41794(csa_tree_add_190_195_groupi_n_7375 ,csa_tree_add_190_195_groupi_n_6425 ,csa_tree_add_190_195_groupi_n_6854);
  and csa_tree_add_190_195_groupi_g41795(csa_tree_add_190_195_groupi_n_7373 ,csa_tree_add_190_195_groupi_n_6432 ,csa_tree_add_190_195_groupi_n_6844);
  or csa_tree_add_190_195_groupi_g41796(csa_tree_add_190_195_groupi_n_7372 ,csa_tree_add_190_195_groupi_n_6347 ,csa_tree_add_190_195_groupi_n_6803);
  or csa_tree_add_190_195_groupi_g41797(csa_tree_add_190_195_groupi_n_7370 ,csa_tree_add_190_195_groupi_n_6245 ,csa_tree_add_190_195_groupi_n_6883);
  and csa_tree_add_190_195_groupi_g41798(csa_tree_add_190_195_groupi_n_7368 ,csa_tree_add_190_195_groupi_n_6528 ,csa_tree_add_190_195_groupi_n_6894);
  and csa_tree_add_190_195_groupi_g41799(csa_tree_add_190_195_groupi_n_7366 ,csa_tree_add_190_195_groupi_n_6234 ,csa_tree_add_190_195_groupi_n_6800);
  and csa_tree_add_190_195_groupi_g41800(csa_tree_add_190_195_groupi_n_7364 ,csa_tree_add_190_195_groupi_n_6482 ,csa_tree_add_190_195_groupi_n_6801);
  or csa_tree_add_190_195_groupi_g41801(csa_tree_add_190_195_groupi_n_7363 ,csa_tree_add_190_195_groupi_n_5738 ,csa_tree_add_190_195_groupi_n_6842);
  and csa_tree_add_190_195_groupi_g41802(csa_tree_add_190_195_groupi_n_7362 ,csa_tree_add_190_195_groupi_n_6540 ,csa_tree_add_190_195_groupi_n_6898);
  and csa_tree_add_190_195_groupi_g41803(csa_tree_add_190_195_groupi_n_7359 ,csa_tree_add_190_195_groupi_n_6423 ,csa_tree_add_190_195_groupi_n_6864);
  and csa_tree_add_190_195_groupi_g41804(csa_tree_add_190_195_groupi_n_7358 ,csa_tree_add_190_195_groupi_n_6529 ,csa_tree_add_190_195_groupi_n_6827);
  or csa_tree_add_190_195_groupi_g41805(csa_tree_add_190_195_groupi_n_7356 ,csa_tree_add_190_195_groupi_n_6484 ,csa_tree_add_190_195_groupi_n_6870);
  and csa_tree_add_190_195_groupi_g41806(csa_tree_add_190_195_groupi_n_7354 ,csa_tree_add_190_195_groupi_n_6338 ,csa_tree_add_190_195_groupi_n_6835);
  and csa_tree_add_190_195_groupi_g41807(csa_tree_add_190_195_groupi_n_7353 ,csa_tree_add_190_195_groupi_n_6538 ,csa_tree_add_190_195_groupi_n_6897);
  or csa_tree_add_190_195_groupi_g41808(csa_tree_add_190_195_groupi_n_7352 ,csa_tree_add_190_195_groupi_n_6411 ,csa_tree_add_190_195_groupi_n_6859);
  or csa_tree_add_190_195_groupi_g41809(csa_tree_add_190_195_groupi_n_7351 ,csa_tree_add_190_195_groupi_n_5679 ,csa_tree_add_190_195_groupi_n_6796);
  or csa_tree_add_190_195_groupi_g41810(csa_tree_add_190_195_groupi_n_7350 ,csa_tree_add_190_195_groupi_n_6409 ,csa_tree_add_190_195_groupi_n_6855);
  or csa_tree_add_190_195_groupi_g41811(csa_tree_add_190_195_groupi_n_7347 ,csa_tree_add_190_195_groupi_n_6206 ,csa_tree_add_190_195_groupi_n_6795);
  and csa_tree_add_190_195_groupi_g41812(csa_tree_add_190_195_groupi_n_7346 ,csa_tree_add_190_195_groupi_n_6205 ,csa_tree_add_190_195_groupi_n_6794);
  or csa_tree_add_190_195_groupi_g41813(csa_tree_add_190_195_groupi_n_7343 ,csa_tree_add_190_195_groupi_n_5766 ,csa_tree_add_190_195_groupi_n_6860);
  and csa_tree_add_190_195_groupi_g41814(csa_tree_add_190_195_groupi_n_7342 ,csa_tree_add_190_195_groupi_n_6427 ,csa_tree_add_190_195_groupi_n_6825);
  and csa_tree_add_190_195_groupi_g41815(csa_tree_add_190_195_groupi_n_7341 ,csa_tree_add_190_195_groupi_n_6158 ,csa_tree_add_190_195_groupi_n_6856);
  or csa_tree_add_190_195_groupi_g41816(csa_tree_add_190_195_groupi_n_7339 ,csa_tree_add_190_195_groupi_n_5697 ,csa_tree_add_190_195_groupi_n_6822);
  and csa_tree_add_190_195_groupi_g41817(csa_tree_add_190_195_groupi_n_7338 ,csa_tree_add_190_195_groupi_n_6553 ,csa_tree_add_190_195_groupi_n_6826);
  and csa_tree_add_190_195_groupi_g41818(csa_tree_add_190_195_groupi_n_7336 ,csa_tree_add_190_195_groupi_n_6554 ,csa_tree_add_190_195_groupi_n_6828);
  or csa_tree_add_190_195_groupi_g41819(csa_tree_add_190_195_groupi_n_7334 ,csa_tree_add_190_195_groupi_n_6112 ,csa_tree_add_190_195_groupi_n_6808);
  or csa_tree_add_190_195_groupi_g41820(csa_tree_add_190_195_groupi_n_7332 ,csa_tree_add_190_195_groupi_n_95 ,csa_tree_add_190_195_groupi_n_6818);
  and csa_tree_add_190_195_groupi_g41821(csa_tree_add_190_195_groupi_n_7330 ,csa_tree_add_190_195_groupi_n_6544 ,csa_tree_add_190_195_groupi_n_6853);
  and csa_tree_add_190_195_groupi_g41822(csa_tree_add_190_195_groupi_n_7328 ,csa_tree_add_190_195_groupi_n_6473 ,csa_tree_add_190_195_groupi_n_6876);
  or csa_tree_add_190_195_groupi_g41823(csa_tree_add_190_195_groupi_n_7327 ,csa_tree_add_190_195_groupi_n_6346 ,csa_tree_add_190_195_groupi_n_6802);
  and csa_tree_add_190_195_groupi_g41824(csa_tree_add_190_195_groupi_n_7325 ,csa_tree_add_190_195_groupi_n_6568 ,csa_tree_add_190_195_groupi_n_6832);
  or csa_tree_add_190_195_groupi_g41825(csa_tree_add_190_195_groupi_n_7323 ,csa_tree_add_190_195_groupi_n_6534 ,csa_tree_add_190_195_groupi_n_6895);
  and csa_tree_add_190_195_groupi_g41826(csa_tree_add_190_195_groupi_n_7320 ,csa_tree_add_190_195_groupi_n_6156 ,csa_tree_add_190_195_groupi_n_6834);
  and csa_tree_add_190_195_groupi_g41827(csa_tree_add_190_195_groupi_n_7318 ,csa_tree_add_190_195_groupi_n_6460 ,csa_tree_add_190_195_groupi_n_6816);
  and csa_tree_add_190_195_groupi_g41828(csa_tree_add_190_195_groupi_n_7317 ,csa_tree_add_190_195_groupi_n_5832 ,csa_tree_add_190_195_groupi_n_6899);
  and csa_tree_add_190_195_groupi_g41829(csa_tree_add_190_195_groupi_n_7316 ,csa_tree_add_190_195_groupi_n_6157 ,csa_tree_add_190_195_groupi_n_6836);
  or csa_tree_add_190_195_groupi_g41830(csa_tree_add_190_195_groupi_n_7315 ,csa_tree_add_190_195_groupi_n_6383 ,csa_tree_add_190_195_groupi_n_6815);
  and csa_tree_add_190_195_groupi_g41831(csa_tree_add_190_195_groupi_n_7314 ,csa_tree_add_190_195_groupi_n_6514 ,csa_tree_add_190_195_groupi_n_6888);
  or csa_tree_add_190_195_groupi_g41832(csa_tree_add_190_195_groupi_n_7313 ,csa_tree_add_190_195_groupi_n_6097 ,csa_tree_add_190_195_groupi_n_6872);
  or csa_tree_add_190_195_groupi_g41833(csa_tree_add_190_195_groupi_n_7312 ,csa_tree_add_190_195_groupi_n_6481 ,csa_tree_add_190_195_groupi_n_6879);
  or csa_tree_add_190_195_groupi_g41834(csa_tree_add_190_195_groupi_n_7309 ,csa_tree_add_190_195_groupi_n_6233 ,csa_tree_add_190_195_groupi_n_6723);
  and csa_tree_add_190_195_groupi_g41835(csa_tree_add_190_195_groupi_n_7308 ,csa_tree_add_190_195_groupi_n_6519 ,csa_tree_add_190_195_groupi_n_6812);
  and csa_tree_add_190_195_groupi_g41836(csa_tree_add_190_195_groupi_n_7306 ,csa_tree_add_190_195_groupi_n_6559 ,csa_tree_add_190_195_groupi_n_6901);
  and csa_tree_add_190_195_groupi_g41837(csa_tree_add_190_195_groupi_n_7305 ,csa_tree_add_190_195_groupi_n_6133 ,csa_tree_add_190_195_groupi_n_6892);
  or csa_tree_add_190_195_groupi_g41838(csa_tree_add_190_195_groupi_n_7303 ,csa_tree_add_190_195_groupi_n_6450 ,csa_tree_add_190_195_groupi_n_6869);
  not csa_tree_add_190_195_groupi_g41839(csa_tree_add_190_195_groupi_n_7230 ,csa_tree_add_190_195_groupi_n_7229);
  not csa_tree_add_190_195_groupi_g41841(csa_tree_add_190_195_groupi_n_7220 ,csa_tree_add_190_195_groupi_n_73);
  not csa_tree_add_190_195_groupi_g41842(csa_tree_add_190_195_groupi_n_7219 ,csa_tree_add_190_195_groupi_n_7218);
  not csa_tree_add_190_195_groupi_g41843(csa_tree_add_190_195_groupi_n_7217 ,csa_tree_add_190_195_groupi_n_7216);
  not csa_tree_add_190_195_groupi_g41844(csa_tree_add_190_195_groupi_n_7208 ,csa_tree_add_190_195_groupi_n_7207);
  not csa_tree_add_190_195_groupi_g41845(csa_tree_add_190_195_groupi_n_7206 ,csa_tree_add_190_195_groupi_n_7205);
  not csa_tree_add_190_195_groupi_g41846(csa_tree_add_190_195_groupi_n_7203 ,csa_tree_add_190_195_groupi_n_7202);
  not csa_tree_add_190_195_groupi_g41848(csa_tree_add_190_195_groupi_n_7192 ,csa_tree_add_190_195_groupi_n_7191);
  not csa_tree_add_190_195_groupi_g41849(csa_tree_add_190_195_groupi_n_7189 ,csa_tree_add_190_195_groupi_n_7188);
  not csa_tree_add_190_195_groupi_g41850(csa_tree_add_190_195_groupi_n_7187 ,csa_tree_add_190_195_groupi_n_7186);
  not csa_tree_add_190_195_groupi_g41851(csa_tree_add_190_195_groupi_n_7185 ,csa_tree_add_190_195_groupi_n_7184);
  not csa_tree_add_190_195_groupi_g41852(csa_tree_add_190_195_groupi_n_7181 ,csa_tree_add_190_195_groupi_n_7180);
  not csa_tree_add_190_195_groupi_g41853(csa_tree_add_190_195_groupi_n_7178 ,csa_tree_add_190_195_groupi_n_7177);
  not csa_tree_add_190_195_groupi_g41854(csa_tree_add_190_195_groupi_n_7175 ,csa_tree_add_190_195_groupi_n_7176);
  not csa_tree_add_190_195_groupi_g41855(csa_tree_add_190_195_groupi_n_7174 ,csa_tree_add_190_195_groupi_n_7173);
  not csa_tree_add_190_195_groupi_g41856(csa_tree_add_190_195_groupi_n_7172 ,csa_tree_add_190_195_groupi_n_7171);
  not csa_tree_add_190_195_groupi_g41857(csa_tree_add_190_195_groupi_n_7169 ,csa_tree_add_190_195_groupi_n_7170);
  not csa_tree_add_190_195_groupi_g41858(csa_tree_add_190_195_groupi_n_7167 ,csa_tree_add_190_195_groupi_n_7168);
  not csa_tree_add_190_195_groupi_g41859(csa_tree_add_190_195_groupi_n_7166 ,csa_tree_add_190_195_groupi_n_7165);
  not csa_tree_add_190_195_groupi_g41860(csa_tree_add_190_195_groupi_n_7164 ,csa_tree_add_190_195_groupi_n_7163);
  not csa_tree_add_190_195_groupi_g41861(csa_tree_add_190_195_groupi_n_7162 ,csa_tree_add_190_195_groupi_n_7161);
  not csa_tree_add_190_195_groupi_g41862(csa_tree_add_190_195_groupi_n_7160 ,csa_tree_add_190_195_groupi_n_7159);
  not csa_tree_add_190_195_groupi_g41863(csa_tree_add_190_195_groupi_n_7157 ,csa_tree_add_190_195_groupi_n_7158);
  not csa_tree_add_190_195_groupi_g41864(csa_tree_add_190_195_groupi_n_7156 ,csa_tree_add_190_195_groupi_n_7155);
  not csa_tree_add_190_195_groupi_g41865(csa_tree_add_190_195_groupi_n_7151 ,csa_tree_add_190_195_groupi_n_21);
  not csa_tree_add_190_195_groupi_g41866(csa_tree_add_190_195_groupi_n_7148 ,csa_tree_add_190_195_groupi_n_7149);
  not csa_tree_add_190_195_groupi_g41867(csa_tree_add_190_195_groupi_n_7145 ,csa_tree_add_190_195_groupi_n_7146);
  not csa_tree_add_190_195_groupi_g41868(csa_tree_add_190_195_groupi_n_7144 ,csa_tree_add_190_195_groupi_n_7143);
  not csa_tree_add_190_195_groupi_g41869(csa_tree_add_190_195_groupi_n_7141 ,csa_tree_add_190_195_groupi_n_7142);
  not csa_tree_add_190_195_groupi_g41870(csa_tree_add_190_195_groupi_n_7139 ,csa_tree_add_190_195_groupi_n_7140);
  not csa_tree_add_190_195_groupi_g41871(csa_tree_add_190_195_groupi_n_7137 ,csa_tree_add_190_195_groupi_n_7136);
  not csa_tree_add_190_195_groupi_g41872(csa_tree_add_190_195_groupi_n_7133 ,csa_tree_add_190_195_groupi_n_7132);
  not csa_tree_add_190_195_groupi_g41873(csa_tree_add_190_195_groupi_n_7131 ,csa_tree_add_190_195_groupi_n_7130);
  not csa_tree_add_190_195_groupi_g41874(csa_tree_add_190_195_groupi_n_7128 ,csa_tree_add_190_195_groupi_n_7129);
  not csa_tree_add_190_195_groupi_g41875(csa_tree_add_190_195_groupi_n_7127 ,csa_tree_add_190_195_groupi_n_7126);
  not csa_tree_add_190_195_groupi_g41876(csa_tree_add_190_195_groupi_n_7125 ,csa_tree_add_190_195_groupi_n_7124);
  not csa_tree_add_190_195_groupi_g41877(csa_tree_add_190_195_groupi_n_7123 ,csa_tree_add_190_195_groupi_n_7122);
  not csa_tree_add_190_195_groupi_g41878(csa_tree_add_190_195_groupi_n_7120 ,csa_tree_add_190_195_groupi_n_7121);
  not csa_tree_add_190_195_groupi_g41879(csa_tree_add_190_195_groupi_n_7118 ,csa_tree_add_190_195_groupi_n_7117);
  not csa_tree_add_190_195_groupi_g41880(csa_tree_add_190_195_groupi_n_7116 ,csa_tree_add_190_195_groupi_n_7115);
  not csa_tree_add_190_195_groupi_g41881(csa_tree_add_190_195_groupi_n_7114 ,csa_tree_add_190_195_groupi_n_7113);
  not csa_tree_add_190_195_groupi_g41882(csa_tree_add_190_195_groupi_n_7112 ,csa_tree_add_190_195_groupi_n_7111);
  not csa_tree_add_190_195_groupi_g41883(csa_tree_add_190_195_groupi_n_7110 ,csa_tree_add_190_195_groupi_n_7109);
  not csa_tree_add_190_195_groupi_g41884(csa_tree_add_190_195_groupi_n_7107 ,csa_tree_add_190_195_groupi_n_7108);
  not csa_tree_add_190_195_groupi_g41885(csa_tree_add_190_195_groupi_n_7104 ,csa_tree_add_190_195_groupi_n_7105);
  not csa_tree_add_190_195_groupi_g41886(csa_tree_add_190_195_groupi_n_7102 ,csa_tree_add_190_195_groupi_n_7103);
  not csa_tree_add_190_195_groupi_g41887(csa_tree_add_190_195_groupi_n_7100 ,csa_tree_add_190_195_groupi_n_7101);
  not csa_tree_add_190_195_groupi_g41888(csa_tree_add_190_195_groupi_n_7099 ,csa_tree_add_190_195_groupi_n_7098);
  not csa_tree_add_190_195_groupi_g41889(csa_tree_add_190_195_groupi_n_7095 ,csa_tree_add_190_195_groupi_n_74);
  not csa_tree_add_190_195_groupi_g41890(csa_tree_add_190_195_groupi_n_7093 ,csa_tree_add_190_195_groupi_n_7092);
  not csa_tree_add_190_195_groupi_g41891(csa_tree_add_190_195_groupi_n_7089 ,csa_tree_add_190_195_groupi_n_7090);
  not csa_tree_add_190_195_groupi_g41892(csa_tree_add_190_195_groupi_n_7087 ,csa_tree_add_190_195_groupi_n_7086);
  not csa_tree_add_190_195_groupi_g41893(csa_tree_add_190_195_groupi_n_7084 ,csa_tree_add_190_195_groupi_n_7085);
  not csa_tree_add_190_195_groupi_g41894(csa_tree_add_190_195_groupi_n_7081 ,csa_tree_add_190_195_groupi_n_7082);
  not csa_tree_add_190_195_groupi_g41895(csa_tree_add_190_195_groupi_n_7079 ,csa_tree_add_190_195_groupi_n_7080);
  not csa_tree_add_190_195_groupi_g41896(csa_tree_add_190_195_groupi_n_7074 ,csa_tree_add_190_195_groupi_n_7075);
  not csa_tree_add_190_195_groupi_g41897(csa_tree_add_190_195_groupi_n_7071 ,csa_tree_add_190_195_groupi_n_7072);
  not csa_tree_add_190_195_groupi_g41898(csa_tree_add_190_195_groupi_n_7069 ,csa_tree_add_190_195_groupi_n_7070);
  not csa_tree_add_190_195_groupi_g41899(csa_tree_add_190_195_groupi_n_7067 ,csa_tree_add_190_195_groupi_n_7066);
  not csa_tree_add_190_195_groupi_g41900(csa_tree_add_190_195_groupi_n_7064 ,csa_tree_add_190_195_groupi_n_7065);
  not csa_tree_add_190_195_groupi_g41901(csa_tree_add_190_195_groupi_n_7062 ,csa_tree_add_190_195_groupi_n_7063);
  and csa_tree_add_190_195_groupi_g41902(csa_tree_add_190_195_groupi_n_7060 ,csa_tree_add_190_195_groupi_n_6351 ,csa_tree_add_190_195_groupi_n_6787);
  or csa_tree_add_190_195_groupi_g41903(csa_tree_add_190_195_groupi_n_7059 ,csa_tree_add_190_195_groupi_n_6906 ,csa_tree_add_190_195_groupi_n_6785);
  and csa_tree_add_190_195_groupi_g41904(csa_tree_add_190_195_groupi_n_7058 ,csa_tree_add_190_195_groupi_n_5687 ,csa_tree_add_190_195_groupi_n_6790);
  or csa_tree_add_190_195_groupi_g41905(csa_tree_add_190_195_groupi_n_7057 ,csa_tree_add_190_195_groupi_n_5199 ,csa_tree_add_190_195_groupi_n_6763);
  nor csa_tree_add_190_195_groupi_g41906(csa_tree_add_190_195_groupi_n_7056 ,csa_tree_add_190_195_groupi_n_5331 ,csa_tree_add_190_195_groupi_n_6953);
  or csa_tree_add_190_195_groupi_g41907(csa_tree_add_190_195_groupi_n_7055 ,csa_tree_add_190_195_groupi_n_5644 ,csa_tree_add_190_195_groupi_n_6779);
  or csa_tree_add_190_195_groupi_g41908(csa_tree_add_190_195_groupi_n_7054 ,csa_tree_add_190_195_groupi_n_4608 ,csa_tree_add_190_195_groupi_n_6772);
  nor csa_tree_add_190_195_groupi_g41909(csa_tree_add_190_195_groupi_n_7053 ,csa_tree_add_190_195_groupi_n_4609 ,csa_tree_add_190_195_groupi_n_6771);
  or csa_tree_add_190_195_groupi_g41910(csa_tree_add_190_195_groupi_n_7052 ,csa_tree_add_190_195_groupi_n_5136 ,csa_tree_add_190_195_groupi_n_6746);
  and csa_tree_add_190_195_groupi_g41911(csa_tree_add_190_195_groupi_n_7051 ,csa_tree_add_190_195_groupi_n_3152 ,csa_tree_add_190_195_groupi_n_6988);
  nor csa_tree_add_190_195_groupi_g41912(csa_tree_add_190_195_groupi_n_7050 ,csa_tree_add_190_195_groupi_n_6575 ,csa_tree_add_190_195_groupi_n_6934);
  or csa_tree_add_190_195_groupi_g41913(csa_tree_add_190_195_groupi_n_7049 ,csa_tree_add_190_195_groupi_n_6574 ,csa_tree_add_190_195_groupi_n_6933);
  and csa_tree_add_190_195_groupi_g41914(csa_tree_add_190_195_groupi_n_7048 ,csa_tree_add_190_195_groupi_n_6992 ,csa_tree_add_190_195_groupi_n_6399);
  or csa_tree_add_190_195_groupi_g41915(csa_tree_add_190_195_groupi_n_7047 ,csa_tree_add_190_195_groupi_n_5818 ,csa_tree_add_190_195_groupi_n_6995);
  and csa_tree_add_190_195_groupi_g41916(csa_tree_add_190_195_groupi_n_7046 ,csa_tree_add_190_195_groupi_n_4877 ,csa_tree_add_190_195_groupi_n_6975);
  nor csa_tree_add_190_195_groupi_g41917(csa_tree_add_190_195_groupi_n_7045 ,csa_tree_add_190_195_groupi_n_6566 ,csa_tree_add_190_195_groupi_n_7016);
  or csa_tree_add_190_195_groupi_g41918(csa_tree_add_190_195_groupi_n_7044 ,csa_tree_add_190_195_groupi_n_6445 ,csa_tree_add_190_195_groupi_n_6990);
  or csa_tree_add_190_195_groupi_g41919(csa_tree_add_190_195_groupi_n_7043 ,csa_tree_add_190_195_groupi_n_3375 ,csa_tree_add_190_195_groupi_n_6984);
  or csa_tree_add_190_195_groupi_g41920(csa_tree_add_190_195_groupi_n_7042 ,csa_tree_add_190_195_groupi_n_7006 ,csa_tree_add_190_195_groupi_n_6173);
  nor csa_tree_add_190_195_groupi_g41921(csa_tree_add_190_195_groupi_n_7041 ,csa_tree_add_190_195_groupi_n_4992 ,csa_tree_add_190_195_groupi_n_6950);
  and csa_tree_add_190_195_groupi_g41922(csa_tree_add_190_195_groupi_n_7040 ,csa_tree_add_190_195_groupi_n_4992 ,csa_tree_add_190_195_groupi_n_6950);
  and csa_tree_add_190_195_groupi_g41923(csa_tree_add_190_195_groupi_n_7039 ,csa_tree_add_190_195_groupi_n_3376 ,csa_tree_add_190_195_groupi_n_6977);
  or csa_tree_add_190_195_groupi_g41924(csa_tree_add_190_195_groupi_n_7038 ,csa_tree_add_190_195_groupi_n_3407 ,csa_tree_add_190_195_groupi_n_7003);
  and csa_tree_add_190_195_groupi_g41925(csa_tree_add_190_195_groupi_n_7037 ,csa_tree_add_190_195_groupi_n_5199 ,csa_tree_add_190_195_groupi_n_6763);
  nor csa_tree_add_190_195_groupi_g41926(csa_tree_add_190_195_groupi_n_7036 ,csa_tree_add_190_195_groupi_n_5839 ,csa_tree_add_190_195_groupi_n_6991);
  and csa_tree_add_190_195_groupi_g41927(csa_tree_add_190_195_groupi_n_7035 ,csa_tree_add_190_195_groupi_n_7011 ,csa_tree_add_190_195_groupi_n_6253);
  xnor csa_tree_add_190_195_groupi_g41928(csa_tree_add_190_195_groupi_n_7034 ,csa_tree_add_190_195_groupi_n_6283 ,csa_tree_add_190_195_groupi_n_5228);
  xnor csa_tree_add_190_195_groupi_g41929(csa_tree_add_190_195_groupi_n_7033 ,csa_tree_add_190_195_groupi_n_6270 ,csa_tree_add_190_195_groupi_n_2016);
  xnor csa_tree_add_190_195_groupi_g41930(csa_tree_add_190_195_groupi_n_7032 ,csa_tree_add_190_195_groupi_n_41 ,csa_tree_add_190_195_groupi_n_5289);
  xnor csa_tree_add_190_195_groupi_g41931(csa_tree_add_190_195_groupi_n_7031 ,csa_tree_add_190_195_groupi_n_6287 ,csa_tree_add_190_195_groupi_n_1941);
  xnor csa_tree_add_190_195_groupi_g41932(csa_tree_add_190_195_groupi_n_7030 ,csa_tree_add_190_195_groupi_n_6289 ,csa_tree_add_190_195_groupi_n_1236);
  xnor csa_tree_add_190_195_groupi_g41933(csa_tree_add_190_195_groupi_n_7029 ,csa_tree_add_190_195_groupi_n_6290 ,csa_tree_add_190_195_groupi_n_5265);
  xnor csa_tree_add_190_195_groupi_g41934(csa_tree_add_190_195_groupi_n_7028 ,csa_tree_add_190_195_groupi_n_27 ,csa_tree_add_190_195_groupi_n_6264);
  xnor csa_tree_add_190_195_groupi_g41935(csa_tree_add_190_195_groupi_n_7027 ,csa_tree_add_190_195_groupi_n_5002 ,csa_tree_add_190_195_groupi_n_6591);
  xnor csa_tree_add_190_195_groupi_g41936(csa_tree_add_190_195_groupi_n_7026 ,csa_tree_add_190_195_groupi_n_4714 ,csa_tree_add_190_195_groupi_n_6587);
  xnor csa_tree_add_190_195_groupi_g41937(csa_tree_add_190_195_groupi_n_7025 ,csa_tree_add_190_195_groupi_n_4935 ,csa_tree_add_190_195_groupi_n_6583);
  xnor csa_tree_add_190_195_groupi_g41938(csa_tree_add_190_195_groupi_n_7024 ,csa_tree_add_190_195_groupi_n_4786 ,csa_tree_add_190_195_groupi_n_6255);
  xnor csa_tree_add_190_195_groupi_g41939(csa_tree_add_190_195_groupi_n_7023 ,csa_tree_add_190_195_groupi_n_4999 ,csa_tree_add_190_195_groupi_n_6581);
  xnor csa_tree_add_190_195_groupi_g41940(csa_tree_add_190_195_groupi_n_7022 ,csa_tree_add_190_195_groupi_n_31 ,csa_tree_add_190_195_groupi_n_6279);
  xnor csa_tree_add_190_195_groupi_g41941(csa_tree_add_190_195_groupi_n_7021 ,csa_tree_add_190_195_groupi_n_5092 ,csa_tree_add_190_195_groupi_n_6578);
  xnor csa_tree_add_190_195_groupi_g41942(csa_tree_add_190_195_groupi_n_7020 ,csa_tree_add_190_195_groupi_n_5017 ,csa_tree_add_190_195_groupi_n_6282);
  xnor csa_tree_add_190_195_groupi_g41944(csa_tree_add_190_195_groupi_n_7019 ,csa_tree_add_190_195_groupi_n_4591 ,csa_tree_add_190_195_groupi_n_6266);
  xnor csa_tree_add_190_195_groupi_g41946(csa_tree_add_190_195_groupi_n_7018 ,csa_tree_add_190_195_groupi_n_4950 ,csa_tree_add_190_195_groupi_n_6262);
  xnor csa_tree_add_190_195_groupi_g41948(csa_tree_add_190_195_groupi_n_7017 ,csa_tree_add_190_195_groupi_n_4901 ,csa_tree_add_190_195_groupi_n_6285);
  and csa_tree_add_190_195_groupi_g41949(csa_tree_add_190_195_groupi_n_7232 ,csa_tree_add_190_195_groupi_n_6335 ,csa_tree_add_190_195_groupi_n_6733);
  xnor csa_tree_add_190_195_groupi_g41950(csa_tree_add_190_195_groupi_n_7231 ,csa_tree_add_190_195_groupi_n_5123 ,csa_tree_add_190_195_groupi_n_6003);
  xnor csa_tree_add_190_195_groupi_g41951(csa_tree_add_190_195_groupi_n_7229 ,csa_tree_add_190_195_groupi_n_5107 ,csa_tree_add_190_195_groupi_n_6044);
  or csa_tree_add_190_195_groupi_g41952(csa_tree_add_190_195_groupi_n_7228 ,csa_tree_add_190_195_groupi_n_6294 ,csa_tree_add_190_195_groupi_n_6738);
  xnor csa_tree_add_190_195_groupi_g41953(csa_tree_add_190_195_groupi_n_7227 ,csa_tree_add_190_195_groupi_n_5992 ,csa_tree_add_190_195_groupi_n_1973);
  and csa_tree_add_190_195_groupi_g41954(csa_tree_add_190_195_groupi_n_7226 ,csa_tree_add_190_195_groupi_n_6392 ,csa_tree_add_190_195_groupi_n_6730);
  xnor csa_tree_add_190_195_groupi_g41955(csa_tree_add_190_195_groupi_n_7225 ,csa_tree_add_190_195_groupi_n_4829 ,csa_tree_add_190_195_groupi_n_6056);
  xnor csa_tree_add_190_195_groupi_g41956(csa_tree_add_190_195_groupi_n_7224 ,csa_tree_add_190_195_groupi_n_4630 ,csa_tree_add_190_195_groupi_n_6030);
  xnor csa_tree_add_190_195_groupi_g41957(csa_tree_add_190_195_groupi_n_7223 ,csa_tree_add_190_195_groupi_n_6039 ,csa_tree_add_190_195_groupi_n_3690);
  and csa_tree_add_190_195_groupi_g41958(csa_tree_add_190_195_groupi_n_7222 ,csa_tree_add_190_195_groupi_n_6314 ,csa_tree_add_190_195_groupi_n_6740);
  xnor csa_tree_add_190_195_groupi_g41959(csa_tree_add_190_195_groupi_n_7221 ,csa_tree_add_190_195_groupi_n_5256 ,csa_tree_add_190_195_groupi_n_6062);
  xnor csa_tree_add_190_195_groupi_g41961(csa_tree_add_190_195_groupi_n_7218 ,csa_tree_add_190_195_groupi_n_6052 ,csa_tree_add_190_195_groupi_n_1074);
  or csa_tree_add_190_195_groupi_g41962(csa_tree_add_190_195_groupi_n_7216 ,csa_tree_add_190_195_groupi_n_3492 ,csa_tree_add_190_195_groupi_n_6748);
  or csa_tree_add_190_195_groupi_g41963(csa_tree_add_190_195_groupi_n_7215 ,csa_tree_add_190_195_groupi_n_5776 ,csa_tree_add_190_195_groupi_n_6728);
  xnor csa_tree_add_190_195_groupi_g41964(csa_tree_add_190_195_groupi_n_7214 ,csa_tree_add_190_195_groupi_n_6024 ,csa_tree_add_190_195_groupi_n_2084);
  xor csa_tree_add_190_195_groupi_g41965(csa_tree_add_190_195_groupi_n_7213 ,csa_tree_add_190_195_groupi_n_6288 ,csa_tree_add_190_195_groupi_n_3908);
  or csa_tree_add_190_195_groupi_g41966(csa_tree_add_190_195_groupi_n_7212 ,csa_tree_add_190_195_groupi_n_6307 ,csa_tree_add_190_195_groupi_n_6727);
  xnor csa_tree_add_190_195_groupi_g41967(csa_tree_add_190_195_groupi_n_7211 ,csa_tree_add_190_195_groupi_n_5146 ,csa_tree_add_190_195_groupi_n_6060);
  or csa_tree_add_190_195_groupi_g41968(csa_tree_add_190_195_groupi_n_7210 ,csa_tree_add_190_195_groupi_n_6183 ,csa_tree_add_190_195_groupi_n_6726);
  xnor csa_tree_add_190_195_groupi_g41969(csa_tree_add_190_195_groupi_n_7209 ,csa_tree_add_190_195_groupi_n_5391 ,csa_tree_add_190_195_groupi_n_6057);
  xnor csa_tree_add_190_195_groupi_g41970(csa_tree_add_190_195_groupi_n_7207 ,csa_tree_add_190_195_groupi_n_5166 ,csa_tree_add_190_195_groupi_n_6017);
  xnor csa_tree_add_190_195_groupi_g41971(csa_tree_add_190_195_groupi_n_7205 ,csa_tree_add_190_195_groupi_n_4800 ,csa_tree_add_190_195_groupi_n_6074);
  xnor csa_tree_add_190_195_groupi_g41972(csa_tree_add_190_195_groupi_n_7204 ,csa_tree_add_190_195_groupi_n_5966 ,csa_tree_add_190_195_groupi_n_6031);
  xnor csa_tree_add_190_195_groupi_g41973(csa_tree_add_190_195_groupi_n_7202 ,csa_tree_add_190_195_groupi_n_3696 ,csa_tree_add_190_195_groupi_n_6000);
  xnor csa_tree_add_190_195_groupi_g41974(csa_tree_add_190_195_groupi_n_7201 ,csa_tree_add_190_195_groupi_n_5148 ,csa_tree_add_190_195_groupi_n_6040);
  xnor csa_tree_add_190_195_groupi_g41975(csa_tree_add_190_195_groupi_n_7200 ,csa_tree_add_190_195_groupi_n_4879 ,csa_tree_add_190_195_groupi_n_6032);
  xnor csa_tree_add_190_195_groupi_g41976(csa_tree_add_190_195_groupi_n_7199 ,csa_tree_add_190_195_groupi_n_5139 ,csa_tree_add_190_195_groupi_n_5991);
  xnor csa_tree_add_190_195_groupi_g41978(csa_tree_add_190_195_groupi_n_7198 ,csa_tree_add_190_195_groupi_n_6584 ,csa_tree_add_190_195_groupi_n_6048);
  xnor csa_tree_add_190_195_groupi_g41980(csa_tree_add_190_195_groupi_n_7197 ,csa_tree_add_190_195_groupi_n_6058 ,csa_tree_add_190_195_groupi_n_1968);
  xnor csa_tree_add_190_195_groupi_g41981(csa_tree_add_190_195_groupi_n_7196 ,csa_tree_add_190_195_groupi_n_4799 ,csa_tree_add_190_195_groupi_n_6063);
  xnor csa_tree_add_190_195_groupi_g41983(csa_tree_add_190_195_groupi_n_7195 ,csa_tree_add_190_195_groupi_n_5984 ,csa_tree_add_190_195_groupi_n_1817);
  or csa_tree_add_190_195_groupi_g41984(csa_tree_add_190_195_groupi_n_7194 ,csa_tree_add_190_195_groupi_n_5627 ,csa_tree_add_190_195_groupi_n_6734);
  xnor csa_tree_add_190_195_groupi_g41985(csa_tree_add_190_195_groupi_n_7193 ,csa_tree_add_190_195_groupi_n_4827 ,csa_tree_add_190_195_groupi_n_6045);
  xnor csa_tree_add_190_195_groupi_g41986(csa_tree_add_190_195_groupi_n_7191 ,csa_tree_add_190_195_groupi_n_5160 ,csa_tree_add_190_195_groupi_n_6013);
  xnor csa_tree_add_190_195_groupi_g41987(csa_tree_add_190_195_groupi_n_7190 ,csa_tree_add_190_195_groupi_n_4679 ,csa_tree_add_190_195_groupi_n_6036);
  xnor csa_tree_add_190_195_groupi_g41988(csa_tree_add_190_195_groupi_n_7188 ,csa_tree_add_190_195_groupi_n_4636 ,csa_tree_add_190_195_groupi_n_6019);
  xnor csa_tree_add_190_195_groupi_g41989(csa_tree_add_190_195_groupi_n_7186 ,csa_tree_add_190_195_groupi_n_4804 ,csa_tree_add_190_195_groupi_n_6023);
  xnor csa_tree_add_190_195_groupi_g41990(csa_tree_add_190_195_groupi_n_7184 ,csa_tree_add_190_195_groupi_n_4837 ,csa_tree_add_190_195_groupi_n_5999);
  xnor csa_tree_add_190_195_groupi_g41991(csa_tree_add_190_195_groupi_n_7183 ,csa_tree_add_190_195_groupi_n_55 ,csa_tree_add_190_195_groupi_n_6016);
  xnor csa_tree_add_190_195_groupi_g41992(csa_tree_add_190_195_groupi_n_7182 ,csa_tree_add_190_195_groupi_n_6034 ,csa_tree_add_190_195_groupi_n_3694);
  xnor csa_tree_add_190_195_groupi_g41993(csa_tree_add_190_195_groupi_n_7180 ,csa_tree_add_190_195_groupi_n_4660 ,csa_tree_add_190_195_groupi_n_6009);
  xnor csa_tree_add_190_195_groupi_g41994(csa_tree_add_190_195_groupi_n_7179 ,csa_tree_add_190_195_groupi_n_4821 ,csa_tree_add_190_195_groupi_n_6007);
  xnor csa_tree_add_190_195_groupi_g41995(csa_tree_add_190_195_groupi_n_7177 ,csa_tree_add_190_195_groupi_n_6041 ,csa_tree_add_190_195_groupi_n_604);
  xnor csa_tree_add_190_195_groupi_g41996(csa_tree_add_190_195_groupi_n_7176 ,csa_tree_add_190_195_groupi_n_5998 ,csa_tree_add_190_195_groupi_n_2210);
  xnor csa_tree_add_190_195_groupi_g41997(csa_tree_add_190_195_groupi_n_7173 ,csa_tree_add_190_195_groupi_n_5011 ,csa_tree_add_190_195_groupi_n_6014);
  xnor csa_tree_add_190_195_groupi_g41998(csa_tree_add_190_195_groupi_n_7171 ,csa_tree_add_190_195_groupi_n_4822 ,csa_tree_add_190_195_groupi_n_6078);
  xnor csa_tree_add_190_195_groupi_g42000(csa_tree_add_190_195_groupi_n_7170 ,csa_tree_add_190_195_groupi_n_4728 ,csa_tree_add_190_195_groupi_n_5997);
  xnor csa_tree_add_190_195_groupi_g42001(csa_tree_add_190_195_groupi_n_7168 ,csa_tree_add_190_195_groupi_n_4683 ,csa_tree_add_190_195_groupi_n_6051);
  xnor csa_tree_add_190_195_groupi_g42002(csa_tree_add_190_195_groupi_n_7165 ,csa_tree_add_190_195_groupi_n_6582 ,csa_tree_add_190_195_groupi_n_5995);
  xnor csa_tree_add_190_195_groupi_g42003(csa_tree_add_190_195_groupi_n_7163 ,csa_tree_add_190_195_groupi_n_4616 ,csa_tree_add_190_195_groupi_n_6042);
  xnor csa_tree_add_190_195_groupi_g42004(csa_tree_add_190_195_groupi_n_7161 ,csa_tree_add_190_195_groupi_n_4588 ,csa_tree_add_190_195_groupi_n_6027);
  xnor csa_tree_add_190_195_groupi_g42005(csa_tree_add_190_195_groupi_n_7159 ,csa_tree_add_190_195_groupi_n_5108 ,csa_tree_add_190_195_groupi_n_6079);
  xnor csa_tree_add_190_195_groupi_g42006(csa_tree_add_190_195_groupi_n_7158 ,csa_tree_add_190_195_groupi_n_4613 ,csa_tree_add_190_195_groupi_n_6072);
  xnor csa_tree_add_190_195_groupi_g42007(csa_tree_add_190_195_groupi_n_7155 ,csa_tree_add_190_195_groupi_n_4917 ,csa_tree_add_190_195_groupi_n_6025);
  xnor csa_tree_add_190_195_groupi_g42008(csa_tree_add_190_195_groupi_n_7154 ,csa_tree_add_190_195_groupi_n_5 ,csa_tree_add_190_195_groupi_n_3846);
  xnor csa_tree_add_190_195_groupi_g42009(csa_tree_add_190_195_groupi_n_7153 ,csa_tree_add_190_195_groupi_n_88 ,csa_tree_add_190_195_groupi_n_2083);
  xnor csa_tree_add_190_195_groupi_g42010(csa_tree_add_190_195_groupi_n_7152 ,csa_tree_add_190_195_groupi_n_6054 ,csa_tree_add_190_195_groupi_n_1848);
  xnor csa_tree_add_190_195_groupi_g42012(csa_tree_add_190_195_groupi_n_7150 ,csa_tree_add_190_195_groupi_n_6020 ,csa_tree_add_190_195_groupi_n_1571);
  xnor csa_tree_add_190_195_groupi_g42013(csa_tree_add_190_195_groupi_n_7149 ,csa_tree_add_190_195_groupi_n_5903 ,csa_tree_add_190_195_groupi_n_6047);
  xnor csa_tree_add_190_195_groupi_g42014(csa_tree_add_190_195_groupi_n_7147 ,csa_tree_add_190_195_groupi_n_5105 ,csa_tree_add_190_195_groupi_n_6082);
  xnor csa_tree_add_190_195_groupi_g42015(csa_tree_add_190_195_groupi_n_7146 ,csa_tree_add_190_195_groupi_n_5987 ,csa_tree_add_190_195_groupi_n_1249);
  xnor csa_tree_add_190_195_groupi_g42016(csa_tree_add_190_195_groupi_n_7143 ,csa_tree_add_190_195_groupi_n_5122 ,csa_tree_add_190_195_groupi_n_6035);
  xnor csa_tree_add_190_195_groupi_g42017(csa_tree_add_190_195_groupi_n_7142 ,csa_tree_add_190_195_groupi_n_4833 ,csa_tree_add_190_195_groupi_n_6021);
  xnor csa_tree_add_190_195_groupi_g42018(csa_tree_add_190_195_groupi_n_7140 ,csa_tree_add_190_195_groupi_n_4796 ,csa_tree_add_190_195_groupi_n_6061);
  xnor csa_tree_add_190_195_groupi_g42019(csa_tree_add_190_195_groupi_n_7138 ,csa_tree_add_190_195_groupi_n_4750 ,csa_tree_add_190_195_groupi_n_6018);
  xnor csa_tree_add_190_195_groupi_g42020(csa_tree_add_190_195_groupi_n_7136 ,csa_tree_add_190_195_groupi_n_6064 ,csa_tree_add_190_195_groupi_n_2215);
  xnor csa_tree_add_190_195_groupi_g42021(csa_tree_add_190_195_groupi_n_7135 ,csa_tree_add_190_195_groupi_n_4758 ,csa_tree_add_190_195_groupi_n_6012);
  xnor csa_tree_add_190_195_groupi_g42022(csa_tree_add_190_195_groupi_n_7134 ,csa_tree_add_190_195_groupi_n_4836 ,csa_tree_add_190_195_groupi_n_6010);
  xnor csa_tree_add_190_195_groupi_g42023(csa_tree_add_190_195_groupi_n_7132 ,csa_tree_add_190_195_groupi_n_4845 ,csa_tree_add_190_195_groupi_n_6015);
  xnor csa_tree_add_190_195_groupi_g42024(csa_tree_add_190_195_groupi_n_7130 ,csa_tree_add_190_195_groupi_n_5134 ,csa_tree_add_190_195_groupi_n_5990);
  xnor csa_tree_add_190_195_groupi_g42025(csa_tree_add_190_195_groupi_n_7129 ,csa_tree_add_190_195_groupi_n_5949 ,csa_tree_add_190_195_groupi_n_6080);
  xnor csa_tree_add_190_195_groupi_g42026(csa_tree_add_190_195_groupi_n_7126 ,csa_tree_add_190_195_groupi_n_5055 ,csa_tree_add_190_195_groupi_n_6037);
  xnor csa_tree_add_190_195_groupi_g42027(csa_tree_add_190_195_groupi_n_7124 ,csa_tree_add_190_195_groupi_n_6592 ,csa_tree_add_190_195_groupi_n_6008);
  xnor csa_tree_add_190_195_groupi_g42028(csa_tree_add_190_195_groupi_n_7122 ,csa_tree_add_190_195_groupi_n_5144 ,csa_tree_add_190_195_groupi_n_6050);
  xnor csa_tree_add_190_195_groupi_g42029(csa_tree_add_190_195_groupi_n_7121 ,csa_tree_add_190_195_groupi_n_6065 ,csa_tree_add_190_195_groupi_n_1673);
  xnor csa_tree_add_190_195_groupi_g42030(csa_tree_add_190_195_groupi_n_7119 ,csa_tree_add_190_195_groupi_n_6046 ,csa_tree_add_190_195_groupi_n_1931);
  xnor csa_tree_add_190_195_groupi_g42031(csa_tree_add_190_195_groupi_n_7117 ,csa_tree_add_190_195_groupi_n_4697 ,csa_tree_add_190_195_groupi_n_6049);
  xnor csa_tree_add_190_195_groupi_g42032(csa_tree_add_190_195_groupi_n_7115 ,csa_tree_add_190_195_groupi_n_4667 ,csa_tree_add_190_195_groupi_n_6005);
  xnor csa_tree_add_190_195_groupi_g42033(csa_tree_add_190_195_groupi_n_7113 ,csa_tree_add_190_195_groupi_n_5418 ,csa_tree_add_190_195_groupi_n_6004);
  xnor csa_tree_add_190_195_groupi_g42034(csa_tree_add_190_195_groupi_n_7111 ,csa_tree_add_190_195_groupi_n_4751 ,csa_tree_add_190_195_groupi_n_6006);
  xnor csa_tree_add_190_195_groupi_g42035(csa_tree_add_190_195_groupi_n_7109 ,csa_tree_add_190_195_groupi_n_5096 ,csa_tree_add_190_195_groupi_n_6081);
  xnor csa_tree_add_190_195_groupi_g42036(csa_tree_add_190_195_groupi_n_7108 ,csa_tree_add_190_195_groupi_n_5985 ,csa_tree_add_190_195_groupi_n_1866);
  xnor csa_tree_add_190_195_groupi_g42037(csa_tree_add_190_195_groupi_n_7106 ,csa_tree_add_190_195_groupi_n_4803 ,csa_tree_add_190_195_groupi_n_6001);
  xnor csa_tree_add_190_195_groupi_g42038(csa_tree_add_190_195_groupi_n_7105 ,csa_tree_add_190_195_groupi_n_4665 ,csa_tree_add_190_195_groupi_n_60);
  xnor csa_tree_add_190_195_groupi_g42039(csa_tree_add_190_195_groupi_n_7103 ,csa_tree_add_190_195_groupi_n_11 ,csa_tree_add_190_195_groupi_n_6043);
  xnor csa_tree_add_190_195_groupi_g42040(csa_tree_add_190_195_groupi_n_7101 ,csa_tree_add_190_195_groupi_n_5595 ,csa_tree_add_190_195_groupi_n_6053);
  xnor csa_tree_add_190_195_groupi_g42041(csa_tree_add_190_195_groupi_n_7098 ,csa_tree_add_190_195_groupi_n_5239 ,csa_tree_add_190_195_groupi_n_5994);
  xnor csa_tree_add_190_195_groupi_g42042(csa_tree_add_190_195_groupi_n_7097 ,csa_tree_add_190_195_groupi_n_5112 ,csa_tree_add_190_195_groupi_n_6086);
  xnor csa_tree_add_190_195_groupi_g42043(csa_tree_add_190_195_groupi_n_7096 ,csa_tree_add_190_195_groupi_n_4748 ,csa_tree_add_190_195_groupi_n_6067);
  xnor csa_tree_add_190_195_groupi_g42045(csa_tree_add_190_195_groupi_n_7094 ,csa_tree_add_190_195_groupi_n_6076 ,csa_tree_add_190_195_groupi_n_1814);
  xnor csa_tree_add_190_195_groupi_g42046(csa_tree_add_190_195_groupi_n_7092 ,csa_tree_add_190_195_groupi_n_5168 ,csa_tree_add_190_195_groupi_n_5989);
  or csa_tree_add_190_195_groupi_g42047(csa_tree_add_190_195_groupi_n_7091 ,csa_tree_add_190_195_groupi_n_6194 ,csa_tree_add_190_195_groupi_n_6752);
  xnor csa_tree_add_190_195_groupi_g42048(csa_tree_add_190_195_groupi_n_7090 ,csa_tree_add_190_195_groupi_n_4615 ,csa_tree_add_190_195_groupi_n_6071);
  xnor csa_tree_add_190_195_groupi_g42049(csa_tree_add_190_195_groupi_n_7088 ,csa_tree_add_190_195_groupi_n_4967 ,csa_tree_add_190_195_groupi_n_6077);
  and csa_tree_add_190_195_groupi_g42050(csa_tree_add_190_195_groupi_n_7086 ,csa_tree_add_190_195_groupi_n_5698 ,csa_tree_add_190_195_groupi_n_6724);
  xnor csa_tree_add_190_195_groupi_g42051(csa_tree_add_190_195_groupi_n_7085 ,csa_tree_add_190_195_groupi_n_5467 ,csa_tree_add_190_195_groupi_n_6069);
  or csa_tree_add_190_195_groupi_g42052(csa_tree_add_190_195_groupi_n_7083 ,csa_tree_add_190_195_groupi_n_6405 ,csa_tree_add_190_195_groupi_n_6725);
  xnor csa_tree_add_190_195_groupi_g42053(csa_tree_add_190_195_groupi_n_7082 ,csa_tree_add_190_195_groupi_n_6073 ,csa_tree_add_190_195_groupi_n_994);
  or csa_tree_add_190_195_groupi_g42054(csa_tree_add_190_195_groupi_n_7080 ,csa_tree_add_190_195_groupi_n_6537 ,csa_tree_add_190_195_groupi_n_6729);
  or csa_tree_add_190_195_groupi_g42055(csa_tree_add_190_195_groupi_n_7078 ,csa_tree_add_190_195_groupi_n_5800 ,csa_tree_add_190_195_groupi_n_6737);
  xnor csa_tree_add_190_195_groupi_g42056(csa_tree_add_190_195_groupi_n_7077 ,csa_tree_add_190_195_groupi_n_6085 ,csa_tree_add_190_195_groupi_n_1849);
  xnor csa_tree_add_190_195_groupi_g42057(csa_tree_add_190_195_groupi_n_7076 ,csa_tree_add_190_195_groupi_n_4841 ,csa_tree_add_190_195_groupi_n_6083);
  xnor csa_tree_add_190_195_groupi_g42058(csa_tree_add_190_195_groupi_n_7075 ,csa_tree_add_190_195_groupi_n_4811 ,csa_tree_add_190_195_groupi_n_6055);
  xnor csa_tree_add_190_195_groupi_g42059(csa_tree_add_190_195_groupi_n_7073 ,csa_tree_add_190_195_groupi_n_5988 ,csa_tree_add_190_195_groupi_n_2083);
  or csa_tree_add_190_195_groupi_g42060(csa_tree_add_190_195_groupi_n_7072 ,csa_tree_add_190_195_groupi_n_6389 ,csa_tree_add_190_195_groupi_n_6739);
  or csa_tree_add_190_195_groupi_g42061(csa_tree_add_190_195_groupi_n_7070 ,csa_tree_add_190_195_groupi_n_6440 ,csa_tree_add_190_195_groupi_n_6741);
  xnor csa_tree_add_190_195_groupi_g42062(csa_tree_add_190_195_groupi_n_7068 ,csa_tree_add_190_195_groupi_n_4826 ,csa_tree_add_190_195_groupi_n_6068);
  or csa_tree_add_190_195_groupi_g42063(csa_tree_add_190_195_groupi_n_7066 ,csa_tree_add_190_195_groupi_n_6090 ,csa_tree_add_190_195_groupi_n_6744);
  xnor csa_tree_add_190_195_groupi_g42064(csa_tree_add_190_195_groupi_n_7065 ,csa_tree_add_190_195_groupi_n_5965 ,csa_tree_add_190_195_groupi_n_6059);
  or csa_tree_add_190_195_groupi_g42065(csa_tree_add_190_195_groupi_n_7063 ,csa_tree_add_190_195_groupi_n_6113 ,csa_tree_add_190_195_groupi_n_6751);
  or csa_tree_add_190_195_groupi_g42066(csa_tree_add_190_195_groupi_n_7061 ,csa_tree_add_190_195_groupi_n_6115 ,csa_tree_add_190_195_groupi_n_6750);
  not csa_tree_add_190_195_groupi_g42067(csa_tree_add_190_195_groupi_n_7015 ,csa_tree_add_190_195_groupi_n_7014);
  not csa_tree_add_190_195_groupi_g42068(csa_tree_add_190_195_groupi_n_7010 ,csa_tree_add_190_195_groupi_n_7009);
  not csa_tree_add_190_195_groupi_g42069(csa_tree_add_190_195_groupi_n_7006 ,csa_tree_add_190_195_groupi_n_7005);
  not csa_tree_add_190_195_groupi_g42071(csa_tree_add_190_195_groupi_n_6999 ,csa_tree_add_190_195_groupi_n_6998);
  not csa_tree_add_190_195_groupi_g42072(csa_tree_add_190_195_groupi_n_6990 ,csa_tree_add_190_195_groupi_n_6989);
  not csa_tree_add_190_195_groupi_g42073(csa_tree_add_190_195_groupi_n_6984 ,csa_tree_add_190_195_groupi_n_6983);
  not csa_tree_add_190_195_groupi_g42074(csa_tree_add_190_195_groupi_n_6967 ,csa_tree_add_190_195_groupi_n_6968);
  not csa_tree_add_190_195_groupi_g42075(csa_tree_add_190_195_groupi_n_6965 ,csa_tree_add_190_195_groupi_n_6966);
  not csa_tree_add_190_195_groupi_g42076(csa_tree_add_190_195_groupi_n_6961 ,csa_tree_add_190_195_groupi_n_6962);
  not csa_tree_add_190_195_groupi_g42077(csa_tree_add_190_195_groupi_n_6959 ,csa_tree_add_190_195_groupi_n_6960);
  not csa_tree_add_190_195_groupi_g42078(csa_tree_add_190_195_groupi_n_6957 ,csa_tree_add_190_195_groupi_n_6958);
  not csa_tree_add_190_195_groupi_g42079(csa_tree_add_190_195_groupi_n_6955 ,csa_tree_add_190_195_groupi_n_6954);
  not csa_tree_add_190_195_groupi_g42080(csa_tree_add_190_195_groupi_n_6953 ,csa_tree_add_190_195_groupi_n_6952);
  not csa_tree_add_190_195_groupi_g42081(csa_tree_add_190_195_groupi_n_6949 ,csa_tree_add_190_195_groupi_n_6948);
  not csa_tree_add_190_195_groupi_g42082(csa_tree_add_190_195_groupi_n_6946 ,csa_tree_add_190_195_groupi_n_6947);
  not csa_tree_add_190_195_groupi_g42083(csa_tree_add_190_195_groupi_n_6944 ,csa_tree_add_190_195_groupi_n_6945);
  not csa_tree_add_190_195_groupi_g42084(csa_tree_add_190_195_groupi_n_6941 ,csa_tree_add_190_195_groupi_n_6942);
  not csa_tree_add_190_195_groupi_g42085(csa_tree_add_190_195_groupi_n_6939 ,csa_tree_add_190_195_groupi_n_6940);
  not csa_tree_add_190_195_groupi_g42086(csa_tree_add_190_195_groupi_n_6937 ,csa_tree_add_190_195_groupi_n_6938);
  not csa_tree_add_190_195_groupi_g42087(csa_tree_add_190_195_groupi_n_6935 ,csa_tree_add_190_195_groupi_n_6936);
  not csa_tree_add_190_195_groupi_g42088(csa_tree_add_190_195_groupi_n_6933 ,csa_tree_add_190_195_groupi_n_6934);
  not csa_tree_add_190_195_groupi_g42089(csa_tree_add_190_195_groupi_n_6930 ,csa_tree_add_190_195_groupi_n_6931);
  not csa_tree_add_190_195_groupi_g42090(csa_tree_add_190_195_groupi_n_6928 ,csa_tree_add_190_195_groupi_n_6929);
  not csa_tree_add_190_195_groupi_g42091(csa_tree_add_190_195_groupi_n_6927 ,csa_tree_add_190_195_groupi_n_6926);
  not csa_tree_add_190_195_groupi_g42092(csa_tree_add_190_195_groupi_n_6924 ,csa_tree_add_190_195_groupi_n_6925);
  not csa_tree_add_190_195_groupi_g42093(csa_tree_add_190_195_groupi_n_6922 ,csa_tree_add_190_195_groupi_n_6923);
  not csa_tree_add_190_195_groupi_g42094(csa_tree_add_190_195_groupi_n_6920 ,csa_tree_add_190_195_groupi_n_6921);
  not csa_tree_add_190_195_groupi_g42096(csa_tree_add_190_195_groupi_n_6917 ,csa_tree_add_190_195_groupi_n_6918);
  not csa_tree_add_190_195_groupi_g42097(csa_tree_add_190_195_groupi_n_6915 ,csa_tree_add_190_195_groupi_n_6916);
  not csa_tree_add_190_195_groupi_g42098(csa_tree_add_190_195_groupi_n_6914 ,csa_tree_add_190_195_groupi_n_6913);
  not csa_tree_add_190_195_groupi_g42099(csa_tree_add_190_195_groupi_n_6911 ,csa_tree_add_190_195_groupi_n_6910);
  not csa_tree_add_190_195_groupi_g42100(csa_tree_add_190_195_groupi_n_6909 ,csa_tree_add_190_195_groupi_n_6908);
  nor csa_tree_add_190_195_groupi_g42101(csa_tree_add_190_195_groupi_n_6907 ,csa_tree_add_190_195_groupi_n_5151 ,csa_tree_add_190_195_groupi_n_6371);
  and csa_tree_add_190_195_groupi_g42102(csa_tree_add_190_195_groupi_n_6906 ,csa_tree_add_190_195_groupi_n_4612 ,csa_tree_add_190_195_groupi_n_6260);
  or csa_tree_add_190_195_groupi_g42103(csa_tree_add_190_195_groupi_n_6905 ,csa_tree_add_190_195_groupi_n_4612 ,csa_tree_add_190_195_groupi_n_6260);
  or csa_tree_add_190_195_groupi_g42104(csa_tree_add_190_195_groupi_n_6904 ,csa_tree_add_190_195_groupi_n_5589 ,csa_tree_add_190_195_groupi_n_6556);
  or csa_tree_add_190_195_groupi_g42105(csa_tree_add_190_195_groupi_n_6903 ,csa_tree_add_190_195_groupi_n_5555 ,csa_tree_add_190_195_groupi_n_6094);
  and csa_tree_add_190_195_groupi_g42106(csa_tree_add_190_195_groupi_n_6902 ,csa_tree_add_190_195_groupi_n_3055 ,csa_tree_add_190_195_groupi_n_6589);
  or csa_tree_add_190_195_groupi_g42107(csa_tree_add_190_195_groupi_n_6901 ,csa_tree_add_190_195_groupi_n_5174 ,csa_tree_add_190_195_groupi_n_6539);
  or csa_tree_add_190_195_groupi_g42108(csa_tree_add_190_195_groupi_n_6900 ,csa_tree_add_190_195_groupi_n_4805 ,csa_tree_add_190_195_groupi_n_6162);
  or csa_tree_add_190_195_groupi_g42109(csa_tree_add_190_195_groupi_n_6899 ,csa_tree_add_190_195_groupi_n_5831 ,csa_tree_add_190_195_groupi_n_6586);
  or csa_tree_add_190_195_groupi_g42110(csa_tree_add_190_195_groupi_n_6898 ,csa_tree_add_190_195_groupi_n_5585 ,csa_tree_add_190_195_groupi_n_94);
  or csa_tree_add_190_195_groupi_g42111(csa_tree_add_190_195_groupi_n_6897 ,csa_tree_add_190_195_groupi_n_5591 ,csa_tree_add_190_195_groupi_n_6536);
  or csa_tree_add_190_195_groupi_g42112(csa_tree_add_190_195_groupi_n_6896 ,csa_tree_add_190_195_groupi_n_4808 ,csa_tree_add_190_195_groupi_n_6126);
  nor csa_tree_add_190_195_groupi_g42113(csa_tree_add_190_195_groupi_n_6895 ,csa_tree_add_190_195_groupi_n_5967 ,csa_tree_add_190_195_groupi_n_6150);
  or csa_tree_add_190_195_groupi_g42114(csa_tree_add_190_195_groupi_n_6894 ,csa_tree_add_190_195_groupi_n_5583 ,csa_tree_add_190_195_groupi_n_6527);
  nor csa_tree_add_190_195_groupi_g42115(csa_tree_add_190_195_groupi_n_6893 ,csa_tree_add_190_195_groupi_n_5125 ,csa_tree_add_190_195_groupi_n_6505);
  or csa_tree_add_190_195_groupi_g42116(csa_tree_add_190_195_groupi_n_6892 ,csa_tree_add_190_195_groupi_n_5552 ,csa_tree_add_190_195_groupi_n_6123);
  or csa_tree_add_190_195_groupi_g42117(csa_tree_add_190_195_groupi_n_6891 ,csa_tree_add_190_195_groupi_n_5596 ,csa_tree_add_190_195_groupi_n_6120);
  and csa_tree_add_190_195_groupi_g42118(csa_tree_add_190_195_groupi_n_6890 ,csa_tree_add_190_195_groupi_n_5121 ,csa_tree_add_190_195_groupi_n_6520);
  or csa_tree_add_190_195_groupi_g42119(csa_tree_add_190_195_groupi_n_6889 ,csa_tree_add_190_195_groupi_n_5580 ,csa_tree_add_190_195_groupi_n_6511);
  or csa_tree_add_190_195_groupi_g42120(csa_tree_add_190_195_groupi_n_6888 ,csa_tree_add_190_195_groupi_n_5592 ,csa_tree_add_190_195_groupi_n_6507);
  and csa_tree_add_190_195_groupi_g42121(csa_tree_add_190_195_groupi_n_6887 ,csa_tree_add_190_195_groupi_n_5236 ,csa_tree_add_190_195_groupi_n_6267);
  nor csa_tree_add_190_195_groupi_g42122(csa_tree_add_190_195_groupi_n_6886 ,csa_tree_add_190_195_groupi_n_5578 ,csa_tree_add_190_195_groupi_n_6498);
  and csa_tree_add_190_195_groupi_g42123(csa_tree_add_190_195_groupi_n_6885 ,csa_tree_add_190_195_groupi_n_5977 ,csa_tree_add_190_195_groupi_n_6493);
  or csa_tree_add_190_195_groupi_g42124(csa_tree_add_190_195_groupi_n_6884 ,csa_tree_add_190_195_groupi_n_5155 ,csa_tree_add_190_195_groupi_n_6490);
  nor csa_tree_add_190_195_groupi_g42125(csa_tree_add_190_195_groupi_n_6883 ,csa_tree_add_190_195_groupi_n_5098 ,csa_tree_add_190_195_groupi_n_6467);
  or csa_tree_add_190_195_groupi_g42126(csa_tree_add_190_195_groupi_n_6882 ,csa_tree_add_190_195_groupi_n_4864 ,csa_tree_add_190_195_groupi_n_6483);
  nor csa_tree_add_190_195_groupi_g42127(csa_tree_add_190_195_groupi_n_6881 ,csa_tree_add_190_195_groupi_n_5602 ,csa_tree_add_190_195_groupi_n_6135);
  or csa_tree_add_190_195_groupi_g42128(csa_tree_add_190_195_groupi_n_6880 ,csa_tree_add_190_195_groupi_n_5079 ,csa_tree_add_190_195_groupi_n_6572);
  nor csa_tree_add_190_195_groupi_g42129(csa_tree_add_190_195_groupi_n_6879 ,csa_tree_add_190_195_groupi_n_5604 ,csa_tree_add_190_195_groupi_n_6476);
  or csa_tree_add_190_195_groupi_g42130(csa_tree_add_190_195_groupi_n_6878 ,csa_tree_add_190_195_groupi_n_5562 ,csa_tree_add_190_195_groupi_n_6480);
  nor csa_tree_add_190_195_groupi_g42131(csa_tree_add_190_195_groupi_n_6877 ,csa_tree_add_190_195_groupi_n_5078 ,csa_tree_add_190_195_groupi_n_6573);
  or csa_tree_add_190_195_groupi_g42132(csa_tree_add_190_195_groupi_n_6876 ,csa_tree_add_190_195_groupi_n_6580 ,csa_tree_add_190_195_groupi_n_6469);
  or csa_tree_add_190_195_groupi_g42133(csa_tree_add_190_195_groupi_n_6875 ,csa_tree_add_190_195_groupi_n_5571 ,csa_tree_add_190_195_groupi_n_6464);
  nor csa_tree_add_190_195_groupi_g42134(csa_tree_add_190_195_groupi_n_6874 ,csa_tree_add_190_195_groupi_n_5897 ,csa_tree_add_190_195_groupi_n_6279);
  or csa_tree_add_190_195_groupi_g42135(csa_tree_add_190_195_groupi_n_6873 ,csa_tree_add_190_195_groupi_n_31 ,csa_tree_add_190_195_groupi_n_85);
  nor csa_tree_add_190_195_groupi_g42136(csa_tree_add_190_195_groupi_n_6872 ,csa_tree_add_190_195_groupi_n_5114 ,csa_tree_add_190_195_groupi_n_6451);
  or csa_tree_add_190_195_groupi_g42137(csa_tree_add_190_195_groupi_n_6871 ,csa_tree_add_190_195_groupi_n_5326 ,csa_tree_add_190_195_groupi_n_6280);
  nor csa_tree_add_190_195_groupi_g42138(csa_tree_add_190_195_groupi_n_6870 ,csa_tree_add_190_195_groupi_n_4844 ,csa_tree_add_190_195_groupi_n_6431);
  and csa_tree_add_190_195_groupi_g42139(csa_tree_add_190_195_groupi_n_6869 ,csa_tree_add_190_195_groupi_n_6285 ,csa_tree_add_190_195_groupi_n_6447);
  nor csa_tree_add_190_195_groupi_g42140(csa_tree_add_190_195_groupi_n_6868 ,csa_tree_add_190_195_groupi_n_4950 ,csa_tree_add_190_195_groupi_n_6261);
  and csa_tree_add_190_195_groupi_g42141(csa_tree_add_190_195_groupi_n_6867 ,csa_tree_add_190_195_groupi_n_5968 ,csa_tree_add_190_195_groupi_n_6438);
  and csa_tree_add_190_195_groupi_g42142(csa_tree_add_190_195_groupi_n_6866 ,csa_tree_add_190_195_groupi_n_5551 ,csa_tree_add_190_195_groupi_n_6433);
  or csa_tree_add_190_195_groupi_g42143(csa_tree_add_190_195_groupi_n_6865 ,csa_tree_add_190_195_groupi_n_4949 ,csa_tree_add_190_195_groupi_n_6262);
  or csa_tree_add_190_195_groupi_g42144(csa_tree_add_190_195_groupi_n_6864 ,csa_tree_add_190_195_groupi_n_5138 ,csa_tree_add_190_195_groupi_n_6416);
  or csa_tree_add_190_195_groupi_g42145(csa_tree_add_190_195_groupi_n_6863 ,csa_tree_add_190_195_groupi_n_5593 ,csa_tree_add_190_195_groupi_n_6413);
  or csa_tree_add_190_195_groupi_g42146(csa_tree_add_190_195_groupi_n_6862 ,csa_tree_add_190_195_groupi_n_14 ,csa_tree_add_190_195_groupi_n_6263);
  or csa_tree_add_190_195_groupi_g42147(csa_tree_add_190_195_groupi_n_6861 ,csa_tree_add_190_195_groupi_n_26 ,csa_tree_add_190_195_groupi_n_6410);
  and csa_tree_add_190_195_groupi_g42148(csa_tree_add_190_195_groupi_n_6860 ,csa_tree_add_190_195_groupi_n_6582 ,csa_tree_add_190_195_groupi_n_5764);
  nor csa_tree_add_190_195_groupi_g42149(csa_tree_add_190_195_groupi_n_6859 ,csa_tree_add_190_195_groupi_n_4871 ,csa_tree_add_190_195_groupi_n_6406);
  nor csa_tree_add_190_195_groupi_g42150(csa_tree_add_190_195_groupi_n_6858 ,csa_tree_add_190_195_groupi_n_5512 ,csa_tree_add_190_195_groupi_n_6264);
  or csa_tree_add_190_195_groupi_g42151(csa_tree_add_190_195_groupi_n_6857 ,csa_tree_add_190_195_groupi_n_5553 ,csa_tree_add_190_195_groupi_n_6560);
  or csa_tree_add_190_195_groupi_g42152(csa_tree_add_190_195_groupi_n_6856 ,csa_tree_add_190_195_groupi_n_5169 ,csa_tree_add_190_195_groupi_n_6200);
  and csa_tree_add_190_195_groupi_g42153(csa_tree_add_190_195_groupi_n_6855 ,csa_tree_add_190_195_groupi_n_5584 ,csa_tree_add_190_195_groupi_n_6396);
  nor csa_tree_add_190_195_groupi_g42154(csa_tree_add_190_195_groupi_n_6854 ,csa_tree_add_190_195_groupi_n_5147 ,csa_tree_add_190_195_groupi_n_6374);
  or csa_tree_add_190_195_groupi_g42155(csa_tree_add_190_195_groupi_n_6853 ,csa_tree_add_190_195_groupi_n_5588 ,csa_tree_add_190_195_groupi_n_6388);
  or csa_tree_add_190_195_groupi_g42156(csa_tree_add_190_195_groupi_n_6852 ,csa_tree_add_190_195_groupi_n_2016 ,csa_tree_add_190_195_groupi_n_6270);
  or csa_tree_add_190_195_groupi_g42157(csa_tree_add_190_195_groupi_n_6851 ,csa_tree_add_190_195_groupi_n_5860 ,csa_tree_add_190_195_groupi_n_6585);
  nor csa_tree_add_190_195_groupi_g42158(csa_tree_add_190_195_groupi_n_6850 ,csa_tree_add_190_195_groupi_n_3516 ,csa_tree_add_190_195_groupi_n_6289);
  or csa_tree_add_190_195_groupi_g42159(csa_tree_add_190_195_groupi_n_6849 ,csa_tree_add_190_195_groupi_n_2041 ,csa_tree_add_190_195_groupi_n_6268);
  and csa_tree_add_190_195_groupi_g42160(csa_tree_add_190_195_groupi_n_6848 ,csa_tree_add_190_195_groupi_n_5326 ,csa_tree_add_190_195_groupi_n_6280);
  or csa_tree_add_190_195_groupi_g42161(csa_tree_add_190_195_groupi_n_6847 ,csa_tree_add_190_195_groupi_n_5321 ,csa_tree_add_190_195_groupi_n_6275);
  or csa_tree_add_190_195_groupi_g42162(csa_tree_add_190_195_groupi_n_6846 ,csa_tree_add_190_195_groupi_n_5171 ,csa_tree_add_190_195_groupi_n_6359);
  and csa_tree_add_190_195_groupi_g42163(csa_tree_add_190_195_groupi_n_6845 ,csa_tree_add_190_195_groupi_n_5321 ,csa_tree_add_190_195_groupi_n_6275);
  or csa_tree_add_190_195_groupi_g42164(csa_tree_add_190_195_groupi_n_6844 ,csa_tree_add_190_195_groupi_n_5173 ,csa_tree_add_190_195_groupi_n_6362);
  nor csa_tree_add_190_195_groupi_g42165(csa_tree_add_190_195_groupi_n_6843 ,csa_tree_add_190_195_groupi_n_6577 ,csa_tree_add_190_195_groupi_n_5473);
  nor csa_tree_add_190_195_groupi_g42166(csa_tree_add_190_195_groupi_n_6842 ,csa_tree_add_190_195_groupi_n_5725 ,csa_tree_add_190_195_groupi_n_6282);
  and csa_tree_add_190_195_groupi_g42167(csa_tree_add_190_195_groupi_n_6841 ,csa_tree_add_190_195_groupi_n_5100 ,csa_tree_add_190_195_groupi_n_6385);
  nor csa_tree_add_190_195_groupi_g42168(csa_tree_add_190_195_groupi_n_6840 ,csa_tree_add_190_195_groupi_n_2627 ,csa_tree_add_190_195_groupi_n_6269);
  and csa_tree_add_190_195_groupi_g42169(csa_tree_add_190_195_groupi_n_6839 ,csa_tree_add_190_195_groupi_n_2016 ,csa_tree_add_190_195_groupi_n_6270);
  and csa_tree_add_190_195_groupi_g42170(csa_tree_add_190_195_groupi_n_6838 ,csa_tree_add_190_195_groupi_n_4846 ,csa_tree_add_190_195_groupi_n_6331);
  and csa_tree_add_190_195_groupi_g42171(csa_tree_add_190_195_groupi_n_6837 ,csa_tree_add_190_195_groupi_n_5609 ,csa_tree_add_190_195_groupi_n_6337);
  or csa_tree_add_190_195_groupi_g42172(csa_tree_add_190_195_groupi_n_6836 ,csa_tree_add_190_195_groupi_n_5556 ,csa_tree_add_190_195_groupi_n_6478);
  or csa_tree_add_190_195_groupi_g42173(csa_tree_add_190_195_groupi_n_6835 ,csa_tree_add_190_195_groupi_n_5573 ,csa_tree_add_190_195_groupi_n_92);
  or csa_tree_add_190_195_groupi_g42174(csa_tree_add_190_195_groupi_n_6834 ,csa_tree_add_190_195_groupi_n_4825 ,csa_tree_add_190_195_groupi_n_6159);
  and csa_tree_add_190_195_groupi_g42175(csa_tree_add_190_195_groupi_n_6833 ,csa_tree_add_190_195_groupi_n_5126 ,csa_tree_add_190_195_groupi_n_6358);
  or csa_tree_add_190_195_groupi_g42176(csa_tree_add_190_195_groupi_n_6832 ,csa_tree_add_190_195_groupi_n_6579 ,csa_tree_add_190_195_groupi_n_6547);
  or csa_tree_add_190_195_groupi_g42177(csa_tree_add_190_195_groupi_n_6831 ,csa_tree_add_190_195_groupi_n_4824 ,csa_tree_add_190_195_groupi_n_6213);
  or csa_tree_add_190_195_groupi_g42178(csa_tree_add_190_195_groupi_n_6830 ,csa_tree_add_190_195_groupi_n_4733 ,csa_tree_add_190_195_groupi_n_6570);
  nor csa_tree_add_190_195_groupi_g42179(csa_tree_add_190_195_groupi_n_6829 ,csa_tree_add_190_195_groupi_n_4734 ,csa_tree_add_190_195_groupi_n_6571);
  or csa_tree_add_190_195_groupi_g42180(csa_tree_add_190_195_groupi_n_6828 ,csa_tree_add_190_195_groupi_n_5120 ,csa_tree_add_190_195_groupi_n_6491);
  or csa_tree_add_190_195_groupi_g42181(csa_tree_add_190_195_groupi_n_6827 ,csa_tree_add_190_195_groupi_n_5570 ,csa_tree_add_190_195_groupi_n_6311);
  or csa_tree_add_190_195_groupi_g42182(csa_tree_add_190_195_groupi_n_6826 ,csa_tree_add_190_195_groupi_n_5559 ,csa_tree_add_190_195_groupi_n_6349);
  or csa_tree_add_190_195_groupi_g42183(csa_tree_add_190_195_groupi_n_6825 ,csa_tree_add_190_195_groupi_n_5567 ,csa_tree_add_190_195_groupi_n_6308);
  or csa_tree_add_190_195_groupi_g42184(csa_tree_add_190_195_groupi_n_6824 ,csa_tree_add_190_195_groupi_n_5587 ,csa_tree_add_190_195_groupi_n_90);
  or csa_tree_add_190_195_groupi_g42185(csa_tree_add_190_195_groupi_n_6823 ,csa_tree_add_190_195_groupi_n_5557 ,csa_tree_add_190_195_groupi_n_6437);
  and csa_tree_add_190_195_groupi_g42186(csa_tree_add_190_195_groupi_n_6822 ,csa_tree_add_190_195_groupi_n_6591 ,csa_tree_add_190_195_groupi_n_5866);
  or csa_tree_add_190_195_groupi_g42187(csa_tree_add_190_195_groupi_n_6821 ,csa_tree_add_190_195_groupi_n_5574 ,csa_tree_add_190_195_groupi_n_6168);
  or csa_tree_add_190_195_groupi_g42188(csa_tree_add_190_195_groupi_n_6820 ,csa_tree_add_190_195_groupi_n_3094 ,csa_tree_add_190_195_groupi_n_6286);
  and csa_tree_add_190_195_groupi_g42189(csa_tree_add_190_195_groupi_n_6819 ,csa_tree_add_190_195_groupi_n_5117 ,csa_tree_add_190_195_groupi_n_6296);
  and csa_tree_add_190_195_groupi_g42190(csa_tree_add_190_195_groupi_n_6818 ,csa_tree_add_190_195_groupi_n_4860 ,csa_tree_add_190_195_groupi_n_6242);
  or csa_tree_add_190_195_groupi_g42191(csa_tree_add_190_195_groupi_n_6817 ,csa_tree_add_190_195_groupi_n_5558 ,csa_tree_add_190_195_groupi_n_6179);
  or csa_tree_add_190_195_groupi_g42192(csa_tree_add_190_195_groupi_n_6816 ,csa_tree_add_190_195_groupi_n_4854 ,csa_tree_add_190_195_groupi_n_6355);
  nor csa_tree_add_190_195_groupi_g42193(csa_tree_add_190_195_groupi_n_6815 ,csa_tree_add_190_195_groupi_n_5569 ,csa_tree_add_190_195_groupi_n_6403);
  or csa_tree_add_190_195_groupi_g42194(csa_tree_add_190_195_groupi_n_6814 ,csa_tree_add_190_195_groupi_n_5111 ,csa_tree_add_190_195_groupi_n_6186);
  or csa_tree_add_190_195_groupi_g42195(csa_tree_add_190_195_groupi_n_6813 ,csa_tree_add_190_195_groupi_n_5568 ,csa_tree_add_190_195_groupi_n_6378);
  or csa_tree_add_190_195_groupi_g42196(csa_tree_add_190_195_groupi_n_6812 ,csa_tree_add_190_195_groupi_n_4817 ,csa_tree_add_190_195_groupi_n_6104);
  and csa_tree_add_190_195_groupi_g42197(csa_tree_add_190_195_groupi_n_6811 ,csa_tree_add_190_195_groupi_n_2803 ,csa_tree_add_190_195_groupi_n_6288);
  or csa_tree_add_190_195_groupi_g42198(csa_tree_add_190_195_groupi_n_6810 ,csa_tree_add_190_195_groupi_n_5572 ,csa_tree_add_190_195_groupi_n_6563);
  or csa_tree_add_190_195_groupi_g42199(csa_tree_add_190_195_groupi_n_6809 ,csa_tree_add_190_195_groupi_n_5236 ,csa_tree_add_190_195_groupi_n_6267);
  and csa_tree_add_190_195_groupi_g42200(csa_tree_add_190_195_groupi_n_6808 ,csa_tree_add_190_195_groupi_n_4855 ,csa_tree_add_190_195_groupi_n_6459);
  or csa_tree_add_190_195_groupi_g42201(csa_tree_add_190_195_groupi_n_6807 ,csa_tree_add_190_195_groupi_n_6576 ,csa_tree_add_190_195_groupi_n_5474);
  or csa_tree_add_190_195_groupi_g42202(csa_tree_add_190_195_groupi_n_6806 ,csa_tree_add_190_195_groupi_n_5158 ,csa_tree_add_190_195_groupi_n_6209);
  and csa_tree_add_190_195_groupi_g42203(csa_tree_add_190_195_groupi_n_6805 ,csa_tree_add_190_195_groupi_n_4870 ,csa_tree_add_190_195_groupi_n_6461);
  or csa_tree_add_190_195_groupi_g42204(csa_tree_add_190_195_groupi_n_6804 ,csa_tree_add_190_195_groupi_n_6284 ,csa_tree_add_190_195_groupi_n_6182);
  and csa_tree_add_190_195_groupi_g42205(csa_tree_add_190_195_groupi_n_6803 ,csa_tree_add_190_195_groupi_n_16 ,csa_tree_add_190_195_groupi_n_6223);
  and csa_tree_add_190_195_groupi_g42206(csa_tree_add_190_195_groupi_n_6802 ,csa_tree_add_190_195_groupi_n_5969 ,csa_tree_add_190_195_groupi_n_6181);
  or csa_tree_add_190_195_groupi_g42207(csa_tree_add_190_195_groupi_n_6801 ,csa_tree_add_190_195_groupi_n_5565 ,csa_tree_add_190_195_groupi_n_6226);
  or csa_tree_add_190_195_groupi_g42208(csa_tree_add_190_195_groupi_n_6800 ,csa_tree_add_190_195_groupi_n_5566 ,csa_tree_add_190_195_groupi_n_6172);
  or csa_tree_add_190_195_groupi_g42209(csa_tree_add_190_195_groupi_n_6799 ,csa_tree_add_190_195_groupi_n_4816 ,csa_tree_add_190_195_groupi_n_6220);
  or csa_tree_add_190_195_groupi_g42210(csa_tree_add_190_195_groupi_n_6798 ,csa_tree_add_190_195_groupi_n_5563 ,csa_tree_add_190_195_groupi_n_91);
  or csa_tree_add_190_195_groupi_g42211(csa_tree_add_190_195_groupi_n_6797 ,csa_tree_add_190_195_groupi_n_4838 ,csa_tree_add_190_195_groupi_n_6144);
  and csa_tree_add_190_195_groupi_g42212(csa_tree_add_190_195_groupi_n_6796 ,csa_tree_add_190_195_groupi_n_6592 ,csa_tree_add_190_195_groupi_n_5671);
  nor csa_tree_add_190_195_groupi_g42213(csa_tree_add_190_195_groupi_n_6795 ,csa_tree_add_190_195_groupi_n_5560 ,csa_tree_add_190_195_groupi_n_6203);
  or csa_tree_add_190_195_groupi_g42214(csa_tree_add_190_195_groupi_n_6794 ,csa_tree_add_190_195_groupi_n_5554 ,csa_tree_add_190_195_groupi_n_6541);
  or csa_tree_add_190_195_groupi_g42215(csa_tree_add_190_195_groupi_n_6793 ,csa_tree_add_190_195_groupi_n_5608 ,csa_tree_add_190_195_groupi_n_6198);
  and csa_tree_add_190_195_groupi_g42216(csa_tree_add_190_195_groupi_n_6792 ,csa_tree_add_190_195_groupi_n_5167 ,csa_tree_add_190_195_groupi_n_6488);
  and csa_tree_add_190_195_groupi_g42217(csa_tree_add_190_195_groupi_n_7016 ,csa_tree_add_190_195_groupi_n_5655 ,csa_tree_add_190_195_groupi_n_6354);
  or csa_tree_add_190_195_groupi_g42218(csa_tree_add_190_195_groupi_n_7014 ,csa_tree_add_190_195_groupi_n_5630 ,csa_tree_add_190_195_groupi_n_6367);
  or csa_tree_add_190_195_groupi_g42219(csa_tree_add_190_195_groupi_n_7013 ,csa_tree_add_190_195_groupi_n_5734 ,csa_tree_add_190_195_groupi_n_6363);
  or csa_tree_add_190_195_groupi_g42220(csa_tree_add_190_195_groupi_n_7012 ,csa_tree_add_190_195_groupi_n_5709 ,csa_tree_add_190_195_groupi_n_6297);
  or csa_tree_add_190_195_groupi_g42221(csa_tree_add_190_195_groupi_n_7011 ,csa_tree_add_190_195_groupi_n_5769 ,csa_tree_add_190_195_groupi_n_6415);
  or csa_tree_add_190_195_groupi_g42222(csa_tree_add_190_195_groupi_n_7009 ,csa_tree_add_190_195_groupi_n_3427 ,csa_tree_add_190_195_groupi_n_6145);
  or csa_tree_add_190_195_groupi_g42223(csa_tree_add_190_195_groupi_n_7008 ,csa_tree_add_190_195_groupi_n_2751 ,csa_tree_add_190_195_groupi_n_6542);
  or csa_tree_add_190_195_groupi_g42224(csa_tree_add_190_195_groupi_n_7007 ,csa_tree_add_190_195_groupi_n_3422 ,csa_tree_add_190_195_groupi_n_6293);
  or csa_tree_add_190_195_groupi_g42225(csa_tree_add_190_195_groupi_n_7005 ,csa_tree_add_190_195_groupi_n_5631 ,csa_tree_add_190_195_groupi_n_6174);
  or csa_tree_add_190_195_groupi_g42226(csa_tree_add_190_195_groupi_n_7004 ,csa_tree_add_190_195_groupi_n_2945 ,csa_tree_add_190_195_groupi_n_6486);
  and csa_tree_add_190_195_groupi_g42227(csa_tree_add_190_195_groupi_n_7003 ,csa_tree_add_190_195_groupi_n_5854 ,csa_tree_add_190_195_groupi_n_6352);
  and csa_tree_add_190_195_groupi_g42228(csa_tree_add_190_195_groupi_n_7002 ,csa_tree_add_190_195_groupi_n_5694 ,csa_tree_add_190_195_groupi_n_6224);
  or csa_tree_add_190_195_groupi_g42229(csa_tree_add_190_195_groupi_n_7001 ,csa_tree_add_190_195_groupi_n_5813 ,csa_tree_add_190_195_groupi_n_6485);
  and csa_tree_add_190_195_groupi_g42230(csa_tree_add_190_195_groupi_n_7000 ,csa_tree_add_190_195_groupi_n_5785 ,csa_tree_add_190_195_groupi_n_6318);
  or csa_tree_add_190_195_groupi_g42231(csa_tree_add_190_195_groupi_n_6998 ,csa_tree_add_190_195_groupi_n_5781 ,csa_tree_add_190_195_groupi_n_6489);
  and csa_tree_add_190_195_groupi_g42232(csa_tree_add_190_195_groupi_n_6997 ,csa_tree_add_190_195_groupi_n_5789 ,csa_tree_add_190_195_groupi_n_6472);
  and csa_tree_add_190_195_groupi_g42233(csa_tree_add_190_195_groupi_n_6996 ,csa_tree_add_190_195_groupi_n_5665 ,csa_tree_add_190_195_groupi_n_6252);
  and csa_tree_add_190_195_groupi_g42234(csa_tree_add_190_195_groupi_n_6995 ,csa_tree_add_190_195_groupi_n_5763 ,csa_tree_add_190_195_groupi_n_6404);
  or csa_tree_add_190_195_groupi_g42235(csa_tree_add_190_195_groupi_n_6994 ,csa_tree_add_190_195_groupi_n_3567 ,csa_tree_add_190_195_groupi_n_6377);
  or csa_tree_add_190_195_groupi_g42236(csa_tree_add_190_195_groupi_n_6993 ,csa_tree_add_190_195_groupi_n_5727 ,csa_tree_add_190_195_groupi_n_6343);
  or csa_tree_add_190_195_groupi_g42237(csa_tree_add_190_195_groupi_n_6992 ,csa_tree_add_190_195_groupi_n_3634 ,csa_tree_add_190_195_groupi_n_6400);
  and csa_tree_add_190_195_groupi_g42238(csa_tree_add_190_195_groupi_n_6991 ,csa_tree_add_190_195_groupi_n_5837 ,csa_tree_add_190_195_groupi_n_6550);
  or csa_tree_add_190_195_groupi_g42239(csa_tree_add_190_195_groupi_n_6989 ,csa_tree_add_190_195_groupi_n_5858 ,csa_tree_add_190_195_groupi_n_6147);
  or csa_tree_add_190_195_groupi_g42240(csa_tree_add_190_195_groupi_n_6988 ,csa_tree_add_190_195_groupi_n_5856 ,csa_tree_add_190_195_groupi_n_6165);
  and csa_tree_add_190_195_groupi_g42241(csa_tree_add_190_195_groupi_n_6987 ,csa_tree_add_190_195_groupi_n_5752 ,csa_tree_add_190_195_groupi_n_6390);
  and csa_tree_add_190_195_groupi_g42242(csa_tree_add_190_195_groupi_n_6986 ,csa_tree_add_190_195_groupi_n_5805 ,csa_tree_add_190_195_groupi_n_6501);
  and csa_tree_add_190_195_groupi_g42243(csa_tree_add_190_195_groupi_n_6985 ,csa_tree_add_190_195_groupi_n_5863 ,csa_tree_add_190_195_groupi_n_6333);
  or csa_tree_add_190_195_groupi_g42244(csa_tree_add_190_195_groupi_n_6983 ,csa_tree_add_190_195_groupi_n_5826 ,csa_tree_add_190_195_groupi_n_6532);
  and csa_tree_add_190_195_groupi_g42245(csa_tree_add_190_195_groupi_n_6982 ,csa_tree_add_190_195_groupi_n_5841 ,csa_tree_add_190_195_groupi_n_6153);
  and csa_tree_add_190_195_groupi_g42246(csa_tree_add_190_195_groupi_n_6981 ,csa_tree_add_190_195_groupi_n_3378 ,csa_tree_add_190_195_groupi_n_6497);
  and csa_tree_add_190_195_groupi_g42247(csa_tree_add_190_195_groupi_n_6980 ,csa_tree_add_190_195_groupi_n_5620 ,csa_tree_add_190_195_groupi_n_6219);
  and csa_tree_add_190_195_groupi_g42248(csa_tree_add_190_195_groupi_n_6979 ,csa_tree_add_190_195_groupi_n_5726 ,csa_tree_add_190_195_groupi_n_6316);
  or csa_tree_add_190_195_groupi_g42249(csa_tree_add_190_195_groupi_n_6978 ,csa_tree_add_190_195_groupi_n_3021 ,csa_tree_add_190_195_groupi_n_6142);
  or csa_tree_add_190_195_groupi_g42250(csa_tree_add_190_195_groupi_n_6977 ,csa_tree_add_190_195_groupi_n_5859 ,csa_tree_add_190_195_groupi_n_6184);
  and csa_tree_add_190_195_groupi_g42251(csa_tree_add_190_195_groupi_n_6976 ,csa_tree_add_190_195_groupi_n_5801 ,csa_tree_add_190_195_groupi_n_6375);
  or csa_tree_add_190_195_groupi_g42252(csa_tree_add_190_195_groupi_n_6975 ,csa_tree_add_190_195_groupi_n_5822 ,csa_tree_add_190_195_groupi_n_6246);
  or csa_tree_add_190_195_groupi_g42253(csa_tree_add_190_195_groupi_n_6974 ,csa_tree_add_190_195_groupi_n_3100 ,csa_tree_add_190_195_groupi_n_6533);
  or csa_tree_add_190_195_groupi_g42254(csa_tree_add_190_195_groupi_n_6973 ,csa_tree_add_190_195_groupi_n_5711 ,csa_tree_add_190_195_groupi_n_6546);
  and csa_tree_add_190_195_groupi_g42255(csa_tree_add_190_195_groupi_n_6972 ,csa_tree_add_190_195_groupi_n_5852 ,csa_tree_add_190_195_groupi_n_6306);
  and csa_tree_add_190_195_groupi_g42256(csa_tree_add_190_195_groupi_n_6971 ,csa_tree_add_190_195_groupi_n_5613 ,csa_tree_add_190_195_groupi_n_6248);
  and csa_tree_add_190_195_groupi_g42257(csa_tree_add_190_195_groupi_n_6970 ,csa_tree_add_190_195_groupi_n_5637 ,csa_tree_add_190_195_groupi_n_6552);
  or csa_tree_add_190_195_groupi_g42258(csa_tree_add_190_195_groupi_n_6969 ,csa_tree_add_190_195_groupi_n_5691 ,csa_tree_add_190_195_groupi_n_6249);
  or csa_tree_add_190_195_groupi_g42259(csa_tree_add_190_195_groupi_n_6968 ,csa_tree_add_190_195_groupi_n_2757 ,csa_tree_add_190_195_groupi_n_6558);
  and csa_tree_add_190_195_groupi_g42260(csa_tree_add_190_195_groupi_n_6966 ,csa_tree_add_190_195_groupi_n_5682 ,csa_tree_add_190_195_groupi_n_6176);
  or csa_tree_add_190_195_groupi_g42261(csa_tree_add_190_195_groupi_n_6964 ,csa_tree_add_190_195_groupi_n_5668 ,csa_tree_add_190_195_groupi_n_6241);
  and csa_tree_add_190_195_groupi_g42262(csa_tree_add_190_195_groupi_n_6963 ,csa_tree_add_190_195_groupi_n_3017 ,csa_tree_add_190_195_groupi_n_6225);
  or csa_tree_add_190_195_groupi_g42263(csa_tree_add_190_195_groupi_n_6962 ,csa_tree_add_190_195_groupi_n_5695 ,csa_tree_add_190_195_groupi_n_6453);
  and csa_tree_add_190_195_groupi_g42264(csa_tree_add_190_195_groupi_n_6960 ,csa_tree_add_190_195_groupi_n_5703 ,csa_tree_add_190_195_groupi_n_6292);
  and csa_tree_add_190_195_groupi_g42265(csa_tree_add_190_195_groupi_n_6958 ,csa_tree_add_190_195_groupi_n_5701 ,csa_tree_add_190_195_groupi_n_6295);
  and csa_tree_add_190_195_groupi_g42266(csa_tree_add_190_195_groupi_n_6956 ,csa_tree_add_190_195_groupi_n_5707 ,csa_tree_add_190_195_groupi_n_6510);
  or csa_tree_add_190_195_groupi_g42267(csa_tree_add_190_195_groupi_n_6954 ,csa_tree_add_190_195_groupi_n_5705 ,csa_tree_add_190_195_groupi_n_6247);
  and csa_tree_add_190_195_groupi_g42268(csa_tree_add_190_195_groupi_n_6952 ,csa_tree_add_190_195_groupi_n_2837 ,csa_tree_add_190_195_groupi_n_6166);
  or csa_tree_add_190_195_groupi_g42269(csa_tree_add_190_195_groupi_n_6951 ,csa_tree_add_190_195_groupi_n_5714 ,csa_tree_add_190_195_groupi_n_6301);
  and csa_tree_add_190_195_groupi_g42270(csa_tree_add_190_195_groupi_n_6950 ,csa_tree_add_190_195_groupi_n_3655 ,csa_tree_add_190_195_groupi_n_6309);
  or csa_tree_add_190_195_groupi_g42271(csa_tree_add_190_195_groupi_n_6948 ,csa_tree_add_190_195_groupi_n_5740 ,csa_tree_add_190_195_groupi_n_6327);
  or csa_tree_add_190_195_groupi_g42272(csa_tree_add_190_195_groupi_n_6947 ,csa_tree_add_190_195_groupi_n_4873 ,csa_tree_add_190_195_groupi_n_6334);
  and csa_tree_add_190_195_groupi_g42273(csa_tree_add_190_195_groupi_n_6945 ,csa_tree_add_190_195_groupi_n_3715 ,csa_tree_add_190_195_groupi_n_6320);
  or csa_tree_add_190_195_groupi_g42274(csa_tree_add_190_195_groupi_n_6943 ,csa_tree_add_190_195_groupi_n_5775 ,csa_tree_add_190_195_groupi_n_6117);
  or csa_tree_add_190_195_groupi_g42275(csa_tree_add_190_195_groupi_n_6942 ,csa_tree_add_190_195_groupi_n_5723 ,csa_tree_add_190_195_groupi_n_6336);
  or csa_tree_add_190_195_groupi_g42276(csa_tree_add_190_195_groupi_n_6940 ,csa_tree_add_190_195_groupi_n_5690 ,csa_tree_add_190_195_groupi_n_6341);
  and csa_tree_add_190_195_groupi_g42277(csa_tree_add_190_195_groupi_n_6938 ,csa_tree_add_190_195_groupi_n_5754 ,csa_tree_add_190_195_groupi_n_6391);
  and csa_tree_add_190_195_groupi_g42278(csa_tree_add_190_195_groupi_n_6936 ,csa_tree_add_190_195_groupi_n_5767 ,csa_tree_add_190_195_groupi_n_6442);
  or csa_tree_add_190_195_groupi_g42279(csa_tree_add_190_195_groupi_n_6934 ,csa_tree_add_190_195_groupi_n_3643 ,csa_tree_add_190_195_groupi_n_6454);
  or csa_tree_add_190_195_groupi_g42280(csa_tree_add_190_195_groupi_n_6932 ,csa_tree_add_190_195_groupi_n_5756 ,csa_tree_add_190_195_groupi_n_6118);
  or csa_tree_add_190_195_groupi_g42281(csa_tree_add_190_195_groupi_n_6931 ,csa_tree_add_190_195_groupi_n_3064 ,csa_tree_add_190_195_groupi_n_6414);
  or csa_tree_add_190_195_groupi_g42282(csa_tree_add_190_195_groupi_n_6929 ,csa_tree_add_190_195_groupi_n_2930 ,csa_tree_add_190_195_groupi_n_6430);
  or csa_tree_add_190_195_groupi_g42283(csa_tree_add_190_195_groupi_n_6926 ,csa_tree_add_190_195_groupi_n_5862 ,csa_tree_add_190_195_groupi_n_6350);
  or csa_tree_add_190_195_groupi_g42284(csa_tree_add_190_195_groupi_n_6925 ,csa_tree_add_190_195_groupi_n_2754 ,csa_tree_add_190_195_groupi_n_6468);
  or csa_tree_add_190_195_groupi_g42285(csa_tree_add_190_195_groupi_n_6923 ,csa_tree_add_190_195_groupi_n_5657 ,csa_tree_add_190_195_groupi_n_6140);
  and csa_tree_add_190_195_groupi_g42286(csa_tree_add_190_195_groupi_n_6921 ,csa_tree_add_190_195_groupi_n_5678 ,csa_tree_add_190_195_groupi_n_6189);
  and csa_tree_add_190_195_groupi_g42287(csa_tree_add_190_195_groupi_n_6919 ,csa_tree_add_190_195_groupi_n_5792 ,csa_tree_add_190_195_groupi_n_6479);
  or csa_tree_add_190_195_groupi_g42288(csa_tree_add_190_195_groupi_n_6918 ,csa_tree_add_190_195_groupi_n_5807 ,csa_tree_add_190_195_groupi_n_6506);
  or csa_tree_add_190_195_groupi_g42289(csa_tree_add_190_195_groupi_n_6916 ,csa_tree_add_190_195_groupi_n_5850 ,csa_tree_add_190_195_groupi_n_6522);
  or csa_tree_add_190_195_groupi_g42290(csa_tree_add_190_195_groupi_n_6913 ,csa_tree_add_190_195_groupi_n_3007 ,csa_tree_add_190_195_groupi_n_6524);
  or csa_tree_add_190_195_groupi_g42291(csa_tree_add_190_195_groupi_n_6912 ,csa_tree_add_190_195_groupi_n_3044 ,csa_tree_add_190_195_groupi_n_6531);
  or csa_tree_add_190_195_groupi_g42292(csa_tree_add_190_195_groupi_n_6910 ,csa_tree_add_190_195_groupi_n_5663 ,csa_tree_add_190_195_groupi_n_6555);
  or csa_tree_add_190_195_groupi_g42293(csa_tree_add_190_195_groupi_n_6908 ,csa_tree_add_190_195_groupi_n_5748 ,csa_tree_add_190_195_groupi_n_6187);
  not csa_tree_add_190_195_groupi_g42294(csa_tree_add_190_195_groupi_n_6785 ,csa_tree_add_190_195_groupi_n_6784);
  not csa_tree_add_190_195_groupi_g42295(csa_tree_add_190_195_groupi_n_6774 ,csa_tree_add_190_195_groupi_n_6773);
  not csa_tree_add_190_195_groupi_g42296(csa_tree_add_190_195_groupi_n_6772 ,csa_tree_add_190_195_groupi_n_6771);
  not csa_tree_add_190_195_groupi_g42297(csa_tree_add_190_195_groupi_n_6769 ,csa_tree_add_190_195_groupi_n_6770);
  not csa_tree_add_190_195_groupi_g42298(csa_tree_add_190_195_groupi_n_6767 ,csa_tree_add_190_195_groupi_n_6766);
  not csa_tree_add_190_195_groupi_g42299(csa_tree_add_190_195_groupi_n_6765 ,csa_tree_add_190_195_groupi_n_6764);
  not csa_tree_add_190_195_groupi_g42300(csa_tree_add_190_195_groupi_n_6761 ,csa_tree_add_190_195_groupi_n_6762);
  not csa_tree_add_190_195_groupi_g42301(csa_tree_add_190_195_groupi_n_6760 ,csa_tree_add_190_195_groupi_n_6759);
  not csa_tree_add_190_195_groupi_g42302(csa_tree_add_190_195_groupi_n_6758 ,csa_tree_add_190_195_groupi_n_35);
  not csa_tree_add_190_195_groupi_g42303(csa_tree_add_190_195_groupi_n_6755 ,csa_tree_add_190_195_groupi_n_6756);
  not csa_tree_add_190_195_groupi_g42304(csa_tree_add_190_195_groupi_n_6753 ,csa_tree_add_190_195_groupi_n_6754);
  and csa_tree_add_190_195_groupi_g42305(csa_tree_add_190_195_groupi_n_6752 ,csa_tree_add_190_195_groupi_n_4872 ,csa_tree_add_190_195_groupi_n_6192);
  and csa_tree_add_190_195_groupi_g42306(csa_tree_add_190_195_groupi_n_6751 ,csa_tree_add_190_195_groupi_n_49 ,csa_tree_add_190_195_groupi_n_6110);
  nor csa_tree_add_190_195_groupi_g42307(csa_tree_add_190_195_groupi_n_6750 ,csa_tree_add_190_195_groupi_n_5600 ,csa_tree_add_190_195_groupi_n_6107);
  nor csa_tree_add_190_195_groupi_g42308(csa_tree_add_190_195_groupi_n_6749 ,csa_tree_add_190_195_groupi_n_5598 ,csa_tree_add_190_195_groupi_n_6215);
  and csa_tree_add_190_195_groupi_g42309(csa_tree_add_190_195_groupi_n_6748 ,csa_tree_add_190_195_groupi_n_3507 ,csa_tree_add_190_195_groupi_n_6287);
  or csa_tree_add_190_195_groupi_g42310(csa_tree_add_190_195_groupi_n_6747 ,csa_tree_add_190_195_groupi_n_5181 ,csa_tree_add_190_195_groupi_n_6273);
  nor csa_tree_add_190_195_groupi_g42311(csa_tree_add_190_195_groupi_n_6746 ,csa_tree_add_190_195_groupi_n_5180 ,csa_tree_add_190_195_groupi_n_6274);
  or csa_tree_add_190_195_groupi_g42312(csa_tree_add_190_195_groupi_n_6745 ,csa_tree_add_190_195_groupi_n_5579 ,csa_tree_add_190_195_groupi_n_6455);
  and csa_tree_add_190_195_groupi_g42313(csa_tree_add_190_195_groupi_n_6744 ,csa_tree_add_190_195_groupi_n_4820 ,csa_tree_add_190_195_groupi_n_6091);
  nor csa_tree_add_190_195_groupi_g42314(csa_tree_add_190_195_groupi_n_6743 ,csa_tree_add_190_195_groupi_n_4634 ,csa_tree_add_190_195_groupi_n_6281);
  and csa_tree_add_190_195_groupi_g42315(csa_tree_add_190_195_groupi_n_6742 ,csa_tree_add_190_195_groupi_n_4634 ,csa_tree_add_190_195_groupi_n_6281);
  and csa_tree_add_190_195_groupi_g42316(csa_tree_add_190_195_groupi_n_6741 ,csa_tree_add_190_195_groupi_n_5103 ,csa_tree_add_190_195_groupi_n_6332);
  or csa_tree_add_190_195_groupi_g42317(csa_tree_add_190_195_groupi_n_6740 ,csa_tree_add_190_195_groupi_n_5976 ,csa_tree_add_190_195_groupi_n_6313);
  nor csa_tree_add_190_195_groupi_g42318(csa_tree_add_190_195_groupi_n_6739 ,csa_tree_add_190_195_groupi_n_4798 ,csa_tree_add_190_195_groupi_n_6429);
  nor csa_tree_add_190_195_groupi_g42319(csa_tree_add_190_195_groupi_n_6738 ,csa_tree_add_190_195_groupi_n_4859 ,csa_tree_add_190_195_groupi_n_6291);
  and csa_tree_add_190_195_groupi_g42320(csa_tree_add_190_195_groupi_n_6737 ,csa_tree_add_190_195_groupi_n_6578 ,csa_tree_add_190_195_groupi_n_5795);
  and csa_tree_add_190_195_groupi_g42321(csa_tree_add_190_195_groupi_n_6736 ,csa_tree_add_190_195_groupi_n_4591 ,csa_tree_add_190_195_groupi_n_6266);
  or csa_tree_add_190_195_groupi_g42322(csa_tree_add_190_195_groupi_n_6735 ,csa_tree_add_190_195_groupi_n_4591 ,csa_tree_add_190_195_groupi_n_6266);
  and csa_tree_add_190_195_groupi_g42323(csa_tree_add_190_195_groupi_n_6734 ,csa_tree_add_190_195_groupi_n_6583 ,csa_tree_add_190_195_groupi_n_5626);
  or csa_tree_add_190_195_groupi_g42324(csa_tree_add_190_195_groupi_n_6733 ,csa_tree_add_190_195_groupi_n_5156 ,csa_tree_add_190_195_groupi_n_6302);
  or csa_tree_add_190_195_groupi_g42325(csa_tree_add_190_195_groupi_n_6732 ,csa_tree_add_190_195_groupi_n_4786 ,csa_tree_add_190_195_groupi_n_6254);
  nor csa_tree_add_190_195_groupi_g42326(csa_tree_add_190_195_groupi_n_6731 ,csa_tree_add_190_195_groupi_n_4785 ,csa_tree_add_190_195_groupi_n_6255);
  or csa_tree_add_190_195_groupi_g42327(csa_tree_add_190_195_groupi_n_6730 ,csa_tree_add_190_195_groupi_n_41 ,csa_tree_add_190_195_groupi_n_6251);
  nor csa_tree_add_190_195_groupi_g42328(csa_tree_add_190_195_groupi_n_6729 ,csa_tree_add_190_195_groupi_n_5129 ,csa_tree_add_190_195_groupi_n_6518);
  nor csa_tree_add_190_195_groupi_g42329(csa_tree_add_190_195_groupi_n_6728 ,csa_tree_add_190_195_groupi_n_5774 ,csa_tree_add_190_195_groupi_n_6581);
  nor csa_tree_add_190_195_groupi_g42330(csa_tree_add_190_195_groupi_n_6727 ,csa_tree_add_190_195_groupi_n_5165 ,csa_tree_add_190_195_groupi_n_6421);
  and csa_tree_add_190_195_groupi_g42331(csa_tree_add_190_195_groupi_n_6726 ,csa_tree_add_190_195_groupi_n_5127 ,csa_tree_add_190_195_groupi_n_6214);
  nor csa_tree_add_190_195_groupi_g42332(csa_tree_add_190_195_groupi_n_6725 ,csa_tree_add_190_195_groupi_n_5131 ,csa_tree_add_190_195_groupi_n_6402);
  or csa_tree_add_190_195_groupi_g42333(csa_tree_add_190_195_groupi_n_6724 ,csa_tree_add_190_195_groupi_n_6588 ,csa_tree_add_190_195_groupi_n_5730);
  and csa_tree_add_190_195_groupi_g42334(csa_tree_add_190_195_groupi_n_6723 ,csa_tree_add_190_195_groupi_n_6290 ,csa_tree_add_190_195_groupi_n_6230);
  xnor csa_tree_add_190_195_groupi_g42335(csa_tree_add_190_195_groupi_n_6722 ,csa_tree_add_190_195_groupi_n_5233 ,csa_tree_add_190_195_groupi_n_5462);
  xnor csa_tree_add_190_195_groupi_g42336(csa_tree_add_190_195_groupi_n_6721 ,csa_tree_add_190_195_groupi_n_5597 ,csa_tree_add_190_195_groupi_n_1188);
  xnor csa_tree_add_190_195_groupi_g42337(csa_tree_add_190_195_groupi_n_6720 ,csa_tree_add_190_195_groupi_n_5238 ,csa_tree_add_190_195_groupi_n_5210);
  xor csa_tree_add_190_195_groupi_g42338(csa_tree_add_190_195_groupi_n_6719 ,csa_tree_add_190_195_groupi_n_5967 ,csa_tree_add_190_195_groupi_n_5960);
  xnor csa_tree_add_190_195_groupi_g42339(csa_tree_add_190_195_groupi_n_6718 ,csa_tree_add_190_195_groupi_n_5888 ,csa_tree_add_190_195_groupi_n_5542);
  xnor csa_tree_add_190_195_groupi_g42340(csa_tree_add_190_195_groupi_n_6717 ,csa_tree_add_190_195_groupi_n_76 ,csa_tree_add_190_195_groupi_n_6);
  xnor csa_tree_add_190_195_groupi_g42341(csa_tree_add_190_195_groupi_n_6716 ,csa_tree_add_190_195_groupi_n_5572 ,csa_tree_add_190_195_groupi_n_5275);
  xnor csa_tree_add_190_195_groupi_g42342(csa_tree_add_190_195_groupi_n_6715 ,csa_tree_add_190_195_groupi_n_5282 ,csa_tree_add_190_195_groupi_n_5270);
  xnor csa_tree_add_190_195_groupi_g42343(csa_tree_add_190_195_groupi_n_6714 ,csa_tree_add_190_195_groupi_n_5062 ,csa_tree_add_190_195_groupi_n_5540);
  xnor csa_tree_add_190_195_groupi_g42344(csa_tree_add_190_195_groupi_n_6713 ,csa_tree_add_190_195_groupi_n_9 ,csa_tree_add_190_195_groupi_n_5889);
  xnor csa_tree_add_190_195_groupi_g42345(csa_tree_add_190_195_groupi_n_6712 ,csa_tree_add_190_195_groupi_n_5980 ,csa_tree_add_190_195_groupi_n_2056);
  xnor csa_tree_add_190_195_groupi_g42346(csa_tree_add_190_195_groupi_n_6711 ,csa_tree_add_190_195_groupi_n_5908 ,csa_tree_add_190_195_groupi_n_5929);
  xnor csa_tree_add_190_195_groupi_g42347(csa_tree_add_190_195_groupi_n_6710 ,csa_tree_add_190_195_groupi_n_5566 ,csa_tree_add_190_195_groupi_n_5444);
  xnor csa_tree_add_190_195_groupi_g42348(csa_tree_add_190_195_groupi_n_6709 ,csa_tree_add_190_195_groupi_n_5488 ,csa_tree_add_190_195_groupi_n_5599);
  xnor csa_tree_add_190_195_groupi_g42349(csa_tree_add_190_195_groupi_n_6708 ,csa_tree_add_190_195_groupi_n_5205 ,csa_tree_add_190_195_groupi_n_1801);
  xnor csa_tree_add_190_195_groupi_g42350(csa_tree_add_190_195_groupi_n_6707 ,csa_tree_add_190_195_groupi_n_5312 ,csa_tree_add_190_195_groupi_n_29);
  xnor csa_tree_add_190_195_groupi_g42351(csa_tree_add_190_195_groupi_n_6706 ,csa_tree_add_190_195_groupi_n_5036 ,csa_tree_add_190_195_groupi_n_5220);
  xnor csa_tree_add_190_195_groupi_g42352(csa_tree_add_190_195_groupi_n_6705 ,csa_tree_add_190_195_groupi_n_5342 ,csa_tree_add_190_195_groupi_n_5584);
  xnor csa_tree_add_190_195_groupi_g42353(csa_tree_add_190_195_groupi_n_6704 ,csa_tree_add_190_195_groupi_n_5310 ,csa_tree_add_190_195_groupi_n_5899);
  xnor csa_tree_add_190_195_groupi_g42354(csa_tree_add_190_195_groupi_n_6703 ,csa_tree_add_190_195_groupi_n_5322 ,csa_tree_add_190_195_groupi_n_5257);
  xnor csa_tree_add_190_195_groupi_g42355(csa_tree_add_190_195_groupi_n_6702 ,csa_tree_add_190_195_groupi_n_5020 ,csa_tree_add_190_195_groupi_n_38);
  xnor csa_tree_add_190_195_groupi_g42356(csa_tree_add_190_195_groupi_n_6701 ,csa_tree_add_190_195_groupi_n_5570 ,csa_tree_add_190_195_groupi_n_5307);
  xor csa_tree_add_190_195_groupi_g42357(csa_tree_add_190_195_groupi_n_6700 ,csa_tree_add_190_195_groupi_n_5235 ,csa_tree_add_190_195_groupi_n_5120);
  xnor csa_tree_add_190_195_groupi_g42358(csa_tree_add_190_195_groupi_n_6699 ,csa_tree_add_190_195_groupi_n_5590 ,csa_tree_add_190_195_groupi_n_1848);
  xor csa_tree_add_190_195_groupi_g42360(csa_tree_add_190_195_groupi_n_6698 ,csa_tree_add_190_195_groupi_n_5596 ,csa_tree_add_190_195_groupi_n_5203);
  xor csa_tree_add_190_195_groupi_g42361(csa_tree_add_190_195_groupi_n_6697 ,csa_tree_add_190_195_groupi_n_5297 ,csa_tree_add_190_195_groupi_n_4805);
  xnor csa_tree_add_190_195_groupi_g42362(csa_tree_add_190_195_groupi_n_6696 ,csa_tree_add_190_195_groupi_n_5187 ,csa_tree_add_190_195_groupi_n_5478);
  xnor csa_tree_add_190_195_groupi_g42363(csa_tree_add_190_195_groupi_n_6695 ,csa_tree_add_190_195_groupi_n_5431 ,csa_tree_add_190_195_groupi_n_5900);
  xnor csa_tree_add_190_195_groupi_g42364(csa_tree_add_190_195_groupi_n_6694 ,csa_tree_add_190_195_groupi_n_5100 ,csa_tree_add_190_195_groupi_n_5296);
  xnor csa_tree_add_190_195_groupi_g42365(csa_tree_add_190_195_groupi_n_6693 ,csa_tree_add_190_195_groupi_n_5274 ,csa_tree_add_190_195_groupi_n_5344);
  xnor csa_tree_add_190_195_groupi_g42366(csa_tree_add_190_195_groupi_n_6692 ,csa_tree_add_190_195_groupi_n_5362 ,csa_tree_add_190_195_groupi_n_5551);
  xnor csa_tree_add_190_195_groupi_g42367(csa_tree_add_190_195_groupi_n_6691 ,csa_tree_add_190_195_groupi_n_5206 ,csa_tree_add_190_195_groupi_n_1845);
  xnor csa_tree_add_190_195_groupi_g42368(csa_tree_add_190_195_groupi_n_6690 ,csa_tree_add_190_195_groupi_n_5573 ,csa_tree_add_190_195_groupi_n_5422);
  xnor csa_tree_add_190_195_groupi_g42369(csa_tree_add_190_195_groupi_n_6689 ,csa_tree_add_190_195_groupi_n_5610 ,csa_tree_add_190_195_groupi_n_1864);
  xnor csa_tree_add_190_195_groupi_g42370(csa_tree_add_190_195_groupi_n_6688 ,csa_tree_add_190_195_groupi_n_71 ,csa_tree_add_190_195_groupi_n_5191);
  xnor csa_tree_add_190_195_groupi_g42371(csa_tree_add_190_195_groupi_n_6687 ,csa_tree_add_190_195_groupi_n_5318 ,csa_tree_add_190_195_groupi_n_5480);
  xnor csa_tree_add_190_195_groupi_g42372(csa_tree_add_190_195_groupi_n_6686 ,csa_tree_add_190_195_groupi_n_5568 ,csa_tree_add_190_195_groupi_n_5285);
  xnor csa_tree_add_190_195_groupi_g42373(csa_tree_add_190_195_groupi_n_6685 ,csa_tree_add_190_195_groupi_n_5364 ,csa_tree_add_190_195_groupi_n_5338);
  xnor csa_tree_add_190_195_groupi_g42374(csa_tree_add_190_195_groupi_n_6684 ,csa_tree_add_190_195_groupi_n_5325 ,csa_tree_add_190_195_groupi_n_5530);
  xnor csa_tree_add_190_195_groupi_g42375(csa_tree_add_190_195_groupi_n_6683 ,csa_tree_add_190_195_groupi_n_4696 ,csa_tree_add_190_195_groupi_n_5499);
  xnor csa_tree_add_190_195_groupi_g42376(csa_tree_add_190_195_groupi_n_6682 ,csa_tree_add_190_195_groupi_n_4561 ,csa_tree_add_190_195_groupi_n_5580);
  xnor csa_tree_add_190_195_groupi_g42377(csa_tree_add_190_195_groupi_n_6681 ,csa_tree_add_190_195_groupi_n_5255 ,csa_tree_add_190_195_groupi_n_5942);
  xnor csa_tree_add_190_195_groupi_g42378(csa_tree_add_190_195_groupi_n_6680 ,csa_tree_add_190_195_groupi_n_5367 ,csa_tree_add_190_195_groupi_n_5356);
  xnor csa_tree_add_190_195_groupi_g42379(csa_tree_add_190_195_groupi_n_6679 ,csa_tree_add_190_195_groupi_n_5581 ,csa_tree_add_190_195_groupi_n_1865);
  xnor csa_tree_add_190_195_groupi_g42380(csa_tree_add_190_195_groupi_n_6678 ,csa_tree_add_190_195_groupi_n_5345 ,csa_tree_add_190_195_groupi_n_80);
  xor csa_tree_add_190_195_groupi_g42381(csa_tree_add_190_195_groupi_n_6677 ,csa_tree_add_190_195_groupi_n_5201 ,csa_tree_add_190_195_groupi_n_4808);
  xnor csa_tree_add_190_195_groupi_g42382(csa_tree_add_190_195_groupi_n_6676 ,csa_tree_add_190_195_groupi_n_5585 ,csa_tree_add_190_195_groupi_n_37);
  xnor csa_tree_add_190_195_groupi_g42383(csa_tree_add_190_195_groupi_n_6675 ,csa_tree_add_190_195_groupi_n_42 ,csa_tree_add_190_195_groupi_n_5490);
  xnor csa_tree_add_190_195_groupi_g42384(csa_tree_add_190_195_groupi_n_6674 ,csa_tree_add_190_195_groupi_n_5567 ,csa_tree_add_190_195_groupi_n_5373);
  xnor csa_tree_add_190_195_groupi_g42385(csa_tree_add_190_195_groupi_n_6673 ,csa_tree_add_190_195_groupi_n_5347 ,csa_tree_add_190_195_groupi_n_5881);
  xnor csa_tree_add_190_195_groupi_g42386(csa_tree_add_190_195_groupi_n_6672 ,csa_tree_add_190_195_groupi_n_5277 ,csa_tree_add_190_195_groupi_n_5948);
  xnor csa_tree_add_190_195_groupi_g42387(csa_tree_add_190_195_groupi_n_6671 ,csa_tree_add_190_195_groupi_n_5576 ,csa_tree_add_190_195_groupi_n_1930);
  xnor csa_tree_add_190_195_groupi_g42388(csa_tree_add_190_195_groupi_n_6670 ,csa_tree_add_190_195_groupi_n_5611 ,csa_tree_add_190_195_groupi_n_1929);
  xnor csa_tree_add_190_195_groupi_g42389(csa_tree_add_190_195_groupi_n_6669 ,csa_tree_add_190_195_groupi_n_59 ,csa_tree_add_190_195_groupi_n_1137);
  xnor csa_tree_add_190_195_groupi_g42390(csa_tree_add_190_195_groupi_n_6668 ,csa_tree_add_190_195_groupi_n_5369 ,csa_tree_add_190_195_groupi_n_5902);
  xnor csa_tree_add_190_195_groupi_g42391(csa_tree_add_190_195_groupi_n_6667 ,csa_tree_add_190_195_groupi_n_5315 ,csa_tree_add_190_195_groupi_n_5472);
  xnor csa_tree_add_190_195_groupi_g42392(csa_tree_add_190_195_groupi_n_6666 ,csa_tree_add_190_195_groupi_n_5298 ,csa_tree_add_190_195_groupi_n_8);
  xnor csa_tree_add_190_195_groupi_g42393(csa_tree_add_190_195_groupi_n_6665 ,csa_tree_add_190_195_groupi_n_61 ,csa_tree_add_190_195_groupi_n_5476);
  xnor csa_tree_add_190_195_groupi_g42394(csa_tree_add_190_195_groupi_n_6664 ,csa_tree_add_190_195_groupi_n_10 ,csa_tree_add_190_195_groupi_n_5425);
  xnor csa_tree_add_190_195_groupi_g42395(csa_tree_add_190_195_groupi_n_6663 ,csa_tree_add_190_195_groupi_n_5575 ,csa_tree_add_190_195_groupi_n_1813);
  xnor csa_tree_add_190_195_groupi_g42396(csa_tree_add_190_195_groupi_n_6662 ,csa_tree_add_190_195_groupi_n_5970 ,csa_tree_add_190_195_groupi_n_1872);
  xnor csa_tree_add_190_195_groupi_g42397(csa_tree_add_190_195_groupi_n_6661 ,csa_tree_add_190_195_groupi_n_4860 ,csa_tree_add_190_195_groupi_n_5286);
  xnor csa_tree_add_190_195_groupi_g42398(csa_tree_add_190_195_groupi_n_6660 ,csa_tree_add_190_195_groupi_n_5569 ,csa_tree_add_190_195_groupi_n_5292);
  xnor csa_tree_add_190_195_groupi_g42399(csa_tree_add_190_195_groupi_n_6659 ,csa_tree_add_190_195_groupi_n_5351 ,csa_tree_add_190_195_groupi_n_5494);
  xnor csa_tree_add_190_195_groupi_g42400(csa_tree_add_190_195_groupi_n_6658 ,csa_tree_add_190_195_groupi_n_5268 ,csa_tree_add_190_195_groupi_n_5421);
  xnor csa_tree_add_190_195_groupi_g42401(csa_tree_add_190_195_groupi_n_6657 ,csa_tree_add_190_195_groupi_n_5167 ,csa_tree_add_190_195_groupi_n_5329);
  xnor csa_tree_add_190_195_groupi_g42402(csa_tree_add_190_195_groupi_n_6656 ,csa_tree_add_190_195_groupi_n_5982 ,csa_tree_add_190_195_groupi_n_1089);
  xnor csa_tree_add_190_195_groupi_g42403(csa_tree_add_190_195_groupi_n_6655 ,csa_tree_add_190_195_groupi_n_5571 ,csa_tree_add_190_195_groupi_n_5905);
  xnor csa_tree_add_190_195_groupi_g42404(csa_tree_add_190_195_groupi_n_6654 ,csa_tree_add_190_195_groupi_n_5244 ,csa_tree_add_190_195_groupi_n_5550);
  xnor csa_tree_add_190_195_groupi_g42405(csa_tree_add_190_195_groupi_n_6653 ,csa_tree_add_190_195_groupi_n_5214 ,csa_tree_add_190_195_groupi_n_5548);
  xnor csa_tree_add_190_195_groupi_g42406(csa_tree_add_190_195_groupi_n_6652 ,csa_tree_add_190_195_groupi_n_5399 ,csa_tree_add_190_195_groupi_n_5869);
  xnor csa_tree_add_190_195_groupi_g42407(csa_tree_add_190_195_groupi_n_6651 ,csa_tree_add_190_195_groupi_n_5574 ,csa_tree_add_190_195_groupi_n_5198);
  xnor csa_tree_add_190_195_groupi_g42408(csa_tree_add_190_195_groupi_n_6650 ,csa_tree_add_190_195_groupi_n_5562 ,csa_tree_add_190_195_groupi_n_5520);
  xnor csa_tree_add_190_195_groupi_g42409(csa_tree_add_190_195_groupi_n_6649 ,csa_tree_add_190_195_groupi_n_4855 ,csa_tree_add_190_195_groupi_n_5401);
  xnor csa_tree_add_190_195_groupi_g42410(csa_tree_add_190_195_groupi_n_6648 ,csa_tree_add_190_195_groupi_n_4846 ,csa_tree_add_190_195_groupi_n_5449);
  xnor csa_tree_add_190_195_groupi_g42411(csa_tree_add_190_195_groupi_n_6647 ,csa_tree_add_190_195_groupi_n_5060 ,csa_tree_add_190_195_groupi_n_5910);
  xnor csa_tree_add_190_195_groupi_g42412(csa_tree_add_190_195_groupi_n_6646 ,csa_tree_add_190_195_groupi_n_5560 ,csa_tree_add_190_195_groupi_n_28);
  xnor csa_tree_add_190_195_groupi_g42413(csa_tree_add_190_195_groupi_n_6645 ,csa_tree_add_190_195_groupi_n_5555 ,csa_tree_add_190_195_groupi_n_5920);
  xnor csa_tree_add_190_195_groupi_g42414(csa_tree_add_190_195_groupi_n_6644 ,csa_tree_add_190_195_groupi_n_5563 ,csa_tree_add_190_195_groupi_n_5916);
  xnor csa_tree_add_190_195_groupi_g42415(csa_tree_add_190_195_groupi_n_6643 ,csa_tree_add_190_195_groupi_n_5248 ,csa_tree_add_190_195_groupi_n_5516);
  xnor csa_tree_add_190_195_groupi_g42416(csa_tree_add_190_195_groupi_n_6642 ,csa_tree_add_190_195_groupi_n_5280 ,csa_tree_add_190_195_groupi_n_5959);
  xnor csa_tree_add_190_195_groupi_g42417(csa_tree_add_190_195_groupi_n_6641 ,csa_tree_add_190_195_groupi_n_5024 ,csa_tree_add_190_195_groupi_n_5360);
  xnor csa_tree_add_190_195_groupi_g42418(csa_tree_add_190_195_groupi_n_6640 ,csa_tree_add_190_195_groupi_n_5022 ,csa_tree_add_190_195_groupi_n_5232);
  xnor csa_tree_add_190_195_groupi_g42419(csa_tree_add_190_195_groupi_n_6639 ,csa_tree_add_190_195_groupi_n_5212 ,csa_tree_add_190_195_groupi_n_4115);
  xnor csa_tree_add_190_195_groupi_g42420(csa_tree_add_190_195_groupi_n_6638 ,csa_tree_add_190_195_groupi_n_4661 ,csa_tree_add_190_195_groupi_n_5240);
  xor csa_tree_add_190_195_groupi_g42421(csa_tree_add_190_195_groupi_n_6637 ,csa_tree_add_190_195_groupi_n_5299 ,csa_tree_add_190_195_groupi_n_4824);
  xnor csa_tree_add_190_195_groupi_g42422(csa_tree_add_190_195_groupi_n_6636 ,csa_tree_add_190_195_groupi_n_5975 ,csa_tree_add_190_195_groupi_n_5294);
  xnor csa_tree_add_190_195_groupi_g42423(csa_tree_add_190_195_groupi_n_6635 ,csa_tree_add_190_195_groupi_n_5407 ,csa_tree_add_190_195_groupi_n_5591);
  xnor csa_tree_add_190_195_groupi_g42424(csa_tree_add_190_195_groupi_n_6634 ,csa_tree_add_190_195_groupi_n_5380 ,csa_tree_add_190_195_groupi_n_5155);
  xnor csa_tree_add_190_195_groupi_g42425(csa_tree_add_190_195_groupi_n_6633 ,csa_tree_add_190_195_groupi_n_5374 ,csa_tree_add_190_195_groupi_n_4694);
  xnor csa_tree_add_190_195_groupi_g42426(csa_tree_add_190_195_groupi_n_6632 ,csa_tree_add_190_195_groupi_n_4738 ,csa_tree_add_190_195_groupi_n_5461);
  xnor csa_tree_add_190_195_groupi_g42427(csa_tree_add_190_195_groupi_n_6631 ,csa_tree_add_190_195_groupi_n_5375 ,csa_tree_add_190_195_groupi_n_4787);
  xnor csa_tree_add_190_195_groupi_g42429(csa_tree_add_190_195_groupi_n_6630 ,csa_tree_add_190_195_groupi_n_4682 ,csa_tree_add_190_195_groupi_n_5459);
  xnor csa_tree_add_190_195_groupi_g42430(csa_tree_add_190_195_groupi_n_6629 ,csa_tree_add_190_195_groupi_n_5164 ,csa_tree_add_190_195_groupi_n_5394);
  xnor csa_tree_add_190_195_groupi_g42431(csa_tree_add_190_195_groupi_n_6628 ,csa_tree_add_190_195_groupi_n_4707 ,csa_tree_add_190_195_groupi_n_5207);
  xnor csa_tree_add_190_195_groupi_g42432(csa_tree_add_190_195_groupi_n_6627 ,csa_tree_add_190_195_groupi_n_4650 ,csa_tree_add_190_195_groupi_n_5416);
  xnor csa_tree_add_190_195_groupi_g42433(csa_tree_add_190_195_groupi_n_6626 ,csa_tree_add_190_195_groupi_n_4586 ,csa_tree_add_190_195_groupi_n_5973);
  xnor csa_tree_add_190_195_groupi_g42434(csa_tree_add_190_195_groupi_n_6625 ,csa_tree_add_190_195_groupi_n_4858 ,csa_tree_add_190_195_groupi_n_5313);
  xor csa_tree_add_190_195_groupi_g42435(csa_tree_add_190_195_groupi_n_6624 ,csa_tree_add_190_195_groupi_n_5114 ,csa_tree_add_190_195_groupi_n_54);
  xnor csa_tree_add_190_195_groupi_g42437(csa_tree_add_190_195_groupi_n_6623 ,csa_tree_add_190_195_groupi_n_5464 ,csa_tree_add_190_195_groupi_n_5509);
  xnor csa_tree_add_190_195_groupi_g42439(csa_tree_add_190_195_groupi_n_6622 ,csa_tree_add_190_195_groupi_n_5320 ,csa_tree_add_190_195_groupi_n_1234);
  xnor csa_tree_add_190_195_groupi_g42440(csa_tree_add_190_195_groupi_n_6621 ,csa_tree_add_190_195_groupi_n_5302 ,csa_tree_add_190_195_groupi_n_5217);
  xnor csa_tree_add_190_195_groupi_g42441(csa_tree_add_190_195_groupi_n_6620 ,csa_tree_add_190_195_groupi_n_4960 ,csa_tree_add_190_195_groupi_n_5907);
  xnor csa_tree_add_190_195_groupi_g42442(csa_tree_add_190_195_groupi_n_6619 ,csa_tree_add_190_195_groupi_n_5545 ,csa_tree_add_190_195_groupi_n_5470);
  xnor csa_tree_add_190_195_groupi_g42443(csa_tree_add_190_195_groupi_n_6618 ,csa_tree_add_190_195_groupi_n_5554 ,csa_tree_add_190_195_groupi_n_5242);
  xnor csa_tree_add_190_195_groupi_g42444(csa_tree_add_190_195_groupi_n_6617 ,csa_tree_add_190_195_groupi_n_5511 ,csa_tree_add_190_195_groupi_n_5446);
  xnor csa_tree_add_190_195_groupi_g42445(csa_tree_add_190_195_groupi_n_6616 ,csa_tree_add_190_195_groupi_n_5873 ,csa_tree_add_190_195_groupi_n_5415);
  xnor csa_tree_add_190_195_groupi_g42446(csa_tree_add_190_195_groupi_n_6615 ,csa_tree_add_190_195_groupi_n_5466 ,csa_tree_add_190_195_groupi_n_5465);
  xnor csa_tree_add_190_195_groupi_g42447(csa_tree_add_190_195_groupi_n_6614 ,csa_tree_add_190_195_groupi_n_5181 ,csa_tree_add_190_195_groupi_n_5136);
  xnor csa_tree_add_190_195_groupi_g42448(csa_tree_add_190_195_groupi_n_6613 ,csa_tree_add_190_195_groupi_n_5938 ,csa_tree_add_190_195_groupi_n_5469);
  xnor csa_tree_add_190_195_groupi_g42449(csa_tree_add_190_195_groupi_n_6612 ,csa_tree_add_190_195_groupi_n_5565 ,csa_tree_add_190_195_groupi_n_5260);
  xnor csa_tree_add_190_195_groupi_g42450(csa_tree_add_190_195_groupi_n_6611 ,csa_tree_add_190_195_groupi_n_5612 ,csa_tree_add_190_195_groupi_n_1750);
  xnor csa_tree_add_190_195_groupi_g42451(csa_tree_add_190_195_groupi_n_6610 ,csa_tree_add_190_195_groupi_n_5397 ,csa_tree_add_190_195_groupi_n_5398);
  xnor csa_tree_add_190_195_groupi_g42452(csa_tree_add_190_195_groupi_n_6609 ,csa_tree_add_190_195_groupi_n_5336 ,csa_tree_add_190_195_groupi_n_5443);
  xnor csa_tree_add_190_195_groupi_g42453(csa_tree_add_190_195_groupi_n_6608 ,csa_tree_add_190_195_groupi_n_5524 ,csa_tree_add_190_195_groupi_n_5519);
  xor csa_tree_add_190_195_groupi_g42454(csa_tree_add_190_195_groupi_n_6607 ,csa_tree_add_190_195_groupi_n_5147 ,csa_tree_add_190_195_groupi_n_5876);
  xnor csa_tree_add_190_195_groupi_g42455(csa_tree_add_190_195_groupi_n_6606 ,csa_tree_add_190_195_groupi_n_5924 ,csa_tree_add_190_195_groupi_n_5951);
  xnor csa_tree_add_190_195_groupi_g42456(csa_tree_add_190_195_groupi_n_6605 ,csa_tree_add_190_195_groupi_n_5126 ,csa_tree_add_190_195_groupi_n_5522);
  xnor csa_tree_add_190_195_groupi_g42457(csa_tree_add_190_195_groupi_n_6604 ,csa_tree_add_190_195_groupi_n_4954 ,csa_tree_add_190_195_groupi_n_5937);
  xnor csa_tree_add_190_195_groupi_g42458(csa_tree_add_190_195_groupi_n_6603 ,csa_tree_add_190_195_groupi_n_5946 ,csa_tree_add_190_195_groupi_n_5977);
  xor csa_tree_add_190_195_groupi_g42459(csa_tree_add_190_195_groupi_n_6602 ,csa_tree_add_190_195_groupi_n_5125 ,csa_tree_add_190_195_groupi_n_17);
  xnor csa_tree_add_190_195_groupi_g42460(csa_tree_add_190_195_groupi_n_6601 ,csa_tree_add_190_195_groupi_n_5592 ,csa_tree_add_190_195_groupi_n_5218);
  xor csa_tree_add_190_195_groupi_g42461(csa_tree_add_190_195_groupi_n_6600 ,csa_tree_add_190_195_groupi_n_5604 ,csa_tree_add_190_195_groupi_n_5917);
  xnor csa_tree_add_190_195_groupi_g42462(csa_tree_add_190_195_groupi_n_6599 ,csa_tree_add_190_195_groupi_n_5979 ,csa_tree_add_190_195_groupi_n_1968);
  xnor csa_tree_add_190_195_groupi_g42463(csa_tree_add_190_195_groupi_n_6598 ,csa_tree_add_190_195_groupi_n_5328 ,csa_tree_add_190_195_groupi_n_5169);
  xnor csa_tree_add_190_195_groupi_g42464(csa_tree_add_190_195_groupi_n_6597 ,csa_tree_add_190_195_groupi_n_5427 ,csa_tree_add_190_195_groupi_n_5202);
  xnor csa_tree_add_190_195_groupi_g42465(csa_tree_add_190_195_groupi_n_6596 ,csa_tree_add_190_195_groupi_n_5603 ,csa_tree_add_190_195_groupi_n_493);
  xnor csa_tree_add_190_195_groupi_g42466(csa_tree_add_190_195_groupi_n_6595 ,csa_tree_add_190_195_groupi_n_4927 ,csa_tree_add_190_195_groupi_n_5912);
  xnor csa_tree_add_190_195_groupi_g42467(csa_tree_add_190_195_groupi_n_6594 ,csa_tree_add_190_195_groupi_n_5423 ,csa_tree_add_190_195_groupi_n_5589);
  xnor csa_tree_add_190_195_groupi_g42469(csa_tree_add_190_195_groupi_n_6593 ,csa_tree_add_190_195_groupi_n_48 ,csa_tree_add_190_195_groupi_n_5578);
  or csa_tree_add_190_195_groupi_g42470(csa_tree_add_190_195_groupi_n_6791 ,csa_tree_add_190_195_groupi_n_5824 ,csa_tree_add_190_195_groupi_n_6152);
  or csa_tree_add_190_195_groupi_g42471(csa_tree_add_190_195_groupi_n_6790 ,csa_tree_add_190_195_groupi_n_3410 ,csa_tree_add_190_195_groupi_n_6114);
  xnor csa_tree_add_190_195_groupi_g42472(csa_tree_add_190_195_groupi_n_6789 ,csa_tree_add_190_195_groupi_n_5178 ,csa_tree_add_190_195_groupi_n_417);
  xnor csa_tree_add_190_195_groupi_g42473(csa_tree_add_190_195_groupi_n_6788 ,csa_tree_add_190_195_groupi_n_5577 ,csa_tree_add_190_195_groupi_n_4137);
  xnor csa_tree_add_190_195_groupi_g42474(csa_tree_add_190_195_groupi_n_6787 ,csa_tree_add_190_195_groupi_n_5594 ,csa_tree_add_190_195_groupi_n_3910);
  xnor csa_tree_add_190_195_groupi_g42475(csa_tree_add_190_195_groupi_n_6786 ,csa_tree_add_190_195_groupi_n_5605 ,csa_tree_add_190_195_groupi_n_3754);
  or csa_tree_add_190_195_groupi_g42476(csa_tree_add_190_195_groupi_n_6784 ,csa_tree_add_190_195_groupi_n_5650 ,csa_tree_add_190_195_groupi_n_6125);
  or csa_tree_add_190_195_groupi_g42477(csa_tree_add_190_195_groupi_n_6783 ,csa_tree_add_190_195_groupi_n_5670 ,csa_tree_add_190_195_groupi_n_6477);
  xnor csa_tree_add_190_195_groupi_g42478(csa_tree_add_190_195_groupi_n_6782 ,csa_tree_add_190_195_groupi_n_5175 ,csa_tree_add_190_195_groupi_n_1934);
  xnor csa_tree_add_190_195_groupi_g42479(csa_tree_add_190_195_groupi_n_6781 ,csa_tree_add_190_195_groupi_n_5972 ,csa_tree_add_190_195_groupi_n_3794);
  xnor csa_tree_add_190_195_groupi_g42480(csa_tree_add_190_195_groupi_n_6780 ,csa_tree_add_190_195_groupi_n_5981 ,csa_tree_add_190_195_groupi_n_39);
  and csa_tree_add_190_195_groupi_g42481(csa_tree_add_190_195_groupi_n_6779 ,csa_tree_add_190_195_groupi_n_5643 ,csa_tree_add_190_195_groupi_n_6105);
  and csa_tree_add_190_195_groupi_g42482(csa_tree_add_190_195_groupi_n_6778 ,csa_tree_add_190_195_groupi_n_5622 ,csa_tree_add_190_195_groupi_n_6155);
  and csa_tree_add_190_195_groupi_g42483(csa_tree_add_190_195_groupi_n_6777 ,csa_tree_add_190_195_groupi_n_3027 ,csa_tree_add_190_195_groupi_n_6517);
  xnor csa_tree_add_190_195_groupi_g42484(csa_tree_add_190_195_groupi_n_6776 ,csa_tree_add_190_195_groupi_n_5177 ,csa_tree_add_190_195_groupi_n_2064);
  or csa_tree_add_190_195_groupi_g42485(csa_tree_add_190_195_groupi_n_6775 ,csa_tree_add_190_195_groupi_n_5636 ,csa_tree_add_190_195_groupi_n_6092);
  or csa_tree_add_190_195_groupi_g42486(csa_tree_add_190_195_groupi_n_6773 ,csa_tree_add_190_195_groupi_n_5811 ,csa_tree_add_190_195_groupi_n_6119);
  or csa_tree_add_190_195_groupi_g42487(csa_tree_add_190_195_groupi_n_6771 ,csa_tree_add_190_195_groupi_n_5640 ,csa_tree_add_190_195_groupi_n_6099);
  or csa_tree_add_190_195_groupi_g42488(csa_tree_add_190_195_groupi_n_6770 ,csa_tree_add_190_195_groupi_n_5619 ,csa_tree_add_190_195_groupi_n_6088);
  or csa_tree_add_190_195_groupi_g42489(csa_tree_add_190_195_groupi_n_6768 ,csa_tree_add_190_195_groupi_n_5634 ,csa_tree_add_190_195_groupi_n_6089);
  or csa_tree_add_190_195_groupi_g42490(csa_tree_add_190_195_groupi_n_6766 ,csa_tree_add_190_195_groupi_n_5848 ,csa_tree_add_190_195_groupi_n_6146);
  and csa_tree_add_190_195_groupi_g42491(csa_tree_add_190_195_groupi_n_6764 ,csa_tree_add_190_195_groupi_n_5780 ,csa_tree_add_190_195_groupi_n_6149);
  xnor csa_tree_add_190_195_groupi_g42492(csa_tree_add_190_195_groupi_n_6763 ,csa_tree_add_190_195_groupi_n_5564 ,csa_tree_add_190_195_groupi_n_3815);
  or csa_tree_add_190_195_groupi_g42493(csa_tree_add_190_195_groupi_n_6762 ,csa_tree_add_190_195_groupi_n_5614 ,csa_tree_add_190_195_groupi_n_6127);
  and csa_tree_add_190_195_groupi_g42494(csa_tree_add_190_195_groupi_n_6759 ,csa_tree_add_190_195_groupi_n_5749 ,csa_tree_add_190_195_groupi_n_6231);
  xnor csa_tree_add_190_195_groupi_g42496(csa_tree_add_190_195_groupi_n_6757 ,csa_tree_add_190_195_groupi_n_5561 ,csa_tree_add_190_195_groupi_n_5176);
  or csa_tree_add_190_195_groupi_g42497(csa_tree_add_190_195_groupi_n_6756 ,csa_tree_add_190_195_groupi_n_5716 ,csa_tree_add_190_195_groupi_n_6121);
  xnor csa_tree_add_190_195_groupi_g42498(csa_tree_add_190_195_groupi_n_6754 ,csa_tree_add_190_195_groupi_n_5601 ,csa_tree_add_190_195_groupi_n_4044);
  not csa_tree_add_190_195_groupi_g42499(csa_tree_add_190_195_groupi_n_6588 ,csa_tree_add_190_195_groupi_n_6587);
  not csa_tree_add_190_195_groupi_g42501(csa_tree_add_190_195_groupi_n_6585 ,csa_tree_add_190_195_groupi_n_6584);
  not csa_tree_add_190_195_groupi_g42503(csa_tree_add_190_195_groupi_n_6576 ,csa_tree_add_190_195_groupi_n_6577);
  not csa_tree_add_190_195_groupi_g42504(csa_tree_add_190_195_groupi_n_6574 ,csa_tree_add_190_195_groupi_n_6575);
  not csa_tree_add_190_195_groupi_g42505(csa_tree_add_190_195_groupi_n_6572 ,csa_tree_add_190_195_groupi_n_6573);
  not csa_tree_add_190_195_groupi_g42506(csa_tree_add_190_195_groupi_n_6570 ,csa_tree_add_190_195_groupi_n_6571);
  or csa_tree_add_190_195_groupi_g42507(csa_tree_add_190_195_groupi_n_6569 ,csa_tree_add_190_195_groupi_n_5280 ,csa_tree_add_190_195_groupi_n_5958);
  or csa_tree_add_190_195_groupi_g42508(csa_tree_add_190_195_groupi_n_6568 ,csa_tree_add_190_195_groupi_n_1944 ,csa_tree_add_190_195_groupi_n_5534);
  nor csa_tree_add_190_195_groupi_g42509(csa_tree_add_190_195_groupi_n_6567 ,csa_tree_add_190_195_groupi_n_2503 ,csa_tree_add_190_195_groupi_n_5278);
  and csa_tree_add_190_195_groupi_g42510(csa_tree_add_190_195_groupi_n_6566 ,csa_tree_add_190_195_groupi_n_1460 ,csa_tree_add_190_195_groupi_n_5278);
  or csa_tree_add_190_195_groupi_g42511(csa_tree_add_190_195_groupi_n_6565 ,csa_tree_add_190_195_groupi_n_2152 ,csa_tree_add_190_195_groupi_n_5370);
  or csa_tree_add_190_195_groupi_g42512(csa_tree_add_190_195_groupi_n_6564 ,csa_tree_add_190_195_groupi_n_715 ,csa_tree_add_190_195_groupi_n_5275);
  and csa_tree_add_190_195_groupi_g42513(csa_tree_add_190_195_groupi_n_6563 ,csa_tree_add_190_195_groupi_n_715 ,csa_tree_add_190_195_groupi_n_5275);
  nor csa_tree_add_190_195_groupi_g42514(csa_tree_add_190_195_groupi_n_6562 ,csa_tree_add_190_195_groupi_n_2604 ,csa_tree_add_190_195_groupi_n_5371);
  or csa_tree_add_190_195_groupi_g42515(csa_tree_add_190_195_groupi_n_6561 ,csa_tree_add_190_195_groupi_n_718 ,csa_tree_add_190_195_groupi_n_5206);
  and csa_tree_add_190_195_groupi_g42516(csa_tree_add_190_195_groupi_n_6560 ,csa_tree_add_190_195_groupi_n_718 ,csa_tree_add_190_195_groupi_n_5206);
  or csa_tree_add_190_195_groupi_g42517(csa_tree_add_190_195_groupi_n_6559 ,csa_tree_add_190_195_groupi_n_4886 ,csa_tree_add_190_195_groupi_n_5418);
  nor csa_tree_add_190_195_groupi_g42518(csa_tree_add_190_195_groupi_n_6558 ,csa_tree_add_190_195_groupi_n_3120 ,csa_tree_add_190_195_groupi_n_5590);
  or csa_tree_add_190_195_groupi_g42519(csa_tree_add_190_195_groupi_n_6557 ,csa_tree_add_190_195_groupi_n_1098 ,csa_tree_add_190_195_groupi_n_5423);
  and csa_tree_add_190_195_groupi_g42520(csa_tree_add_190_195_groupi_n_6556 ,csa_tree_add_190_195_groupi_n_1099 ,csa_tree_add_190_195_groupi_n_5423);
  nor csa_tree_add_190_195_groupi_g42521(csa_tree_add_190_195_groupi_n_6555 ,csa_tree_add_190_195_groupi_n_5105 ,csa_tree_add_190_195_groupi_n_5846);
  or csa_tree_add_190_195_groupi_g42522(csa_tree_add_190_195_groupi_n_6554 ,csa_tree_add_190_195_groupi_n_4745 ,csa_tree_add_190_195_groupi_n_5235);
  or csa_tree_add_190_195_groupi_g42523(csa_tree_add_190_195_groupi_n_6553 ,csa_tree_add_190_195_groupi_n_2402 ,csa_tree_add_190_195_groupi_n_5431);
  or csa_tree_add_190_195_groupi_g42524(csa_tree_add_190_195_groupi_n_6552 ,csa_tree_add_190_195_groupi_n_5166 ,csa_tree_add_190_195_groupi_n_5638);
  nor csa_tree_add_190_195_groupi_g42525(csa_tree_add_190_195_groupi_n_6551 ,csa_tree_add_190_195_groupi_n_4127 ,csa_tree_add_190_195_groupi_n_5521);
  or csa_tree_add_190_195_groupi_g42526(csa_tree_add_190_195_groupi_n_6550 ,csa_tree_add_190_195_groupi_n_5161 ,csa_tree_add_190_195_groupi_n_5838);
  or csa_tree_add_190_195_groupi_g42527(csa_tree_add_190_195_groupi_n_6549 ,csa_tree_add_190_195_groupi_n_4651 ,csa_tree_add_190_195_groupi_n_5416);
  and csa_tree_add_190_195_groupi_g42528(csa_tree_add_190_195_groupi_n_6548 ,csa_tree_add_190_195_groupi_n_17 ,csa_tree_add_190_195_groupi_n_5877);
  nor csa_tree_add_190_195_groupi_g42529(csa_tree_add_190_195_groupi_n_6547 ,csa_tree_add_190_195_groupi_n_2690 ,csa_tree_add_190_195_groupi_n_70);
  nor csa_tree_add_190_195_groupi_g42530(csa_tree_add_190_195_groupi_n_6546 ,csa_tree_add_190_195_groupi_n_5148 ,csa_tree_add_190_195_groupi_n_5843);
  or csa_tree_add_190_195_groupi_g42531(csa_tree_add_190_195_groupi_n_6545 ,csa_tree_add_190_195_groupi_n_4759 ,csa_tree_add_190_195_groupi_n_5452);
  or csa_tree_add_190_195_groupi_g42532(csa_tree_add_190_195_groupi_n_6544 ,csa_tree_add_190_195_groupi_n_5035 ,csa_tree_add_190_195_groupi_n_5219);
  and csa_tree_add_190_195_groupi_g42533(csa_tree_add_190_195_groupi_n_6543 ,csa_tree_add_190_195_groupi_n_4759 ,csa_tree_add_190_195_groupi_n_5452);
  and csa_tree_add_190_195_groupi_g42534(csa_tree_add_190_195_groupi_n_6542 ,csa_tree_add_190_195_groupi_n_3025 ,csa_tree_add_190_195_groupi_n_5612);
  and csa_tree_add_190_195_groupi_g42535(csa_tree_add_190_195_groupi_n_6541 ,csa_tree_add_190_195_groupi_n_5243 ,csa_tree_add_190_195_groupi_n_5242);
  or csa_tree_add_190_195_groupi_g42536(csa_tree_add_190_195_groupi_n_6540 ,csa_tree_add_190_195_groupi_n_2403 ,csa_tree_add_190_195_groupi_n_5411);
  and csa_tree_add_190_195_groupi_g42537(csa_tree_add_190_195_groupi_n_6539 ,csa_tree_add_190_195_groupi_n_4886 ,csa_tree_add_190_195_groupi_n_5418);
  or csa_tree_add_190_195_groupi_g42539(csa_tree_add_190_195_groupi_n_6538 ,csa_tree_add_190_195_groupi_n_5408 ,csa_tree_add_190_195_groupi_n_5407);
  nor csa_tree_add_190_195_groupi_g42540(csa_tree_add_190_195_groupi_n_6537 ,csa_tree_add_190_195_groupi_n_5870 ,csa_tree_add_190_195_groupi_n_5399);
  and csa_tree_add_190_195_groupi_g42541(csa_tree_add_190_195_groupi_n_6536 ,csa_tree_add_190_195_groupi_n_5408 ,csa_tree_add_190_195_groupi_n_5407);
  or csa_tree_add_190_195_groupi_g42542(csa_tree_add_190_195_groupi_n_6535 ,csa_tree_add_190_195_groupi_n_5282 ,csa_tree_add_190_195_groupi_n_5270);
  and csa_tree_add_190_195_groupi_g42543(csa_tree_add_190_195_groupi_n_6534 ,csa_tree_add_190_195_groupi_n_5962 ,csa_tree_add_190_195_groupi_n_5960);
  and csa_tree_add_190_195_groupi_g42544(csa_tree_add_190_195_groupi_n_6533 ,csa_tree_add_190_195_groupi_n_3081 ,csa_tree_add_190_195_groupi_n_5979);
  nor csa_tree_add_190_195_groupi_g42545(csa_tree_add_190_195_groupi_n_6532 ,csa_tree_add_190_195_groupi_n_5135 ,csa_tree_add_190_195_groupi_n_5825);
  and csa_tree_add_190_195_groupi_g42546(csa_tree_add_190_195_groupi_n_6531 ,csa_tree_add_190_195_groupi_n_3252 ,csa_tree_add_190_195_groupi_n_5978);
  nor csa_tree_add_190_195_groupi_g42547(csa_tree_add_190_195_groupi_n_6530 ,csa_tree_add_190_195_groupi_n_5544 ,csa_tree_add_190_195_groupi_n_20);
  or csa_tree_add_190_195_groupi_g42548(csa_tree_add_190_195_groupi_n_6529 ,csa_tree_add_190_195_groupi_n_5413 ,csa_tree_add_190_195_groupi_n_5307);
  or csa_tree_add_190_195_groupi_g42549(csa_tree_add_190_195_groupi_n_6528 ,csa_tree_add_190_195_groupi_n_5398 ,csa_tree_add_190_195_groupi_n_5397);
  and csa_tree_add_190_195_groupi_g42550(csa_tree_add_190_195_groupi_n_6527 ,csa_tree_add_190_195_groupi_n_5398 ,csa_tree_add_190_195_groupi_n_5397);
  or csa_tree_add_190_195_groupi_g42551(csa_tree_add_190_195_groupi_n_6526 ,csa_tree_add_190_195_groupi_n_4976 ,csa_tree_add_190_195_groupi_n_5952);
  nor csa_tree_add_190_195_groupi_g42552(csa_tree_add_190_195_groupi_n_6525 ,csa_tree_add_190_195_groupi_n_4977 ,csa_tree_add_190_195_groupi_n_5953);
  nor csa_tree_add_190_195_groupi_g42553(csa_tree_add_190_195_groupi_n_6524 ,csa_tree_add_190_195_groupi_n_3072 ,csa_tree_add_190_195_groupi_n_5582);
  nor csa_tree_add_190_195_groupi_g42554(csa_tree_add_190_195_groupi_n_6523 ,csa_tree_add_190_195_groupi_n_5393 ,csa_tree_add_190_195_groupi_n_5392);
  nor csa_tree_add_190_195_groupi_g42555(csa_tree_add_190_195_groupi_n_6522 ,csa_tree_add_190_195_groupi_n_5128 ,csa_tree_add_190_195_groupi_n_5849);
  and csa_tree_add_190_195_groupi_g42556(csa_tree_add_190_195_groupi_n_6521 ,csa_tree_add_190_195_groupi_n_5393 ,csa_tree_add_190_195_groupi_n_5392);
  or csa_tree_add_190_195_groupi_g42557(csa_tree_add_190_195_groupi_n_6520 ,csa_tree_add_190_195_groupi_n_4981 ,csa_tree_add_190_195_groupi_n_5390);
  or csa_tree_add_190_195_groupi_g42558(csa_tree_add_190_195_groupi_n_6519 ,csa_tree_add_190_195_groupi_n_5923 ,csa_tree_add_190_195_groupi_n_5950);
  and csa_tree_add_190_195_groupi_g42559(csa_tree_add_190_195_groupi_n_6518 ,csa_tree_add_190_195_groupi_n_5870 ,csa_tree_add_190_195_groupi_n_5399);
  or csa_tree_add_190_195_groupi_g42560(csa_tree_add_190_195_groupi_n_6517 ,csa_tree_add_190_195_groupi_n_2921 ,csa_tree_add_190_195_groupi_n_5581);
  or csa_tree_add_190_195_groupi_g42561(csa_tree_add_190_195_groupi_n_6516 ,csa_tree_add_190_195_groupi_n_5389 ,csa_tree_add_190_195_groupi_n_5388);
  and csa_tree_add_190_195_groupi_g42562(csa_tree_add_190_195_groupi_n_6515 ,csa_tree_add_190_195_groupi_n_5389 ,csa_tree_add_190_195_groupi_n_5388);
  or csa_tree_add_190_195_groupi_g42563(csa_tree_add_190_195_groupi_n_6514 ,csa_tree_add_190_195_groupi_n_5218 ,csa_tree_add_190_195_groupi_n_5385);
  nor csa_tree_add_190_195_groupi_g42564(csa_tree_add_190_195_groupi_n_6513 ,csa_tree_add_190_195_groupi_n_4765 ,csa_tree_add_190_195_groupi_n_5386);
  or csa_tree_add_190_195_groupi_g42565(csa_tree_add_190_195_groupi_n_6512 ,csa_tree_add_190_195_groupi_n_4560 ,csa_tree_add_190_195_groupi_n_5943);
  nor csa_tree_add_190_195_groupi_g42566(csa_tree_add_190_195_groupi_n_6511 ,csa_tree_add_190_195_groupi_n_4561 ,csa_tree_add_190_195_groupi_n_5944);
  or csa_tree_add_190_195_groupi_g42567(csa_tree_add_190_195_groupi_n_6510 ,csa_tree_add_190_195_groupi_n_4843 ,csa_tree_add_190_195_groupi_n_5758);
  or csa_tree_add_190_195_groupi_g42568(csa_tree_add_190_195_groupi_n_6509 ,csa_tree_add_190_195_groupi_n_5255 ,csa_tree_add_190_195_groupi_n_5941);
  nor csa_tree_add_190_195_groupi_g42569(csa_tree_add_190_195_groupi_n_6508 ,csa_tree_add_190_195_groupi_n_5254 ,csa_tree_add_190_195_groupi_n_5942);
  and csa_tree_add_190_195_groupi_g42570(csa_tree_add_190_195_groupi_n_6507 ,csa_tree_add_190_195_groupi_n_5218 ,csa_tree_add_190_195_groupi_n_5385);
  nor csa_tree_add_190_195_groupi_g42571(csa_tree_add_190_195_groupi_n_6506 ,csa_tree_add_190_195_groupi_n_5163 ,csa_tree_add_190_195_groupi_n_5742);
  nor csa_tree_add_190_195_groupi_g42572(csa_tree_add_190_195_groupi_n_6505 ,csa_tree_add_190_195_groupi_n_17 ,csa_tree_add_190_195_groupi_n_5877);
  or csa_tree_add_190_195_groupi_g42573(csa_tree_add_190_195_groupi_n_6504 ,csa_tree_add_190_195_groupi_n_5380 ,csa_tree_add_190_195_groupi_n_5379);
  or csa_tree_add_190_195_groupi_g42574(csa_tree_add_190_195_groupi_n_6503 ,csa_tree_add_190_195_groupi_n_4953 ,csa_tree_add_190_195_groupi_n_5936);
  nor csa_tree_add_190_195_groupi_g42575(csa_tree_add_190_195_groupi_n_6502 ,csa_tree_add_190_195_groupi_n_4954 ,csa_tree_add_190_195_groupi_n_5937);
  or csa_tree_add_190_195_groupi_g42576(csa_tree_add_190_195_groupi_n_6501 ,csa_tree_add_190_195_groupi_n_5153 ,csa_tree_add_190_195_groupi_n_5804);
  nor csa_tree_add_190_195_groupi_g42577(csa_tree_add_190_195_groupi_n_6500 ,csa_tree_add_190_195_groupi_n_5334 ,csa_tree_add_190_195_groupi_n_5935);
  nor csa_tree_add_190_195_groupi_g42578(csa_tree_add_190_195_groupi_n_6499 ,csa_tree_add_190_195_groupi_n_5933 ,csa_tree_add_190_195_groupi_n_48);
  and csa_tree_add_190_195_groupi_g42579(csa_tree_add_190_195_groupi_n_6498 ,csa_tree_add_190_195_groupi_n_5933 ,csa_tree_add_190_195_groupi_n_48);
  or csa_tree_add_190_195_groupi_g42580(csa_tree_add_190_195_groupi_n_6497 ,csa_tree_add_190_195_groupi_n_3356 ,csa_tree_add_190_195_groupi_n_5981);
  nor csa_tree_add_190_195_groupi_g42581(csa_tree_add_190_195_groupi_n_6496 ,csa_tree_add_190_195_groupi_n_5930 ,csa_tree_add_190_195_groupi_n_58);
  or csa_tree_add_190_195_groupi_g42582(csa_tree_add_190_195_groupi_n_6495 ,csa_tree_add_190_195_groupi_n_5931 ,csa_tree_add_190_195_groupi_n_5376);
  nor csa_tree_add_190_195_groupi_g42583(csa_tree_add_190_195_groupi_n_6494 ,csa_tree_add_190_195_groupi_n_5945 ,csa_tree_add_190_195_groupi_n_24);
  or csa_tree_add_190_195_groupi_g42584(csa_tree_add_190_195_groupi_n_6493 ,csa_tree_add_190_195_groupi_n_5946 ,csa_tree_add_190_195_groupi_n_5447);
  or csa_tree_add_190_195_groupi_g42585(csa_tree_add_190_195_groupi_n_6492 ,csa_tree_add_190_195_groupi_n_5233 ,csa_tree_add_190_195_groupi_n_5463);
  nor csa_tree_add_190_195_groupi_g42586(csa_tree_add_190_195_groupi_n_6491 ,csa_tree_add_190_195_groupi_n_4746 ,csa_tree_add_190_195_groupi_n_5234);
  and csa_tree_add_190_195_groupi_g42587(csa_tree_add_190_195_groupi_n_6490 ,csa_tree_add_190_195_groupi_n_5380 ,csa_tree_add_190_195_groupi_n_5379);
  and csa_tree_add_190_195_groupi_g42588(csa_tree_add_190_195_groupi_n_6489 ,csa_tree_add_190_195_groupi_n_4800 ,csa_tree_add_190_195_groupi_n_5783);
  or csa_tree_add_190_195_groupi_g42589(csa_tree_add_190_195_groupi_n_6488 ,csa_tree_add_190_195_groupi_n_2398 ,csa_tree_add_190_195_groupi_n_5546);
  and csa_tree_add_190_195_groupi_g42590(csa_tree_add_190_195_groupi_n_6487 ,csa_tree_add_190_195_groupi_n_5282 ,csa_tree_add_190_195_groupi_n_5270);
  and csa_tree_add_190_195_groupi_g42591(csa_tree_add_190_195_groupi_n_6486 ,csa_tree_add_190_195_groupi_n_2942 ,csa_tree_add_190_195_groupi_n_5982);
  and csa_tree_add_190_195_groupi_g42592(csa_tree_add_190_195_groupi_n_6485 ,csa_tree_add_190_195_groupi_n_5654 ,csa_tree_add_190_195_groupi_n_5966);
  and csa_tree_add_190_195_groupi_g42593(csa_tree_add_190_195_groupi_n_6484 ,csa_tree_add_190_195_groupi_n_5080 ,csa_tree_add_190_195_groupi_n_5903);
  and csa_tree_add_190_195_groupi_g42594(csa_tree_add_190_195_groupi_n_6483 ,csa_tree_add_190_195_groupi_n_4694 ,csa_tree_add_190_195_groupi_n_5374);
  or csa_tree_add_190_195_groupi_g42595(csa_tree_add_190_195_groupi_n_6482 ,csa_tree_add_190_195_groupi_n_5260 ,csa_tree_add_190_195_groupi_n_5259);
  and csa_tree_add_190_195_groupi_g42596(csa_tree_add_190_195_groupi_n_6481 ,csa_tree_add_190_195_groupi_n_5918 ,csa_tree_add_190_195_groupi_n_5917);
  nor csa_tree_add_190_195_groupi_g42597(csa_tree_add_190_195_groupi_n_6480 ,csa_tree_add_190_195_groupi_n_1312 ,csa_tree_add_190_195_groupi_n_18);
  or csa_tree_add_190_195_groupi_g42598(csa_tree_add_190_195_groupi_n_6479 ,csa_tree_add_190_195_groupi_n_4823 ,csa_tree_add_190_195_groupi_n_5791);
  nor csa_tree_add_190_195_groupi_g42599(csa_tree_add_190_195_groupi_n_6478 ,csa_tree_add_190_195_groupi_n_5191 ,csa_tree_add_190_195_groupi_n_5432);
  nor csa_tree_add_190_195_groupi_g42600(csa_tree_add_190_195_groupi_n_6477 ,csa_tree_add_190_195_groupi_n_4847 ,csa_tree_add_190_195_groupi_n_5674);
  nor csa_tree_add_190_195_groupi_g42601(csa_tree_add_190_195_groupi_n_6476 ,csa_tree_add_190_195_groupi_n_5918 ,csa_tree_add_190_195_groupi_n_5917);
  or csa_tree_add_190_195_groupi_g42602(csa_tree_add_190_195_groupi_n_6475 ,csa_tree_add_190_195_groupi_n_5261 ,csa_tree_add_190_195_groupi_n_5914);
  nor csa_tree_add_190_195_groupi_g42603(csa_tree_add_190_195_groupi_n_6474 ,csa_tree_add_190_195_groupi_n_5262 ,csa_tree_add_190_195_groupi_n_5915);
  or csa_tree_add_190_195_groupi_g42604(csa_tree_add_190_195_groupi_n_6473 ,csa_tree_add_190_195_groupi_n_4926 ,csa_tree_add_190_195_groupi_n_5911);
  or csa_tree_add_190_195_groupi_g42605(csa_tree_add_190_195_groupi_n_6472 ,csa_tree_add_190_195_groupi_n_5109 ,csa_tree_add_190_195_groupi_n_5788);
  or csa_tree_add_190_195_groupi_g42606(csa_tree_add_190_195_groupi_n_6471 ,csa_tree_add_190_195_groupi_n_4990 ,csa_tree_add_190_195_groupi_n_5284);
  or csa_tree_add_190_195_groupi_g42607(csa_tree_add_190_195_groupi_n_6470 ,csa_tree_add_190_195_groupi_n_5060 ,csa_tree_add_190_195_groupi_n_5909);
  nor csa_tree_add_190_195_groupi_g42608(csa_tree_add_190_195_groupi_n_6469 ,csa_tree_add_190_195_groupi_n_4927 ,csa_tree_add_190_195_groupi_n_5912);
  and csa_tree_add_190_195_groupi_g42609(csa_tree_add_190_195_groupi_n_6468 ,csa_tree_add_190_195_groupi_n_2870 ,csa_tree_add_190_195_groupi_n_5972);
  nor csa_tree_add_190_195_groupi_g42610(csa_tree_add_190_195_groupi_n_6467 ,csa_tree_add_190_195_groupi_n_4918 ,csa_tree_add_190_195_groupi_n_5949);
  and csa_tree_add_190_195_groupi_g42611(csa_tree_add_190_195_groupi_n_6466 ,csa_tree_add_190_195_groupi_n_5266 ,csa_tree_add_190_195_groupi_n_5311);
  or csa_tree_add_190_195_groupi_g42612(csa_tree_add_190_195_groupi_n_6465 ,csa_tree_add_190_195_groupi_n_5369 ,csa_tree_add_190_195_groupi_n_5901);
  nor csa_tree_add_190_195_groupi_g42613(csa_tree_add_190_195_groupi_n_6464 ,csa_tree_add_190_195_groupi_n_4133 ,csa_tree_add_190_195_groupi_n_5905);
  nor csa_tree_add_190_195_groupi_g42614(csa_tree_add_190_195_groupi_n_6463 ,csa_tree_add_190_195_groupi_n_5368 ,csa_tree_add_190_195_groupi_n_5902);
  or csa_tree_add_190_195_groupi_g42615(csa_tree_add_190_195_groupi_n_6462 ,csa_tree_add_190_195_groupi_n_5898 ,csa_tree_add_190_195_groupi_n_5310);
  or csa_tree_add_190_195_groupi_g42616(csa_tree_add_190_195_groupi_n_6461 ,csa_tree_add_190_195_groupi_n_4708 ,csa_tree_add_190_195_groupi_n_5207);
  or csa_tree_add_190_195_groupi_g42617(csa_tree_add_190_195_groupi_n_6460 ,csa_tree_add_190_195_groupi_n_4787 ,csa_tree_add_190_195_groupi_n_5375);
  or csa_tree_add_190_195_groupi_g42618(csa_tree_add_190_195_groupi_n_6459 ,csa_tree_add_190_195_groupi_n_4618 ,csa_tree_add_190_195_groupi_n_5402);
  or csa_tree_add_190_195_groupi_g42620(csa_tree_add_190_195_groupi_n_6458 ,csa_tree_add_190_195_groupi_n_4134 ,csa_tree_add_190_195_groupi_n_5904);
  and csa_tree_add_190_195_groupi_g42621(csa_tree_add_190_195_groupi_n_6457 ,csa_tree_add_190_195_groupi_n_5298 ,csa_tree_add_190_195_groupi_n_5396);
  nor csa_tree_add_190_195_groupi_g42622(csa_tree_add_190_195_groupi_n_6456 ,csa_tree_add_190_195_groupi_n_5059 ,csa_tree_add_190_195_groupi_n_5910);
  nor csa_tree_add_190_195_groupi_g42623(csa_tree_add_190_195_groupi_n_6455 ,csa_tree_add_190_195_groupi_n_5899 ,csa_tree_add_190_195_groupi_n_5309);
  and csa_tree_add_190_195_groupi_g42624(csa_tree_add_190_195_groupi_n_6454 ,csa_tree_add_190_195_groupi_n_3665 ,csa_tree_add_190_195_groupi_n_5980);
  and csa_tree_add_190_195_groupi_g42625(csa_tree_add_190_195_groupi_n_6453 ,csa_tree_add_190_195_groupi_n_4812 ,csa_tree_add_190_195_groupi_n_5693);
  or csa_tree_add_190_195_groupi_g42626(csa_tree_add_190_195_groupi_n_6452 ,csa_tree_add_190_195_groupi_n_5023 ,csa_tree_add_190_195_groupi_n_5360);
  nor csa_tree_add_190_195_groupi_g42627(csa_tree_add_190_195_groupi_n_6451 ,csa_tree_add_190_195_groupi_n_54 ,csa_tree_add_190_195_groupi_n_5896);
  nor csa_tree_add_190_195_groupi_g42628(csa_tree_add_190_195_groupi_n_6450 ,csa_tree_add_190_195_groupi_n_4900 ,csa_tree_add_190_195_groupi_n_5456);
  nor csa_tree_add_190_195_groupi_g42629(csa_tree_add_190_195_groupi_n_6449 ,csa_tree_add_190_195_groupi_n_5024 ,csa_tree_add_190_195_groupi_n_5359);
  nor csa_tree_add_190_195_groupi_g42630(csa_tree_add_190_195_groupi_n_6448 ,csa_tree_add_190_195_groupi_n_5274 ,csa_tree_add_190_195_groupi_n_5343);
  or csa_tree_add_190_195_groupi_g42631(csa_tree_add_190_195_groupi_n_6447 ,csa_tree_add_190_195_groupi_n_4901 ,csa_tree_add_190_195_groupi_n_5455);
  or csa_tree_add_190_195_groupi_g42632(csa_tree_add_190_195_groupi_n_6446 ,csa_tree_add_190_195_groupi_n_5884 ,csa_tree_add_190_195_groupi_n_5878);
  nor csa_tree_add_190_195_groupi_g42633(csa_tree_add_190_195_groupi_n_6445 ,csa_tree_add_190_195_groupi_n_4966 ,csa_tree_add_190_195_groupi_n_5215);
  nor csa_tree_add_190_195_groupi_g42634(csa_tree_add_190_195_groupi_n_6444 ,csa_tree_add_190_195_groupi_n_4570 ,csa_tree_add_190_195_groupi_n_5514);
  nor csa_tree_add_190_195_groupi_g42635(csa_tree_add_190_195_groupi_n_6443 ,csa_tree_add_190_195_groupi_n_5886 ,csa_tree_add_190_195_groupi_n_5362);
  or csa_tree_add_190_195_groupi_g42636(csa_tree_add_190_195_groupi_n_6442 ,csa_tree_add_190_195_groupi_n_4828 ,csa_tree_add_190_195_groupi_n_5696);
  or csa_tree_add_190_195_groupi_g42637(csa_tree_add_190_195_groupi_n_6441 ,csa_tree_add_190_195_groupi_n_5273 ,csa_tree_add_190_195_groupi_n_5344);
  nor csa_tree_add_190_195_groupi_g42638(csa_tree_add_190_195_groupi_n_6440 ,csa_tree_add_190_195_groupi_n_5337 ,csa_tree_add_190_195_groupi_n_5364);
  and csa_tree_add_190_195_groupi_g42639(csa_tree_add_190_195_groupi_n_6439 ,csa_tree_add_190_195_groupi_n_5442 ,csa_tree_add_190_195_groupi_n_5414);
  or csa_tree_add_190_195_groupi_g42640(csa_tree_add_190_195_groupi_n_6438 ,csa_tree_add_190_195_groupi_n_9 ,csa_tree_add_190_195_groupi_n_5889);
  and csa_tree_add_190_195_groupi_g42641(csa_tree_add_190_195_groupi_n_6437 ,csa_tree_add_190_195_groupi_n_29 ,csa_tree_add_190_195_groupi_n_5312);
  nor csa_tree_add_190_195_groupi_g42642(csa_tree_add_190_195_groupi_n_6436 ,csa_tree_add_190_195_groupi_n_5358 ,csa_tree_add_190_195_groupi_n_5882);
  or csa_tree_add_190_195_groupi_g42643(csa_tree_add_190_195_groupi_n_6435 ,csa_tree_add_190_195_groupi_n_5357 ,csa_tree_add_190_195_groupi_n_5883);
  or csa_tree_add_190_195_groupi_g42644(csa_tree_add_190_195_groupi_n_6434 ,csa_tree_add_190_195_groupi_n_5356 ,csa_tree_add_190_195_groupi_n_5367);
  or csa_tree_add_190_195_groupi_g42645(csa_tree_add_190_195_groupi_n_6433 ,csa_tree_add_190_195_groupi_n_5887 ,csa_tree_add_190_195_groupi_n_5361);
  or csa_tree_add_190_195_groupi_g42646(csa_tree_add_190_195_groupi_n_6432 ,csa_tree_add_190_195_groupi_n_1362 ,csa_tree_add_190_195_groupi_n_5204);
  nor csa_tree_add_190_195_groupi_g42647(csa_tree_add_190_195_groupi_n_6431 ,csa_tree_add_190_195_groupi_n_5080 ,csa_tree_add_190_195_groupi_n_5903);
  and csa_tree_add_190_195_groupi_g42648(csa_tree_add_190_195_groupi_n_6430 ,csa_tree_add_190_195_groupi_n_3575 ,csa_tree_add_190_195_groupi_n_5594);
  and csa_tree_add_190_195_groupi_g42649(csa_tree_add_190_195_groupi_n_6429 ,csa_tree_add_190_195_groupi_n_4756 ,csa_tree_add_190_195_groupi_n_5239);
  nor csa_tree_add_190_195_groupi_g42650(csa_tree_add_190_195_groupi_n_6428 ,csa_tree_add_190_195_groupi_n_5353 ,csa_tree_add_190_195_groupi_n_5352);
  or csa_tree_add_190_195_groupi_g42651(csa_tree_add_190_195_groupi_n_6427 ,csa_tree_add_190_195_groupi_n_5377 ,csa_tree_add_190_195_groupi_n_5372);
  and csa_tree_add_190_195_groupi_g42652(csa_tree_add_190_195_groupi_n_6426 ,csa_tree_add_190_195_groupi_n_5353 ,csa_tree_add_190_195_groupi_n_5352);
  and csa_tree_add_190_195_groupi_g42653(csa_tree_add_190_195_groupi_n_6425 ,csa_tree_add_190_195_groupi_n_5961 ,csa_tree_add_190_195_groupi_n_5876);
  and csa_tree_add_190_195_groupi_g42654(csa_tree_add_190_195_groupi_n_6424 ,csa_tree_add_190_195_groupi_n_5356 ,csa_tree_add_190_195_groupi_n_5367);
  or csa_tree_add_190_195_groupi_g42655(csa_tree_add_190_195_groupi_n_6423 ,csa_tree_add_190_195_groupi_n_4987 ,csa_tree_add_190_195_groupi_n_5256);
  or csa_tree_add_190_195_groupi_g42656(csa_tree_add_190_195_groupi_n_6422 ,csa_tree_add_190_195_groupi_n_5350 ,csa_tree_add_190_195_groupi_n_5348);
  and csa_tree_add_190_195_groupi_g42657(csa_tree_add_190_195_groupi_n_6421 ,csa_tree_add_190_195_groupi_n_5395 ,csa_tree_add_190_195_groupi_n_5349);
  or csa_tree_add_190_195_groupi_g42658(csa_tree_add_190_195_groupi_n_6420 ,csa_tree_add_190_195_groupi_n_5412 ,csa_tree_add_190_195_groupi_n_5405);
  nor csa_tree_add_190_195_groupi_g42659(csa_tree_add_190_195_groupi_n_6419 ,csa_tree_add_190_195_groupi_n_5880 ,csa_tree_add_190_195_groupi_n_5347);
  and csa_tree_add_190_195_groupi_g42660(csa_tree_add_190_195_groupi_n_6418 ,csa_tree_add_190_195_groupi_n_5350 ,csa_tree_add_190_195_groupi_n_5348);
  or csa_tree_add_190_195_groupi_g42661(csa_tree_add_190_195_groupi_n_6417 ,csa_tree_add_190_195_groupi_n_80 ,csa_tree_add_190_195_groupi_n_5345);
  and csa_tree_add_190_195_groupi_g42662(csa_tree_add_190_195_groupi_n_6416 ,csa_tree_add_190_195_groupi_n_4987 ,csa_tree_add_190_195_groupi_n_5256);
  and csa_tree_add_190_195_groupi_g42663(csa_tree_add_190_195_groupi_n_6415 ,csa_tree_add_190_195_groupi_n_5102 ,csa_tree_add_190_195_groupi_n_5768);
  nor csa_tree_add_190_195_groupi_g42664(csa_tree_add_190_195_groupi_n_6414 ,csa_tree_add_190_195_groupi_n_2834 ,csa_tree_add_190_195_groupi_n_5576);
  and csa_tree_add_190_195_groupi_g42665(csa_tree_add_190_195_groupi_n_6413 ,csa_tree_add_190_195_groupi_n_80 ,csa_tree_add_190_195_groupi_n_5345);
  or csa_tree_add_190_195_groupi_g42666(csa_tree_add_190_195_groupi_n_6412 ,csa_tree_add_190_195_groupi_n_4695 ,csa_tree_add_190_195_groupi_n_5498);
  and csa_tree_add_190_195_groupi_g42667(csa_tree_add_190_195_groupi_n_6411 ,csa_tree_add_190_195_groupi_n_4979 ,csa_tree_add_190_195_groupi_n_11);
  nor csa_tree_add_190_195_groupi_g42668(csa_tree_add_190_195_groupi_n_6410 ,csa_tree_add_190_195_groupi_n_4114 ,csa_tree_add_190_195_groupi_n_5212);
  nor csa_tree_add_190_195_groupi_g42669(csa_tree_add_190_195_groupi_n_6409 ,csa_tree_add_190_195_groupi_n_5342 ,csa_tree_add_190_195_groupi_n_5871);
  and csa_tree_add_190_195_groupi_g42670(csa_tree_add_190_195_groupi_n_6408 ,csa_tree_add_190_195_groupi_n_5873 ,csa_tree_add_190_195_groupi_n_5415);
  or csa_tree_add_190_195_groupi_g42671(csa_tree_add_190_195_groupi_n_6407 ,csa_tree_add_190_195_groupi_n_4959 ,csa_tree_add_190_195_groupi_n_5906);
  nor csa_tree_add_190_195_groupi_g42672(csa_tree_add_190_195_groupi_n_6406 ,csa_tree_add_190_195_groupi_n_4979 ,csa_tree_add_190_195_groupi_n_11);
  nor csa_tree_add_190_195_groupi_g42673(csa_tree_add_190_195_groupi_n_6405 ,csa_tree_add_190_195_groupi_n_4705 ,csa_tree_add_190_195_groupi_n_5875);
  or csa_tree_add_190_195_groupi_g42674(csa_tree_add_190_195_groupi_n_6404 ,csa_tree_add_190_195_groupi_n_5762 ,csa_tree_add_190_195_groupi_n_5974);
  nor csa_tree_add_190_195_groupi_g42675(csa_tree_add_190_195_groupi_n_6403 ,csa_tree_add_190_195_groupi_n_4686 ,csa_tree_add_190_195_groupi_n_5292);
  and csa_tree_add_190_195_groupi_g42676(csa_tree_add_190_195_groupi_n_6402 ,csa_tree_add_190_195_groupi_n_4705 ,csa_tree_add_190_195_groupi_n_5875);
  nor csa_tree_add_190_195_groupi_g42677(csa_tree_add_190_195_groupi_n_6401 ,csa_tree_add_190_195_groupi_n_5481 ,csa_tree_add_190_195_groupi_n_5340);
  and csa_tree_add_190_195_groupi_g42678(csa_tree_add_190_195_groupi_n_6400 ,csa_tree_add_190_195_groupi_n_3646 ,csa_tree_add_190_195_groupi_n_5575);
  or csa_tree_add_190_195_groupi_g42679(csa_tree_add_190_195_groupi_n_6399 ,csa_tree_add_190_195_groupi_n_5482 ,csa_tree_add_190_195_groupi_n_5339);
  or csa_tree_add_190_195_groupi_g42680(csa_tree_add_190_195_groupi_n_6398 ,csa_tree_add_190_195_groupi_n_5351 ,csa_tree_add_190_195_groupi_n_5495);
  or csa_tree_add_190_195_groupi_g42681(csa_tree_add_190_195_groupi_n_6397 ,csa_tree_add_190_195_groupi_n_5443 ,csa_tree_add_190_195_groupi_n_5336);
  or csa_tree_add_190_195_groupi_g42682(csa_tree_add_190_195_groupi_n_6396 ,csa_tree_add_190_195_groupi_n_5341 ,csa_tree_add_190_195_groupi_n_5872);
  nor csa_tree_add_190_195_groupi_g42683(csa_tree_add_190_195_groupi_n_6395 ,csa_tree_add_190_195_groupi_n_5873 ,csa_tree_add_190_195_groupi_n_5415);
  or csa_tree_add_190_195_groupi_g42684(csa_tree_add_190_195_groupi_n_6394 ,csa_tree_add_190_195_groupi_n_5543 ,csa_tree_add_190_195_groupi_n_5308);
  nor csa_tree_add_190_195_groupi_g42685(csa_tree_add_190_195_groupi_n_6393 ,csa_tree_add_190_195_groupi_n_5381 ,csa_tree_add_190_195_groupi_n_75);
  or csa_tree_add_190_195_groupi_g42686(csa_tree_add_190_195_groupi_n_6392 ,csa_tree_add_190_195_groupi_n_4784 ,csa_tree_add_190_195_groupi_n_5289);
  or csa_tree_add_190_195_groupi_g42687(csa_tree_add_190_195_groupi_n_6391 ,csa_tree_add_190_195_groupi_n_5142 ,csa_tree_add_190_195_groupi_n_5753);
  or csa_tree_add_190_195_groupi_g42688(csa_tree_add_190_195_groupi_n_6390 ,csa_tree_add_190_195_groupi_n_5143 ,csa_tree_add_190_195_groupi_n_5751);
  nor csa_tree_add_190_195_groupi_g42689(csa_tree_add_190_195_groupi_n_6389 ,csa_tree_add_190_195_groupi_n_4756 ,csa_tree_add_190_195_groupi_n_5239);
  nor csa_tree_add_190_195_groupi_g42690(csa_tree_add_190_195_groupi_n_6388 ,csa_tree_add_190_195_groupi_n_5036 ,csa_tree_add_190_195_groupi_n_5220);
  or csa_tree_add_190_195_groupi_g42691(csa_tree_add_190_195_groupi_n_6387 ,csa_tree_add_190_195_groupi_n_5229 ,csa_tree_add_190_195_groupi_n_5230);
  or csa_tree_add_190_195_groupi_g42692(csa_tree_add_190_195_groupi_n_6386 ,csa_tree_add_190_195_groupi_n_4662 ,csa_tree_add_190_195_groupi_n_5240);
  or csa_tree_add_190_195_groupi_g42693(csa_tree_add_190_195_groupi_n_6385 ,csa_tree_add_190_195_groupi_n_5184 ,csa_tree_add_190_195_groupi_n_5295);
  or csa_tree_add_190_195_groupi_g42694(csa_tree_add_190_195_groupi_n_6384 ,csa_tree_add_190_195_groupi_n_1386 ,csa_tree_add_190_195_groupi_n_5919);
  and csa_tree_add_190_195_groupi_g42695(csa_tree_add_190_195_groupi_n_6383 ,csa_tree_add_190_195_groupi_n_4686 ,csa_tree_add_190_195_groupi_n_5292);
  or csa_tree_add_190_195_groupi_g42696(csa_tree_add_190_195_groupi_n_6382 ,csa_tree_add_190_195_groupi_n_5335 ,csa_tree_add_190_195_groupi_n_5934);
  or csa_tree_add_190_195_groupi_g42697(csa_tree_add_190_195_groupi_n_6381 ,csa_tree_add_190_195_groupi_n_5442 ,csa_tree_add_190_195_groupi_n_5414);
  or csa_tree_add_190_195_groupi_g42698(csa_tree_add_190_195_groupi_n_6380 ,csa_tree_add_190_195_groupi_n_4904 ,csa_tree_add_190_195_groupi_n_5892);
  nor csa_tree_add_190_195_groupi_g42699(csa_tree_add_190_195_groupi_n_6379 ,csa_tree_add_190_195_groupi_n_5410 ,csa_tree_add_190_195_groupi_n_5300);
  nor csa_tree_add_190_195_groupi_g42700(csa_tree_add_190_195_groupi_n_6378 ,csa_tree_add_190_195_groupi_n_4991 ,csa_tree_add_190_195_groupi_n_5285);
  and csa_tree_add_190_195_groupi_g42701(csa_tree_add_190_195_groupi_n_6377 ,csa_tree_add_190_195_groupi_n_3562 ,csa_tree_add_190_195_groupi_n_5611);
  or csa_tree_add_190_195_groupi_g42702(csa_tree_add_190_195_groupi_n_6376 ,csa_tree_add_190_195_groupi_n_4922 ,csa_tree_add_190_195_groupi_n_5921);
  or csa_tree_add_190_195_groupi_g42703(csa_tree_add_190_195_groupi_n_6375 ,csa_tree_add_190_195_groupi_n_5149 ,csa_tree_add_190_195_groupi_n_5743);
  nor csa_tree_add_190_195_groupi_g42704(csa_tree_add_190_195_groupi_n_6374 ,csa_tree_add_190_195_groupi_n_5961 ,csa_tree_add_190_195_groupi_n_5876);
  and csa_tree_add_190_195_groupi_g42705(csa_tree_add_190_195_groupi_n_6373 ,csa_tree_add_190_195_groupi_n_5464 ,csa_tree_add_190_195_groupi_n_5509);
  nor csa_tree_add_190_195_groupi_g42706(csa_tree_add_190_195_groupi_n_6372 ,csa_tree_add_190_195_groupi_n_4921 ,csa_tree_add_190_195_groupi_n_5922);
  nor csa_tree_add_190_195_groupi_g42707(csa_tree_add_190_195_groupi_n_6371 ,csa_tree_add_190_195_groupi_n_5464 ,csa_tree_add_190_195_groupi_n_5509);
  nor csa_tree_add_190_195_groupi_g42708(csa_tree_add_190_195_groupi_n_6370 ,csa_tree_add_190_195_groupi_n_5529 ,csa_tree_add_190_195_groupi_n_5325);
  or csa_tree_add_190_195_groupi_g42709(csa_tree_add_190_195_groupi_n_6369 ,csa_tree_add_190_195_groupi_n_5530 ,csa_tree_add_190_195_groupi_n_5324);
  and csa_tree_add_190_195_groupi_g42710(csa_tree_add_190_195_groupi_n_6368 ,csa_tree_add_190_195_groupi_n_4628 ,csa_tree_add_190_195_groupi_n_5323);
  and csa_tree_add_190_195_groupi_g42711(csa_tree_add_190_195_groupi_n_6367 ,csa_tree_add_190_195_groupi_n_4869 ,csa_tree_add_190_195_groupi_n_5629);
  or csa_tree_add_190_195_groupi_g42712(csa_tree_add_190_195_groupi_n_6366 ,csa_tree_add_190_195_groupi_n_4898 ,csa_tree_add_190_195_groupi_n_5429);
  or csa_tree_add_190_195_groupi_g42713(csa_tree_add_190_195_groupi_n_6365 ,csa_tree_add_190_195_groupi_n_4569 ,csa_tree_add_190_195_groupi_n_5468);
  or csa_tree_add_190_195_groupi_g42714(csa_tree_add_190_195_groupi_n_6364 ,csa_tree_add_190_195_groupi_n_4892 ,csa_tree_add_190_195_groupi_n_5485);
  nor csa_tree_add_190_195_groupi_g42715(csa_tree_add_190_195_groupi_n_6363 ,csa_tree_add_190_195_groupi_n_5099 ,csa_tree_add_190_195_groupi_n_5733);
  nor csa_tree_add_190_195_groupi_g42716(csa_tree_add_190_195_groupi_n_6362 ,csa_tree_add_190_195_groupi_n_954 ,csa_tree_add_190_195_groupi_n_5205);
  nor csa_tree_add_190_195_groupi_g42717(csa_tree_add_190_195_groupi_n_6361 ,csa_tree_add_190_195_groupi_n_4919 ,csa_tree_add_190_195_groupi_n_5183);
  or csa_tree_add_190_195_groupi_g42718(csa_tree_add_190_195_groupi_n_6360 ,csa_tree_add_190_195_groupi_n_688 ,csa_tree_add_190_195_groupi_n_5319);
  nor csa_tree_add_190_195_groupi_g42719(csa_tree_add_190_195_groupi_n_6359 ,csa_tree_add_190_195_groupi_n_378 ,csa_tree_add_190_195_groupi_n_5320);
  or csa_tree_add_190_195_groupi_g42720(csa_tree_add_190_195_groupi_n_6358 ,csa_tree_add_190_195_groupi_n_4126 ,csa_tree_add_190_195_groupi_n_5522);
  and csa_tree_add_190_195_groupi_g42721(csa_tree_add_190_195_groupi_n_6357 ,csa_tree_add_190_195_groupi_n_6 ,csa_tree_add_190_195_groupi_n_76);
  and csa_tree_add_190_195_groupi_g42722(csa_tree_add_190_195_groupi_n_6356 ,csa_tree_add_190_195_groupi_n_1188 ,csa_tree_add_190_195_groupi_n_5504);
  and csa_tree_add_190_195_groupi_g42723(csa_tree_add_190_195_groupi_n_6355 ,csa_tree_add_190_195_groupi_n_4787 ,csa_tree_add_190_195_groupi_n_5375);
  or csa_tree_add_190_195_groupi_g42724(csa_tree_add_190_195_groupi_n_6354 ,csa_tree_add_190_195_groupi_n_5139 ,csa_tree_add_190_195_groupi_n_5737);
  nor csa_tree_add_190_195_groupi_g42725(csa_tree_add_190_195_groupi_n_6353 ,csa_tree_add_190_195_groupi_n_5479 ,csa_tree_add_190_195_groupi_n_5318);
  or csa_tree_add_190_195_groupi_g42726(csa_tree_add_190_195_groupi_n_6352 ,csa_tree_add_190_195_groupi_n_5107 ,csa_tree_add_190_195_groupi_n_5853);
  or csa_tree_add_190_195_groupi_g42727(csa_tree_add_190_195_groupi_n_6351 ,csa_tree_add_190_195_groupi_n_5480 ,csa_tree_add_190_195_groupi_n_5317);
  nor csa_tree_add_190_195_groupi_g42728(csa_tree_add_190_195_groupi_n_6350 ,csa_tree_add_190_195_groupi_n_4852 ,csa_tree_add_190_195_groupi_n_5861);
  nor csa_tree_add_190_195_groupi_g42729(csa_tree_add_190_195_groupi_n_6349 ,csa_tree_add_190_195_groupi_n_1311 ,csa_tree_add_190_195_groupi_n_5430);
  or csa_tree_add_190_195_groupi_g42730(csa_tree_add_190_195_groupi_n_6348 ,csa_tree_add_190_195_groupi_n_5472 ,csa_tree_add_190_195_groupi_n_5316);
  nor csa_tree_add_190_195_groupi_g42731(csa_tree_add_190_195_groupi_n_6347 ,csa_tree_add_190_195_groupi_n_5947 ,csa_tree_add_190_195_groupi_n_5277);
  and csa_tree_add_190_195_groupi_g42732(csa_tree_add_190_195_groupi_n_6346 ,csa_tree_add_190_195_groupi_n_5888 ,csa_tree_add_190_195_groupi_n_5542);
  nor csa_tree_add_190_195_groupi_g42733(csa_tree_add_190_195_groupi_n_6345 ,csa_tree_add_190_195_groupi_n_4565 ,csa_tree_add_190_195_groupi_n_5448);
  nor csa_tree_add_190_195_groupi_g42734(csa_tree_add_190_195_groupi_n_6344 ,csa_tree_add_190_195_groupi_n_4696 ,csa_tree_add_190_195_groupi_n_5499);
  and csa_tree_add_190_195_groupi_g42735(csa_tree_add_190_195_groupi_n_6343 ,csa_tree_add_190_195_groupi_n_5134 ,csa_tree_add_190_195_groupi_n_5836);
  nor csa_tree_add_190_195_groupi_g42736(csa_tree_add_190_195_groupi_n_6342 ,csa_tree_add_190_195_groupi_n_5437 ,csa_tree_add_190_195_groupi_n_5223);
  and csa_tree_add_190_195_groupi_g42737(csa_tree_add_190_195_groupi_n_6341 ,csa_tree_add_190_195_groupi_n_5168 ,csa_tree_add_190_195_groupi_n_5724);
  or csa_tree_add_190_195_groupi_g42738(csa_tree_add_190_195_groupi_n_6340 ,csa_tree_add_190_195_groupi_n_5438 ,csa_tree_add_190_195_groupi_n_5222);
  nor csa_tree_add_190_195_groupi_g42739(csa_tree_add_190_195_groupi_n_6339 ,csa_tree_add_190_195_groupi_n_5424 ,csa_tree_add_190_195_groupi_n_10);
  or csa_tree_add_190_195_groupi_g42740(csa_tree_add_190_195_groupi_n_6338 ,csa_tree_add_190_195_groupi_n_2399 ,csa_tree_add_190_195_groupi_n_5269);
  or csa_tree_add_190_195_groupi_g42741(csa_tree_add_190_195_groupi_n_6337 ,csa_tree_add_190_195_groupi_n_5425 ,csa_tree_add_190_195_groupi_n_5305);
  and csa_tree_add_190_195_groupi_g42742(csa_tree_add_190_195_groupi_n_6336 ,csa_tree_add_190_195_groupi_n_4833 ,csa_tree_add_190_195_groupi_n_5722);
  or csa_tree_add_190_195_groupi_g42744(csa_tree_add_190_195_groupi_n_6335 ,csa_tree_add_190_195_groupi_n_5021 ,csa_tree_add_190_195_groupi_n_5232);
  and csa_tree_add_190_195_groupi_g42745(csa_tree_add_190_195_groupi_n_6334 ,csa_tree_add_190_195_groupi_n_4580 ,csa_tree_add_190_195_groupi_n_5561);
  or csa_tree_add_190_195_groupi_g42746(csa_tree_add_190_195_groupi_n_6333 ,csa_tree_add_190_195_groupi_n_5119 ,csa_tree_add_190_195_groupi_n_5700);
  or csa_tree_add_190_195_groupi_g42747(csa_tree_add_190_195_groupi_n_6332 ,csa_tree_add_190_195_groupi_n_5338 ,csa_tree_add_190_195_groupi_n_5363);
  or csa_tree_add_190_195_groupi_g42749(csa_tree_add_190_195_groupi_n_6331 ,csa_tree_add_190_195_groupi_n_4564 ,csa_tree_add_190_195_groupi_n_5449);
  or csa_tree_add_190_195_groupi_g42750(csa_tree_add_190_195_groupi_n_6330 ,csa_tree_add_190_195_groupi_n_5908 ,csa_tree_add_190_195_groupi_n_5929);
  and csa_tree_add_190_195_groupi_g42751(csa_tree_add_190_195_groupi_n_6329 ,csa_tree_add_190_195_groupi_n_4892 ,csa_tree_add_190_195_groupi_n_5485);
  nor csa_tree_add_190_195_groupi_g42752(csa_tree_add_190_195_groupi_n_6328 ,csa_tree_add_190_195_groupi_n_81 ,csa_tree_add_190_195_groupi_n_5406);
  nor csa_tree_add_190_195_groupi_g42753(csa_tree_add_190_195_groupi_n_6327 ,csa_tree_add_190_195_groupi_n_4813 ,csa_tree_add_190_195_groupi_n_5720);
  nor csa_tree_add_190_195_groupi_g42754(csa_tree_add_190_195_groupi_n_6326 ,csa_tree_add_190_195_groupi_n_5298 ,csa_tree_add_190_195_groupi_n_5396);
  and csa_tree_add_190_195_groupi_g42755(csa_tree_add_190_195_groupi_n_6325 ,csa_tree_add_190_195_groupi_n_5217 ,csa_tree_add_190_195_groupi_n_5302);
  or csa_tree_add_190_195_groupi_g42756(csa_tree_add_190_195_groupi_n_6324 ,csa_tree_add_190_195_groupi_n_2396 ,csa_tree_add_190_195_groupi_n_5322);
  or csa_tree_add_190_195_groupi_g42757(csa_tree_add_190_195_groupi_n_6323 ,csa_tree_add_190_195_groupi_n_2395 ,csa_tree_add_190_195_groupi_n_5237);
  nor csa_tree_add_190_195_groupi_g42758(csa_tree_add_190_195_groupi_n_6322 ,csa_tree_add_190_195_groupi_n_4980 ,csa_tree_add_190_195_groupi_n_5391);
  or csa_tree_add_190_195_groupi_g42759(csa_tree_add_190_195_groupi_n_6321 ,csa_tree_add_190_195_groupi_n_6 ,csa_tree_add_190_195_groupi_n_76);
  or csa_tree_add_190_195_groupi_g42760(csa_tree_add_190_195_groupi_n_6320 ,csa_tree_add_190_195_groupi_n_3712 ,csa_tree_add_190_195_groupi_n_5577);
  and csa_tree_add_190_195_groupi_g42761(csa_tree_add_190_195_groupi_n_6319 ,csa_tree_add_190_195_groupi_n_554 ,csa_tree_add_190_195_groupi_n_5241);
  or csa_tree_add_190_195_groupi_g42763(csa_tree_add_190_195_groupi_n_6318 ,csa_tree_add_190_195_groupi_n_4866 ,csa_tree_add_190_195_groupi_n_5677);
  or csa_tree_add_190_195_groupi_g42764(csa_tree_add_190_195_groupi_n_6317 ,csa_tree_add_190_195_groupi_n_5263 ,csa_tree_add_190_195_groupi_n_5297);
  or csa_tree_add_190_195_groupi_g42765(csa_tree_add_190_195_groupi_n_6316 ,csa_tree_add_190_195_groupi_n_4841 ,csa_tree_add_190_195_groupi_n_5660);
  nor csa_tree_add_190_195_groupi_g42766(csa_tree_add_190_195_groupi_n_6315 ,csa_tree_add_190_195_groupi_n_4752 ,csa_tree_add_190_195_groupi_n_5246);
  or csa_tree_add_190_195_groupi_g42767(csa_tree_add_190_195_groupi_n_6314 ,csa_tree_add_190_195_groupi_n_4620 ,csa_tree_add_190_195_groupi_n_5294);
  nor csa_tree_add_190_195_groupi_g42768(csa_tree_add_190_195_groupi_n_6313 ,csa_tree_add_190_195_groupi_n_4621 ,csa_tree_add_190_195_groupi_n_5293);
  nor csa_tree_add_190_195_groupi_g42769(csa_tree_add_190_195_groupi_n_6312 ,csa_tree_add_190_195_groupi_n_5383 ,csa_tree_add_190_195_groupi_n_5291);
  nor csa_tree_add_190_195_groupi_g42770(csa_tree_add_190_195_groupi_n_6311 ,csa_tree_add_190_195_groupi_n_32 ,csa_tree_add_190_195_groupi_n_5306);
  or csa_tree_add_190_195_groupi_g42771(csa_tree_add_190_195_groupi_n_6310 ,csa_tree_add_190_195_groupi_n_5384 ,csa_tree_add_190_195_groupi_n_5290);
  or csa_tree_add_190_195_groupi_g42772(csa_tree_add_190_195_groupi_n_6309 ,csa_tree_add_190_195_groupi_n_3651 ,csa_tree_add_190_195_groupi_n_5971);
  nor csa_tree_add_190_195_groupi_g42773(csa_tree_add_190_195_groupi_n_6308 ,csa_tree_add_190_195_groupi_n_5378 ,csa_tree_add_190_195_groupi_n_5373);
  nor csa_tree_add_190_195_groupi_g42774(csa_tree_add_190_195_groupi_n_6307 ,csa_tree_add_190_195_groupi_n_5395 ,csa_tree_add_190_195_groupi_n_5349);
  or csa_tree_add_190_195_groupi_g42775(csa_tree_add_190_195_groupi_n_6306 ,csa_tree_add_190_195_groupi_n_5101 ,csa_tree_add_190_195_groupi_n_5851);
  nor csa_tree_add_190_195_groupi_g42776(csa_tree_add_190_195_groupi_n_6305 ,csa_tree_add_190_195_groupi_n_5185 ,csa_tree_add_190_195_groupi_n_5296);
  nor csa_tree_add_190_195_groupi_g42777(csa_tree_add_190_195_groupi_n_6304 ,csa_tree_add_190_195_groupi_n_5279 ,csa_tree_add_190_195_groupi_n_5959);
  and csa_tree_add_190_195_groupi_g42778(csa_tree_add_190_195_groupi_n_6303 ,csa_tree_add_190_195_groupi_n_9 ,csa_tree_add_190_195_groupi_n_5889);
  nor csa_tree_add_190_195_groupi_g42779(csa_tree_add_190_195_groupi_n_6302 ,csa_tree_add_190_195_groupi_n_5022 ,csa_tree_add_190_195_groupi_n_5231);
  and csa_tree_add_190_195_groupi_g42780(csa_tree_add_190_195_groupi_n_6301 ,csa_tree_add_190_195_groupi_n_5097 ,csa_tree_add_190_195_groupi_n_5712);
  nor csa_tree_add_190_195_groupi_g42781(csa_tree_add_190_195_groupi_n_6300 ,csa_tree_add_190_195_groupi_n_5094 ,csa_tree_add_190_195_groupi_n_5956);
  or csa_tree_add_190_195_groupi_g42782(csa_tree_add_190_195_groupi_n_6299 ,csa_tree_add_190_195_groupi_n_4706 ,csa_tree_add_190_195_groupi_n_5288);
  and csa_tree_add_190_195_groupi_g42783(csa_tree_add_190_195_groupi_n_6298 ,csa_tree_add_190_195_groupi_n_483 ,csa_tree_add_190_195_groupi_n_5513);
  nor csa_tree_add_190_195_groupi_g42784(csa_tree_add_190_195_groupi_n_6297 ,csa_tree_add_190_195_groupi_n_5115 ,csa_tree_add_190_195_groupi_n_5708);
  or csa_tree_add_190_195_groupi_g42785(csa_tree_add_190_195_groupi_n_6296 ,csa_tree_add_190_195_groupi_n_398 ,csa_tree_add_190_195_groupi_n_5513);
  or csa_tree_add_190_195_groupi_g42786(csa_tree_add_190_195_groupi_n_6295 ,csa_tree_add_190_195_groupi_n_4850 ,csa_tree_add_190_195_groupi_n_5686);
  nor csa_tree_add_190_195_groupi_g42787(csa_tree_add_190_195_groupi_n_6294 ,csa_tree_add_190_195_groupi_n_4566 ,csa_tree_add_190_195_groupi_n_5314);
  and csa_tree_add_190_195_groupi_g42788(csa_tree_add_190_195_groupi_n_6293 ,csa_tree_add_190_195_groupi_n_3436 ,csa_tree_add_190_195_groupi_n_5610);
  or csa_tree_add_190_195_groupi_g42789(csa_tree_add_190_195_groupi_n_6292 ,csa_tree_add_190_195_groupi_n_4857 ,csa_tree_add_190_195_groupi_n_5819);
  and csa_tree_add_190_195_groupi_g42790(csa_tree_add_190_195_groupi_n_6291 ,csa_tree_add_190_195_groupi_n_4566 ,csa_tree_add_190_195_groupi_n_5314);
  or csa_tree_add_190_195_groupi_g42791(csa_tree_add_190_195_groupi_n_6592 ,csa_tree_add_190_195_groupi_n_3601 ,csa_tree_add_190_195_groupi_n_5652);
  or csa_tree_add_190_195_groupi_g42792(csa_tree_add_190_195_groupi_n_6591 ,csa_tree_add_190_195_groupi_n_3369 ,csa_tree_add_190_195_groupi_n_5713);
  and csa_tree_add_190_195_groupi_g42793(csa_tree_add_190_195_groupi_n_6590 ,csa_tree_add_190_195_groupi_n_3160 ,csa_tree_add_190_195_groupi_n_5718);
  or csa_tree_add_190_195_groupi_g42794(csa_tree_add_190_195_groupi_n_6589 ,csa_tree_add_190_195_groupi_n_4324 ,csa_tree_add_190_195_groupi_n_5833);
  or csa_tree_add_190_195_groupi_g42795(csa_tree_add_190_195_groupi_n_6587 ,csa_tree_add_190_195_groupi_n_2986 ,csa_tree_add_190_195_groupi_n_5731);
  and csa_tree_add_190_195_groupi_g42796(csa_tree_add_190_195_groupi_n_6586 ,csa_tree_add_190_195_groupi_n_4244 ,csa_tree_add_190_195_groupi_n_5830);
  or csa_tree_add_190_195_groupi_g42797(csa_tree_add_190_195_groupi_n_6584 ,csa_tree_add_190_195_groupi_n_2972 ,csa_tree_add_190_195_groupi_n_5745);
  or csa_tree_add_190_195_groupi_g42798(csa_tree_add_190_195_groupi_n_6583 ,csa_tree_add_190_195_groupi_n_3189 ,csa_tree_add_190_195_groupi_n_5828);
  or csa_tree_add_190_195_groupi_g42799(csa_tree_add_190_195_groupi_n_6582 ,csa_tree_add_190_195_groupi_n_2946 ,csa_tree_add_190_195_groupi_n_5765);
  and csa_tree_add_190_195_groupi_g42800(csa_tree_add_190_195_groupi_n_6581 ,csa_tree_add_190_195_groupi_n_4394 ,csa_tree_add_190_195_groupi_n_5772);
  and csa_tree_add_190_195_groupi_g42801(csa_tree_add_190_195_groupi_n_6580 ,csa_tree_add_190_195_groupi_n_2916 ,csa_tree_add_190_195_groupi_n_5757);
  and csa_tree_add_190_195_groupi_g42802(csa_tree_add_190_195_groupi_n_6579 ,csa_tree_add_190_195_groupi_n_3550 ,csa_tree_add_190_195_groupi_n_5675);
  or csa_tree_add_190_195_groupi_g42803(csa_tree_add_190_195_groupi_n_6578 ,csa_tree_add_190_195_groupi_n_3339 ,csa_tree_add_190_195_groupi_n_5797);
  and csa_tree_add_190_195_groupi_g42804(csa_tree_add_190_195_groupi_n_6577 ,csa_tree_add_190_195_groupi_n_3425 ,csa_tree_add_190_195_groupi_n_5732);
  or csa_tree_add_190_195_groupi_g42805(csa_tree_add_190_195_groupi_n_6575 ,csa_tree_add_190_195_groupi_n_3309 ,csa_tree_add_190_195_groupi_n_5761);
  or csa_tree_add_190_195_groupi_g42806(csa_tree_add_190_195_groupi_n_6573 ,csa_tree_add_190_195_groupi_n_3637 ,csa_tree_add_190_195_groupi_n_5790);
  or csa_tree_add_190_195_groupi_g42807(csa_tree_add_190_195_groupi_n_6571 ,csa_tree_add_190_195_groupi_n_3251 ,csa_tree_add_190_195_groupi_n_5719);
  not csa_tree_add_190_195_groupi_g42808(csa_tree_add_190_195_groupi_n_6286 ,csa_tree_add_190_195_groupi_n_5);
  not csa_tree_add_190_195_groupi_g42809(csa_tree_add_190_195_groupi_n_6284 ,csa_tree_add_190_195_groupi_n_6283);
  not csa_tree_add_190_195_groupi_g42810(csa_tree_add_190_195_groupi_n_6279 ,csa_tree_add_190_195_groupi_n_85);
  not csa_tree_add_190_195_groupi_g42811(csa_tree_add_190_195_groupi_n_6277 ,csa_tree_add_190_195_groupi_n_6278);
  not csa_tree_add_190_195_groupi_g42812(csa_tree_add_190_195_groupi_n_6273 ,csa_tree_add_190_195_groupi_n_6274);
  not csa_tree_add_190_195_groupi_g42813(csa_tree_add_190_195_groupi_n_6271 ,csa_tree_add_190_195_groupi_n_6272);
  not csa_tree_add_190_195_groupi_g42814(csa_tree_add_190_195_groupi_n_6268 ,csa_tree_add_190_195_groupi_n_6269);
  not csa_tree_add_190_195_groupi_g42815(csa_tree_add_190_195_groupi_n_6263 ,csa_tree_add_190_195_groupi_n_6264);
  not csa_tree_add_190_195_groupi_g42816(csa_tree_add_190_195_groupi_n_6261 ,csa_tree_add_190_195_groupi_n_6262);
  not csa_tree_add_190_195_groupi_g42817(csa_tree_add_190_195_groupi_n_6258 ,csa_tree_add_190_195_groupi_n_6259);
  not csa_tree_add_190_195_groupi_g42818(csa_tree_add_190_195_groupi_n_6256 ,csa_tree_add_190_195_groupi_n_6257);
  not csa_tree_add_190_195_groupi_g42819(csa_tree_add_190_195_groupi_n_6254 ,csa_tree_add_190_195_groupi_n_6255);
  or csa_tree_add_190_195_groupi_g42820(csa_tree_add_190_195_groupi_n_6253 ,csa_tree_add_190_195_groupi_n_5881 ,csa_tree_add_190_195_groupi_n_5346);
  or csa_tree_add_190_195_groupi_g42821(csa_tree_add_190_195_groupi_n_6252 ,csa_tree_add_190_195_groupi_n_4840 ,csa_tree_add_190_195_groupi_n_5676);
  and csa_tree_add_190_195_groupi_g42822(csa_tree_add_190_195_groupi_n_6251 ,csa_tree_add_190_195_groupi_n_4784 ,csa_tree_add_190_195_groupi_n_5289);
  and csa_tree_add_190_195_groupi_g42823(csa_tree_add_190_195_groupi_n_6250 ,csa_tree_add_190_195_groupi_n_5433 ,csa_tree_add_190_195_groupi_n_5253);
  and csa_tree_add_190_195_groupi_g42824(csa_tree_add_190_195_groupi_n_6249 ,csa_tree_add_190_195_groupi_n_4826 ,csa_tree_add_190_195_groupi_n_5835);
  or csa_tree_add_190_195_groupi_g42825(csa_tree_add_190_195_groupi_n_6248 ,csa_tree_add_190_195_groupi_n_4839 ,csa_tree_add_190_195_groupi_n_5617);
  nor csa_tree_add_190_195_groupi_g42826(csa_tree_add_190_195_groupi_n_6247 ,csa_tree_add_190_195_groupi_n_5122 ,csa_tree_add_190_195_groupi_n_5809);
  and csa_tree_add_190_195_groupi_g42827(csa_tree_add_190_195_groupi_n_6246 ,csa_tree_add_190_195_groupi_n_5146 ,csa_tree_add_190_195_groupi_n_5799);
  and csa_tree_add_190_195_groupi_g42828(csa_tree_add_190_195_groupi_n_6245 ,csa_tree_add_190_195_groupi_n_4918 ,csa_tree_add_190_195_groupi_n_5949);
  or csa_tree_add_190_195_groupi_g42829(csa_tree_add_190_195_groupi_n_6244 ,csa_tree_add_190_195_groupi_n_5433 ,csa_tree_add_190_195_groupi_n_5253);
  or csa_tree_add_190_195_groupi_g42830(csa_tree_add_190_195_groupi_n_6243 ,csa_tree_add_190_195_groupi_n_5516 ,csa_tree_add_190_195_groupi_n_5247);
  or csa_tree_add_190_195_groupi_g42831(csa_tree_add_190_195_groupi_n_6242 ,csa_tree_add_190_195_groupi_n_2397 ,csa_tree_add_190_195_groupi_n_5541);
  and csa_tree_add_190_195_groupi_g42832(csa_tree_add_190_195_groupi_n_6241 ,csa_tree_add_190_195_groupi_n_4811 ,csa_tree_add_190_195_groupi_n_5666);
  and csa_tree_add_190_195_groupi_g42833(csa_tree_add_190_195_groupi_n_6240 ,csa_tree_add_190_195_groupi_n_5443 ,csa_tree_add_190_195_groupi_n_5336);
  and csa_tree_add_190_195_groupi_g42834(csa_tree_add_190_195_groupi_n_6239 ,csa_tree_add_190_195_groupi_n_4570 ,csa_tree_add_190_195_groupi_n_5514);
  or csa_tree_add_190_195_groupi_g42835(csa_tree_add_190_195_groupi_n_6238 ,csa_tree_add_190_195_groupi_n_4694 ,csa_tree_add_190_195_groupi_n_5374);
  nor csa_tree_add_190_195_groupi_g42836(csa_tree_add_190_195_groupi_n_6237 ,csa_tree_add_190_195_groupi_n_5420 ,csa_tree_add_190_195_groupi_n_5268);
  and csa_tree_add_190_195_groupi_g42837(csa_tree_add_190_195_groupi_n_6236 ,csa_tree_add_190_195_groupi_n_196 ,csa_tree_add_190_195_groupi_n_5283);
  and csa_tree_add_190_195_groupi_g42838(csa_tree_add_190_195_groupi_n_6235 ,csa_tree_add_190_195_groupi_n_4708 ,csa_tree_add_190_195_groupi_n_5207);
  or csa_tree_add_190_195_groupi_g42839(csa_tree_add_190_195_groupi_n_6234 ,csa_tree_add_190_195_groupi_n_5444 ,csa_tree_add_190_195_groupi_n_5225);
  nor csa_tree_add_190_195_groupi_g42840(csa_tree_add_190_195_groupi_n_6233 ,csa_tree_add_190_195_groupi_n_4760 ,csa_tree_add_190_195_groupi_n_5265);
  or csa_tree_add_190_195_groupi_g42841(csa_tree_add_190_195_groupi_n_6232 ,csa_tree_add_190_195_groupi_n_4628 ,csa_tree_add_190_195_groupi_n_5323);
  or csa_tree_add_190_195_groupi_g42842(csa_tree_add_190_195_groupi_n_6231 ,csa_tree_add_190_195_groupi_n_5144 ,csa_tree_add_190_195_groupi_n_5744);
  or csa_tree_add_190_195_groupi_g42843(csa_tree_add_190_195_groupi_n_6230 ,csa_tree_add_190_195_groupi_n_4761 ,csa_tree_add_190_195_groupi_n_5264);
  or csa_tree_add_190_195_groupi_g42844(csa_tree_add_190_195_groupi_n_6229 ,csa_tree_add_190_195_groupi_n_463 ,csa_tree_add_190_195_groupi_n_5241);
  nor csa_tree_add_190_195_groupi_g42845(csa_tree_add_190_195_groupi_n_6228 ,csa_tree_add_190_195_groupi_n_5266 ,csa_tree_add_190_195_groupi_n_5311);
  and csa_tree_add_190_195_groupi_g42846(csa_tree_add_190_195_groupi_n_6227 ,csa_tree_add_190_195_groupi_n_4752 ,csa_tree_add_190_195_groupi_n_5246);
  and csa_tree_add_190_195_groupi_g42847(csa_tree_add_190_195_groupi_n_6226 ,csa_tree_add_190_195_groupi_n_5260 ,csa_tree_add_190_195_groupi_n_5259);
  or csa_tree_add_190_195_groupi_g42848(csa_tree_add_190_195_groupi_n_6225 ,csa_tree_add_190_195_groupi_n_2899 ,csa_tree_add_190_195_groupi_n_5564);
  or csa_tree_add_190_195_groupi_g42849(csa_tree_add_190_195_groupi_n_6224 ,csa_tree_add_190_195_groupi_n_5124 ,csa_tree_add_190_195_groupi_n_5692);
  or csa_tree_add_190_195_groupi_g42850(csa_tree_add_190_195_groupi_n_6223 ,csa_tree_add_190_195_groupi_n_5948 ,csa_tree_add_190_195_groupi_n_5276);
  nor csa_tree_add_190_195_groupi_g42851(csa_tree_add_190_195_groupi_n_6222 ,csa_tree_add_190_195_groupi_n_4906 ,csa_tree_add_190_195_groupi_n_5893);
  nor csa_tree_add_190_195_groupi_g42852(csa_tree_add_190_195_groupi_n_6221 ,csa_tree_add_190_195_groupi_n_5545 ,csa_tree_add_190_195_groupi_n_5470);
  and csa_tree_add_190_195_groupi_g42853(csa_tree_add_190_195_groupi_n_6220 ,csa_tree_add_190_195_groupi_n_4904 ,csa_tree_add_190_195_groupi_n_5892);
  or csa_tree_add_190_195_groupi_g42854(csa_tree_add_190_195_groupi_n_6219 ,csa_tree_add_190_195_groupi_n_4845 ,csa_tree_add_190_195_groupi_n_5618);
  and csa_tree_add_190_195_groupi_g42855(csa_tree_add_190_195_groupi_n_6218 ,csa_tree_add_190_195_groupi_n_5233 ,csa_tree_add_190_195_groupi_n_5463);
  or csa_tree_add_190_195_groupi_g42856(csa_tree_add_190_195_groupi_n_6217 ,csa_tree_add_190_195_groupi_n_2404 ,csa_tree_add_190_195_groupi_n_5252);
  or csa_tree_add_190_195_groupi_g42857(csa_tree_add_190_195_groupi_n_6216 ,csa_tree_add_190_195_groupi_n_4905 ,csa_tree_add_190_195_groupi_n_5894);
  nor csa_tree_add_190_195_groupi_g42858(csa_tree_add_190_195_groupi_n_6215 ,csa_tree_add_190_195_groupi_n_1189 ,csa_tree_add_190_195_groupi_n_5504);
  or csa_tree_add_190_195_groupi_g42859(csa_tree_add_190_195_groupi_n_6214 ,csa_tree_add_190_195_groupi_n_4737 ,csa_tree_add_190_195_groupi_n_5461);
  and csa_tree_add_190_195_groupi_g42860(csa_tree_add_190_195_groupi_n_6213 ,csa_tree_add_190_195_groupi_n_4978 ,csa_tree_add_190_195_groupi_n_5299);
  nor csa_tree_add_190_195_groupi_g42861(csa_tree_add_190_195_groupi_n_6212 ,csa_tree_add_190_195_groupi_n_5515 ,csa_tree_add_190_195_groupi_n_5248);
  or csa_tree_add_190_195_groupi_g42862(csa_tree_add_190_195_groupi_n_6211 ,csa_tree_add_190_195_groupi_n_5197 ,csa_tree_add_190_195_groupi_n_5527);
  and csa_tree_add_190_195_groupi_g42863(csa_tree_add_190_195_groupi_n_6210 ,csa_tree_add_190_195_groupi_n_5472 ,csa_tree_add_190_195_groupi_n_5316);
  and csa_tree_add_190_195_groupi_g42864(csa_tree_add_190_195_groupi_n_6209 ,csa_tree_add_190_195_groupi_n_4651 ,csa_tree_add_190_195_groupi_n_5416);
  or csa_tree_add_190_195_groupi_g42865(csa_tree_add_190_195_groupi_n_6208 ,csa_tree_add_190_195_groupi_n_5436 ,csa_tree_add_190_195_groupi_n_5224);
  or csa_tree_add_190_195_groupi_g42866(csa_tree_add_190_195_groupi_n_6207 ,csa_tree_add_190_195_groupi_n_2401 ,csa_tree_add_190_195_groupi_n_5244);
  and csa_tree_add_190_195_groupi_g42867(csa_tree_add_190_195_groupi_n_6206 ,csa_tree_add_190_195_groupi_n_28 ,csa_tree_add_190_195_groupi_n_5549);
  or csa_tree_add_190_195_groupi_g42869(csa_tree_add_190_195_groupi_n_6205 ,csa_tree_add_190_195_groupi_n_5243 ,csa_tree_add_190_195_groupi_n_5242);
  or csa_tree_add_190_195_groupi_g42870(csa_tree_add_190_195_groupi_n_6204 ,csa_tree_add_190_195_groupi_n_5434 ,csa_tree_add_190_195_groupi_n_5533);
  nor csa_tree_add_190_195_groupi_g42871(csa_tree_add_190_195_groupi_n_6203 ,csa_tree_add_190_195_groupi_n_28 ,csa_tree_add_190_195_groupi_n_5549);
  or csa_tree_add_190_195_groupi_g42872(csa_tree_add_190_195_groupi_n_6202 ,csa_tree_add_190_195_groupi_n_1330 ,csa_tree_add_190_195_groupi_n_5211);
  or csa_tree_add_190_195_groupi_g42873(csa_tree_add_190_195_groupi_n_6201 ,csa_tree_add_190_195_groupi_n_5421 ,csa_tree_add_190_195_groupi_n_5267);
  nor csa_tree_add_190_195_groupi_g42874(csa_tree_add_190_195_groupi_n_6200 ,csa_tree_add_190_195_groupi_n_4640 ,csa_tree_add_190_195_groupi_n_5327);
  or csa_tree_add_190_195_groupi_g42875(csa_tree_add_190_195_groupi_n_6199 ,csa_tree_add_190_195_groupi_n_2400 ,csa_tree_add_190_195_groupi_n_5517);
  and csa_tree_add_190_195_groupi_g42876(csa_tree_add_190_195_groupi_n_6198 ,csa_tree_add_190_195_groupi_n_4662 ,csa_tree_add_190_195_groupi_n_5240);
  nor csa_tree_add_190_195_groupi_g42877(csa_tree_add_190_195_groupi_n_6197 ,csa_tree_add_190_195_groupi_n_5526 ,csa_tree_add_190_195_groupi_n_5221);
  and csa_tree_add_190_195_groupi_g42878(csa_tree_add_190_195_groupi_n_6196 ,csa_tree_add_190_195_groupi_n_4898 ,csa_tree_add_190_195_groupi_n_5429);
  and csa_tree_add_190_195_groupi_g42879(csa_tree_add_190_195_groupi_n_6195 ,csa_tree_add_190_195_groupi_n_5351 ,csa_tree_add_190_195_groupi_n_5495);
  nor csa_tree_add_190_195_groupi_g42880(csa_tree_add_190_195_groupi_n_6194 ,csa_tree_add_190_195_groupi_n_5214 ,csa_tree_add_190_195_groupi_n_5547);
  or csa_tree_add_190_195_groupi_g42881(csa_tree_add_190_195_groupi_n_6193 ,csa_tree_add_190_195_groupi_n_4711 ,csa_tree_add_190_195_groupi_n_5272);
  or csa_tree_add_190_195_groupi_g42882(csa_tree_add_190_195_groupi_n_6192 ,csa_tree_add_190_195_groupi_n_5213 ,csa_tree_add_190_195_groupi_n_5548);
  and csa_tree_add_190_195_groupi_g42883(csa_tree_add_190_195_groupi_n_6191 ,csa_tree_add_190_195_groupi_n_5908 ,csa_tree_add_190_195_groupi_n_5929);
  or csa_tree_add_190_195_groupi_g42884(csa_tree_add_190_195_groupi_n_6190 ,csa_tree_add_190_195_groupi_n_5217 ,csa_tree_add_190_195_groupi_n_5302);
  or csa_tree_add_190_195_groupi_g42885(csa_tree_add_190_195_groupi_n_6189 ,csa_tree_add_190_195_groupi_n_5113 ,csa_tree_add_190_195_groupi_n_5615);
  nor csa_tree_add_190_195_groupi_g42886(csa_tree_add_190_195_groupi_n_6188 ,csa_tree_add_190_195_groupi_n_4712 ,csa_tree_add_190_195_groupi_n_5271);
  and csa_tree_add_190_195_groupi_g42887(csa_tree_add_190_195_groupi_n_6187 ,csa_tree_add_190_195_groupi_n_5152 ,csa_tree_add_190_195_groupi_n_5664);
  nor csa_tree_add_190_195_groupi_g42888(csa_tree_add_190_195_groupi_n_6186 ,csa_tree_add_190_195_groupi_n_4960 ,csa_tree_add_190_195_groupi_n_5907);
  or csa_tree_add_190_195_groupi_g42889(csa_tree_add_190_195_groupi_n_6185 ,csa_tree_add_190_195_groupi_n_900 ,csa_tree_add_190_195_groupi_n_5283);
  and csa_tree_add_190_195_groupi_g42890(csa_tree_add_190_195_groupi_n_6184 ,csa_tree_add_190_195_groupi_n_4829 ,csa_tree_add_190_195_groupi_n_5864);
  nor csa_tree_add_190_195_groupi_g42891(csa_tree_add_190_195_groupi_n_6183 ,csa_tree_add_190_195_groupi_n_4738 ,csa_tree_add_190_195_groupi_n_5460);
  and csa_tree_add_190_195_groupi_g42892(csa_tree_add_190_195_groupi_n_6182 ,csa_tree_add_190_195_groupi_n_5229 ,csa_tree_add_190_195_groupi_n_5230);
  or csa_tree_add_190_195_groupi_g42893(csa_tree_add_190_195_groupi_n_6181 ,csa_tree_add_190_195_groupi_n_5888 ,csa_tree_add_190_195_groupi_n_5542);
  or csa_tree_add_190_195_groupi_g42894(csa_tree_add_190_195_groupi_n_6180 ,csa_tree_add_190_195_groupi_n_5061 ,csa_tree_add_190_195_groupi_n_5539);
  nor csa_tree_add_190_195_groupi_g42895(csa_tree_add_190_195_groupi_n_6179 ,csa_tree_add_190_195_groupi_n_5062 ,csa_tree_add_190_195_groupi_n_5540);
  or csa_tree_add_190_195_groupi_g42896(csa_tree_add_190_195_groupi_n_6178 ,csa_tree_add_190_195_groupi_n_5510 ,csa_tree_add_190_195_groupi_n_5445);
  or csa_tree_add_190_195_groupi_g42897(csa_tree_add_190_195_groupi_n_6177 ,csa_tree_add_190_195_groupi_n_5441 ,csa_tree_add_190_195_groupi_n_5537);
  or csa_tree_add_190_195_groupi_g42898(csa_tree_add_190_195_groupi_n_6176 ,csa_tree_add_190_195_groupi_n_5112 ,csa_tree_add_190_195_groupi_n_5667);
  nor csa_tree_add_190_195_groupi_g42899(csa_tree_add_190_195_groupi_n_6175 ,csa_tree_add_190_195_groupi_n_5511 ,csa_tree_add_190_195_groupi_n_5446);
  and csa_tree_add_190_195_groupi_g42900(csa_tree_add_190_195_groupi_n_6174 ,csa_tree_add_190_195_groupi_n_5160 ,csa_tree_add_190_195_groupi_n_5628);
  nor csa_tree_add_190_195_groupi_g42901(csa_tree_add_190_195_groupi_n_6173 ,csa_tree_add_190_195_groupi_n_5440 ,csa_tree_add_190_195_groupi_n_5538);
  and csa_tree_add_190_195_groupi_g42902(csa_tree_add_190_195_groupi_n_6172 ,csa_tree_add_190_195_groupi_n_5444 ,csa_tree_add_190_195_groupi_n_5225);
  and csa_tree_add_190_195_groupi_g42903(csa_tree_add_190_195_groupi_n_6171 ,csa_tree_add_190_195_groupi_n_5436 ,csa_tree_add_190_195_groupi_n_5224);
  and csa_tree_add_190_195_groupi_g42904(csa_tree_add_190_195_groupi_n_6170 ,csa_tree_add_190_195_groupi_n_4676 ,csa_tree_add_190_195_groupi_n_5258);
  or csa_tree_add_190_195_groupi_g42905(csa_tree_add_190_195_groupi_n_6169 ,csa_tree_add_190_195_groupi_n_5525 ,csa_tree_add_190_195_groupi_n_66);
  nor csa_tree_add_190_195_groupi_g42906(csa_tree_add_190_195_groupi_n_6168 ,csa_tree_add_190_195_groupi_n_5198 ,csa_tree_add_190_195_groupi_n_5528);
  or csa_tree_add_190_195_groupi_g42907(csa_tree_add_190_195_groupi_n_6167 ,csa_tree_add_190_195_groupi_n_29 ,csa_tree_add_190_195_groupi_n_5312);
  or csa_tree_add_190_195_groupi_g42908(csa_tree_add_190_195_groupi_n_6166 ,csa_tree_add_190_195_groupi_n_2897 ,csa_tree_add_190_195_groupi_n_5606);
  and csa_tree_add_190_195_groupi_g42910(csa_tree_add_190_195_groupi_n_6165 ,csa_tree_add_190_195_groupi_n_4827 ,csa_tree_add_190_195_groupi_n_5855);
  nor csa_tree_add_190_195_groupi_g42911(csa_tree_add_190_195_groupi_n_6164 ,csa_tree_add_190_195_groupi_n_5435 ,csa_tree_add_190_195_groupi_n_5532);
  or csa_tree_add_190_195_groupi_g42912(csa_tree_add_190_195_groupi_n_6163 ,csa_tree_add_190_195_groupi_n_4764 ,csa_tree_add_190_195_groupi_n_5387);
  and csa_tree_add_190_195_groupi_g42913(csa_tree_add_190_195_groupi_n_6162 ,csa_tree_add_190_195_groupi_n_5263 ,csa_tree_add_190_195_groupi_n_5297);
  or csa_tree_add_190_195_groupi_g42914(csa_tree_add_190_195_groupi_n_6161 ,csa_tree_add_190_195_groupi_n_5409 ,csa_tree_add_190_195_groupi_n_5301);
  and csa_tree_add_190_195_groupi_g42915(csa_tree_add_190_195_groupi_n_6160 ,csa_tree_add_190_195_groupi_n_4706 ,csa_tree_add_190_195_groupi_n_5288);
  nor csa_tree_add_190_195_groupi_g42916(csa_tree_add_190_195_groupi_n_6159 ,csa_tree_add_190_195_groupi_n_5524 ,csa_tree_add_190_195_groupi_n_5519);
  or csa_tree_add_190_195_groupi_g42917(csa_tree_add_190_195_groupi_n_6158 ,csa_tree_add_190_195_groupi_n_4639 ,csa_tree_add_190_195_groupi_n_5328);
  or csa_tree_add_190_195_groupi_g42918(csa_tree_add_190_195_groupi_n_6157 ,csa_tree_add_190_195_groupi_n_5190 ,csa_tree_add_190_195_groupi_n_71);
  or csa_tree_add_190_195_groupi_g42919(csa_tree_add_190_195_groupi_n_6156 ,csa_tree_add_190_195_groupi_n_5523 ,csa_tree_add_190_195_groupi_n_5518);
  or csa_tree_add_190_195_groupi_g42920(csa_tree_add_190_195_groupi_n_6155 ,csa_tree_add_190_195_groupi_n_4832 ,csa_tree_add_190_195_groupi_n_5645);
  or csa_tree_add_190_195_groupi_g42921(csa_tree_add_190_195_groupi_n_6154 ,csa_tree_add_190_195_groupi_n_4965 ,csa_tree_add_190_195_groupi_n_5216);
  or csa_tree_add_190_195_groupi_g42922(csa_tree_add_190_195_groupi_n_6153 ,csa_tree_add_190_195_groupi_n_5672 ,csa_tree_add_190_195_groupi_n_5965);
  nor csa_tree_add_190_195_groupi_g42923(csa_tree_add_190_195_groupi_n_6152 ,csa_tree_add_190_195_groupi_n_5132 ,csa_tree_add_190_195_groupi_n_5820);
  nor csa_tree_add_190_195_groupi_g42924(csa_tree_add_190_195_groupi_n_6151 ,csa_tree_add_190_195_groupi_n_1313 ,csa_tree_add_190_195_groupi_n_5238);
  nor csa_tree_add_190_195_groupi_g42925(csa_tree_add_190_195_groupi_n_6150 ,csa_tree_add_190_195_groupi_n_5962 ,csa_tree_add_190_195_groupi_n_5960);
  or csa_tree_add_190_195_groupi_g42926(csa_tree_add_190_195_groupi_n_6149 ,csa_tree_add_190_195_groupi_n_5116 ,csa_tree_add_190_195_groupi_n_5779);
  or csa_tree_add_190_195_groupi_g42927(csa_tree_add_190_195_groupi_n_6148 ,csa_tree_add_190_195_groupi_n_4676 ,csa_tree_add_190_195_groupi_n_5258);
  and csa_tree_add_190_195_groupi_g42928(csa_tree_add_190_195_groupi_n_6147 ,csa_tree_add_190_195_groupi_n_4799 ,csa_tree_add_190_195_groupi_n_5857);
  nor csa_tree_add_190_195_groupi_g42929(csa_tree_add_190_195_groupi_n_6146 ,csa_tree_add_190_195_groupi_n_4862 ,csa_tree_add_190_195_groupi_n_5847);
  and csa_tree_add_190_195_groupi_g42930(csa_tree_add_190_195_groupi_n_6145 ,csa_tree_add_190_195_groupi_n_3451 ,csa_tree_add_190_195_groupi_n_59);
  and csa_tree_add_190_195_groupi_g42931(csa_tree_add_190_195_groupi_n_6144 ,csa_tree_add_190_195_groupi_n_4569 ,csa_tree_add_190_195_groupi_n_5468);
  or csa_tree_add_190_195_groupi_g42932(csa_tree_add_190_195_groupi_n_6143 ,csa_tree_add_190_195_groupi_n_4135 ,csa_tree_add_190_195_groupi_n_5203);
  and csa_tree_add_190_195_groupi_g42933(csa_tree_add_190_195_groupi_n_6142 ,csa_tree_add_190_195_groupi_n_3070 ,csa_tree_add_190_195_groupi_n_5603);
  nor csa_tree_add_190_195_groupi_g42934(csa_tree_add_190_195_groupi_n_6141 ,csa_tree_add_190_195_groupi_n_4658 ,csa_tree_add_190_195_groupi_n_5458);
  nor csa_tree_add_190_195_groupi_g42935(csa_tree_add_190_195_groupi_n_6140 ,csa_tree_add_190_195_groupi_n_4810 ,csa_tree_add_190_195_groupi_n_5656);
  or csa_tree_add_190_195_groupi_g42936(csa_tree_add_190_195_groupi_n_6139 ,csa_tree_add_190_195_groupi_n_4659 ,csa_tree_add_190_195_groupi_n_5457);
  or csa_tree_add_190_195_groupi_g42937(csa_tree_add_190_195_groupi_n_6138 ,csa_tree_add_190_195_groupi_n_5068 ,csa_tree_add_190_195_groupi_n_5500);
  and csa_tree_add_190_195_groupi_g42938(csa_tree_add_190_195_groupi_n_6137 ,csa_tree_add_190_195_groupi_n_228 ,csa_tree_add_190_195_groupi_n_5895);
  or csa_tree_add_190_195_groupi_g42939(csa_tree_add_190_195_groupi_n_6136 ,csa_tree_add_190_195_groupi_n_5505 ,csa_tree_add_190_195_groupi_n_5502);
  nor csa_tree_add_190_195_groupi_g42940(csa_tree_add_190_195_groupi_n_6135 ,csa_tree_add_190_195_groupi_n_262 ,csa_tree_add_190_195_groupi_n_5895);
  nor csa_tree_add_190_195_groupi_g42941(csa_tree_add_190_195_groupi_n_6134 ,csa_tree_add_190_195_groupi_n_5506 ,csa_tree_add_190_195_groupi_n_5503);
  or csa_tree_add_190_195_groupi_g42942(csa_tree_add_190_195_groupi_n_6133 ,csa_tree_add_190_195_groupi_n_5202 ,csa_tree_add_190_195_groupi_n_5427);
  nor csa_tree_add_190_195_groupi_g42943(csa_tree_add_190_195_groupi_n_6132 ,csa_tree_add_190_195_groupi_n_5069 ,csa_tree_add_190_195_groupi_n_5501);
  or csa_tree_add_190_195_groupi_g42944(csa_tree_add_190_195_groupi_n_6131 ,csa_tree_add_190_195_groupi_n_77 ,csa_tree_add_190_195_groupi_n_5428);
  or csa_tree_add_190_195_groupi_g42945(csa_tree_add_190_195_groupi_n_6130 ,csa_tree_add_190_195_groupi_n_5419 ,csa_tree_add_190_195_groupi_n_5201);
  or csa_tree_add_190_195_groupi_g42946(csa_tree_add_190_195_groupi_n_6129 ,csa_tree_add_190_195_groupi_n_4648 ,csa_tree_add_190_195_groupi_n_5496);
  nor csa_tree_add_190_195_groupi_g42947(csa_tree_add_190_195_groupi_n_6128 ,csa_tree_add_190_195_groupi_n_4649 ,csa_tree_add_190_195_groupi_n_5497);
  and csa_tree_add_190_195_groupi_g42948(csa_tree_add_190_195_groupi_n_6127 ,csa_tree_add_190_195_groupi_n_4821 ,csa_tree_add_190_195_groupi_n_5621);
  and csa_tree_add_190_195_groupi_g42949(csa_tree_add_190_195_groupi_n_6126 ,csa_tree_add_190_195_groupi_n_5419 ,csa_tree_add_190_195_groupi_n_5201);
  nor csa_tree_add_190_195_groupi_g42950(csa_tree_add_190_195_groupi_n_6125 ,csa_tree_add_190_195_groupi_n_4837 ,csa_tree_add_190_195_groupi_n_5649);
  and csa_tree_add_190_195_groupi_g42951(csa_tree_add_190_195_groupi_n_6124 ,csa_tree_add_190_195_groupi_n_5545 ,csa_tree_add_190_195_groupi_n_5470);
  and csa_tree_add_190_195_groupi_g42952(csa_tree_add_190_195_groupi_n_6123 ,csa_tree_add_190_195_groupi_n_5202 ,csa_tree_add_190_195_groupi_n_5427);
  or csa_tree_add_190_195_groupi_g42953(csa_tree_add_190_195_groupi_n_6122 ,csa_tree_add_190_195_groupi_n_4920 ,csa_tree_add_190_195_groupi_n_5182);
  and csa_tree_add_190_195_groupi_g42954(csa_tree_add_190_195_groupi_n_6121 ,csa_tree_add_190_195_groupi_n_4865 ,csa_tree_add_190_195_groupi_n_5782);
  and csa_tree_add_190_195_groupi_g42955(csa_tree_add_190_195_groupi_n_6120 ,csa_tree_add_190_195_groupi_n_4135 ,csa_tree_add_190_195_groupi_n_5203);
  and csa_tree_add_190_195_groupi_g42956(csa_tree_add_190_195_groupi_n_6119 ,csa_tree_add_190_195_groupi_n_5595 ,csa_tree_add_190_195_groupi_n_5840);
  and csa_tree_add_190_195_groupi_g42957(csa_tree_add_190_195_groupi_n_6118 ,csa_tree_add_190_195_groupi_n_4803 ,csa_tree_add_190_195_groupi_n_5777);
  and csa_tree_add_190_195_groupi_g42958(csa_tree_add_190_195_groupi_n_6117 ,csa_tree_add_190_195_groupi_n_4804 ,csa_tree_add_190_195_groupi_n_5641);
  or csa_tree_add_190_195_groupi_g42959(csa_tree_add_190_195_groupi_n_6116 ,csa_tree_add_190_195_groupi_n_5093 ,csa_tree_add_190_195_groupi_n_5957);
  and csa_tree_add_190_195_groupi_g42960(csa_tree_add_190_195_groupi_n_6115 ,csa_tree_add_190_195_groupi_n_5491 ,csa_tree_add_190_195_groupi_n_5488);
  and csa_tree_add_190_195_groupi_g42961(csa_tree_add_190_195_groupi_n_6114 ,csa_tree_add_190_195_groupi_n_3414 ,csa_tree_add_190_195_groupi_n_5601);
  nor csa_tree_add_190_195_groupi_g42962(csa_tree_add_190_195_groupi_n_6113 ,csa_tree_add_190_195_groupi_n_5489 ,csa_tree_add_190_195_groupi_n_42);
  and csa_tree_add_190_195_groupi_g42963(csa_tree_add_190_195_groupi_n_6112 ,csa_tree_add_190_195_groupi_n_4618 ,csa_tree_add_190_195_groupi_n_5402);
  nor csa_tree_add_190_195_groupi_g42964(csa_tree_add_190_195_groupi_n_6111 ,csa_tree_add_190_195_groupi_n_5885 ,csa_tree_add_190_195_groupi_n_5879);
  or csa_tree_add_190_195_groupi_g42965(csa_tree_add_190_195_groupi_n_6110 ,csa_tree_add_190_195_groupi_n_5490 ,csa_tree_add_190_195_groupi_n_5194);
  or csa_tree_add_190_195_groupi_g42966(csa_tree_add_190_195_groupi_n_6109 ,csa_tree_add_190_195_groupi_n_5483 ,csa_tree_add_190_195_groupi_n_5189);
  nor csa_tree_add_190_195_groupi_g42967(csa_tree_add_190_195_groupi_n_6108 ,csa_tree_add_190_195_groupi_n_5484 ,csa_tree_add_190_195_groupi_n_5188);
  nor csa_tree_add_190_195_groupi_g42968(csa_tree_add_190_195_groupi_n_6107 ,csa_tree_add_190_195_groupi_n_5491 ,csa_tree_add_190_195_groupi_n_5488);
  or csa_tree_add_190_195_groupi_g42969(csa_tree_add_190_195_groupi_n_6106 ,csa_tree_add_190_195_groupi_n_4978 ,csa_tree_add_190_195_groupi_n_5299);
  or csa_tree_add_190_195_groupi_g42970(csa_tree_add_190_195_groupi_n_6105 ,csa_tree_add_190_195_groupi_n_4801 ,csa_tree_add_190_195_groupi_n_5642);
  nor csa_tree_add_190_195_groupi_g42971(csa_tree_add_190_195_groupi_n_6104 ,csa_tree_add_190_195_groupi_n_5924 ,csa_tree_add_190_195_groupi_n_5951);
  nor csa_tree_add_190_195_groupi_g42972(csa_tree_add_190_195_groupi_n_6103 ,csa_tree_add_190_195_groupi_n_5477 ,csa_tree_add_190_195_groupi_n_5187);
  or csa_tree_add_190_195_groupi_g42973(csa_tree_add_190_195_groupi_n_6102 ,csa_tree_add_190_195_groupi_n_5475 ,csa_tree_add_190_195_groupi_n_5426);
  or csa_tree_add_190_195_groupi_g42974(csa_tree_add_190_195_groupi_n_6101 ,csa_tree_add_190_195_groupi_n_5478 ,csa_tree_add_190_195_groupi_n_5186);
  nor csa_tree_add_190_195_groupi_g42975(csa_tree_add_190_195_groupi_n_6100 ,csa_tree_add_190_195_groupi_n_61 ,csa_tree_add_190_195_groupi_n_5476);
  and csa_tree_add_190_195_groupi_g42976(csa_tree_add_190_195_groupi_n_6099 ,csa_tree_add_190_195_groupi_n_38 ,csa_tree_add_190_195_groupi_n_5639);
  and csa_tree_add_190_195_groupi_g42977(csa_tree_add_190_195_groupi_n_6098 ,csa_tree_add_190_195_groupi_n_5938 ,csa_tree_add_190_195_groupi_n_5469);
  and csa_tree_add_190_195_groupi_g42978(csa_tree_add_190_195_groupi_n_6097 ,csa_tree_add_190_195_groupi_n_54 ,csa_tree_add_190_195_groupi_n_5896);
  nor csa_tree_add_190_195_groupi_g42979(csa_tree_add_190_195_groupi_n_6096 ,csa_tree_add_190_195_groupi_n_5938 ,csa_tree_add_190_195_groupi_n_5469);
  and csa_tree_add_190_195_groupi_g42980(csa_tree_add_190_195_groupi_n_6095 ,csa_tree_add_190_195_groupi_n_5466 ,csa_tree_add_190_195_groupi_n_5465);
  nor csa_tree_add_190_195_groupi_g42981(csa_tree_add_190_195_groupi_n_6094 ,csa_tree_add_190_195_groupi_n_1928 ,csa_tree_add_190_195_groupi_n_5920);
  nor csa_tree_add_190_195_groupi_g42982(csa_tree_add_190_195_groupi_n_6093 ,csa_tree_add_190_195_groupi_n_5466 ,csa_tree_add_190_195_groupi_n_5465);
  nor csa_tree_add_190_195_groupi_g42983(csa_tree_add_190_195_groupi_n_6092 ,csa_tree_add_190_195_groupi_n_4831 ,csa_tree_add_190_195_groupi_n_5635);
  or csa_tree_add_190_195_groupi_g42984(csa_tree_add_190_195_groupi_n_6091 ,csa_tree_add_190_195_groupi_n_4682 ,csa_tree_add_190_195_groupi_n_5459);
  and csa_tree_add_190_195_groupi_g42985(csa_tree_add_190_195_groupi_n_6090 ,csa_tree_add_190_195_groupi_n_4682 ,csa_tree_add_190_195_groupi_n_5459);
  nor csa_tree_add_190_195_groupi_g42986(csa_tree_add_190_195_groupi_n_6089 ,csa_tree_add_190_195_groupi_n_4802 ,csa_tree_add_190_195_groupi_n_5633);
  and csa_tree_add_190_195_groupi_g42987(csa_tree_add_190_195_groupi_n_6088 ,csa_tree_add_190_195_groupi_n_4836 ,csa_tree_add_190_195_groupi_n_5616);
  xnor csa_tree_add_190_195_groupi_g42988(csa_tree_add_190_195_groupi_n_6087 ,csa_tree_add_190_195_groupi_n_3699 ,csa_tree_add_190_195_groupi_n_5086);
  xnor csa_tree_add_190_195_groupi_g42989(csa_tree_add_190_195_groupi_n_6086 ,csa_tree_add_190_195_groupi_n_4731 ,csa_tree_add_190_195_groupi_n_4720);
  xor csa_tree_add_190_195_groupi_g42990(csa_tree_add_190_195_groupi_n_6085 ,csa_tree_add_190_195_groupi_n_5119 ,csa_tree_add_190_195_groupi_n_5053);
  xnor csa_tree_add_190_195_groupi_g42991(csa_tree_add_190_195_groupi_n_6084 ,csa_tree_add_190_195_groupi_n_4642 ,csa_tree_add_190_195_groupi_n_1961);
  xnor csa_tree_add_190_195_groupi_g42992(csa_tree_add_190_195_groupi_n_6083 ,csa_tree_add_190_195_groupi_n_4653 ,csa_tree_add_190_195_groupi_n_5009);
  xnor csa_tree_add_190_195_groupi_g42993(csa_tree_add_190_195_groupi_n_6082 ,csa_tree_add_190_195_groupi_n_4689 ,csa_tree_add_190_195_groupi_n_4881);
  xor csa_tree_add_190_195_groupi_g42994(csa_tree_add_190_195_groupi_n_6081 ,csa_tree_add_190_195_groupi_n_5149 ,csa_tree_add_190_195_groupi_n_4924);
  xor csa_tree_add_190_195_groupi_g42995(csa_tree_add_190_195_groupi_n_6080 ,csa_tree_add_190_195_groupi_n_5098 ,csa_tree_add_190_195_groupi_n_4918);
  xnor csa_tree_add_190_195_groupi_g42996(csa_tree_add_190_195_groupi_n_6079 ,csa_tree_add_190_195_groupi_n_5067 ,csa_tree_add_190_195_groupi_n_1741);
  xnor csa_tree_add_190_195_groupi_g42997(csa_tree_add_190_195_groupi_n_6078 ,csa_tree_add_190_195_groupi_n_4595 ,csa_tree_add_190_195_groupi_n_5084);
  xor csa_tree_add_190_195_groupi_g42998(csa_tree_add_190_195_groupi_n_6077 ,csa_tree_add_190_195_groupi_n_5128 ,csa_tree_add_190_195_groupi_n_1846);
  xnor csa_tree_add_190_195_groupi_g42999(csa_tree_add_190_195_groupi_n_6076 ,csa_tree_add_190_195_groupi_n_5106 ,csa_tree_add_190_195_groupi_n_1156);
  xnor csa_tree_add_190_195_groupi_g43000(csa_tree_add_190_195_groupi_n_6075 ,csa_tree_add_190_195_groupi_n_5014 ,csa_tree_add_190_195_groupi_n_5029);
  xnor csa_tree_add_190_195_groupi_g43001(csa_tree_add_190_195_groupi_n_6074 ,csa_tree_add_190_195_groupi_n_5004 ,csa_tree_add_190_195_groupi_n_1811);
  xnor csa_tree_add_190_195_groupi_g43002(csa_tree_add_190_195_groupi_n_6073 ,csa_tree_add_190_195_groupi_n_5140 ,csa_tree_add_190_195_groupi_n_1095);
  xor csa_tree_add_190_195_groupi_g43003(csa_tree_add_190_195_groupi_n_6072 ,csa_tree_add_190_195_groupi_n_4617 ,csa_tree_add_190_195_groupi_n_4850);
  xnor csa_tree_add_190_195_groupi_g43004(csa_tree_add_190_195_groupi_n_6071 ,csa_tree_add_190_195_groupi_n_4801 ,csa_tree_add_190_195_groupi_n_960);
  xnor csa_tree_add_190_195_groupi_g43005(csa_tree_add_190_195_groupi_n_6070 ,csa_tree_add_190_195_groupi_n_4693 ,csa_tree_add_190_195_groupi_n_4685);
  xor csa_tree_add_190_195_groupi_g43006(csa_tree_add_190_195_groupi_n_6069 ,csa_tree_add_190_195_groupi_n_4838 ,csa_tree_add_190_195_groupi_n_4569);
  xnor csa_tree_add_190_195_groupi_g43007(csa_tree_add_190_195_groupi_n_6068 ,csa_tree_add_190_195_groupi_n_4563 ,csa_tree_add_190_195_groupi_n_4741);
  xnor csa_tree_add_190_195_groupi_g43008(csa_tree_add_190_195_groupi_n_6067 ,csa_tree_add_190_195_groupi_n_5097 ,csa_tree_add_190_195_groupi_n_4743);
  xnor csa_tree_add_190_195_groupi_g43009(csa_tree_add_190_195_groupi_n_6066 ,csa_tree_add_190_195_groupi_n_5133 ,csa_tree_add_190_195_groupi_n_2055);
  xor csa_tree_add_190_195_groupi_g43010(csa_tree_add_190_195_groupi_n_6065 ,csa_tree_add_190_195_groupi_n_4908 ,csa_tree_add_190_195_groupi_n_5161);
  xor csa_tree_add_190_195_groupi_g43011(csa_tree_add_190_195_groupi_n_6064 ,csa_tree_add_190_195_groupi_n_4928 ,csa_tree_add_190_195_groupi_n_5143);
  xnor csa_tree_add_190_195_groupi_g43012(csa_tree_add_190_195_groupi_n_6063 ,csa_tree_add_190_195_groupi_n_5071 ,csa_tree_add_190_195_groupi_n_1812);
  xor csa_tree_add_190_195_groupi_g43013(csa_tree_add_190_195_groupi_n_6062 ,csa_tree_add_190_195_groupi_n_5138 ,csa_tree_add_190_195_groupi_n_4987);
  xnor csa_tree_add_190_195_groupi_g43014(csa_tree_add_190_195_groupi_n_6061 ,csa_tree_add_190_195_groupi_n_5007 ,csa_tree_add_190_195_groupi_n_4828);
  xnor csa_tree_add_190_195_groupi_g43015(csa_tree_add_190_195_groupi_n_6060 ,csa_tree_add_190_195_groupi_n_4896 ,csa_tree_add_190_195_groupi_n_3695);
  xnor csa_tree_add_190_195_groupi_g43016(csa_tree_add_190_195_groupi_n_6059 ,csa_tree_add_190_195_groupi_n_4996 ,csa_tree_add_190_195_groupi_n_1866);
  xnor csa_tree_add_190_195_groupi_g43017(csa_tree_add_190_195_groupi_n_6058 ,csa_tree_add_190_195_groupi_n_4806 ,csa_tree_add_190_195_groupi_n_561);
  xnor csa_tree_add_190_195_groupi_g43018(csa_tree_add_190_195_groupi_n_6057 ,csa_tree_add_190_195_groupi_n_5121 ,csa_tree_add_190_195_groupi_n_4981);
  xnor csa_tree_add_190_195_groupi_g43019(csa_tree_add_190_195_groupi_n_6056 ,csa_tree_add_190_195_groupi_n_5045 ,in56[11]);
  xnor csa_tree_add_190_195_groupi_g43020(csa_tree_add_190_195_groupi_n_6055 ,csa_tree_add_190_195_groupi_n_4597 ,csa_tree_add_190_195_groupi_n_4736);
  xnor csa_tree_add_190_195_groupi_g43021(csa_tree_add_190_195_groupi_n_6054 ,csa_tree_add_190_195_groupi_n_5102 ,csa_tree_add_190_195_groupi_n_4985);
  xnor csa_tree_add_190_195_groupi_g43022(csa_tree_add_190_195_groupi_n_6053 ,csa_tree_add_190_195_groupi_n_4775 ,csa_tree_add_190_195_groupi_n_4773);
  xnor csa_tree_add_190_195_groupi_g43023(csa_tree_add_190_195_groupi_n_6052 ,csa_tree_add_190_195_groupi_n_5172 ,csa_tree_add_190_195_groupi_n_1969);
  xnor csa_tree_add_190_195_groupi_g43024(csa_tree_add_190_195_groupi_n_6051 ,csa_tree_add_190_195_groupi_n_4809 ,csa_tree_add_190_195_groupi_n_5025);
  xnor csa_tree_add_190_195_groupi_g43025(csa_tree_add_190_195_groupi_n_6050 ,csa_tree_add_190_195_groupi_n_4969 ,csa_tree_add_190_195_groupi_n_4943);
  xnor csa_tree_add_190_195_groupi_g43026(csa_tree_add_190_195_groupi_n_6049 ,csa_tree_add_190_195_groupi_n_4757 ,csa_tree_add_190_195_groupi_n_4813);
  xnor csa_tree_add_190_195_groupi_g43027(csa_tree_add_190_195_groupi_n_6048 ,csa_tree_add_190_195_groupi_n_4941 ,csa_tree_add_190_195_groupi_n_1944);
  xor csa_tree_add_190_195_groupi_g43028(csa_tree_add_190_195_groupi_n_6047 ,csa_tree_add_190_195_groupi_n_4844 ,csa_tree_add_190_195_groupi_n_5080);
  xnor csa_tree_add_190_195_groupi_g43029(csa_tree_add_190_195_groupi_n_6046 ,csa_tree_add_190_195_groupi_n_4815 ,csa_tree_add_190_195_groupi_n_1928);
  xnor csa_tree_add_190_195_groupi_g43030(csa_tree_add_190_195_groupi_n_6045 ,csa_tree_add_190_195_groupi_n_5064 ,in56[9]);
  xnor csa_tree_add_190_195_groupi_g43031(csa_tree_add_190_195_groupi_n_6044 ,csa_tree_add_190_195_groupi_n_4948 ,in56[10]);
  xnor csa_tree_add_190_195_groupi_g43032(csa_tree_add_190_195_groupi_n_6043 ,csa_tree_add_190_195_groupi_n_4871 ,csa_tree_add_190_195_groupi_n_4979);
  xnor csa_tree_add_190_195_groupi_g43033(csa_tree_add_190_195_groupi_n_6042 ,csa_tree_add_190_195_groupi_n_4619 ,csa_tree_add_190_195_groupi_n_4802);
  xnor csa_tree_add_190_195_groupi_g43034(csa_tree_add_190_195_groupi_n_6041 ,csa_tree_add_190_195_groupi_n_5150 ,csa_tree_add_190_195_groupi_n_2210);
  xnor csa_tree_add_190_195_groupi_g43035(csa_tree_add_190_195_groupi_n_6040 ,csa_tree_add_190_195_groupi_n_4739 ,in60[14]);
  xnor csa_tree_add_190_195_groupi_g43036(csa_tree_add_190_195_groupi_n_6039 ,csa_tree_add_190_195_groupi_n_4909 ,csa_tree_add_190_195_groupi_n_4869);
  xnor csa_tree_add_190_195_groupi_g43037(csa_tree_add_190_195_groupi_n_6038 ,csa_tree_add_190_195_groupi_n_4831 ,csa_tree_add_190_195_groupi_n_5003);
  xnor csa_tree_add_190_195_groupi_g43038(csa_tree_add_190_195_groupi_n_6037 ,csa_tree_add_190_195_groupi_n_4673 ,csa_tree_add_190_195_groupi_n_4843);
  xnor csa_tree_add_190_195_groupi_g43039(csa_tree_add_190_195_groupi_n_6036 ,csa_tree_add_190_195_groupi_n_4839 ,csa_tree_add_190_195_groupi_n_4681);
  xnor csa_tree_add_190_195_groupi_g43040(csa_tree_add_190_195_groupi_n_6035 ,csa_tree_add_190_195_groupi_n_4729 ,csa_tree_add_190_195_groupi_n_5065);
  xnor csa_tree_add_190_195_groupi_g43041(csa_tree_add_190_195_groupi_n_6034 ,csa_tree_add_190_195_groupi_n_5154 ,csa_tree_add_190_195_groupi_n_2089);
  xnor csa_tree_add_190_195_groupi_g43042(csa_tree_add_190_195_groupi_n_6033 ,csa_tree_add_190_195_groupi_n_4584 ,csa_tree_add_190_195_groupi_n_5027);
  xnor csa_tree_add_190_195_groupi_g43043(csa_tree_add_190_195_groupi_n_6032 ,csa_tree_add_190_195_groupi_n_5132 ,csa_tree_add_190_195_groupi_n_4958);
  xnor csa_tree_add_190_195_groupi_g43044(csa_tree_add_190_195_groupi_n_6031 ,csa_tree_add_190_195_groupi_n_5089 ,csa_tree_add_190_195_groupi_n_1965);
  xor csa_tree_add_190_195_groupi_g43045(csa_tree_add_190_195_groupi_n_6030 ,csa_tree_add_190_195_groupi_n_4866 ,csa_tree_add_190_195_groupi_n_4710);
  xnor csa_tree_add_190_195_groupi_g43046(csa_tree_add_190_195_groupi_n_6029 ,csa_tree_add_190_195_groupi_n_5116 ,csa_tree_add_190_195_groupi_n_5032);
  xnor csa_tree_add_190_195_groupi_g43047(csa_tree_add_190_195_groupi_n_6028 ,csa_tree_add_190_195_groupi_n_5047 ,csa_tree_add_190_195_groupi_n_4937);
  xnor csa_tree_add_190_195_groupi_g43048(csa_tree_add_190_195_groupi_n_6027 ,csa_tree_add_190_195_groupi_n_5075 ,csa_tree_add_190_195_groupi_n_5152);
  xnor csa_tree_add_190_195_groupi_g43049(csa_tree_add_190_195_groupi_n_6026 ,csa_tree_add_190_195_groupi_n_4882 ,csa_tree_add_190_195_groupi_n_4883);
  xnor csa_tree_add_190_195_groupi_g43050(csa_tree_add_190_195_groupi_n_6025 ,csa_tree_add_190_195_groupi_n_4862 ,csa_tree_add_190_195_groupi_n_1293);
  xnor csa_tree_add_190_195_groupi_g43051(csa_tree_add_190_195_groupi_n_6024 ,csa_tree_add_190_195_groupi_n_5012 ,csa_tree_add_190_195_groupi_n_5142);
  xnor csa_tree_add_190_195_groupi_g43052(csa_tree_add_190_195_groupi_n_6023 ,csa_tree_add_190_195_groupi_n_4668 ,csa_tree_add_190_195_groupi_n_4647);
  xor csa_tree_add_190_195_groupi_g43053(csa_tree_add_190_195_groupi_n_6022 ,csa_tree_add_190_195_groupi_n_5135 ,csa_tree_add_190_195_groupi_n_4955);
  xnor csa_tree_add_190_195_groupi_g43055(csa_tree_add_190_195_groupi_n_6021 ,csa_tree_add_190_195_groupi_n_4644 ,csa_tree_add_190_195_groupi_n_4732);
  xnor csa_tree_add_190_195_groupi_g43056(csa_tree_add_190_195_groupi_n_6020 ,csa_tree_add_190_195_groupi_n_5099 ,csa_tree_add_190_195_groupi_n_5090);
  xnor csa_tree_add_190_195_groupi_g43057(csa_tree_add_190_195_groupi_n_6019 ,csa_tree_add_190_195_groupi_n_4638 ,csa_tree_add_190_195_groupi_n_4865);
  xnor csa_tree_add_190_195_groupi_g43058(csa_tree_add_190_195_groupi_n_6018 ,csa_tree_add_190_195_groupi_n_4812 ,csa_tree_add_190_195_groupi_n_4726);
  xnor csa_tree_add_190_195_groupi_g43059(csa_tree_add_190_195_groupi_n_6017 ,csa_tree_add_190_195_groupi_n_4887 ,csa_tree_add_190_195_groupi_n_1159);
  xor csa_tree_add_190_195_groupi_g43060(csa_tree_add_190_195_groupi_n_6016 ,csa_tree_add_190_195_groupi_n_4904 ,csa_tree_add_190_195_groupi_n_4816);
  xnor csa_tree_add_190_195_groupi_g43061(csa_tree_add_190_195_groupi_n_6015 ,csa_tree_add_190_195_groupi_n_4778 ,csa_tree_add_190_195_groupi_n_3693);
  xnor csa_tree_add_190_195_groupi_g43062(csa_tree_add_190_195_groupi_n_6014 ,csa_tree_add_190_195_groupi_n_5153 ,csa_tree_add_190_195_groupi_n_2153);
  xnor csa_tree_add_190_195_groupi_g43063(csa_tree_add_190_195_groupi_n_6013 ,csa_tree_add_190_195_groupi_n_4885 ,csa_tree_add_190_195_groupi_n_1354);
  xnor csa_tree_add_190_195_groupi_g43064(csa_tree_add_190_195_groupi_n_6012 ,csa_tree_add_190_195_groupi_n_4852 ,csa_tree_add_190_195_groupi_n_1903);
  xnor csa_tree_add_190_195_groupi_g43065(csa_tree_add_190_195_groupi_n_6011 ,csa_tree_add_190_195_groupi_n_4118 ,csa_tree_add_190_195_groupi_n_4834);
  xnor csa_tree_add_190_195_groupi_g43066(csa_tree_add_190_195_groupi_n_6010 ,csa_tree_add_190_195_groupi_n_4670 ,csa_tree_add_190_195_groupi_n_4781);
  xnor csa_tree_add_190_195_groupi_g43067(csa_tree_add_190_195_groupi_n_6009 ,csa_tree_add_190_195_groupi_n_4677 ,csa_tree_add_190_195_groupi_n_4840);
  xnor csa_tree_add_190_195_groupi_g43068(csa_tree_add_190_195_groupi_n_6008 ,csa_tree_add_190_195_groupi_n_4769 ,csa_tree_add_190_195_groupi_n_4890);
  xnor csa_tree_add_190_195_groupi_g43069(csa_tree_add_190_195_groupi_n_6007 ,csa_tree_add_190_195_groupi_n_4722 ,csa_tree_add_190_195_groupi_n_4939);
  xnor csa_tree_add_190_195_groupi_g43070(csa_tree_add_190_195_groupi_n_6006 ,csa_tree_add_190_195_groupi_n_5163 ,csa_tree_add_190_195_groupi_n_4894);
  xnor csa_tree_add_190_195_groupi_g43071(csa_tree_add_190_195_groupi_n_6005 ,csa_tree_add_190_195_groupi_n_5113 ,csa_tree_add_190_195_groupi_n_4964);
  xor csa_tree_add_190_195_groupi_g43072(csa_tree_add_190_195_groupi_n_6004 ,csa_tree_add_190_195_groupi_n_4886 ,csa_tree_add_190_195_groupi_n_5174);
  xnor csa_tree_add_190_195_groupi_g43073(csa_tree_add_190_195_groupi_n_6003 ,csa_tree_add_190_195_groupi_n_4702 ,csa_tree_add_190_195_groupi_n_1930);
  xnor csa_tree_add_190_195_groupi_g43074(csa_tree_add_190_195_groupi_n_6002 ,csa_tree_add_190_195_groupi_n_4646 ,csa_tree_add_190_195_groupi_n_4590);
  xnor csa_tree_add_190_195_groupi_g43075(csa_tree_add_190_195_groupi_n_6001 ,csa_tree_add_190_195_groupi_n_4715 ,csa_tree_add_190_195_groupi_n_895);
  xnor csa_tree_add_190_195_groupi_g43076(csa_tree_add_190_195_groupi_n_6000 ,csa_tree_add_190_195_groupi_n_3697 ,csa_tree_add_190_195_groupi_n_4851);
  xnor csa_tree_add_190_195_groupi_g43077(csa_tree_add_190_195_groupi_n_5999 ,csa_tree_add_190_195_groupi_n_4643 ,csa_tree_add_190_195_groupi_n_4691);
  xor csa_tree_add_190_195_groupi_g43078(csa_tree_add_190_195_groupi_n_5998 ,csa_tree_add_190_195_groupi_n_5115 ,csa_tree_add_190_195_groupi_n_5056);
  xnor csa_tree_add_190_195_groupi_g43079(csa_tree_add_190_195_groupi_n_5997 ,csa_tree_add_190_195_groupi_n_4688 ,csa_tree_add_190_195_groupi_n_4857);
  xnor csa_tree_add_190_195_groupi_g43080(csa_tree_add_190_195_groupi_n_5996 ,csa_tree_add_190_195_groupi_n_4793 ,csa_tree_add_190_195_groupi_n_4593);
  xnor csa_tree_add_190_195_groupi_g43081(csa_tree_add_190_195_groupi_n_5995 ,csa_tree_add_190_195_groupi_n_4744 ,csa_tree_add_190_195_groupi_n_4794);
  xnor csa_tree_add_190_195_groupi_g43082(csa_tree_add_190_195_groupi_n_5994 ,csa_tree_add_190_195_groupi_n_4756 ,csa_tree_add_190_195_groupi_n_4798);
  xnor csa_tree_add_190_195_groupi_g43083(csa_tree_add_190_195_groupi_n_5993 ,csa_tree_add_190_195_groupi_n_4986 ,csa_tree_add_190_195_groupi_n_5087);
  xnor csa_tree_add_190_195_groupi_g43084(csa_tree_add_190_195_groupi_n_5992 ,csa_tree_add_190_195_groupi_n_5137 ,csa_tree_add_190_195_groupi_n_1277);
  xnor csa_tree_add_190_195_groupi_g43085(csa_tree_add_190_195_groupi_n_5991 ,csa_tree_add_190_195_groupi_n_4117 ,csa_tree_add_190_195_groupi_n_4913);
  xnor csa_tree_add_190_195_groupi_g43086(csa_tree_add_190_195_groupi_n_5990 ,csa_tree_add_190_195_groupi_n_4776 ,csa_tree_add_190_195_groupi_n_4899);
  xnor csa_tree_add_190_195_groupi_g43087(csa_tree_add_190_195_groupi_n_5989 ,csa_tree_add_190_195_groupi_n_5018 ,csa_tree_add_190_195_groupi_n_4753);
  xnor csa_tree_add_190_195_groupi_g43088(csa_tree_add_190_195_groupi_n_5988 ,csa_tree_add_190_195_groupi_n_4861 ,csa_tree_add_190_195_groupi_n_976);
  xnor csa_tree_add_190_195_groupi_g43089(csa_tree_add_190_195_groupi_n_5987 ,csa_tree_add_190_195_groupi_n_4867 ,csa_tree_add_190_195_groupi_n_1751);
  xnor csa_tree_add_190_195_groupi_g43091(csa_tree_add_190_195_groupi_n_5986 ,csa_tree_add_190_195_groupi_n_4848 ,csa_tree_add_190_195_groupi_n_1988);
  xnor csa_tree_add_190_195_groupi_g43092(csa_tree_add_190_195_groupi_n_5985 ,csa_tree_add_190_195_groupi_n_4807 ,csa_tree_add_190_195_groupi_n_1760);
  xor csa_tree_add_190_195_groupi_g43093(csa_tree_add_190_195_groupi_n_5984 ,csa_tree_add_190_195_groupi_n_5101 ,csa_tree_add_190_195_groupi_n_4767);
  or csa_tree_add_190_195_groupi_g43094(csa_tree_add_190_195_groupi_n_6290 ,csa_tree_add_190_195_groupi_n_3180 ,csa_tree_add_190_195_groupi_n_5683);
  and csa_tree_add_190_195_groupi_g43095(csa_tree_add_190_195_groupi_n_6289 ,csa_tree_add_190_195_groupi_n_3353 ,csa_tree_add_190_195_groupi_n_5632);
  xnor csa_tree_add_190_195_groupi_g43096(csa_tree_add_190_195_groupi_n_6288 ,csa_tree_add_190_195_groupi_n_4574 ,csa_tree_add_190_195_groupi_n_2091);
  xnor csa_tree_add_190_195_groupi_g43097(csa_tree_add_190_195_groupi_n_6287 ,csa_tree_add_190_195_groupi_n_4575 ,csa_tree_add_190_195_groupi_n_592);
  or csa_tree_add_190_195_groupi_g43099(csa_tree_add_190_195_groupi_n_6285 ,csa_tree_add_190_195_groupi_n_4356 ,csa_tree_add_190_195_groupi_n_5778);
  or csa_tree_add_190_195_groupi_g43100(csa_tree_add_190_195_groupi_n_6283 ,csa_tree_add_190_195_groupi_n_3214 ,csa_tree_add_190_195_groupi_n_5681);
  and csa_tree_add_190_195_groupi_g43101(csa_tree_add_190_195_groupi_n_6282 ,csa_tree_add_190_195_groupi_n_4578 ,csa_tree_add_190_195_groupi_n_5625);
  and csa_tree_add_190_195_groupi_g43103(csa_tree_add_190_195_groupi_n_6281 ,csa_tree_add_190_195_groupi_n_2766 ,csa_tree_add_190_195_groupi_n_5648);
  xnor csa_tree_add_190_195_groupi_g43104(csa_tree_add_190_195_groupi_n_6280 ,csa_tree_add_190_195_groupi_n_5130 ,csa_tree_add_190_195_groupi_n_3881);
  xnor csa_tree_add_190_195_groupi_g43106(csa_tree_add_190_195_groupi_n_6278 ,csa_tree_add_190_195_groupi_n_4818 ,csa_tree_add_190_195_groupi_n_3813);
  xnor csa_tree_add_190_195_groupi_g43107(csa_tree_add_190_195_groupi_n_6276 ,csa_tree_add_190_195_groupi_n_3203 ,csa_tree_add_190_195_groupi_n_4849);
  xnor csa_tree_add_190_195_groupi_g43108(csa_tree_add_190_195_groupi_n_6275 ,csa_tree_add_190_195_groupi_n_5104 ,csa_tree_add_190_195_groupi_n_3936);
  xnor csa_tree_add_190_195_groupi_g43109(csa_tree_add_190_195_groupi_n_6274 ,csa_tree_add_190_195_groupi_n_5145 ,csa_tree_add_190_195_groupi_n_3882);
  xnor csa_tree_add_190_195_groupi_g43110(csa_tree_add_190_195_groupi_n_6272 ,csa_tree_add_190_195_groupi_n_4120 ,csa_tree_add_190_195_groupi_n_4856);
  or csa_tree_add_190_195_groupi_g43111(csa_tree_add_190_195_groupi_n_6270 ,csa_tree_add_190_195_groupi_n_4392 ,csa_tree_add_190_195_groupi_n_5680);
  or csa_tree_add_190_195_groupi_g43112(csa_tree_add_190_195_groupi_n_6269 ,csa_tree_add_190_195_groupi_n_2854 ,csa_tree_add_190_195_groupi_n_5823);
  xnor csa_tree_add_190_195_groupi_g43113(csa_tree_add_190_195_groupi_n_6267 ,csa_tree_add_190_195_groupi_n_5162 ,csa_tree_add_190_195_groupi_n_3895);
  or csa_tree_add_190_195_groupi_g43114(csa_tree_add_190_195_groupi_n_6266 ,csa_tree_add_190_195_groupi_n_3020 ,csa_tree_add_190_195_groupi_n_5806);
  xor csa_tree_add_190_195_groupi_g43115(csa_tree_add_190_195_groupi_n_6265 ,csa_tree_add_190_195_groupi_n_4797 ,csa_tree_add_190_195_groupi_n_3769);
  xnor csa_tree_add_190_195_groupi_g43116(csa_tree_add_190_195_groupi_n_6264 ,csa_tree_add_190_195_groupi_n_4842 ,csa_tree_add_190_195_groupi_n_4098);
  and csa_tree_add_190_195_groupi_g43117(csa_tree_add_190_195_groupi_n_6262 ,csa_tree_add_190_195_groupi_n_2977 ,csa_tree_add_190_195_groupi_n_5659);
  and csa_tree_add_190_195_groupi_g43118(csa_tree_add_190_195_groupi_n_6260 ,csa_tree_add_190_195_groupi_n_3629 ,csa_tree_add_190_195_groupi_n_5651);
  xnor csa_tree_add_190_195_groupi_g43119(csa_tree_add_190_195_groupi_n_6259 ,csa_tree_add_190_195_groupi_n_4830 ,csa_tree_add_190_195_groupi_n_3855);
  xnor csa_tree_add_190_195_groupi_g43120(csa_tree_add_190_195_groupi_n_6257 ,csa_tree_add_190_195_groupi_n_5141 ,csa_tree_add_190_195_groupi_n_3918);
  xnor csa_tree_add_190_195_groupi_g43121(csa_tree_add_190_195_groupi_n_6255 ,csa_tree_add_190_195_groupi_n_5118 ,csa_tree_add_190_195_groupi_n_4571);
  not csa_tree_add_190_195_groupi_g43123(csa_tree_add_190_195_groupi_n_5976 ,csa_tree_add_190_195_groupi_n_5975);
  not csa_tree_add_190_195_groupi_g43124(csa_tree_add_190_195_groupi_n_5974 ,csa_tree_add_190_195_groupi_n_5973);
  not csa_tree_add_190_195_groupi_g43125(csa_tree_add_190_195_groupi_n_5971 ,csa_tree_add_190_195_groupi_n_5970);
  not csa_tree_add_190_195_groupi_g43126(csa_tree_add_190_195_groupi_n_5963 ,csa_tree_add_190_195_groupi_n_5964);
  not csa_tree_add_190_195_groupi_g43127(csa_tree_add_190_195_groupi_n_5958 ,csa_tree_add_190_195_groupi_n_5959);
  not csa_tree_add_190_195_groupi_g43128(csa_tree_add_190_195_groupi_n_5956 ,csa_tree_add_190_195_groupi_n_5957);
  not csa_tree_add_190_195_groupi_g43129(csa_tree_add_190_195_groupi_n_5955 ,csa_tree_add_190_195_groupi_n_50);
  not csa_tree_add_190_195_groupi_g43130(csa_tree_add_190_195_groupi_n_5954 ,csa_tree_add_190_195_groupi_n_65);
  not csa_tree_add_190_195_groupi_g43131(csa_tree_add_190_195_groupi_n_5952 ,csa_tree_add_190_195_groupi_n_5953);
  not csa_tree_add_190_195_groupi_g43132(csa_tree_add_190_195_groupi_n_5950 ,csa_tree_add_190_195_groupi_n_5951);
  not csa_tree_add_190_195_groupi_g43133(csa_tree_add_190_195_groupi_n_5947 ,csa_tree_add_190_195_groupi_n_5948);
  not csa_tree_add_190_195_groupi_g43134(csa_tree_add_190_195_groupi_n_5945 ,csa_tree_add_190_195_groupi_n_5946);
  not csa_tree_add_190_195_groupi_g43135(csa_tree_add_190_195_groupi_n_5943 ,csa_tree_add_190_195_groupi_n_5944);
  not csa_tree_add_190_195_groupi_g43136(csa_tree_add_190_195_groupi_n_5941 ,csa_tree_add_190_195_groupi_n_5942);
  not csa_tree_add_190_195_groupi_g43137(csa_tree_add_190_195_groupi_n_5939 ,csa_tree_add_190_195_groupi_n_5940);
  not csa_tree_add_190_195_groupi_g43138(csa_tree_add_190_195_groupi_n_5936 ,csa_tree_add_190_195_groupi_n_5937);
  not csa_tree_add_190_195_groupi_g43139(csa_tree_add_190_195_groupi_n_5934 ,csa_tree_add_190_195_groupi_n_5935);
  not csa_tree_add_190_195_groupi_g43140(csa_tree_add_190_195_groupi_n_5933 ,csa_tree_add_190_195_groupi_n_5932);
  not csa_tree_add_190_195_groupi_g43141(csa_tree_add_190_195_groupi_n_5930 ,csa_tree_add_190_195_groupi_n_5931);
  not csa_tree_add_190_195_groupi_g43142(csa_tree_add_190_195_groupi_n_5927 ,csa_tree_add_190_195_groupi_n_5928);
  not csa_tree_add_190_195_groupi_g43143(csa_tree_add_190_195_groupi_n_5925 ,csa_tree_add_190_195_groupi_n_5926);
  not csa_tree_add_190_195_groupi_g43144(csa_tree_add_190_195_groupi_n_5923 ,csa_tree_add_190_195_groupi_n_5924);
  not csa_tree_add_190_195_groupi_g43145(csa_tree_add_190_195_groupi_n_5921 ,csa_tree_add_190_195_groupi_n_5922);
  not csa_tree_add_190_195_groupi_g43146(csa_tree_add_190_195_groupi_n_5919 ,csa_tree_add_190_195_groupi_n_5920);
  not csa_tree_add_190_195_groupi_g43148(csa_tree_add_190_195_groupi_n_5914 ,csa_tree_add_190_195_groupi_n_5915);
  not csa_tree_add_190_195_groupi_g43149(csa_tree_add_190_195_groupi_n_5913 ,csa_tree_add_190_195_groupi_n_53);
  not csa_tree_add_190_195_groupi_g43150(csa_tree_add_190_195_groupi_n_5911 ,csa_tree_add_190_195_groupi_n_5912);
  not csa_tree_add_190_195_groupi_g43151(csa_tree_add_190_195_groupi_n_5909 ,csa_tree_add_190_195_groupi_n_5910);
  not csa_tree_add_190_195_groupi_g43152(csa_tree_add_190_195_groupi_n_5906 ,csa_tree_add_190_195_groupi_n_5907);
  not csa_tree_add_190_195_groupi_g43154(csa_tree_add_190_195_groupi_n_5904 ,csa_tree_add_190_195_groupi_n_5905);
  not csa_tree_add_190_195_groupi_g43155(csa_tree_add_190_195_groupi_n_5901 ,csa_tree_add_190_195_groupi_n_5902);
  not csa_tree_add_190_195_groupi_g43157(csa_tree_add_190_195_groupi_n_5898 ,csa_tree_add_190_195_groupi_n_5899);
  not csa_tree_add_190_195_groupi_g43158(csa_tree_add_190_195_groupi_n_5897 ,csa_tree_add_190_195_groupi_n_31);
  not csa_tree_add_190_195_groupi_g43159(csa_tree_add_190_195_groupi_n_5893 ,csa_tree_add_190_195_groupi_n_5894);
  not csa_tree_add_190_195_groupi_g43160(csa_tree_add_190_195_groupi_n_5892 ,csa_tree_add_190_195_groupi_n_55);
  not csa_tree_add_190_195_groupi_g43161(csa_tree_add_190_195_groupi_n_5891 ,csa_tree_add_190_195_groupi_n_5890);
  not csa_tree_add_190_195_groupi_g43162(csa_tree_add_190_195_groupi_n_5886 ,csa_tree_add_190_195_groupi_n_5887);
  not csa_tree_add_190_195_groupi_g43163(csa_tree_add_190_195_groupi_n_5884 ,csa_tree_add_190_195_groupi_n_5885);
  not csa_tree_add_190_195_groupi_g43164(csa_tree_add_190_195_groupi_n_5882 ,csa_tree_add_190_195_groupi_n_5883);
  not csa_tree_add_190_195_groupi_g43165(csa_tree_add_190_195_groupi_n_5880 ,csa_tree_add_190_195_groupi_n_5881);
  not csa_tree_add_190_195_groupi_g43166(csa_tree_add_190_195_groupi_n_5878 ,csa_tree_add_190_195_groupi_n_5879);
  not csa_tree_add_190_195_groupi_g43167(csa_tree_add_190_195_groupi_n_5875 ,csa_tree_add_190_195_groupi_n_5874);
  not csa_tree_add_190_195_groupi_g43168(csa_tree_add_190_195_groupi_n_5871 ,csa_tree_add_190_195_groupi_n_5872);
  not csa_tree_add_190_195_groupi_g43169(csa_tree_add_190_195_groupi_n_5870 ,csa_tree_add_190_195_groupi_n_5869);
  not csa_tree_add_190_195_groupi_g43170(csa_tree_add_190_195_groupi_n_5867 ,csa_tree_add_190_195_groupi_n_5868);
  or csa_tree_add_190_195_groupi_g43171(csa_tree_add_190_195_groupi_n_5866 ,csa_tree_add_190_195_groupi_n_4582 ,csa_tree_add_190_195_groupi_n_5001);
  or csa_tree_add_190_195_groupi_g43172(csa_tree_add_190_195_groupi_n_5865 ,csa_tree_add_190_195_groupi_n_1944 ,csa_tree_add_190_195_groupi_n_4940);
  or csa_tree_add_190_195_groupi_g43173(csa_tree_add_190_195_groupi_n_5864 ,csa_tree_add_190_195_groupi_n_2721 ,csa_tree_add_190_195_groupi_n_5045);
  or csa_tree_add_190_195_groupi_g43174(csa_tree_add_190_195_groupi_n_5863 ,csa_tree_add_190_195_groupi_n_1849 ,csa_tree_add_190_195_groupi_n_5052);
  nor csa_tree_add_190_195_groupi_g43175(csa_tree_add_190_195_groupi_n_5862 ,csa_tree_add_190_195_groupi_n_2535 ,csa_tree_add_190_195_groupi_n_4758);
  and csa_tree_add_190_195_groupi_g43176(csa_tree_add_190_195_groupi_n_5861 ,csa_tree_add_190_195_groupi_n_2535 ,csa_tree_add_190_195_groupi_n_4758);
  nor csa_tree_add_190_195_groupi_g43177(csa_tree_add_190_195_groupi_n_5860 ,csa_tree_add_190_195_groupi_n_2690 ,csa_tree_add_190_195_groupi_n_4941);
  nor csa_tree_add_190_195_groupi_g43178(csa_tree_add_190_195_groupi_n_5859 ,in56[11] ,csa_tree_add_190_195_groupi_n_5044);
  nor csa_tree_add_190_195_groupi_g43179(csa_tree_add_190_195_groupi_n_5858 ,csa_tree_add_190_195_groupi_n_2527 ,csa_tree_add_190_195_groupi_n_5071);
  or csa_tree_add_190_195_groupi_g43180(csa_tree_add_190_195_groupi_n_5857 ,csa_tree_add_190_195_groupi_n_1812 ,csa_tree_add_190_195_groupi_n_5070);
  nor csa_tree_add_190_195_groupi_g43181(csa_tree_add_190_195_groupi_n_5856 ,in56[9] ,csa_tree_add_190_195_groupi_n_5063);
  or csa_tree_add_190_195_groupi_g43182(csa_tree_add_190_195_groupi_n_5855 ,csa_tree_add_190_195_groupi_n_2556 ,csa_tree_add_190_195_groupi_n_5064);
  or csa_tree_add_190_195_groupi_g43183(csa_tree_add_190_195_groupi_n_5854 ,in56[10] ,csa_tree_add_190_195_groupi_n_4947);
  nor csa_tree_add_190_195_groupi_g43184(csa_tree_add_190_195_groupi_n_5853 ,csa_tree_add_190_195_groupi_n_2563 ,csa_tree_add_190_195_groupi_n_4948);
  or csa_tree_add_190_195_groupi_g43185(csa_tree_add_190_195_groupi_n_5852 ,csa_tree_add_190_195_groupi_n_1817 ,csa_tree_add_190_195_groupi_n_4766);
  nor csa_tree_add_190_195_groupi_g43186(csa_tree_add_190_195_groupi_n_5851 ,csa_tree_add_190_195_groupi_n_2674 ,csa_tree_add_190_195_groupi_n_4767);
  nor csa_tree_add_190_195_groupi_g43187(csa_tree_add_190_195_groupi_n_5850 ,csa_tree_add_190_195_groupi_n_2648 ,csa_tree_add_190_195_groupi_n_4967);
  and csa_tree_add_190_195_groupi_g43188(csa_tree_add_190_195_groupi_n_5849 ,csa_tree_add_190_195_groupi_n_1390 ,csa_tree_add_190_195_groupi_n_4967);
  nor csa_tree_add_190_195_groupi_g43189(csa_tree_add_190_195_groupi_n_5848 ,csa_tree_add_190_195_groupi_n_1546 ,csa_tree_add_190_195_groupi_n_4917);
  and csa_tree_add_190_195_groupi_g43190(csa_tree_add_190_195_groupi_n_5847 ,csa_tree_add_190_195_groupi_n_731 ,csa_tree_add_190_195_groupi_n_4917);
  nor csa_tree_add_190_195_groupi_g43191(csa_tree_add_190_195_groupi_n_5846 ,csa_tree_add_190_195_groupi_n_4689 ,csa_tree_add_190_195_groupi_n_4881);
  nor csa_tree_add_190_195_groupi_g43192(csa_tree_add_190_195_groupi_n_5845 ,csa_tree_add_190_195_groupi_n_4882 ,csa_tree_add_190_195_groupi_n_4883);
  and csa_tree_add_190_195_groupi_g43193(csa_tree_add_190_195_groupi_n_5844 ,csa_tree_add_190_195_groupi_n_4897 ,csa_tree_add_190_195_groupi_n_4916);
  and csa_tree_add_190_195_groupi_g43194(csa_tree_add_190_195_groupi_n_5843 ,csa_tree_add_190_195_groupi_n_2726 ,csa_tree_add_190_195_groupi_n_4739);
  nor csa_tree_add_190_195_groupi_g43195(csa_tree_add_190_195_groupi_n_5842 ,csa_tree_add_190_195_groupi_n_4989 ,csa_tree_add_190_195_groupi_n_4907);
  or csa_tree_add_190_195_groupi_g43196(csa_tree_add_190_195_groupi_n_5841 ,csa_tree_add_190_195_groupi_n_2683 ,csa_tree_add_190_195_groupi_n_4995);
  or csa_tree_add_190_195_groupi_g43197(csa_tree_add_190_195_groupi_n_5840 ,csa_tree_add_190_195_groupi_n_4775 ,csa_tree_add_190_195_groupi_n_4772);
  and csa_tree_add_190_195_groupi_g43198(csa_tree_add_190_195_groupi_n_5839 ,csa_tree_add_190_195_groupi_n_4989 ,csa_tree_add_190_195_groupi_n_4907);
  and csa_tree_add_190_195_groupi_g43199(csa_tree_add_190_195_groupi_n_5838 ,csa_tree_add_190_195_groupi_n_1673 ,csa_tree_add_190_195_groupi_n_4908);
  or csa_tree_add_190_195_groupi_g43200(csa_tree_add_190_195_groupi_n_5837 ,csa_tree_add_190_195_groupi_n_1673 ,csa_tree_add_190_195_groupi_n_4908);
  or csa_tree_add_190_195_groupi_g43201(csa_tree_add_190_195_groupi_n_5836 ,csa_tree_add_190_195_groupi_n_4776 ,csa_tree_add_190_195_groupi_n_4899);
  or csa_tree_add_190_195_groupi_g43202(csa_tree_add_190_195_groupi_n_5835 ,csa_tree_add_190_195_groupi_n_4562 ,csa_tree_add_190_195_groupi_n_4741);
  or csa_tree_add_190_195_groupi_g43203(csa_tree_add_190_195_groupi_n_5834 ,csa_tree_add_190_195_groupi_n_4897 ,csa_tree_add_190_195_groupi_n_4916);
  and csa_tree_add_190_195_groupi_g43204(csa_tree_add_190_195_groupi_n_5833 ,csa_tree_add_190_195_groupi_n_4322 ,csa_tree_add_190_195_groupi_n_4851);
  or csa_tree_add_190_195_groupi_g43205(csa_tree_add_190_195_groupi_n_5832 ,csa_tree_add_190_195_groupi_n_2532 ,csa_tree_add_190_195_groupi_n_5030);
  nor csa_tree_add_190_195_groupi_g43206(csa_tree_add_190_195_groupi_n_5831 ,csa_tree_add_190_195_groupi_n_1945 ,csa_tree_add_190_195_groupi_n_5031);
  or csa_tree_add_190_195_groupi_g43207(csa_tree_add_190_195_groupi_n_5830 ,csa_tree_add_190_195_groupi_n_4195 ,csa_tree_add_190_195_groupi_n_5154);
  or csa_tree_add_190_195_groupi_g43208(csa_tree_add_190_195_groupi_n_5829 ,csa_tree_add_190_195_groupi_n_5048 ,csa_tree_add_190_195_groupi_n_4945);
  nor csa_tree_add_190_195_groupi_g43209(csa_tree_add_190_195_groupi_n_5828 ,csa_tree_add_190_195_groupi_n_2827 ,csa_tree_add_190_195_groupi_n_5141);
  nor csa_tree_add_190_195_groupi_g43210(csa_tree_add_190_195_groupi_n_5827 ,csa_tree_add_190_195_groupi_n_5049 ,csa_tree_add_190_195_groupi_n_4946);
  and csa_tree_add_190_195_groupi_g43211(csa_tree_add_190_195_groupi_n_5826 ,csa_tree_add_190_195_groupi_n_607 ,csa_tree_add_190_195_groupi_n_4955);
  nor csa_tree_add_190_195_groupi_g43212(csa_tree_add_190_195_groupi_n_5825 ,csa_tree_add_190_195_groupi_n_425 ,csa_tree_add_190_195_groupi_n_4955);
  nor csa_tree_add_190_195_groupi_g43213(csa_tree_add_190_195_groupi_n_5824 ,csa_tree_add_190_195_groupi_n_4880 ,csa_tree_add_190_195_groupi_n_4958);
  and csa_tree_add_190_195_groupi_g43214(csa_tree_add_190_195_groupi_n_5823 ,csa_tree_add_190_195_groupi_n_3611 ,csa_tree_add_190_195_groupi_n_4815);
  nor csa_tree_add_190_195_groupi_g43215(csa_tree_add_190_195_groupi_n_5822 ,csa_tree_add_190_195_groupi_n_2394 ,csa_tree_add_190_195_groupi_n_4896);
  nor csa_tree_add_190_195_groupi_g43216(csa_tree_add_190_195_groupi_n_5821 ,csa_tree_add_190_195_groupi_n_4903 ,csa_tree_add_190_195_groupi_n_4780);
  and csa_tree_add_190_195_groupi_g43217(csa_tree_add_190_195_groupi_n_5820 ,csa_tree_add_190_195_groupi_n_4880 ,csa_tree_add_190_195_groupi_n_4958);
  nor csa_tree_add_190_195_groupi_g43218(csa_tree_add_190_195_groupi_n_5819 ,csa_tree_add_190_195_groupi_n_4728 ,csa_tree_add_190_195_groupi_n_4687);
  nor csa_tree_add_190_195_groupi_g43219(csa_tree_add_190_195_groupi_n_5818 ,csa_tree_add_190_195_groupi_n_4973 ,csa_tree_add_190_195_groupi_n_4970);
  or csa_tree_add_190_195_groupi_g43220(csa_tree_add_190_195_groupi_n_5817 ,csa_tree_add_190_195_groupi_n_4975 ,csa_tree_add_190_195_groupi_n_4703);
  or csa_tree_add_190_195_groupi_g43221(csa_tree_add_190_195_groupi_n_5816 ,csa_tree_add_190_195_groupi_n_4723 ,csa_tree_add_190_195_groupi_n_4631);
  or csa_tree_add_190_195_groupi_g43222(csa_tree_add_190_195_groupi_n_5815 ,csa_tree_add_190_195_groupi_n_4606 ,csa_tree_add_190_195_groupi_n_4600);
  and csa_tree_add_190_195_groupi_g43223(csa_tree_add_190_195_groupi_n_5814 ,csa_tree_add_190_195_groupi_n_1041 ,csa_tree_add_190_195_groupi_n_5005);
  nor csa_tree_add_190_195_groupi_g43224(csa_tree_add_190_195_groupi_n_5813 ,csa_tree_add_190_195_groupi_n_1501 ,csa_tree_add_190_195_groupi_n_5089);
  nor csa_tree_add_190_195_groupi_g43225(csa_tree_add_190_195_groupi_n_5812 ,csa_tree_add_190_195_groupi_n_1041 ,csa_tree_add_190_195_groupi_n_5005);
  nor csa_tree_add_190_195_groupi_g43226(csa_tree_add_190_195_groupi_n_5811 ,csa_tree_add_190_195_groupi_n_4774 ,csa_tree_add_190_195_groupi_n_4773);
  or csa_tree_add_190_195_groupi_g43227(csa_tree_add_190_195_groupi_n_5810 ,csa_tree_add_190_195_groupi_n_5013 ,csa_tree_add_190_195_groupi_n_5029);
  nor csa_tree_add_190_195_groupi_g43228(csa_tree_add_190_195_groupi_n_5809 ,csa_tree_add_190_195_groupi_n_4729 ,csa_tree_add_190_195_groupi_n_5065);
  nor csa_tree_add_190_195_groupi_g43229(csa_tree_add_190_195_groupi_n_5808 ,csa_tree_add_190_195_groupi_n_5014 ,csa_tree_add_190_195_groupi_n_5028);
  and csa_tree_add_190_195_groupi_g43230(csa_tree_add_190_195_groupi_n_5807 ,csa_tree_add_190_195_groupi_n_4751 ,csa_tree_add_190_195_groupi_n_4894);
  nor csa_tree_add_190_195_groupi_g43231(csa_tree_add_190_195_groupi_n_5806 ,csa_tree_add_190_195_groupi_n_2838 ,csa_tree_add_190_195_groupi_n_5106);
  or csa_tree_add_190_195_groupi_g43232(csa_tree_add_190_195_groupi_n_5805 ,csa_tree_add_190_195_groupi_n_1438 ,csa_tree_add_190_195_groupi_n_5010);
  nor csa_tree_add_190_195_groupi_g43233(csa_tree_add_190_195_groupi_n_5804 ,csa_tree_add_190_195_groupi_n_2153 ,csa_tree_add_190_195_groupi_n_5011);
  nor csa_tree_add_190_195_groupi_g43234(csa_tree_add_190_195_groupi_n_5803 ,csa_tree_add_190_195_groupi_n_5042 ,csa_tree_add_190_195_groupi_n_5077);
  nor csa_tree_add_190_195_groupi_g43235(csa_tree_add_190_195_groupi_n_5802 ,csa_tree_add_190_195_groupi_n_4607 ,csa_tree_add_190_195_groupi_n_4601);
  or csa_tree_add_190_195_groupi_g43236(csa_tree_add_190_195_groupi_n_5801 ,csa_tree_add_190_195_groupi_n_5096 ,csa_tree_add_190_195_groupi_n_4923);
  nor csa_tree_add_190_195_groupi_g43237(csa_tree_add_190_195_groupi_n_5800 ,csa_tree_add_190_195_groupi_n_5081 ,csa_tree_add_190_195_groupi_n_5092);
  or csa_tree_add_190_195_groupi_g43238(csa_tree_add_190_195_groupi_n_5799 ,csa_tree_add_190_195_groupi_n_1351 ,csa_tree_add_190_195_groupi_n_4895);
  or csa_tree_add_190_195_groupi_g43239(csa_tree_add_190_195_groupi_n_5798 ,csa_tree_add_190_195_groupi_n_4645 ,csa_tree_add_190_195_groupi_n_4590);
  and csa_tree_add_190_195_groupi_g43240(csa_tree_add_190_195_groupi_n_5797 ,csa_tree_add_190_195_groupi_n_3368 ,csa_tree_add_190_195_groupi_n_5137);
  nor csa_tree_add_190_195_groupi_g43241(csa_tree_add_190_195_groupi_n_5796 ,csa_tree_add_190_195_groupi_n_4771 ,csa_tree_add_190_195_groupi_n_4930);
  or csa_tree_add_190_195_groupi_g43242(csa_tree_add_190_195_groupi_n_5795 ,csa_tree_add_190_195_groupi_n_5082 ,csa_tree_add_190_195_groupi_n_5091);
  nor csa_tree_add_190_195_groupi_g43243(csa_tree_add_190_195_groupi_n_5794 ,csa_tree_add_190_195_groupi_n_4656 ,csa_tree_add_190_195_groupi_n_4791);
  or csa_tree_add_190_195_groupi_g43244(csa_tree_add_190_195_groupi_n_5793 ,csa_tree_add_190_195_groupi_n_4986 ,csa_tree_add_190_195_groupi_n_5087);
  or csa_tree_add_190_195_groupi_g43245(csa_tree_add_190_195_groupi_n_5792 ,csa_tree_add_190_195_groupi_n_4594 ,csa_tree_add_190_195_groupi_n_5083);
  nor csa_tree_add_190_195_groupi_g43246(csa_tree_add_190_195_groupi_n_5791 ,csa_tree_add_190_195_groupi_n_4595 ,csa_tree_add_190_195_groupi_n_5084);
  and csa_tree_add_190_195_groupi_g43247(csa_tree_add_190_195_groupi_n_5790 ,csa_tree_add_190_195_groupi_n_3625 ,csa_tree_add_190_195_groupi_n_5104);
  or csa_tree_add_190_195_groupi_g43248(csa_tree_add_190_195_groupi_n_5789 ,csa_tree_add_190_195_groupi_n_2498 ,csa_tree_add_190_195_groupi_n_5066);
  nor csa_tree_add_190_195_groupi_g43249(csa_tree_add_190_195_groupi_n_5788 ,csa_tree_add_190_195_groupi_n_792 ,csa_tree_add_190_195_groupi_n_5067);
  nor csa_tree_add_190_195_groupi_g43250(csa_tree_add_190_195_groupi_n_5787 ,csa_tree_add_190_195_groupi_n_1961 ,csa_tree_add_190_195_groupi_n_4642);
  or csa_tree_add_190_195_groupi_g43251(csa_tree_add_190_195_groupi_n_5786 ,csa_tree_add_190_195_groupi_n_4699 ,csa_tree_add_190_195_groupi_n_4624);
  or csa_tree_add_190_195_groupi_g43252(csa_tree_add_190_195_groupi_n_5785 ,csa_tree_add_190_195_groupi_n_4709 ,csa_tree_add_190_195_groupi_n_4629);
  or csa_tree_add_190_195_groupi_g43253(csa_tree_add_190_195_groupi_n_5784 ,csa_tree_add_190_195_groupi_n_5043 ,csa_tree_add_190_195_groupi_n_5076);
  or csa_tree_add_190_195_groupi_g43254(csa_tree_add_190_195_groupi_n_5783 ,csa_tree_add_190_195_groupi_n_1811 ,csa_tree_add_190_195_groupi_n_5004);
  or csa_tree_add_190_195_groupi_g43255(csa_tree_add_190_195_groupi_n_5782 ,csa_tree_add_190_195_groupi_n_4637 ,csa_tree_add_190_195_groupi_n_4636);
  and csa_tree_add_190_195_groupi_g43256(csa_tree_add_190_195_groupi_n_5781 ,csa_tree_add_190_195_groupi_n_1811 ,csa_tree_add_190_195_groupi_n_5004);
  or csa_tree_add_190_195_groupi_g43257(csa_tree_add_190_195_groupi_n_5780 ,csa_tree_add_190_195_groupi_n_723 ,csa_tree_add_190_195_groupi_n_5032);
  and csa_tree_add_190_195_groupi_g43258(csa_tree_add_190_195_groupi_n_5779 ,csa_tree_add_190_195_groupi_n_723 ,csa_tree_add_190_195_groupi_n_5032);
  and csa_tree_add_190_195_groupi_g43259(csa_tree_add_190_195_groupi_n_5778 ,csa_tree_add_190_195_groupi_n_4354 ,csa_tree_add_190_195_groupi_n_5118);
  or csa_tree_add_190_195_groupi_g43260(csa_tree_add_190_195_groupi_n_5777 ,csa_tree_add_190_195_groupi_n_243 ,csa_tree_add_190_195_groupi_n_4715);
  nor csa_tree_add_190_195_groupi_g43261(csa_tree_add_190_195_groupi_n_5776 ,csa_tree_add_190_195_groupi_n_5000 ,csa_tree_add_190_195_groupi_n_4893);
  and csa_tree_add_190_195_groupi_g43262(csa_tree_add_190_195_groupi_n_5775 ,csa_tree_add_190_195_groupi_n_4668 ,csa_tree_add_190_195_groupi_n_4647);
  and csa_tree_add_190_195_groupi_g43263(csa_tree_add_190_195_groupi_n_5774 ,csa_tree_add_190_195_groupi_n_5000 ,csa_tree_add_190_195_groupi_n_4893);
  or csa_tree_add_190_195_groupi_g43264(csa_tree_add_190_195_groupi_n_5773 ,csa_tree_add_190_195_groupi_n_4997 ,csa_tree_add_190_195_groupi_n_4993);
  or csa_tree_add_190_195_groupi_g43265(csa_tree_add_190_195_groupi_n_5772 ,csa_tree_add_190_195_groupi_n_4395 ,csa_tree_add_190_195_groupi_n_5159);
  nor csa_tree_add_190_195_groupi_g43266(csa_tree_add_190_195_groupi_n_5771 ,csa_tree_add_190_195_groupi_n_4998 ,csa_tree_add_190_195_groupi_n_4994);
  and csa_tree_add_190_195_groupi_g43267(csa_tree_add_190_195_groupi_n_5770 ,csa_tree_add_190_195_groupi_n_4986 ,csa_tree_add_190_195_groupi_n_5087);
  nor csa_tree_add_190_195_groupi_g43268(csa_tree_add_190_195_groupi_n_5769 ,csa_tree_add_190_195_groupi_n_1848 ,csa_tree_add_190_195_groupi_n_4985);
  or csa_tree_add_190_195_groupi_g43269(csa_tree_add_190_195_groupi_n_5768 ,csa_tree_add_190_195_groupi_n_2688 ,csa_tree_add_190_195_groupi_n_4984);
  or csa_tree_add_190_195_groupi_g43270(csa_tree_add_190_195_groupi_n_5767 ,csa_tree_add_190_195_groupi_n_5006 ,csa_tree_add_190_195_groupi_n_4796);
  and csa_tree_add_190_195_groupi_g43271(csa_tree_add_190_195_groupi_n_5766 ,csa_tree_add_190_195_groupi_n_4744 ,csa_tree_add_190_195_groupi_n_4794);
  nor csa_tree_add_190_195_groupi_g43272(csa_tree_add_190_195_groupi_n_5765 ,csa_tree_add_190_195_groupi_n_3107 ,csa_tree_add_190_195_groupi_n_5130);
  or csa_tree_add_190_195_groupi_g43273(csa_tree_add_190_195_groupi_n_5764 ,csa_tree_add_190_195_groupi_n_4744 ,csa_tree_add_190_195_groupi_n_4794);
  or csa_tree_add_190_195_groupi_g43274(csa_tree_add_190_195_groupi_n_5763 ,csa_tree_add_190_195_groupi_n_942 ,csa_tree_add_190_195_groupi_n_4585);
  nor csa_tree_add_190_195_groupi_g43275(csa_tree_add_190_195_groupi_n_5762 ,csa_tree_add_190_195_groupi_n_2465 ,csa_tree_add_190_195_groupi_n_4586);
  and csa_tree_add_190_195_groupi_g43276(csa_tree_add_190_195_groupi_n_5761 ,csa_tree_add_190_195_groupi_n_3367 ,csa_tree_add_190_195_groupi_n_5133);
  nor csa_tree_add_190_195_groupi_g43277(csa_tree_add_190_195_groupi_n_5760 ,csa_tree_add_190_195_groupi_n_4724 ,csa_tree_add_190_195_groupi_n_4632);
  nor csa_tree_add_190_195_groupi_g43278(csa_tree_add_190_195_groupi_n_5759 ,csa_tree_add_190_195_groupi_n_4718 ,csa_tree_add_190_195_groupi_n_4983);
  nor csa_tree_add_190_195_groupi_g43279(csa_tree_add_190_195_groupi_n_5758 ,csa_tree_add_190_195_groupi_n_4673 ,csa_tree_add_190_195_groupi_n_5054);
  or csa_tree_add_190_195_groupi_g43280(csa_tree_add_190_195_groupi_n_5757 ,csa_tree_add_190_195_groupi_n_3038 ,csa_tree_add_190_195_groupi_n_5140);
  and csa_tree_add_190_195_groupi_g43281(csa_tree_add_190_195_groupi_n_5756 ,csa_tree_add_190_195_groupi_n_1200 ,csa_tree_add_190_195_groupi_n_4715);
  or csa_tree_add_190_195_groupi_g43282(csa_tree_add_190_195_groupi_n_5755 ,csa_tree_add_190_195_groupi_n_4770 ,csa_tree_add_190_195_groupi_n_4929);
  or csa_tree_add_190_195_groupi_g43283(csa_tree_add_190_195_groupi_n_5754 ,csa_tree_add_190_195_groupi_n_2084 ,csa_tree_add_190_195_groupi_n_5012);
  and csa_tree_add_190_195_groupi_g43284(csa_tree_add_190_195_groupi_n_5753 ,csa_tree_add_190_195_groupi_n_2084 ,csa_tree_add_190_195_groupi_n_5012);
  or csa_tree_add_190_195_groupi_g43285(csa_tree_add_190_195_groupi_n_5752 ,csa_tree_add_190_195_groupi_n_2215 ,csa_tree_add_190_195_groupi_n_4928);
  and csa_tree_add_190_195_groupi_g43286(csa_tree_add_190_195_groupi_n_5751 ,csa_tree_add_190_195_groupi_n_2215 ,csa_tree_add_190_195_groupi_n_4928);
  or csa_tree_add_190_195_groupi_g43287(csa_tree_add_190_195_groupi_n_5750 ,csa_tree_add_190_195_groupi_n_4792 ,csa_tree_add_190_195_groupi_n_4592);
  or csa_tree_add_190_195_groupi_g43288(csa_tree_add_190_195_groupi_n_5749 ,csa_tree_add_190_195_groupi_n_4968 ,csa_tree_add_190_195_groupi_n_4943);
  nor csa_tree_add_190_195_groupi_g43289(csa_tree_add_190_195_groupi_n_5748 ,csa_tree_add_190_195_groupi_n_4588 ,csa_tree_add_190_195_groupi_n_5075);
  or csa_tree_add_190_195_groupi_g43290(csa_tree_add_190_195_groupi_n_5747 ,csa_tree_add_190_195_groupi_n_4902 ,csa_tree_add_190_195_groupi_n_4779);
  nor csa_tree_add_190_195_groupi_g43291(csa_tree_add_190_195_groupi_n_5746 ,csa_tree_add_190_195_groupi_n_4793 ,csa_tree_add_190_195_groupi_n_4593);
  and csa_tree_add_190_195_groupi_g43292(csa_tree_add_190_195_groupi_n_5745 ,csa_tree_add_190_195_groupi_n_2775 ,csa_tree_add_190_195_groupi_n_5145);
  nor csa_tree_add_190_195_groupi_g43293(csa_tree_add_190_195_groupi_n_5744 ,csa_tree_add_190_195_groupi_n_4969 ,csa_tree_add_190_195_groupi_n_4942);
  nor csa_tree_add_190_195_groupi_g43294(csa_tree_add_190_195_groupi_n_5743 ,csa_tree_add_190_195_groupi_n_5095 ,csa_tree_add_190_195_groupi_n_4924);
  nor csa_tree_add_190_195_groupi_g43295(csa_tree_add_190_195_groupi_n_5742 ,csa_tree_add_190_195_groupi_n_4751 ,csa_tree_add_190_195_groupi_n_4894);
  and csa_tree_add_190_195_groupi_g43296(csa_tree_add_190_195_groupi_n_5741 ,csa_tree_add_190_195_groupi_n_4882 ,csa_tree_add_190_195_groupi_n_4883);
  and csa_tree_add_190_195_groupi_g43297(csa_tree_add_190_195_groupi_n_5740 ,csa_tree_add_190_195_groupi_n_4697 ,csa_tree_add_190_195_groupi_n_4757);
  nor csa_tree_add_190_195_groupi_g43298(csa_tree_add_190_195_groupi_n_5739 ,csa_tree_add_190_195_groupi_n_4603 ,csa_tree_add_190_195_groupi_n_4961);
  and csa_tree_add_190_195_groupi_g43299(csa_tree_add_190_195_groupi_n_5738 ,csa_tree_add_190_195_groupi_n_5017 ,csa_tree_add_190_195_groupi_n_4944);
  nor csa_tree_add_190_195_groupi_g43300(csa_tree_add_190_195_groupi_n_5737 ,csa_tree_add_190_195_groupi_n_4117 ,csa_tree_add_190_195_groupi_n_4913);
  nor csa_tree_add_190_195_groupi_g43301(csa_tree_add_190_195_groupi_n_5736 ,csa_tree_add_190_195_groupi_n_4692 ,csa_tree_add_190_195_groupi_n_4685);
  nor csa_tree_add_190_195_groupi_g43302(csa_tree_add_190_195_groupi_n_5735 ,csa_tree_add_190_195_groupi_n_4974 ,csa_tree_add_190_195_groupi_n_4704);
  nor csa_tree_add_190_195_groupi_g43303(csa_tree_add_190_195_groupi_n_5734 ,csa_tree_add_190_195_groupi_n_713 ,csa_tree_add_190_195_groupi_n_5090);
  and csa_tree_add_190_195_groupi_g43304(csa_tree_add_190_195_groupi_n_5733 ,csa_tree_add_190_195_groupi_n_712 ,csa_tree_add_190_195_groupi_n_5090);
  or csa_tree_add_190_195_groupi_g43305(csa_tree_add_190_195_groupi_n_5732 ,csa_tree_add_190_195_groupi_n_3402 ,csa_tree_add_190_195_groupi_n_5172);
  nor csa_tree_add_190_195_groupi_g43306(csa_tree_add_190_195_groupi_n_5731 ,csa_tree_add_190_195_groupi_n_2872 ,csa_tree_add_190_195_groupi_n_5162);
  nor csa_tree_add_190_195_groupi_g43307(csa_tree_add_190_195_groupi_n_5730 ,csa_tree_add_190_195_groupi_n_4755 ,csa_tree_add_190_195_groupi_n_4713);
  or csa_tree_add_190_195_groupi_g43308(csa_tree_add_190_195_groupi_n_5729 ,csa_tree_add_190_195_groupi_n_4657 ,csa_tree_add_190_195_groupi_n_4790);
  nor csa_tree_add_190_195_groupi_g43309(csa_tree_add_190_195_groupi_n_5728 ,csa_tree_add_190_195_groupi_n_4698 ,csa_tree_add_190_195_groupi_n_4625);
  and csa_tree_add_190_195_groupi_g43310(csa_tree_add_190_195_groupi_n_5727 ,csa_tree_add_190_195_groupi_n_4776 ,csa_tree_add_190_195_groupi_n_4899);
  or csa_tree_add_190_195_groupi_g43311(csa_tree_add_190_195_groupi_n_5726 ,csa_tree_add_190_195_groupi_n_4652 ,csa_tree_add_190_195_groupi_n_5008);
  nor csa_tree_add_190_195_groupi_g43312(csa_tree_add_190_195_groupi_n_5725 ,csa_tree_add_190_195_groupi_n_5017 ,csa_tree_add_190_195_groupi_n_4944);
  or csa_tree_add_190_195_groupi_g43313(csa_tree_add_190_195_groupi_n_5724 ,csa_tree_add_190_195_groupi_n_5018 ,csa_tree_add_190_195_groupi_n_4753);
  and csa_tree_add_190_195_groupi_g43314(csa_tree_add_190_195_groupi_n_5723 ,csa_tree_add_190_195_groupi_n_4644 ,csa_tree_add_190_195_groupi_n_4732);
  or csa_tree_add_190_195_groupi_g43315(csa_tree_add_190_195_groupi_n_5722 ,csa_tree_add_190_195_groupi_n_4644 ,csa_tree_add_190_195_groupi_n_4732);
  or csa_tree_add_190_195_groupi_g43316(csa_tree_add_190_195_groupi_n_5721 ,csa_tree_add_190_195_groupi_n_2462 ,csa_tree_add_190_195_groupi_n_4641);
  nor csa_tree_add_190_195_groupi_g43317(csa_tree_add_190_195_groupi_n_5720 ,csa_tree_add_190_195_groupi_n_4697 ,csa_tree_add_190_195_groupi_n_4757);
  and csa_tree_add_190_195_groupi_g43318(csa_tree_add_190_195_groupi_n_5719 ,csa_tree_add_190_195_groupi_n_2855 ,csa_tree_add_190_195_groupi_n_4797);
  or csa_tree_add_190_195_groupi_g43319(csa_tree_add_190_195_groupi_n_5718 ,csa_tree_add_190_195_groupi_n_2789 ,csa_tree_add_190_195_groupi_n_4868);
  or csa_tree_add_190_195_groupi_g43320(csa_tree_add_190_195_groupi_n_5717 ,csa_tree_add_190_195_groupi_n_4910 ,csa_tree_add_190_195_groupi_n_4598);
  nor csa_tree_add_190_195_groupi_g43321(csa_tree_add_190_195_groupi_n_5716 ,csa_tree_add_190_195_groupi_n_4638 ,csa_tree_add_190_195_groupi_n_4635);
  and csa_tree_add_190_195_groupi_g43322(csa_tree_add_190_195_groupi_n_5715 ,csa_tree_add_190_195_groupi_n_4716 ,csa_tree_add_190_195_groupi_n_5039);
  nor csa_tree_add_190_195_groupi_g43323(csa_tree_add_190_195_groupi_n_5714 ,csa_tree_add_190_195_groupi_n_4747 ,csa_tree_add_190_195_groupi_n_4743);
  and csa_tree_add_190_195_groupi_g43324(csa_tree_add_190_195_groupi_n_5713 ,csa_tree_add_190_195_groupi_n_3372 ,csa_tree_add_190_195_groupi_n_4861);
  or csa_tree_add_190_195_groupi_g43325(csa_tree_add_190_195_groupi_n_5712 ,csa_tree_add_190_195_groupi_n_4748 ,csa_tree_add_190_195_groupi_n_4742);
  nor csa_tree_add_190_195_groupi_g43326(csa_tree_add_190_195_groupi_n_5711 ,csa_tree_add_190_195_groupi_n_2726 ,csa_tree_add_190_195_groupi_n_4739);
  nor csa_tree_add_190_195_groupi_g43327(csa_tree_add_190_195_groupi_n_5710 ,csa_tree_add_190_195_groupi_n_5015 ,csa_tree_add_190_195_groupi_n_5034);
  and csa_tree_add_190_195_groupi_g43328(csa_tree_add_190_195_groupi_n_5709 ,csa_tree_add_190_195_groupi_n_2210 ,csa_tree_add_190_195_groupi_n_5056);
  nor csa_tree_add_190_195_groupi_g43329(csa_tree_add_190_195_groupi_n_5708 ,csa_tree_add_190_195_groupi_n_2210 ,csa_tree_add_190_195_groupi_n_5056);
  or csa_tree_add_190_195_groupi_g43330(csa_tree_add_190_195_groupi_n_5707 ,csa_tree_add_190_195_groupi_n_4672 ,csa_tree_add_190_195_groupi_n_5055);
  or csa_tree_add_190_195_groupi_g43331(csa_tree_add_190_195_groupi_n_5706 ,csa_tree_add_190_195_groupi_n_5047 ,csa_tree_add_190_195_groupi_n_4936);
  and csa_tree_add_190_195_groupi_g43332(csa_tree_add_190_195_groupi_n_5705 ,csa_tree_add_190_195_groupi_n_4729 ,csa_tree_add_190_195_groupi_n_5065);
  or csa_tree_add_190_195_groupi_g43333(csa_tree_add_190_195_groupi_n_5704 ,csa_tree_add_190_195_groupi_n_5016 ,csa_tree_add_190_195_groupi_n_5033);
  or csa_tree_add_190_195_groupi_g43334(csa_tree_add_190_195_groupi_n_5703 ,csa_tree_add_190_195_groupi_n_4727 ,csa_tree_add_190_195_groupi_n_4688);
  nor csa_tree_add_190_195_groupi_g43335(csa_tree_add_190_195_groupi_n_5702 ,csa_tree_add_190_195_groupi_n_4583 ,csa_tree_add_190_195_groupi_n_5027);
  or csa_tree_add_190_195_groupi_g43336(csa_tree_add_190_195_groupi_n_5701 ,csa_tree_add_190_195_groupi_n_4617 ,csa_tree_add_190_195_groupi_n_4613);
  nor csa_tree_add_190_195_groupi_g43337(csa_tree_add_190_195_groupi_n_5700 ,csa_tree_add_190_195_groupi_n_2682 ,csa_tree_add_190_195_groupi_n_5053);
  or csa_tree_add_190_195_groupi_g43338(csa_tree_add_190_195_groupi_n_5699 ,csa_tree_add_190_195_groupi_n_4602 ,csa_tree_add_190_195_groupi_n_4962);
  or csa_tree_add_190_195_groupi_g43339(csa_tree_add_190_195_groupi_n_5698 ,csa_tree_add_190_195_groupi_n_4754 ,csa_tree_add_190_195_groupi_n_4714);
  nor csa_tree_add_190_195_groupi_g43340(csa_tree_add_190_195_groupi_n_5697 ,csa_tree_add_190_195_groupi_n_4581 ,csa_tree_add_190_195_groupi_n_5002);
  nor csa_tree_add_190_195_groupi_g43341(csa_tree_add_190_195_groupi_n_5696 ,csa_tree_add_190_195_groupi_n_5007 ,csa_tree_add_190_195_groupi_n_4795);
  nor csa_tree_add_190_195_groupi_g43342(csa_tree_add_190_195_groupi_n_5695 ,csa_tree_add_190_195_groupi_n_4726 ,csa_tree_add_190_195_groupi_n_4749);
  or csa_tree_add_190_195_groupi_g43343(csa_tree_add_190_195_groupi_n_5694 ,csa_tree_add_190_195_groupi_n_1930 ,csa_tree_add_190_195_groupi_n_4701);
  or csa_tree_add_190_195_groupi_g43344(csa_tree_add_190_195_groupi_n_5693 ,csa_tree_add_190_195_groupi_n_4725 ,csa_tree_add_190_195_groupi_n_4750);
  nor csa_tree_add_190_195_groupi_g43345(csa_tree_add_190_195_groupi_n_5692 ,csa_tree_add_190_195_groupi_n_2616 ,csa_tree_add_190_195_groupi_n_4702);
  nor csa_tree_add_190_195_groupi_g43346(csa_tree_add_190_195_groupi_n_5691 ,csa_tree_add_190_195_groupi_n_4563 ,csa_tree_add_190_195_groupi_n_4740);
  and csa_tree_add_190_195_groupi_g43347(csa_tree_add_190_195_groupi_n_5690 ,csa_tree_add_190_195_groupi_n_5018 ,csa_tree_add_190_195_groupi_n_4753);
  nor csa_tree_add_190_195_groupi_g43348(csa_tree_add_190_195_groupi_n_5689 ,csa_tree_add_190_195_groupi_n_4911 ,csa_tree_add_190_195_groupi_n_4599);
  and csa_tree_add_190_195_groupi_g43349(csa_tree_add_190_195_groupi_n_5688 ,csa_tree_add_190_195_groupi_n_4690 ,csa_tree_add_190_195_groupi_n_4925);
  or csa_tree_add_190_195_groupi_g43350(csa_tree_add_190_195_groupi_n_5687 ,csa_tree_add_190_195_groupi_n_4626 ,csa_tree_add_190_195_groupi_n_4623);
  and csa_tree_add_190_195_groupi_g43351(csa_tree_add_190_195_groupi_n_5686 ,csa_tree_add_190_195_groupi_n_4617 ,csa_tree_add_190_195_groupi_n_4613);
  nor csa_tree_add_190_195_groupi_g43352(csa_tree_add_190_195_groupi_n_5685 ,csa_tree_add_190_195_groupi_n_4716 ,csa_tree_add_190_195_groupi_n_5039);
  or csa_tree_add_190_195_groupi_g43353(csa_tree_add_190_195_groupi_n_5684 ,csa_tree_add_190_195_groupi_n_4717 ,csa_tree_add_190_195_groupi_n_4982);
  nor csa_tree_add_190_195_groupi_g43354(csa_tree_add_190_195_groupi_n_5683 ,csa_tree_add_190_195_groupi_n_3300 ,csa_tree_add_190_195_groupi_n_4830);
  or csa_tree_add_190_195_groupi_g43355(csa_tree_add_190_195_groupi_n_5682 ,csa_tree_add_190_195_groupi_n_4730 ,csa_tree_add_190_195_groupi_n_4719);
  and csa_tree_add_190_195_groupi_g43356(csa_tree_add_190_195_groupi_n_5681 ,csa_tree_add_190_195_groupi_n_3220 ,csa_tree_add_190_195_groupi_n_4856);
  and csa_tree_add_190_195_groupi_g43357(csa_tree_add_190_195_groupi_n_5680 ,csa_tree_add_190_195_groupi_n_4393 ,csa_tree_add_190_195_groupi_n_4848);
  nor csa_tree_add_190_195_groupi_g43358(csa_tree_add_190_195_groupi_n_5679 ,csa_tree_add_190_195_groupi_n_4769 ,csa_tree_add_190_195_groupi_n_4889);
  or csa_tree_add_190_195_groupi_g43359(csa_tree_add_190_195_groupi_n_5678 ,csa_tree_add_190_195_groupi_n_4963 ,csa_tree_add_190_195_groupi_n_4667);
  nor csa_tree_add_190_195_groupi_g43360(csa_tree_add_190_195_groupi_n_5677 ,csa_tree_add_190_195_groupi_n_4710 ,csa_tree_add_190_195_groupi_n_4630);
  and csa_tree_add_190_195_groupi_g43361(csa_tree_add_190_195_groupi_n_5676 ,csa_tree_add_190_195_groupi_n_4660 ,csa_tree_add_190_195_groupi_n_4677);
  or csa_tree_add_190_195_groupi_g43362(csa_tree_add_190_195_groupi_n_5675 ,csa_tree_add_190_195_groupi_n_3686 ,csa_tree_add_190_195_groupi_n_4819);
  nor csa_tree_add_190_195_groupi_g43363(csa_tree_add_190_195_groupi_n_5674 ,csa_tree_add_190_195_groupi_n_1303 ,csa_tree_add_190_195_groupi_n_4665);
  or csa_tree_add_190_195_groupi_g43364(csa_tree_add_190_195_groupi_n_5673 ,csa_tree_add_190_195_groupi_n_4690 ,csa_tree_add_190_195_groupi_n_4925);
  nor csa_tree_add_190_195_groupi_g43365(csa_tree_add_190_195_groupi_n_5672 ,csa_tree_add_190_195_groupi_n_1866 ,csa_tree_add_190_195_groupi_n_4996);
  or csa_tree_add_190_195_groupi_g43366(csa_tree_add_190_195_groupi_n_5671 ,csa_tree_add_190_195_groupi_n_4768 ,csa_tree_add_190_195_groupi_n_4890);
  and csa_tree_add_190_195_groupi_g43367(csa_tree_add_190_195_groupi_n_5670 ,csa_tree_add_190_195_groupi_n_506 ,csa_tree_add_190_195_groupi_n_4665);
  or csa_tree_add_190_195_groupi_g43368(csa_tree_add_190_195_groupi_n_5669 ,csa_tree_add_190_195_groupi_n_4693 ,csa_tree_add_190_195_groupi_n_4684);
  nor csa_tree_add_190_195_groupi_g43369(csa_tree_add_190_195_groupi_n_5668 ,csa_tree_add_190_195_groupi_n_4596 ,csa_tree_add_190_195_groupi_n_4736);
  nor csa_tree_add_190_195_groupi_g43370(csa_tree_add_190_195_groupi_n_5667 ,csa_tree_add_190_195_groupi_n_4731 ,csa_tree_add_190_195_groupi_n_4720);
  or csa_tree_add_190_195_groupi_g43371(csa_tree_add_190_195_groupi_n_5666 ,csa_tree_add_190_195_groupi_n_4597 ,csa_tree_add_190_195_groupi_n_4735);
  or csa_tree_add_190_195_groupi_g43372(csa_tree_add_190_195_groupi_n_5665 ,csa_tree_add_190_195_groupi_n_4660 ,csa_tree_add_190_195_groupi_n_4677);
  or csa_tree_add_190_195_groupi_g43373(csa_tree_add_190_195_groupi_n_5664 ,csa_tree_add_190_195_groupi_n_4587 ,csa_tree_add_190_195_groupi_n_5074);
  and csa_tree_add_190_195_groupi_g43374(csa_tree_add_190_195_groupi_n_5663 ,csa_tree_add_190_195_groupi_n_4689 ,csa_tree_add_190_195_groupi_n_4881);
  or csa_tree_add_190_195_groupi_g43375(csa_tree_add_190_195_groupi_n_5662 ,csa_tree_add_190_195_groupi_n_4972 ,csa_tree_add_190_195_groupi_n_4971);
  and csa_tree_add_190_195_groupi_g43376(csa_tree_add_190_195_groupi_n_5661 ,csa_tree_add_190_195_groupi_n_4671 ,csa_tree_add_190_195_groupi_n_4669);
  nor csa_tree_add_190_195_groupi_g43377(csa_tree_add_190_195_groupi_n_5660 ,csa_tree_add_190_195_groupi_n_4653 ,csa_tree_add_190_195_groupi_n_5009);
  or csa_tree_add_190_195_groupi_g43378(csa_tree_add_190_195_groupi_n_5659 ,csa_tree_add_190_195_groupi_n_3091 ,csa_tree_add_190_195_groupi_n_4814);
  or csa_tree_add_190_195_groupi_g43379(csa_tree_add_190_195_groupi_n_5658 ,csa_tree_add_190_195_groupi_n_4671 ,csa_tree_add_190_195_groupi_n_4669);
  and csa_tree_add_190_195_groupi_g43380(csa_tree_add_190_195_groupi_n_5657 ,csa_tree_add_190_195_groupi_n_4683 ,csa_tree_add_190_195_groupi_n_5025);
  nor csa_tree_add_190_195_groupi_g43381(csa_tree_add_190_195_groupi_n_5656 ,csa_tree_add_190_195_groupi_n_4683 ,csa_tree_add_190_195_groupi_n_5025);
  or csa_tree_add_190_195_groupi_g43382(csa_tree_add_190_195_groupi_n_5655 ,csa_tree_add_190_195_groupi_n_4116 ,csa_tree_add_190_195_groupi_n_4912);
  or csa_tree_add_190_195_groupi_g43383(csa_tree_add_190_195_groupi_n_5654 ,csa_tree_add_190_195_groupi_n_1965 ,csa_tree_add_190_195_groupi_n_5088);
  nor csa_tree_add_190_195_groupi_g43384(csa_tree_add_190_195_groupi_n_5653 ,csa_tree_add_190_195_groupi_n_4646 ,csa_tree_add_190_195_groupi_n_4589);
  and csa_tree_add_190_195_groupi_g43385(csa_tree_add_190_195_groupi_n_5652 ,csa_tree_add_190_195_groupi_n_3535 ,csa_tree_add_190_195_groupi_n_4842);
  or csa_tree_add_190_195_groupi_g43386(csa_tree_add_190_195_groupi_n_5651 ,csa_tree_add_190_195_groupi_n_3654 ,csa_tree_add_190_195_groupi_n_4807);
  and csa_tree_add_190_195_groupi_g43387(csa_tree_add_190_195_groupi_n_5650 ,csa_tree_add_190_195_groupi_n_4643 ,csa_tree_add_190_195_groupi_n_4691);
  nor csa_tree_add_190_195_groupi_g43388(csa_tree_add_190_195_groupi_n_5649 ,csa_tree_add_190_195_groupi_n_4643 ,csa_tree_add_190_195_groupi_n_4691);
  or csa_tree_add_190_195_groupi_g43389(csa_tree_add_190_195_groupi_n_5648 ,csa_tree_add_190_195_groupi_n_3179 ,csa_tree_add_190_195_groupi_n_4806);
  or csa_tree_add_190_195_groupi_g43390(csa_tree_add_190_195_groupi_n_5647 ,csa_tree_add_190_195_groupi_n_4584 ,csa_tree_add_190_195_groupi_n_5026);
  nor csa_tree_add_190_195_groupi_g43391(csa_tree_add_190_195_groupi_n_5646 ,csa_tree_add_190_195_groupi_n_4627 ,csa_tree_add_190_195_groupi_n_4622);
  nor csa_tree_add_190_195_groupi_g43392(csa_tree_add_190_195_groupi_n_5645 ,csa_tree_add_190_195_groupi_n_3698 ,csa_tree_add_190_195_groupi_n_5086);
  nor csa_tree_add_190_195_groupi_g43393(csa_tree_add_190_195_groupi_n_5644 ,csa_tree_add_190_195_groupi_n_5046 ,csa_tree_add_190_195_groupi_n_4937);
  or csa_tree_add_190_195_groupi_g43394(csa_tree_add_190_195_groupi_n_5643 ,csa_tree_add_190_195_groupi_n_1401 ,csa_tree_add_190_195_groupi_n_4614);
  nor csa_tree_add_190_195_groupi_g43395(csa_tree_add_190_195_groupi_n_5642 ,csa_tree_add_190_195_groupi_n_387 ,csa_tree_add_190_195_groupi_n_4615);
  or csa_tree_add_190_195_groupi_g43396(csa_tree_add_190_195_groupi_n_5641 ,csa_tree_add_190_195_groupi_n_4668 ,csa_tree_add_190_195_groupi_n_4647);
  nor csa_tree_add_190_195_groupi_g43397(csa_tree_add_190_195_groupi_n_5640 ,csa_tree_add_190_195_groupi_n_5020 ,csa_tree_add_190_195_groupi_n_4605);
  or csa_tree_add_190_195_groupi_g43398(csa_tree_add_190_195_groupi_n_5639 ,csa_tree_add_190_195_groupi_n_5019 ,csa_tree_add_190_195_groupi_n_4604);
  and csa_tree_add_190_195_groupi_g43399(csa_tree_add_190_195_groupi_n_5638 ,csa_tree_add_190_195_groupi_n_832 ,csa_tree_add_190_195_groupi_n_4887);
  or csa_tree_add_190_195_groupi_g43400(csa_tree_add_190_195_groupi_n_5637 ,csa_tree_add_190_195_groupi_n_978 ,csa_tree_add_190_195_groupi_n_4887);
  and csa_tree_add_190_195_groupi_g43401(csa_tree_add_190_195_groupi_n_5636 ,csa_tree_add_190_195_groupi_n_625 ,csa_tree_add_190_195_groupi_n_5003);
  nor csa_tree_add_190_195_groupi_g43402(csa_tree_add_190_195_groupi_n_5635 ,csa_tree_add_190_195_groupi_n_582 ,csa_tree_add_190_195_groupi_n_5003);
  and csa_tree_add_190_195_groupi_g43403(csa_tree_add_190_195_groupi_n_5634 ,csa_tree_add_190_195_groupi_n_4619 ,csa_tree_add_190_195_groupi_n_4616);
  nor csa_tree_add_190_195_groupi_g43404(csa_tree_add_190_195_groupi_n_5633 ,csa_tree_add_190_195_groupi_n_4619 ,csa_tree_add_190_195_groupi_n_4616);
  or csa_tree_add_190_195_groupi_g43405(csa_tree_add_190_195_groupi_n_5632 ,csa_tree_add_190_195_groupi_n_3345 ,csa_tree_add_190_195_groupi_n_5150);
  nor csa_tree_add_190_195_groupi_g43406(csa_tree_add_190_195_groupi_n_5631 ,csa_tree_add_190_195_groupi_n_3202 ,csa_tree_add_190_195_groupi_n_4885);
  and csa_tree_add_190_195_groupi_g43407(csa_tree_add_190_195_groupi_n_5630 ,csa_tree_add_190_195_groupi_n_3691 ,csa_tree_add_190_195_groupi_n_4909);
  or csa_tree_add_190_195_groupi_g43408(csa_tree_add_190_195_groupi_n_5629 ,csa_tree_add_190_195_groupi_n_1314 ,csa_tree_add_190_195_groupi_n_4909);
  or csa_tree_add_190_195_groupi_g43409(csa_tree_add_190_195_groupi_n_5628 ,csa_tree_add_190_195_groupi_n_2393 ,csa_tree_add_190_195_groupi_n_4884);
  nor csa_tree_add_190_195_groupi_g43410(csa_tree_add_190_195_groupi_n_5627 ,csa_tree_add_190_195_groupi_n_4933 ,csa_tree_add_190_195_groupi_n_4935);
  or csa_tree_add_190_195_groupi_g43411(csa_tree_add_190_195_groupi_n_5626 ,csa_tree_add_190_195_groupi_n_4932 ,csa_tree_add_190_195_groupi_n_4934);
  or csa_tree_add_190_195_groupi_g43412(csa_tree_add_190_195_groupi_n_5625 ,csa_tree_add_190_195_groupi_n_4576 ,csa_tree_add_190_195_groupi_n_4835);
  nor csa_tree_add_190_195_groupi_g43413(csa_tree_add_190_195_groupi_n_5624 ,csa_tree_add_190_195_groupi_n_5051 ,csa_tree_add_190_195_groupi_n_4952);
  or csa_tree_add_190_195_groupi_g43414(csa_tree_add_190_195_groupi_n_5623 ,csa_tree_add_190_195_groupi_n_5050 ,csa_tree_add_190_195_groupi_n_4951);
  or csa_tree_add_190_195_groupi_g43415(csa_tree_add_190_195_groupi_n_5622 ,csa_tree_add_190_195_groupi_n_3699 ,csa_tree_add_190_195_groupi_n_5085);
  or csa_tree_add_190_195_groupi_g43416(csa_tree_add_190_195_groupi_n_5621 ,csa_tree_add_190_195_groupi_n_4721 ,csa_tree_add_190_195_groupi_n_4939);
  or csa_tree_add_190_195_groupi_g43417(csa_tree_add_190_195_groupi_n_5620 ,csa_tree_add_190_195_groupi_n_3693 ,csa_tree_add_190_195_groupi_n_4777);
  and csa_tree_add_190_195_groupi_g43418(csa_tree_add_190_195_groupi_n_5619 ,csa_tree_add_190_195_groupi_n_4670 ,csa_tree_add_190_195_groupi_n_4781);
  nor csa_tree_add_190_195_groupi_g43419(csa_tree_add_190_195_groupi_n_5618 ,csa_tree_add_190_195_groupi_n_3692 ,csa_tree_add_190_195_groupi_n_4778);
  nor csa_tree_add_190_195_groupi_g43420(csa_tree_add_190_195_groupi_n_5617 ,csa_tree_add_190_195_groupi_n_4681 ,csa_tree_add_190_195_groupi_n_4679);
  or csa_tree_add_190_195_groupi_g43421(csa_tree_add_190_195_groupi_n_5616 ,csa_tree_add_190_195_groupi_n_4670 ,csa_tree_add_190_195_groupi_n_4781);
  nor csa_tree_add_190_195_groupi_g43422(csa_tree_add_190_195_groupi_n_5615 ,csa_tree_add_190_195_groupi_n_4964 ,csa_tree_add_190_195_groupi_n_4666);
  nor csa_tree_add_190_195_groupi_g43423(csa_tree_add_190_195_groupi_n_5614 ,csa_tree_add_190_195_groupi_n_4722 ,csa_tree_add_190_195_groupi_n_4938);
  or csa_tree_add_190_195_groupi_g43424(csa_tree_add_190_195_groupi_n_5613 ,csa_tree_add_190_195_groupi_n_4680 ,csa_tree_add_190_195_groupi_n_4678);
  and csa_tree_add_190_195_groupi_g43425(csa_tree_add_190_195_groupi_n_5983 ,csa_tree_add_190_195_groupi_n_3204 ,csa_tree_add_190_195_groupi_n_4849);
  xnor csa_tree_add_190_195_groupi_g43426(csa_tree_add_190_195_groupi_n_5982 ,csa_tree_add_190_195_groupi_n_15 ,csa_tree_add_190_195_groupi_n_952);
  and csa_tree_add_190_195_groupi_g43427(csa_tree_add_190_195_groupi_n_5981 ,csa_tree_add_190_195_groupi_n_3684 ,csa_tree_add_190_195_groupi_n_4874);
  xnor csa_tree_add_190_195_groupi_g43428(csa_tree_add_190_195_groupi_n_5980 ,csa_tree_add_190_195_groupi_n_3923 ,csa_tree_add_190_195_groupi_n_1129);
  xnor csa_tree_add_190_195_groupi_g43429(csa_tree_add_190_195_groupi_n_5979 ,csa_tree_add_190_195_groupi_n_3924 ,csa_tree_add_190_195_groupi_n_1838);
  xnor csa_tree_add_190_195_groupi_g43430(csa_tree_add_190_195_groupi_n_5978 ,csa_tree_add_190_195_groupi_n_4026 ,in61[14]);
  xnor csa_tree_add_190_195_groupi_g43431(csa_tree_add_190_195_groupi_n_5977 ,csa_tree_add_190_195_groupi_n_4080 ,csa_tree_add_190_195_groupi_n_1997);
  or csa_tree_add_190_195_groupi_g43432(csa_tree_add_190_195_groupi_n_5975 ,csa_tree_add_190_195_groupi_n_3487 ,csa_tree_add_190_195_groupi_n_4577);
  or csa_tree_add_190_195_groupi_g43433(csa_tree_add_190_195_groupi_n_5973 ,csa_tree_add_190_195_groupi_n_3109 ,csa_tree_add_190_195_groupi_n_4579);
  xnor csa_tree_add_190_195_groupi_g43434(csa_tree_add_190_195_groupi_n_5972 ,csa_tree_add_190_195_groupi_n_3932 ,in59[3]);
  xnor csa_tree_add_190_195_groupi_g43435(csa_tree_add_190_195_groupi_n_5970 ,csa_tree_add_190_195_groupi_n_4140 ,csa_tree_add_190_195_groupi_n_4081);
  xnor csa_tree_add_190_195_groupi_g43436(csa_tree_add_190_195_groupi_n_5969 ,csa_tree_add_190_195_groupi_n_4000 ,csa_tree_add_190_195_groupi_n_1898);
  xnor csa_tree_add_190_195_groupi_g43437(csa_tree_add_190_195_groupi_n_5968 ,csa_tree_add_190_195_groupi_n_3808 ,csa_tree_add_190_195_groupi_n_1158);
  xor csa_tree_add_190_195_groupi_g43438(csa_tree_add_190_195_groupi_n_5967 ,csa_tree_add_190_195_groupi_n_3770 ,csa_tree_add_190_195_groupi_n_1629);
  or csa_tree_add_190_195_groupi_g43439(csa_tree_add_190_195_groupi_n_5966 ,csa_tree_add_190_195_groupi_n_3385 ,csa_tree_add_190_195_groupi_n_4875);
  and csa_tree_add_190_195_groupi_g43440(csa_tree_add_190_195_groupi_n_5965 ,csa_tree_add_190_195_groupi_n_3458 ,csa_tree_add_190_195_groupi_n_4876);
  xnor csa_tree_add_190_195_groupi_g43441(csa_tree_add_190_195_groupi_n_5964 ,csa_tree_add_190_195_groupi_n_3861 ,csa_tree_add_190_195_groupi_n_1081);
  xnor csa_tree_add_190_195_groupi_g43442(csa_tree_add_190_195_groupi_n_5962 ,csa_tree_add_190_195_groupi_n_3765 ,csa_tree_add_190_195_groupi_n_628);
  xnor csa_tree_add_190_195_groupi_g43443(csa_tree_add_190_195_groupi_n_5961 ,csa_tree_add_190_195_groupi_n_3913 ,csa_tree_add_190_195_groupi_n_910);
  xnor csa_tree_add_190_195_groupi_g43444(csa_tree_add_190_195_groupi_n_5960 ,csa_tree_add_190_195_groupi_n_3851 ,csa_tree_add_190_195_groupi_n_1862);
  xnor csa_tree_add_190_195_groupi_g43445(csa_tree_add_190_195_groupi_n_5959 ,csa_tree_add_190_195_groupi_n_4052 ,csa_tree_add_190_195_groupi_n_2006);
  xnor csa_tree_add_190_195_groupi_g43446(csa_tree_add_190_195_groupi_n_5957 ,csa_tree_add_190_195_groupi_n_3821 ,csa_tree_add_190_195_groupi_n_1987);
  xnor csa_tree_add_190_195_groupi_g43449(csa_tree_add_190_195_groupi_n_5953 ,csa_tree_add_190_195_groupi_n_3982 ,csa_tree_add_190_195_groupi_n_2215);
  xnor csa_tree_add_190_195_groupi_g43450(csa_tree_add_190_195_groupi_n_5951 ,csa_tree_add_190_195_groupi_n_3730 ,csa_tree_add_190_195_groupi_n_1120);
  xnor csa_tree_add_190_195_groupi_g43451(csa_tree_add_190_195_groupi_n_5949 ,csa_tree_add_190_195_groupi_n_3887 ,csa_tree_add_190_195_groupi_n_1915);
  xnor csa_tree_add_190_195_groupi_g43452(csa_tree_add_190_195_groupi_n_5948 ,csa_tree_add_190_195_groupi_n_3819 ,csa_tree_add_190_195_groupi_n_898);
  xnor csa_tree_add_190_195_groupi_g43453(csa_tree_add_190_195_groupi_n_5946 ,csa_tree_add_190_195_groupi_n_3811 ,csa_tree_add_190_195_groupi_n_1305);
  xnor csa_tree_add_190_195_groupi_g43454(csa_tree_add_190_195_groupi_n_5944 ,csa_tree_add_190_195_groupi_n_3853 ,in61[4]);
  xnor csa_tree_add_190_195_groupi_g43455(csa_tree_add_190_195_groupi_n_5942 ,csa_tree_add_190_195_groupi_n_4094 ,csa_tree_add_190_195_groupi_n_1039);
  xnor csa_tree_add_190_195_groupi_g43456(csa_tree_add_190_195_groupi_n_5940 ,csa_tree_add_190_195_groupi_n_4035 ,csa_tree_add_190_195_groupi_n_1045);
  xnor csa_tree_add_190_195_groupi_g43457(csa_tree_add_190_195_groupi_n_5938 ,csa_tree_add_190_195_groupi_n_3753 ,csa_tree_add_190_195_groupi_n_2039);
  xnor csa_tree_add_190_195_groupi_g43458(csa_tree_add_190_195_groupi_n_5937 ,csa_tree_add_190_195_groupi_n_4059 ,csa_tree_add_190_195_groupi_n_1993);
  xnor csa_tree_add_190_195_groupi_g43459(csa_tree_add_190_195_groupi_n_5935 ,csa_tree_add_190_195_groupi_n_4064 ,csa_tree_add_190_195_groupi_n_1104);
  xnor csa_tree_add_190_195_groupi_g43460(csa_tree_add_190_195_groupi_n_5932 ,csa_tree_add_190_195_groupi_n_3744 ,csa_tree_add_190_195_groupi_n_1690);
  xnor csa_tree_add_190_195_groupi_g43461(csa_tree_add_190_195_groupi_n_5931 ,csa_tree_add_190_195_groupi_n_3868 ,csa_tree_add_190_195_groupi_n_2052);
  xnor csa_tree_add_190_195_groupi_g43462(csa_tree_add_190_195_groupi_n_5929 ,csa_tree_add_190_195_groupi_n_4109 ,csa_tree_add_190_195_groupi_n_2085);
  xnor csa_tree_add_190_195_groupi_g43463(csa_tree_add_190_195_groupi_n_5928 ,csa_tree_add_190_195_groupi_n_3946 ,csa_tree_add_190_195_groupi_n_1972);
  xnor csa_tree_add_190_195_groupi_g43464(csa_tree_add_190_195_groupi_n_5926 ,csa_tree_add_190_195_groupi_n_3792 ,csa_tree_add_190_195_groupi_n_570);
  xnor csa_tree_add_190_195_groupi_g43465(csa_tree_add_190_195_groupi_n_5924 ,csa_tree_add_190_195_groupi_n_3786 ,csa_tree_add_190_195_groupi_n_1774);
  xnor csa_tree_add_190_195_groupi_g43466(csa_tree_add_190_195_groupi_n_5922 ,csa_tree_add_190_195_groupi_n_3745 ,csa_tree_add_190_195_groupi_n_1287);
  xnor csa_tree_add_190_195_groupi_g43467(csa_tree_add_190_195_groupi_n_5920 ,csa_tree_add_190_195_groupi_n_3825 ,in58[6]);
  xnor csa_tree_add_190_195_groupi_g43468(csa_tree_add_190_195_groupi_n_5918 ,csa_tree_add_190_195_groupi_n_4113 ,csa_tree_add_190_195_groupi_n_1714);
  xnor csa_tree_add_190_195_groupi_g43469(csa_tree_add_190_195_groupi_n_5917 ,csa_tree_add_190_195_groupi_n_3947 ,csa_tree_add_190_195_groupi_n_1584);
  xnor csa_tree_add_190_195_groupi_g43470(csa_tree_add_190_195_groupi_n_5916 ,csa_tree_add_190_195_groupi_n_3779 ,csa_tree_add_190_195_groupi_n_1611);
  xnor csa_tree_add_190_195_groupi_g43471(csa_tree_add_190_195_groupi_n_5915 ,csa_tree_add_190_195_groupi_n_4005 ,csa_tree_add_190_195_groupi_n_1856);
  xnor csa_tree_add_190_195_groupi_g43473(csa_tree_add_190_195_groupi_n_5912 ,csa_tree_add_190_195_groupi_n_4073 ,csa_tree_add_190_195_groupi_n_556);
  xnor csa_tree_add_190_195_groupi_g43474(csa_tree_add_190_195_groupi_n_5910 ,csa_tree_add_190_195_groupi_n_45 ,csa_tree_add_190_195_groupi_n_1689);
  xnor csa_tree_add_190_195_groupi_g43475(csa_tree_add_190_195_groupi_n_5908 ,csa_tree_add_190_195_groupi_n_3969 ,csa_tree_add_190_195_groupi_n_1950);
  xnor csa_tree_add_190_195_groupi_g43476(csa_tree_add_190_195_groupi_n_5907 ,csa_tree_add_190_195_groupi_n_4129 ,csa_tree_add_190_195_groupi_n_1825);
  xnor csa_tree_add_190_195_groupi_g43478(csa_tree_add_190_195_groupi_n_5905 ,csa_tree_add_190_195_groupi_n_3864 ,in61[3]);
  xnor csa_tree_add_190_195_groupi_g43479(csa_tree_add_190_195_groupi_n_5903 ,csa_tree_add_190_195_groupi_n_3750 ,csa_tree_add_190_195_groupi_n_496);
  xnor csa_tree_add_190_195_groupi_g43480(csa_tree_add_190_195_groupi_n_5902 ,csa_tree_add_190_195_groupi_n_4002 ,csa_tree_add_190_195_groupi_n_2119);
  xnor csa_tree_add_190_195_groupi_g43481(csa_tree_add_190_195_groupi_n_5900 ,csa_tree_add_190_195_groupi_n_3768 ,csa_tree_add_190_195_groupi_n_1588);
  xnor csa_tree_add_190_195_groupi_g43482(csa_tree_add_190_195_groupi_n_5899 ,csa_tree_add_190_195_groupi_n_3835 ,in58[8]);
  xnor csa_tree_add_190_195_groupi_g43485(csa_tree_add_190_195_groupi_n_5896 ,csa_tree_add_190_195_groupi_n_33 ,csa_tree_add_190_195_groupi_n_1827);
  xnor csa_tree_add_190_195_groupi_g43486(csa_tree_add_190_195_groupi_n_5895 ,csa_tree_add_190_195_groupi_n_3863 ,csa_tree_add_190_195_groupi_n_466);
  xnor csa_tree_add_190_195_groupi_g43487(csa_tree_add_190_195_groupi_n_5894 ,csa_tree_add_190_195_groupi_n_3872 ,csa_tree_add_190_195_groupi_n_1299);
  xnor csa_tree_add_190_195_groupi_g43489(csa_tree_add_190_195_groupi_n_5890 ,csa_tree_add_190_195_groupi_n_4124 ,csa_tree_add_190_195_groupi_n_2453);
  xnor csa_tree_add_190_195_groupi_g43490(csa_tree_add_190_195_groupi_n_5889 ,csa_tree_add_190_195_groupi_n_3782 ,csa_tree_add_190_195_groupi_n_1920);
  xnor csa_tree_add_190_195_groupi_g43491(csa_tree_add_190_195_groupi_n_5888 ,csa_tree_add_190_195_groupi_n_3789 ,csa_tree_add_190_195_groupi_n_1180);
  xnor csa_tree_add_190_195_groupi_g43492(csa_tree_add_190_195_groupi_n_5887 ,csa_tree_add_190_195_groupi_n_3843 ,csa_tree_add_190_195_groupi_n_473);
  xnor csa_tree_add_190_195_groupi_g43493(csa_tree_add_190_195_groupi_n_5885 ,csa_tree_add_190_195_groupi_n_3916 ,csa_tree_add_190_195_groupi_n_1289);
  xnor csa_tree_add_190_195_groupi_g43494(csa_tree_add_190_195_groupi_n_5883 ,csa_tree_add_190_195_groupi_n_3942 ,csa_tree_add_190_195_groupi_n_1976);
  xnor csa_tree_add_190_195_groupi_g43495(csa_tree_add_190_195_groupi_n_5881 ,csa_tree_add_190_195_groupi_n_3797 ,csa_tree_add_190_195_groupi_n_1710);
  xnor csa_tree_add_190_195_groupi_g43496(csa_tree_add_190_195_groupi_n_5879 ,csa_tree_add_190_195_groupi_n_3978 ,csa_tree_add_190_195_groupi_n_1996);
  xnor csa_tree_add_190_195_groupi_g43497(csa_tree_add_190_195_groupi_n_5877 ,csa_tree_add_190_195_groupi_n_3929 ,csa_tree_add_190_195_groupi_n_1745);
  xnor csa_tree_add_190_195_groupi_g43498(csa_tree_add_190_195_groupi_n_5876 ,csa_tree_add_190_195_groupi_n_3772 ,csa_tree_add_190_195_groupi_n_454);
  xnor csa_tree_add_190_195_groupi_g43499(csa_tree_add_190_195_groupi_n_5874 ,csa_tree_add_190_195_groupi_n_3998 ,csa_tree_add_190_195_groupi_n_2049);
  xnor csa_tree_add_190_195_groupi_g43500(csa_tree_add_190_195_groupi_n_5873 ,csa_tree_add_190_195_groupi_n_3875 ,csa_tree_add_190_195_groupi_n_903);
  xnor csa_tree_add_190_195_groupi_g43501(csa_tree_add_190_195_groupi_n_5872 ,csa_tree_add_190_195_groupi_n_4039 ,csa_tree_add_190_195_groupi_n_867);
  xnor csa_tree_add_190_195_groupi_g43502(csa_tree_add_190_195_groupi_n_5869 ,csa_tree_add_190_195_groupi_n_3931 ,csa_tree_add_190_195_groupi_n_1916);
  xnor csa_tree_add_190_195_groupi_g43503(csa_tree_add_190_195_groupi_n_5868 ,csa_tree_add_190_195_groupi_n_3885 ,csa_tree_add_190_195_groupi_n_1174);
  not csa_tree_add_190_195_groupi_g43504(csa_tree_add_190_195_groupi_n_5608 ,csa_tree_add_190_195_groupi_n_5607);
  not csa_tree_add_190_195_groupi_g43505(csa_tree_add_190_195_groupi_n_5606 ,csa_tree_add_190_195_groupi_n_5605);
  not csa_tree_add_190_195_groupi_g43506(csa_tree_add_190_195_groupi_n_5600 ,csa_tree_add_190_195_groupi_n_5599);
  not csa_tree_add_190_195_groupi_g43507(csa_tree_add_190_195_groupi_n_5598 ,csa_tree_add_190_195_groupi_n_5597);
  not csa_tree_add_190_195_groupi_g43508(csa_tree_add_190_195_groupi_n_5587 ,csa_tree_add_190_195_groupi_n_5586);
  not csa_tree_add_190_195_groupi_g43510(csa_tree_add_190_195_groupi_n_5547 ,csa_tree_add_190_195_groupi_n_5548);
  not csa_tree_add_190_195_groupi_g43512(csa_tree_add_190_195_groupi_n_5543 ,csa_tree_add_190_195_groupi_n_5544);
  not csa_tree_add_190_195_groupi_g43514(csa_tree_add_190_195_groupi_n_5539 ,csa_tree_add_190_195_groupi_n_5540);
  not csa_tree_add_190_195_groupi_g43515(csa_tree_add_190_195_groupi_n_5537 ,csa_tree_add_190_195_groupi_n_5538);
  not csa_tree_add_190_195_groupi_g43516(csa_tree_add_190_195_groupi_n_5535 ,csa_tree_add_190_195_groupi_n_5536);
  not csa_tree_add_190_195_groupi_g43517(csa_tree_add_190_195_groupi_n_5534 ,csa_tree_add_190_195_groupi_n_70);
  not csa_tree_add_190_195_groupi_g43518(csa_tree_add_190_195_groupi_n_5532 ,csa_tree_add_190_195_groupi_n_5533);
  not csa_tree_add_190_195_groupi_g43519(csa_tree_add_190_195_groupi_n_5530 ,csa_tree_add_190_195_groupi_n_5529);
  not csa_tree_add_190_195_groupi_g43520(csa_tree_add_190_195_groupi_n_5527 ,csa_tree_add_190_195_groupi_n_5528);
  not csa_tree_add_190_195_groupi_g43521(csa_tree_add_190_195_groupi_n_5525 ,csa_tree_add_190_195_groupi_n_5526);
  not csa_tree_add_190_195_groupi_g43522(csa_tree_add_190_195_groupi_n_5523 ,csa_tree_add_190_195_groupi_n_5524);
  not csa_tree_add_190_195_groupi_g43523(csa_tree_add_190_195_groupi_n_5521 ,csa_tree_add_190_195_groupi_n_5522);
  not csa_tree_add_190_195_groupi_g43525(csa_tree_add_190_195_groupi_n_5518 ,csa_tree_add_190_195_groupi_n_5519);
  not csa_tree_add_190_195_groupi_g43526(csa_tree_add_190_195_groupi_n_5517 ,csa_tree_add_190_195_groupi_n_18);
  not csa_tree_add_190_195_groupi_g43527(csa_tree_add_190_195_groupi_n_5515 ,csa_tree_add_190_195_groupi_n_5516);
  not csa_tree_add_190_195_groupi_g43528(csa_tree_add_190_195_groupi_n_5512 ,csa_tree_add_190_195_groupi_n_14);
  not csa_tree_add_190_195_groupi_g43529(csa_tree_add_190_195_groupi_n_5510 ,csa_tree_add_190_195_groupi_n_5511);
  not csa_tree_add_190_195_groupi_g43530(csa_tree_add_190_195_groupi_n_5507 ,csa_tree_add_190_195_groupi_n_5508);
  not csa_tree_add_190_195_groupi_g43531(csa_tree_add_190_195_groupi_n_5505 ,csa_tree_add_190_195_groupi_n_5506);
  not csa_tree_add_190_195_groupi_g43532(csa_tree_add_190_195_groupi_n_5502 ,csa_tree_add_190_195_groupi_n_5503);
  not csa_tree_add_190_195_groupi_g43533(csa_tree_add_190_195_groupi_n_5500 ,csa_tree_add_190_195_groupi_n_5501);
  not csa_tree_add_190_195_groupi_g43534(csa_tree_add_190_195_groupi_n_5498 ,csa_tree_add_190_195_groupi_n_5499);
  not csa_tree_add_190_195_groupi_g43535(csa_tree_add_190_195_groupi_n_5496 ,csa_tree_add_190_195_groupi_n_5497);
  not csa_tree_add_190_195_groupi_g43536(csa_tree_add_190_195_groupi_n_5495 ,csa_tree_add_190_195_groupi_n_5494);
  not csa_tree_add_190_195_groupi_g43537(csa_tree_add_190_195_groupi_n_5492 ,csa_tree_add_190_195_groupi_n_5493);
  not csa_tree_add_190_195_groupi_g43538(csa_tree_add_190_195_groupi_n_5489 ,csa_tree_add_190_195_groupi_n_5490);
  not csa_tree_add_190_195_groupi_g43539(csa_tree_add_190_195_groupi_n_5486 ,csa_tree_add_190_195_groupi_n_5487);
  not csa_tree_add_190_195_groupi_g43540(csa_tree_add_190_195_groupi_n_5483 ,csa_tree_add_190_195_groupi_n_5484);
  not csa_tree_add_190_195_groupi_g43541(csa_tree_add_190_195_groupi_n_5481 ,csa_tree_add_190_195_groupi_n_5482);
  not csa_tree_add_190_195_groupi_g43542(csa_tree_add_190_195_groupi_n_5479 ,csa_tree_add_190_195_groupi_n_5480);
  not csa_tree_add_190_195_groupi_g43543(csa_tree_add_190_195_groupi_n_5477 ,csa_tree_add_190_195_groupi_n_5478);
  not csa_tree_add_190_195_groupi_g43544(csa_tree_add_190_195_groupi_n_5475 ,csa_tree_add_190_195_groupi_n_5476);
  not csa_tree_add_190_195_groupi_g43545(csa_tree_add_190_195_groupi_n_5473 ,csa_tree_add_190_195_groupi_n_5474);
  not csa_tree_add_190_195_groupi_g43546(csa_tree_add_190_195_groupi_n_5468 ,csa_tree_add_190_195_groupi_n_5467);
  not csa_tree_add_190_195_groupi_g43547(csa_tree_add_190_195_groupi_n_5463 ,csa_tree_add_190_195_groupi_n_5462);
  not csa_tree_add_190_195_groupi_g43548(csa_tree_add_190_195_groupi_n_5461 ,csa_tree_add_190_195_groupi_n_5460);
  not csa_tree_add_190_195_groupi_g43549(csa_tree_add_190_195_groupi_n_5458 ,csa_tree_add_190_195_groupi_n_5457);
  not csa_tree_add_190_195_groupi_g43550(csa_tree_add_190_195_groupi_n_5456 ,csa_tree_add_190_195_groupi_n_5455);
  not csa_tree_add_190_195_groupi_g43551(csa_tree_add_190_195_groupi_n_5453 ,csa_tree_add_190_195_groupi_n_5454);
  not csa_tree_add_190_195_groupi_g43552(csa_tree_add_190_195_groupi_n_5450 ,csa_tree_add_190_195_groupi_n_5451);
  not csa_tree_add_190_195_groupi_g43553(csa_tree_add_190_195_groupi_n_5448 ,csa_tree_add_190_195_groupi_n_5449);
  not csa_tree_add_190_195_groupi_g43554(csa_tree_add_190_195_groupi_n_5447 ,csa_tree_add_190_195_groupi_n_24);
  not csa_tree_add_190_195_groupi_g43555(csa_tree_add_190_195_groupi_n_5445 ,csa_tree_add_190_195_groupi_n_5446);
  not csa_tree_add_190_195_groupi_g43556(csa_tree_add_190_195_groupi_n_5440 ,csa_tree_add_190_195_groupi_n_5441);
  not csa_tree_add_190_195_groupi_g43557(csa_tree_add_190_195_groupi_n_5439 ,csa_tree_add_190_195_groupi_n_64);
  not csa_tree_add_190_195_groupi_g43558(csa_tree_add_190_195_groupi_n_5437 ,csa_tree_add_190_195_groupi_n_5438);
  not csa_tree_add_190_195_groupi_g43559(csa_tree_add_190_195_groupi_n_5434 ,csa_tree_add_190_195_groupi_n_5435);
  not csa_tree_add_190_195_groupi_g43560(csa_tree_add_190_195_groupi_n_5432 ,csa_tree_add_190_195_groupi_n_71);
  not csa_tree_add_190_195_groupi_g43561(csa_tree_add_190_195_groupi_n_5431 ,csa_tree_add_190_195_groupi_n_5430);
  not csa_tree_add_190_195_groupi_g43562(csa_tree_add_190_195_groupi_n_5428 ,csa_tree_add_190_195_groupi_n_75);
  not csa_tree_add_190_195_groupi_g43563(csa_tree_add_190_195_groupi_n_5426 ,csa_tree_add_190_195_groupi_n_61);
  not csa_tree_add_190_195_groupi_g43564(csa_tree_add_190_195_groupi_n_5424 ,csa_tree_add_190_195_groupi_n_5425);
  not csa_tree_add_190_195_groupi_g43566(csa_tree_add_190_195_groupi_n_5420 ,csa_tree_add_190_195_groupi_n_5421);
  not csa_tree_add_190_195_groupi_g43567(csa_tree_add_190_195_groupi_n_5413 ,csa_tree_add_190_195_groupi_n_32);
  not csa_tree_add_190_195_groupi_g43568(csa_tree_add_190_195_groupi_n_5412 ,csa_tree_add_190_195_groupi_n_81);
  not csa_tree_add_190_195_groupi_g43570(csa_tree_add_190_195_groupi_n_5409 ,csa_tree_add_190_195_groupi_n_5410);
  not csa_tree_add_190_195_groupi_g43571(csa_tree_add_190_195_groupi_n_5405 ,csa_tree_add_190_195_groupi_n_5406);
  not csa_tree_add_190_195_groupi_g43572(csa_tree_add_190_195_groupi_n_5403 ,csa_tree_add_190_195_groupi_n_5404);
  not csa_tree_add_190_195_groupi_g43573(csa_tree_add_190_195_groupi_n_5402 ,csa_tree_add_190_195_groupi_n_5401);
  not csa_tree_add_190_195_groupi_g43574(csa_tree_add_190_195_groupi_n_5396 ,csa_tree_add_190_195_groupi_n_8);
  not csa_tree_add_190_195_groupi_g43575(csa_tree_add_190_195_groupi_n_5395 ,csa_tree_add_190_195_groupi_n_5394);
  not csa_tree_add_190_195_groupi_g43576(csa_tree_add_190_195_groupi_n_5390 ,csa_tree_add_190_195_groupi_n_5391);
  not csa_tree_add_190_195_groupi_g43577(csa_tree_add_190_195_groupi_n_5386 ,csa_tree_add_190_195_groupi_n_5387);
  not csa_tree_add_190_195_groupi_g43578(csa_tree_add_190_195_groupi_n_5383 ,csa_tree_add_190_195_groupi_n_5384);
  not csa_tree_add_190_195_groupi_g43579(csa_tree_add_190_195_groupi_n_5381 ,csa_tree_add_190_195_groupi_n_77);
  not csa_tree_add_190_195_groupi_g43580(csa_tree_add_190_195_groupi_n_5377 ,csa_tree_add_190_195_groupi_n_5378);
  not csa_tree_add_190_195_groupi_g43581(csa_tree_add_190_195_groupi_n_5376 ,csa_tree_add_190_195_groupi_n_58);
  not csa_tree_add_190_195_groupi_g43582(csa_tree_add_190_195_groupi_n_5372 ,csa_tree_add_190_195_groupi_n_5373);
  not csa_tree_add_190_195_groupi_g43583(csa_tree_add_190_195_groupi_n_5370 ,csa_tree_add_190_195_groupi_n_5371);
  not csa_tree_add_190_195_groupi_g43584(csa_tree_add_190_195_groupi_n_5368 ,csa_tree_add_190_195_groupi_n_5369);
  not csa_tree_add_190_195_groupi_g43585(csa_tree_add_190_195_groupi_n_5363 ,csa_tree_add_190_195_groupi_n_5364);
  not csa_tree_add_190_195_groupi_g43586(csa_tree_add_190_195_groupi_n_5361 ,csa_tree_add_190_195_groupi_n_5362);
  not csa_tree_add_190_195_groupi_g43587(csa_tree_add_190_195_groupi_n_5359 ,csa_tree_add_190_195_groupi_n_5360);
  not csa_tree_add_190_195_groupi_g43588(csa_tree_add_190_195_groupi_n_5357 ,csa_tree_add_190_195_groupi_n_5358);
  not csa_tree_add_190_195_groupi_g43589(csa_tree_add_190_195_groupi_n_5354 ,csa_tree_add_190_195_groupi_n_5355);
  not csa_tree_add_190_195_groupi_g43590(csa_tree_add_190_195_groupi_n_5346 ,csa_tree_add_190_195_groupi_n_5347);
  not csa_tree_add_190_195_groupi_g43591(csa_tree_add_190_195_groupi_n_5343 ,csa_tree_add_190_195_groupi_n_5344);
  not csa_tree_add_190_195_groupi_g43592(csa_tree_add_190_195_groupi_n_5341 ,csa_tree_add_190_195_groupi_n_5342);
  not csa_tree_add_190_195_groupi_g43593(csa_tree_add_190_195_groupi_n_5339 ,csa_tree_add_190_195_groupi_n_5340);
  not csa_tree_add_190_195_groupi_g43594(csa_tree_add_190_195_groupi_n_5337 ,csa_tree_add_190_195_groupi_n_5338);
  not csa_tree_add_190_195_groupi_g43595(csa_tree_add_190_195_groupi_n_5334 ,csa_tree_add_190_195_groupi_n_5335);
  not csa_tree_add_190_195_groupi_g43596(csa_tree_add_190_195_groupi_n_5332 ,csa_tree_add_190_195_groupi_n_5333);
  not csa_tree_add_190_195_groupi_g43597(csa_tree_add_190_195_groupi_n_5330 ,csa_tree_add_190_195_groupi_n_5331);
  not csa_tree_add_190_195_groupi_g43599(csa_tree_add_190_195_groupi_n_5327 ,csa_tree_add_190_195_groupi_n_5328);
  not csa_tree_add_190_195_groupi_g43600(csa_tree_add_190_195_groupi_n_5324 ,csa_tree_add_190_195_groupi_n_5325);
  not csa_tree_add_190_195_groupi_g43602(csa_tree_add_190_195_groupi_n_5319 ,csa_tree_add_190_195_groupi_n_5320);
  not csa_tree_add_190_195_groupi_g43603(csa_tree_add_190_195_groupi_n_5317 ,csa_tree_add_190_195_groupi_n_5318);
  not csa_tree_add_190_195_groupi_g43604(csa_tree_add_190_195_groupi_n_5316 ,csa_tree_add_190_195_groupi_n_5315);
  not csa_tree_add_190_195_groupi_g43605(csa_tree_add_190_195_groupi_n_5314 ,csa_tree_add_190_195_groupi_n_5313);
  not csa_tree_add_190_195_groupi_g43606(csa_tree_add_190_195_groupi_n_5309 ,csa_tree_add_190_195_groupi_n_5310);
  not csa_tree_add_190_195_groupi_g43607(csa_tree_add_190_195_groupi_n_5308 ,csa_tree_add_190_195_groupi_n_20);
  not csa_tree_add_190_195_groupi_g43608(csa_tree_add_190_195_groupi_n_5307 ,csa_tree_add_190_195_groupi_n_5306);
  not csa_tree_add_190_195_groupi_g43609(csa_tree_add_190_195_groupi_n_5305 ,csa_tree_add_190_195_groupi_n_10);
  not csa_tree_add_190_195_groupi_g43610(csa_tree_add_190_195_groupi_n_5303 ,csa_tree_add_190_195_groupi_n_5304);
  not csa_tree_add_190_195_groupi_g43611(csa_tree_add_190_195_groupi_n_5300 ,csa_tree_add_190_195_groupi_n_5301);
  not csa_tree_add_190_195_groupi_g43612(csa_tree_add_190_195_groupi_n_5295 ,csa_tree_add_190_195_groupi_n_5296);
  not csa_tree_add_190_195_groupi_g43613(csa_tree_add_190_195_groupi_n_5293 ,csa_tree_add_190_195_groupi_n_5294);
  not csa_tree_add_190_195_groupi_g43614(csa_tree_add_190_195_groupi_n_5290 ,csa_tree_add_190_195_groupi_n_5291);
  not csa_tree_add_190_195_groupi_g43615(csa_tree_add_190_195_groupi_n_5288 ,csa_tree_add_190_195_groupi_n_5287);
  not csa_tree_add_190_195_groupi_g43617(csa_tree_add_190_195_groupi_n_5284 ,csa_tree_add_190_195_groupi_n_5285);
  not csa_tree_add_190_195_groupi_g43618(csa_tree_add_190_195_groupi_n_5279 ,csa_tree_add_190_195_groupi_n_5280);
  not csa_tree_add_190_195_groupi_g43619(csa_tree_add_190_195_groupi_n_5276 ,csa_tree_add_190_195_groupi_n_5277);
  not csa_tree_add_190_195_groupi_g43620(csa_tree_add_190_195_groupi_n_5273 ,csa_tree_add_190_195_groupi_n_5274);
  not csa_tree_add_190_195_groupi_g43621(csa_tree_add_190_195_groupi_n_5271 ,csa_tree_add_190_195_groupi_n_5272);
  not csa_tree_add_190_195_groupi_g43623(csa_tree_add_190_195_groupi_n_5267 ,csa_tree_add_190_195_groupi_n_5268);
  not csa_tree_add_190_195_groupi_g43624(csa_tree_add_190_195_groupi_n_5264 ,csa_tree_add_190_195_groupi_n_5265);
  not csa_tree_add_190_195_groupi_g43625(csa_tree_add_190_195_groupi_n_5261 ,csa_tree_add_190_195_groupi_n_5262);
  not csa_tree_add_190_195_groupi_g43627(csa_tree_add_190_195_groupi_n_5254 ,csa_tree_add_190_195_groupi_n_5255);
  not csa_tree_add_190_195_groupi_g43629(csa_tree_add_190_195_groupi_n_5251 ,csa_tree_add_190_195_groupi_n_56);
  not csa_tree_add_190_195_groupi_g43630(csa_tree_add_190_195_groupi_n_5249 ,csa_tree_add_190_195_groupi_n_5250);
  not csa_tree_add_190_195_groupi_g43631(csa_tree_add_190_195_groupi_n_5247 ,csa_tree_add_190_195_groupi_n_5248);
  not csa_tree_add_190_195_groupi_g43632(csa_tree_add_190_195_groupi_n_5246 ,csa_tree_add_190_195_groupi_n_5245);
  not csa_tree_add_190_195_groupi_g43634(csa_tree_add_190_195_groupi_n_5237 ,csa_tree_add_190_195_groupi_n_5238);
  not csa_tree_add_190_195_groupi_g43635(csa_tree_add_190_195_groupi_n_5235 ,csa_tree_add_190_195_groupi_n_5234);
  not csa_tree_add_190_195_groupi_g43636(csa_tree_add_190_195_groupi_n_5231 ,csa_tree_add_190_195_groupi_n_5232);
  not csa_tree_add_190_195_groupi_g43637(csa_tree_add_190_195_groupi_n_5229 ,csa_tree_add_190_195_groupi_n_5228);
  not csa_tree_add_190_195_groupi_g43638(csa_tree_add_190_195_groupi_n_5226 ,csa_tree_add_190_195_groupi_n_5227);
  not csa_tree_add_190_195_groupi_g43639(csa_tree_add_190_195_groupi_n_5222 ,csa_tree_add_190_195_groupi_n_5223);
  not csa_tree_add_190_195_groupi_g43640(csa_tree_add_190_195_groupi_n_5221 ,csa_tree_add_190_195_groupi_n_66);
  not csa_tree_add_190_195_groupi_g43641(csa_tree_add_190_195_groupi_n_5219 ,csa_tree_add_190_195_groupi_n_5220);
  not csa_tree_add_190_195_groupi_g43642(csa_tree_add_190_195_groupi_n_5215 ,csa_tree_add_190_195_groupi_n_5216);
  not csa_tree_add_190_195_groupi_g43643(csa_tree_add_190_195_groupi_n_5213 ,csa_tree_add_190_195_groupi_n_5214);
  not csa_tree_add_190_195_groupi_g43644(csa_tree_add_190_195_groupi_n_5211 ,csa_tree_add_190_195_groupi_n_5212);
  not csa_tree_add_190_195_groupi_g43646(csa_tree_add_190_195_groupi_n_5208 ,csa_tree_add_190_195_groupi_n_5209);
  not csa_tree_add_190_195_groupi_g43647(csa_tree_add_190_195_groupi_n_5204 ,csa_tree_add_190_195_groupi_n_5205);
  not csa_tree_add_190_195_groupi_g43648(csa_tree_add_190_195_groupi_n_5197 ,csa_tree_add_190_195_groupi_n_5198);
  not csa_tree_add_190_195_groupi_g43649(csa_tree_add_190_195_groupi_n_5195 ,csa_tree_add_190_195_groupi_n_5196);
  not csa_tree_add_190_195_groupi_g43650(csa_tree_add_190_195_groupi_n_5194 ,csa_tree_add_190_195_groupi_n_42);
  not csa_tree_add_190_195_groupi_g43651(csa_tree_add_190_195_groupi_n_5192 ,csa_tree_add_190_195_groupi_n_5193);
  not csa_tree_add_190_195_groupi_g43652(csa_tree_add_190_195_groupi_n_5190 ,csa_tree_add_190_195_groupi_n_5191);
  not csa_tree_add_190_195_groupi_g43653(csa_tree_add_190_195_groupi_n_5188 ,csa_tree_add_190_195_groupi_n_5189);
  not csa_tree_add_190_195_groupi_g43654(csa_tree_add_190_195_groupi_n_5186 ,csa_tree_add_190_195_groupi_n_5187);
  not csa_tree_add_190_195_groupi_g43655(csa_tree_add_190_195_groupi_n_5184 ,csa_tree_add_190_195_groupi_n_5185);
  not csa_tree_add_190_195_groupi_g43656(csa_tree_add_190_195_groupi_n_5182 ,csa_tree_add_190_195_groupi_n_5183);
  not csa_tree_add_190_195_groupi_g43657(csa_tree_add_190_195_groupi_n_5180 ,csa_tree_add_190_195_groupi_n_5181);
  xnor csa_tree_add_190_195_groupi_g43658(csa_tree_add_190_195_groupi_n_5179 ,csa_tree_add_190_195_groupi_n_4141 ,csa_tree_add_190_195_groupi_n_1932);
  xnor csa_tree_add_190_195_groupi_g43659(csa_tree_add_190_195_groupi_n_5178 ,csa_tree_add_190_195_groupi_n_4138 ,csa_tree_add_190_195_groupi_n_1988);
  xnor csa_tree_add_190_195_groupi_g43660(csa_tree_add_190_195_groupi_n_5177 ,csa_tree_add_190_195_groupi_n_4142 ,csa_tree_add_190_195_groupi_n_510);
  xnor csa_tree_add_190_195_groupi_g43661(csa_tree_add_190_195_groupi_n_5176 ,csa_tree_add_190_195_groupi_n_4567 ,csa_tree_add_190_195_groupi_n_1846);
  xnor csa_tree_add_190_195_groupi_g43662(csa_tree_add_190_195_groupi_n_5175 ,csa_tree_add_190_195_groupi_n_4139 ,csa_tree_add_190_195_groupi_n_1994);
  xnor csa_tree_add_190_195_groupi_g43663(csa_tree_add_190_195_groupi_n_5612 ,csa_tree_add_190_195_groupi_n_3838 ,in58[9]);
  xnor csa_tree_add_190_195_groupi_g43664(csa_tree_add_190_195_groupi_n_5611 ,csa_tree_add_190_195_groupi_n_3798 ,in59[2]);
  xnor csa_tree_add_190_195_groupi_g43665(csa_tree_add_190_195_groupi_n_5610 ,csa_tree_add_190_195_groupi_n_3860 ,in58[10]);
  xnor csa_tree_add_190_195_groupi_g43666(csa_tree_add_190_195_groupi_n_5609 ,csa_tree_add_190_195_groupi_n_3974 ,csa_tree_add_190_195_groupi_n_1810);
  xnor csa_tree_add_190_195_groupi_g43668(csa_tree_add_190_195_groupi_n_5607 ,csa_tree_add_190_195_groupi_n_4121 ,csa_tree_add_190_195_groupi_n_1699);
  xnor csa_tree_add_190_195_groupi_g43669(csa_tree_add_190_195_groupi_n_5605 ,csa_tree_add_190_195_groupi_n_3816 ,csa_tree_add_190_195_groupi_n_2153);
  xor csa_tree_add_190_195_groupi_g43670(csa_tree_add_190_195_groupi_n_5604 ,csa_tree_add_190_195_groupi_n_3965 ,csa_tree_add_190_195_groupi_n_1084);
  xnor csa_tree_add_190_195_groupi_g43673(csa_tree_add_190_195_groupi_n_5603 ,csa_tree_add_190_195_groupi_n_3834 ,in58[11]);
  xor csa_tree_add_190_195_groupi_g43674(csa_tree_add_190_195_groupi_n_5602 ,csa_tree_add_190_195_groupi_n_3943 ,csa_tree_add_190_195_groupi_n_1998);
  xnor csa_tree_add_190_195_groupi_g43675(csa_tree_add_190_195_groupi_n_5601 ,csa_tree_add_190_195_groupi_n_3917 ,csa_tree_add_190_195_groupi_n_1824);
  xnor csa_tree_add_190_195_groupi_g43677(csa_tree_add_190_195_groupi_n_5599 ,csa_tree_add_190_195_groupi_n_4034 ,csa_tree_add_190_195_groupi_n_1742);
  xnor csa_tree_add_190_195_groupi_g43678(csa_tree_add_190_195_groupi_n_5597 ,csa_tree_add_190_195_groupi_n_3888 ,csa_tree_add_190_195_groupi_n_607);
  xor csa_tree_add_190_195_groupi_g43679(csa_tree_add_190_195_groupi_n_5596 ,csa_tree_add_190_195_groupi_n_4053 ,in61[15]);
  xnor csa_tree_add_190_195_groupi_g43681(csa_tree_add_190_195_groupi_n_5595 ,csa_tree_add_190_195_groupi_n_270 ,csa_tree_add_190_195_groupi_n_1330);
  xnor csa_tree_add_190_195_groupi_g43682(csa_tree_add_190_195_groupi_n_5594 ,csa_tree_add_190_195_groupi_n_3702 ,csa_tree_add_190_195_groupi_n_3735);
  xnor csa_tree_add_190_195_groupi_g43683(csa_tree_add_190_195_groupi_n_5593 ,csa_tree_add_190_195_groupi_n_4144 ,csa_tree_add_190_195_groupi_n_1964);
  xnor csa_tree_add_190_195_groupi_g43684(csa_tree_add_190_195_groupi_n_5592 ,csa_tree_add_190_195_groupi_n_2 ,csa_tree_add_190_195_groupi_n_1107);
  xnor csa_tree_add_190_195_groupi_g43686(csa_tree_add_190_195_groupi_n_5591 ,csa_tree_add_190_195_groupi_n_4104 ,csa_tree_add_190_195_groupi_n_762);
  xnor csa_tree_add_190_195_groupi_g43687(csa_tree_add_190_195_groupi_n_5590 ,csa_tree_add_190_195_groupi_n_3949 ,in60[5]);
  xnor csa_tree_add_190_195_groupi_g43688(csa_tree_add_190_195_groupi_n_5589 ,csa_tree_add_190_195_groupi_n_3985 ,csa_tree_add_190_195_groupi_n_1978);
  xnor csa_tree_add_190_195_groupi_g43689(csa_tree_add_190_195_groupi_n_5588 ,csa_tree_add_190_195_groupi_n_4122 ,csa_tree_add_190_195_groupi_n_2050);
  xnor csa_tree_add_190_195_groupi_g43690(csa_tree_add_190_195_groupi_n_5586 ,csa_tree_add_190_195_groupi_n_4040 ,csa_tree_add_190_195_groupi_n_1892);
  xnor csa_tree_add_190_195_groupi_g43691(csa_tree_add_190_195_groupi_n_5585 ,csa_tree_add_190_195_groupi_n_3818 ,csa_tree_add_190_195_groupi_n_1161);
  xnor csa_tree_add_190_195_groupi_g43692(csa_tree_add_190_195_groupi_n_5584 ,csa_tree_add_190_195_groupi_n_3958 ,csa_tree_add_190_195_groupi_n_758);
  xnor csa_tree_add_190_195_groupi_g43693(csa_tree_add_190_195_groupi_n_5583 ,csa_tree_add_190_195_groupi_n_3733 ,csa_tree_add_190_195_groupi_n_1688);
  xnor csa_tree_add_190_195_groupi_g43694(csa_tree_add_190_195_groupi_n_5582 ,csa_tree_add_190_195_groupi_n_4015 ,in59[4]);
  xnor csa_tree_add_190_195_groupi_g43695(csa_tree_add_190_195_groupi_n_5581 ,csa_tree_add_190_195_groupi_n_3989 ,in56[12]);
  xnor csa_tree_add_190_195_groupi_g43696(csa_tree_add_190_195_groupi_n_5580 ,csa_tree_add_190_195_groupi_n_4050 ,csa_tree_add_190_195_groupi_n_933);
  xnor csa_tree_add_190_195_groupi_g43697(csa_tree_add_190_195_groupi_n_5579 ,csa_tree_add_190_195_groupi_n_3829 ,in57[8]);
  xnor csa_tree_add_190_195_groupi_g43698(csa_tree_add_190_195_groupi_n_5578 ,csa_tree_add_190_195_groupi_n_4089 ,csa_tree_add_190_195_groupi_n_2053);
  xnor csa_tree_add_190_195_groupi_g43699(csa_tree_add_190_195_groupi_n_5577 ,csa_tree_add_190_195_groupi_n_4020 ,in60[1]);
  xnor csa_tree_add_190_195_groupi_g43700(csa_tree_add_190_195_groupi_n_5576 ,csa_tree_add_190_195_groupi_n_4056 ,csa_tree_add_190_195_groupi_n_1265);
  xnor csa_tree_add_190_195_groupi_g43701(csa_tree_add_190_195_groupi_n_5575 ,csa_tree_add_190_195_groupi_n_4129 ,csa_tree_add_190_195_groupi_n_1978);
  xnor csa_tree_add_190_195_groupi_g43702(csa_tree_add_190_195_groupi_n_5574 ,csa_tree_add_190_195_groupi_n_3751 ,csa_tree_add_190_195_groupi_n_1704);
  xnor csa_tree_add_190_195_groupi_g43703(csa_tree_add_190_195_groupi_n_5573 ,csa_tree_add_190_195_groupi_n_4004 ,csa_tree_add_190_195_groupi_n_1009);
  xnor csa_tree_add_190_195_groupi_g43704(csa_tree_add_190_195_groupi_n_5572 ,csa_tree_add_190_195_groupi_n_3991 ,in59[7]);
  xnor csa_tree_add_190_195_groupi_g43705(csa_tree_add_190_195_groupi_n_5571 ,csa_tree_add_190_195_groupi_n_3856 ,in57[3]);
  xnor csa_tree_add_190_195_groupi_g43706(csa_tree_add_190_195_groupi_n_5570 ,csa_tree_add_190_195_groupi_n_4046 ,csa_tree_add_190_195_groupi_n_1977);
  xnor csa_tree_add_190_195_groupi_g43707(csa_tree_add_190_195_groupi_n_5569 ,csa_tree_add_190_195_groupi_n_4096 ,csa_tree_add_190_195_groupi_n_1704);
  xnor csa_tree_add_190_195_groupi_g43708(csa_tree_add_190_195_groupi_n_5568 ,csa_tree_add_190_195_groupi_n_3747 ,csa_tree_add_190_195_groupi_n_1824);
  xnor csa_tree_add_190_195_groupi_g43709(csa_tree_add_190_195_groupi_n_5567 ,csa_tree_add_190_195_groupi_n_3748 ,csa_tree_add_190_195_groupi_n_1996);
  xnor csa_tree_add_190_195_groupi_g43710(csa_tree_add_190_195_groupi_n_5566 ,csa_tree_add_190_195_groupi_n_3755 ,csa_tree_add_190_195_groupi_n_1920);
  xnor csa_tree_add_190_195_groupi_g43711(csa_tree_add_190_195_groupi_n_5565 ,csa_tree_add_190_195_groupi_n_1 ,csa_tree_add_190_195_groupi_n_1710);
  xnor csa_tree_add_190_195_groupi_g43712(csa_tree_add_190_195_groupi_n_5564 ,csa_tree_add_190_195_groupi_n_3849 ,in57[6]);
  xnor csa_tree_add_190_195_groupi_g43713(csa_tree_add_190_195_groupi_n_5563 ,csa_tree_add_190_195_groupi_n_3899 ,csa_tree_add_190_195_groupi_n_1809);
  xnor csa_tree_add_190_195_groupi_g43714(csa_tree_add_190_195_groupi_n_5562 ,csa_tree_add_190_195_groupi_n_3740 ,csa_tree_add_190_195_groupi_n_1021);
  xnor csa_tree_add_190_195_groupi_g43715(csa_tree_add_190_195_groupi_n_5561 ,csa_tree_add_190_195_groupi_n_4018 ,in56[1]);
  xnor csa_tree_add_190_195_groupi_g43716(csa_tree_add_190_195_groupi_n_5560 ,csa_tree_add_190_195_groupi_n_4033 ,csa_tree_add_190_195_groupi_n_2117);
  xnor csa_tree_add_190_195_groupi_g43717(csa_tree_add_190_195_groupi_n_5559 ,csa_tree_add_190_195_groupi_n_4106 ,csa_tree_add_190_195_groupi_n_1595);
  xnor csa_tree_add_190_195_groupi_g43718(csa_tree_add_190_195_groupi_n_5558 ,csa_tree_add_190_195_groupi_n_4120 ,csa_tree_add_190_195_groupi_n_1911);
  xnor csa_tree_add_190_195_groupi_g43719(csa_tree_add_190_195_groupi_n_5557 ,csa_tree_add_190_195_groupi_n_3966 ,csa_tree_add_190_195_groupi_n_1908);
  xnor csa_tree_add_190_195_groupi_g43720(csa_tree_add_190_195_groupi_n_5556 ,csa_tree_add_190_195_groupi_n_12 ,csa_tree_add_190_195_groupi_n_1963);
  xnor csa_tree_add_190_195_groupi_g43721(csa_tree_add_190_195_groupi_n_5555 ,csa_tree_add_190_195_groupi_n_3842 ,in55[7]);
  xnor csa_tree_add_190_195_groupi_g43722(csa_tree_add_190_195_groupi_n_5554 ,csa_tree_add_190_195_groupi_n_4131 ,csa_tree_add_190_195_groupi_n_1837);
  xnor csa_tree_add_190_195_groupi_g43723(csa_tree_add_190_195_groupi_n_5553 ,csa_tree_add_190_195_groupi_n_3840 ,in57[9]);
  xnor csa_tree_add_190_195_groupi_g43724(csa_tree_add_190_195_groupi_n_5552 ,csa_tree_add_190_195_groupi_n_3771 ,csa_tree_add_190_195_groupi_n_1042);
  xnor csa_tree_add_190_195_groupi_g43725(csa_tree_add_190_195_groupi_n_5551 ,csa_tree_add_190_195_groupi_n_4016 ,csa_tree_add_190_195_groupi_n_1839);
  xnor csa_tree_add_190_195_groupi_g43726(csa_tree_add_190_195_groupi_n_5550 ,csa_tree_add_190_195_groupi_n_3832 ,csa_tree_add_190_195_groupi_n_1891);
  xnor csa_tree_add_190_195_groupi_g43728(csa_tree_add_190_195_groupi_n_5549 ,csa_tree_add_190_195_groupi_n_3776 ,csa_tree_add_190_195_groupi_n_1694);
  xnor csa_tree_add_190_195_groupi_g43729(csa_tree_add_190_195_groupi_n_5548 ,csa_tree_add_190_195_groupi_n_4006 ,csa_tree_add_190_195_groupi_n_800);
  xnor csa_tree_add_190_195_groupi_g43730(csa_tree_add_190_195_groupi_n_5546 ,csa_tree_add_190_195_groupi_n_4024 ,csa_tree_add_190_195_groupi_n_1808);
  xnor csa_tree_add_190_195_groupi_g43731(csa_tree_add_190_195_groupi_n_5545 ,csa_tree_add_190_195_groupi_n_4123 ,csa_tree_add_190_195_groupi_n_522);
  xnor csa_tree_add_190_195_groupi_g43732(csa_tree_add_190_195_groupi_n_5544 ,csa_tree_add_190_195_groupi_n_3784 ,csa_tree_add_190_195_groupi_n_1679);
  xnor csa_tree_add_190_195_groupi_g43733(csa_tree_add_190_195_groupi_n_5542 ,csa_tree_add_190_195_groupi_n_3921 ,csa_tree_add_190_195_groupi_n_1862);
  xnor csa_tree_add_190_195_groupi_g43734(csa_tree_add_190_195_groupi_n_5541 ,csa_tree_add_190_195_groupi_n_4071 ,csa_tree_add_190_195_groupi_n_1897);
  xnor csa_tree_add_190_195_groupi_g43735(csa_tree_add_190_195_groupi_n_5540 ,csa_tree_add_190_195_groupi_n_3925 ,csa_tree_add_190_195_groupi_n_1697);
  xnor csa_tree_add_190_195_groupi_g43736(csa_tree_add_190_195_groupi_n_5538 ,csa_tree_add_190_195_groupi_n_4105 ,csa_tree_add_190_195_groupi_n_1822);
  xnor csa_tree_add_190_195_groupi_g43737(csa_tree_add_190_195_groupi_n_5536 ,csa_tree_add_190_195_groupi_n_3934 ,csa_tree_add_190_195_groupi_n_1904);
  xnor csa_tree_add_190_195_groupi_g43739(csa_tree_add_190_195_groupi_n_5533 ,csa_tree_add_190_195_groupi_n_4084 ,csa_tree_add_190_195_groupi_n_1659);
  xnor csa_tree_add_190_195_groupi_g43740(csa_tree_add_190_195_groupi_n_5531 ,csa_tree_add_190_195_groupi_n_3738 ,csa_tree_add_190_195_groupi_n_2006);
  xnor csa_tree_add_190_195_groupi_g43741(csa_tree_add_190_195_groupi_n_5529 ,csa_tree_add_190_195_groupi_n_3854 ,csa_tree_add_190_195_groupi_n_2708);
  xnor csa_tree_add_190_195_groupi_g43743(csa_tree_add_190_195_groupi_n_5528 ,csa_tree_add_190_195_groupi_n_3820 ,csa_tree_add_190_195_groupi_n_1825);
  xnor csa_tree_add_190_195_groupi_g43744(csa_tree_add_190_195_groupi_n_5526 ,csa_tree_add_190_195_groupi_n_3866 ,csa_tree_add_190_195_groupi_n_1864);
  xnor csa_tree_add_190_195_groupi_g43745(csa_tree_add_190_195_groupi_n_5524 ,csa_tree_add_190_195_groupi_n_3886 ,csa_tree_add_190_195_groupi_n_1297);
  xnor csa_tree_add_190_195_groupi_g43746(csa_tree_add_190_195_groupi_n_5522 ,csa_tree_add_190_195_groupi_n_3830 ,in60[12]);
  xnor csa_tree_add_190_195_groupi_g43747(csa_tree_add_190_195_groupi_n_5520 ,csa_tree_add_190_195_groupi_n_3741 ,csa_tree_add_190_195_groupi_n_802);
  xnor csa_tree_add_190_195_groupi_g43748(csa_tree_add_190_195_groupi_n_5519 ,csa_tree_add_190_195_groupi_n_3912 ,csa_tree_add_190_195_groupi_n_2054);
  xnor csa_tree_add_190_195_groupi_g43750(csa_tree_add_190_195_groupi_n_5516 ,csa_tree_add_190_195_groupi_n_83 ,csa_tree_add_190_195_groupi_n_804);
  xnor csa_tree_add_190_195_groupi_g43751(csa_tree_add_190_195_groupi_n_5514 ,csa_tree_add_190_195_groupi_n_3795 ,csa_tree_add_190_195_groupi_n_1810);
  xnor csa_tree_add_190_195_groupi_g43752(csa_tree_add_190_195_groupi_n_5513 ,csa_tree_add_190_195_groupi_n_3884 ,csa_tree_add_190_195_groupi_n_2153);
  xnor csa_tree_add_190_195_groupi_g43755(csa_tree_add_190_195_groupi_n_5511 ,csa_tree_add_190_195_groupi_n_3731 ,csa_tree_add_190_195_groupi_n_1263);
  xnor csa_tree_add_190_195_groupi_g43756(csa_tree_add_190_195_groupi_n_5509 ,csa_tree_add_190_195_groupi_n_3977 ,csa_tree_add_190_195_groupi_n_1911);
  xnor csa_tree_add_190_195_groupi_g43757(csa_tree_add_190_195_groupi_n_5508 ,csa_tree_add_190_195_groupi_n_4043 ,csa_tree_add_190_195_groupi_n_1814);
  xnor csa_tree_add_190_195_groupi_g43758(csa_tree_add_190_195_groupi_n_5506 ,csa_tree_add_190_195_groupi_n_3927 ,csa_tree_add_190_195_groupi_n_1948);
  xnor csa_tree_add_190_195_groupi_g43759(csa_tree_add_190_195_groupi_n_5504 ,csa_tree_add_190_195_groupi_n_3930 ,csa_tree_add_190_195_groupi_n_1838);
  xnor csa_tree_add_190_195_groupi_g43760(csa_tree_add_190_195_groupi_n_5503 ,csa_tree_add_190_195_groupi_n_3800 ,csa_tree_add_190_195_groupi_n_886);
  xnor csa_tree_add_190_195_groupi_g43761(csa_tree_add_190_195_groupi_n_5501 ,csa_tree_add_190_195_groupi_n_3897 ,csa_tree_add_190_195_groupi_n_2016);
  xnor csa_tree_add_190_195_groupi_g43762(csa_tree_add_190_195_groupi_n_5499 ,csa_tree_add_190_195_groupi_n_3790 ,csa_tree_add_190_195_groupi_n_550);
  xnor csa_tree_add_190_195_groupi_g43763(csa_tree_add_190_195_groupi_n_5497 ,csa_tree_add_190_195_groupi_n_3941 ,csa_tree_add_190_195_groupi_n_1905);
  xnor csa_tree_add_190_195_groupi_g43764(csa_tree_add_190_195_groupi_n_5494 ,csa_tree_add_190_195_groupi_n_3951 ,csa_tree_add_190_195_groupi_n_1675);
  xnor csa_tree_add_190_195_groupi_g43765(csa_tree_add_190_195_groupi_n_5493 ,csa_tree_add_190_195_groupi_n_3898 ,csa_tree_add_190_195_groupi_n_1943);
  xnor csa_tree_add_190_195_groupi_g43766(csa_tree_add_190_195_groupi_n_5491 ,csa_tree_add_190_195_groupi_n_3870 ,csa_tree_add_190_195_groupi_n_981);
  xnor csa_tree_add_190_195_groupi_g43767(csa_tree_add_190_195_groupi_n_5490 ,csa_tree_add_190_195_groupi_n_3828 ,csa_tree_add_190_195_groupi_n_1060);
  xnor csa_tree_add_190_195_groupi_g43768(csa_tree_add_190_195_groupi_n_5488 ,csa_tree_add_190_195_groupi_n_3883 ,csa_tree_add_190_195_groupi_n_1147);
  xnor csa_tree_add_190_195_groupi_g43769(csa_tree_add_190_195_groupi_n_5487 ,csa_tree_add_190_195_groupi_n_4137 ,csa_tree_add_190_195_groupi_n_1665);
  xnor csa_tree_add_190_195_groupi_g43770(csa_tree_add_190_195_groupi_n_5485 ,csa_tree_add_190_195_groupi_n_3963 ,csa_tree_add_190_195_groupi_n_1849);
  xnor csa_tree_add_190_195_groupi_g43771(csa_tree_add_190_195_groupi_n_5484 ,csa_tree_add_190_195_groupi_n_4119 ,csa_tree_add_190_195_groupi_n_2119);
  xnor csa_tree_add_190_195_groupi_g43772(csa_tree_add_190_195_groupi_n_5482 ,csa_tree_add_190_195_groupi_n_3869 ,csa_tree_add_190_195_groupi_n_1297);
  xnor csa_tree_add_190_195_groupi_g43773(csa_tree_add_190_195_groupi_n_5480 ,csa_tree_add_190_195_groupi_n_3911 ,csa_tree_add_190_195_groupi_n_1063);
  xnor csa_tree_add_190_195_groupi_g43774(csa_tree_add_190_195_groupi_n_5478 ,csa_tree_add_190_195_groupi_n_3801 ,csa_tree_add_190_195_groupi_n_2006);
  xnor csa_tree_add_190_195_groupi_g43775(csa_tree_add_190_195_groupi_n_5476 ,csa_tree_add_190_195_groupi_n_3999 ,csa_tree_add_190_195_groupi_n_1224);
  xnor csa_tree_add_190_195_groupi_g43776(csa_tree_add_190_195_groupi_n_5474 ,csa_tree_add_190_195_groupi_n_3926 ,csa_tree_add_190_195_groupi_n_1301);
  xnor csa_tree_add_190_195_groupi_g43777(csa_tree_add_190_195_groupi_n_5472 ,csa_tree_add_190_195_groupi_n_3823 ,csa_tree_add_190_195_groupi_n_1709);
  xnor csa_tree_add_190_195_groupi_g43778(csa_tree_add_190_195_groupi_n_5471 ,csa_tree_add_190_195_groupi_n_4093 ,csa_tree_add_190_195_groupi_n_1780);
  xnor csa_tree_add_190_195_groupi_g43779(csa_tree_add_190_195_groupi_n_5470 ,csa_tree_add_190_195_groupi_n_3873 ,csa_tree_add_190_195_groupi_n_1843);
  xnor csa_tree_add_190_195_groupi_g43780(csa_tree_add_190_195_groupi_n_5469 ,csa_tree_add_190_195_groupi_n_4102 ,csa_tree_add_190_195_groupi_n_985);
  xnor csa_tree_add_190_195_groupi_g43781(csa_tree_add_190_195_groupi_n_5467 ,csa_tree_add_190_195_groupi_n_3877 ,csa_tree_add_190_195_groupi_n_1828);
  xnor csa_tree_add_190_195_groupi_g43782(csa_tree_add_190_195_groupi_n_5466 ,csa_tree_add_190_195_groupi_n_3948 ,csa_tree_add_190_195_groupi_n_1131);
  xnor csa_tree_add_190_195_groupi_g43783(csa_tree_add_190_195_groupi_n_5465 ,csa_tree_add_190_195_groupi_n_4130 ,csa_tree_add_190_195_groupi_n_2118);
  xnor csa_tree_add_190_195_groupi_g43784(csa_tree_add_190_195_groupi_n_5464 ,csa_tree_add_190_195_groupi_n_3756 ,csa_tree_add_190_195_groupi_n_1820);
  xnor csa_tree_add_190_195_groupi_g43785(csa_tree_add_190_195_groupi_n_5462 ,csa_tree_add_190_195_groupi_n_4067 ,csa_tree_add_190_195_groupi_n_1994);
  xnor csa_tree_add_190_195_groupi_g43786(csa_tree_add_190_195_groupi_n_5460 ,csa_tree_add_190_195_groupi_n_4568 ,csa_tree_add_190_195_groupi_n_1840);
  xnor csa_tree_add_190_195_groupi_g43787(csa_tree_add_190_195_groupi_n_5459 ,csa_tree_add_190_195_groupi_n_4145 ,csa_tree_add_190_195_groupi_n_1155);
  xnor csa_tree_add_190_195_groupi_g43788(csa_tree_add_190_195_groupi_n_5457 ,csa_tree_add_190_195_groupi_n_4143 ,csa_tree_add_190_195_groupi_n_1755);
  xnor csa_tree_add_190_195_groupi_g43789(csa_tree_add_190_195_groupi_n_5455 ,csa_tree_add_190_195_groupi_n_3705 ,csa_tree_add_190_195_groupi_n_3960);
  xnor csa_tree_add_190_195_groupi_g43790(csa_tree_add_190_195_groupi_n_5454 ,csa_tree_add_190_195_groupi_n_3871 ,csa_tree_add_190_195_groupi_n_1828);
  xnor csa_tree_add_190_195_groupi_g43791(csa_tree_add_190_195_groupi_n_5452 ,csa_tree_add_190_195_groupi_n_3976 ,csa_tree_add_190_195_groupi_n_583);
  xnor csa_tree_add_190_195_groupi_g43793(csa_tree_add_190_195_groupi_n_5451 ,csa_tree_add_190_195_groupi_n_4058 ,csa_tree_add_190_195_groupi_n_512);
  xnor csa_tree_add_190_195_groupi_g43795(csa_tree_add_190_195_groupi_n_5449 ,csa_tree_add_190_195_groupi_n_3984 ,in56[14]);
  xnor csa_tree_add_190_195_groupi_g43797(csa_tree_add_190_195_groupi_n_5446 ,csa_tree_add_190_195_groupi_n_3806 ,csa_tree_add_190_195_groupi_n_1756);
  xnor csa_tree_add_190_195_groupi_g43798(csa_tree_add_190_195_groupi_n_5444 ,csa_tree_add_190_195_groupi_n_3981 ,csa_tree_add_190_195_groupi_n_541);
  xnor csa_tree_add_190_195_groupi_g43799(csa_tree_add_190_195_groupi_n_5443 ,csa_tree_add_190_195_groupi_n_3971 ,csa_tree_add_190_195_groupi_n_419);
  xnor csa_tree_add_190_195_groupi_g43800(csa_tree_add_190_195_groupi_n_5442 ,csa_tree_add_190_195_groupi_n_4054 ,csa_tree_add_190_195_groupi_n_486);
  xnor csa_tree_add_190_195_groupi_g43801(csa_tree_add_190_195_groupi_n_5441 ,csa_tree_add_190_195_groupi_n_3961 ,csa_tree_add_190_195_groupi_n_1309);
  xnor csa_tree_add_190_195_groupi_g43804(csa_tree_add_190_195_groupi_n_5438 ,csa_tree_add_190_195_groupi_n_3909 ,csa_tree_add_190_195_groupi_n_2001);
  xnor csa_tree_add_190_195_groupi_g43805(csa_tree_add_190_195_groupi_n_5436 ,csa_tree_add_190_195_groupi_n_4045 ,csa_tree_add_190_195_groupi_n_586);
  xnor csa_tree_add_190_195_groupi_g43807(csa_tree_add_190_195_groupi_n_5435 ,csa_tree_add_190_195_groupi_n_4041 ,csa_tree_add_190_195_groupi_n_547);
  xnor csa_tree_add_190_195_groupi_g43808(csa_tree_add_190_195_groupi_n_5433 ,csa_tree_add_190_195_groupi_n_4076 ,csa_tree_add_190_195_groupi_n_1279);
  xnor csa_tree_add_190_195_groupi_g43810(csa_tree_add_190_195_groupi_n_5430 ,csa_tree_add_190_195_groupi_n_4031 ,csa_tree_add_190_195_groupi_n_979);
  xnor csa_tree_add_190_195_groupi_g43811(csa_tree_add_190_195_groupi_n_5429 ,csa_tree_add_190_195_groupi_n_4038 ,csa_tree_add_190_195_groupi_n_577);
  xnor csa_tree_add_190_195_groupi_g43814(csa_tree_add_190_195_groupi_n_5427 ,csa_tree_add_190_195_groupi_n_4030 ,csa_tree_add_190_195_groupi_n_544);
  xnor csa_tree_add_190_195_groupi_g43816(csa_tree_add_190_195_groupi_n_5425 ,csa_tree_add_190_195_groupi_n_3781 ,in61[1]);
  xnor csa_tree_add_190_195_groupi_g43817(csa_tree_add_190_195_groupi_n_5423 ,csa_tree_add_190_195_groupi_n_3996 ,in59[5]);
  xnor csa_tree_add_190_195_groupi_g43818(csa_tree_add_190_195_groupi_n_5422 ,csa_tree_add_190_195_groupi_n_3896 ,csa_tree_add_190_195_groupi_n_1600);
  xnor csa_tree_add_190_195_groupi_g43819(csa_tree_add_190_195_groupi_n_5421 ,csa_tree_add_190_195_groupi_n_3915 ,csa_tree_add_190_195_groupi_n_2088);
  xnor csa_tree_add_190_195_groupi_g43820(csa_tree_add_190_195_groupi_n_5419 ,csa_tree_add_190_195_groupi_n_3848 ,in57[11]);
  xnor csa_tree_add_190_195_groupi_g43821(csa_tree_add_190_195_groupi_n_5418 ,csa_tree_add_190_195_groupi_n_3933 ,csa_tree_add_190_195_groupi_n_1844);
  xnor csa_tree_add_190_195_groupi_g43822(csa_tree_add_190_195_groupi_n_5417 ,csa_tree_add_190_195_groupi_n_3953 ,csa_tree_add_190_195_groupi_n_928);
  xnor csa_tree_add_190_195_groupi_g43823(csa_tree_add_190_195_groupi_n_5416 ,csa_tree_add_190_195_groupi_n_3987 ,csa_tree_add_190_195_groupi_n_1065);
  xnor csa_tree_add_190_195_groupi_g43824(csa_tree_add_190_195_groupi_n_5415 ,csa_tree_add_190_195_groupi_n_3904 ,csa_tree_add_190_195_groupi_n_957);
  xnor csa_tree_add_190_195_groupi_g43825(csa_tree_add_190_195_groupi_n_5414 ,csa_tree_add_190_195_groupi_n_3807 ,csa_tree_add_190_195_groupi_n_2061);
  xnor csa_tree_add_190_195_groupi_g43828(csa_tree_add_190_195_groupi_n_5411 ,csa_tree_add_190_195_groupi_n_4011 ,csa_tree_add_190_195_groupi_n_2058);
  xnor csa_tree_add_190_195_groupi_g43829(csa_tree_add_190_195_groupi_n_5410 ,csa_tree_add_190_195_groupi_n_3783 ,csa_tree_add_190_195_groupi_n_1577);
  xnor csa_tree_add_190_195_groupi_g43830(csa_tree_add_190_195_groupi_n_5408 ,csa_tree_add_190_195_groupi_n_4012 ,csa_tree_add_190_195_groupi_n_1605);
  xnor csa_tree_add_190_195_groupi_g43831(csa_tree_add_190_195_groupi_n_5407 ,csa_tree_add_190_195_groupi_n_4048 ,csa_tree_add_190_195_groupi_n_1685);
  xnor csa_tree_add_190_195_groupi_g43832(csa_tree_add_190_195_groupi_n_5406 ,csa_tree_add_190_195_groupi_n_4075 ,csa_tree_add_190_195_groupi_n_1850);
  xnor csa_tree_add_190_195_groupi_g43833(csa_tree_add_190_195_groupi_n_5404 ,csa_tree_add_190_195_groupi_n_3889 ,csa_tree_add_190_195_groupi_n_1606);
  xnor csa_tree_add_190_195_groupi_g43834(csa_tree_add_190_195_groupi_n_5401 ,csa_tree_add_190_195_groupi_n_3785 ,csa_tree_add_190_195_groupi_n_1974);
  xnor csa_tree_add_190_195_groupi_g43835(csa_tree_add_190_195_groupi_n_5400 ,csa_tree_add_190_195_groupi_n_3787 ,csa_tree_add_190_195_groupi_n_806);
  xnor csa_tree_add_190_195_groupi_g43836(csa_tree_add_190_195_groupi_n_5399 ,csa_tree_add_190_195_groupi_n_4100 ,csa_tree_add_190_195_groupi_n_1927);
  xnor csa_tree_add_190_195_groupi_g43837(csa_tree_add_190_195_groupi_n_5398 ,csa_tree_add_190_195_groupi_n_4125 ,csa_tree_add_190_195_groupi_n_1686);
  xnor csa_tree_add_190_195_groupi_g43838(csa_tree_add_190_195_groupi_n_5397 ,csa_tree_add_190_195_groupi_n_3878 ,csa_tree_add_190_195_groupi_n_1609);
  xnor csa_tree_add_190_195_groupi_g43840(csa_tree_add_190_195_groupi_n_5394 ,csa_tree_add_190_195_groupi_n_3907 ,csa_tree_add_190_195_groupi_n_2210);
  xnor csa_tree_add_190_195_groupi_g43841(csa_tree_add_190_195_groupi_n_5393 ,csa_tree_add_190_195_groupi_n_4101 ,csa_tree_add_190_195_groupi_n_1841);
  xnor csa_tree_add_190_195_groupi_g43842(csa_tree_add_190_195_groupi_n_5392 ,csa_tree_add_190_195_groupi_n_3742 ,csa_tree_add_190_195_groupi_n_1923);
  xnor csa_tree_add_190_195_groupi_g43843(csa_tree_add_190_195_groupi_n_5391 ,csa_tree_add_190_195_groupi_n_0 ,in55[1]);
  xnor csa_tree_add_190_195_groupi_g43845(csa_tree_add_190_195_groupi_n_5389 ,csa_tree_add_190_195_groupi_n_3979 ,csa_tree_add_190_195_groupi_n_1904);
  xnor csa_tree_add_190_195_groupi_g43846(csa_tree_add_190_195_groupi_n_5388 ,csa_tree_add_190_195_groupi_n_3952 ,csa_tree_add_190_195_groupi_n_1056);
  xnor csa_tree_add_190_195_groupi_g43847(csa_tree_add_190_195_groupi_n_5387 ,csa_tree_add_190_195_groupi_n_4128 ,csa_tree_add_190_195_groupi_n_2154);
  xnor csa_tree_add_190_195_groupi_g43848(csa_tree_add_190_195_groupi_n_5385 ,csa_tree_add_190_195_groupi_n_69 ,csa_tree_add_190_195_groupi_n_1915);
  xnor csa_tree_add_190_195_groupi_g43849(csa_tree_add_190_195_groupi_n_5384 ,csa_tree_add_190_195_groupi_n_63 ,csa_tree_add_190_195_groupi_n_2002);
  xnor csa_tree_add_190_195_groupi_g43850(csa_tree_add_190_195_groupi_n_5382 ,csa_tree_add_190_195_groupi_n_3763 ,csa_tree_add_190_195_groupi_n_1715);
  xnor csa_tree_add_190_195_groupi_g43852(csa_tree_add_190_195_groupi_n_5380 ,csa_tree_add_190_195_groupi_n_4090 ,in59[13]);
  xnor csa_tree_add_190_195_groupi_g43854(csa_tree_add_190_195_groupi_n_5379 ,csa_tree_add_190_195_groupi_n_4088 ,in58[13]);
  xnor csa_tree_add_190_195_groupi_g43855(csa_tree_add_190_195_groupi_n_5378 ,csa_tree_add_190_195_groupi_n_3803 ,csa_tree_add_190_195_groupi_n_1993);
  xnor csa_tree_add_190_195_groupi_g43857(csa_tree_add_190_195_groupi_n_5375 ,csa_tree_add_190_195_groupi_n_3857 ,csa_tree_add_190_195_groupi_n_2008);
  xnor csa_tree_add_190_195_groupi_g43858(csa_tree_add_190_195_groupi_n_5374 ,csa_tree_add_190_195_groupi_n_3920 ,csa_tree_add_190_195_groupi_n_1670);
  xnor csa_tree_add_190_195_groupi_g43859(csa_tree_add_190_195_groupi_n_5373 ,csa_tree_add_190_195_groupi_n_3767 ,csa_tree_add_190_195_groupi_n_1889);
  xnor csa_tree_add_190_195_groupi_g43860(csa_tree_add_190_195_groupi_n_5371 ,csa_tree_add_190_195_groupi_n_4124 ,csa_tree_add_190_195_groupi_n_1307);
  xnor csa_tree_add_190_195_groupi_g43861(csa_tree_add_190_195_groupi_n_5369 ,csa_tree_add_190_195_groupi_n_4119 ,csa_tree_add_190_195_groupi_n_1904);
  xnor csa_tree_add_190_195_groupi_g43862(csa_tree_add_190_195_groupi_n_5367 ,csa_tree_add_190_195_groupi_n_3812 ,csa_tree_add_190_195_groupi_n_1638);
  xnor csa_tree_add_190_195_groupi_g43863(csa_tree_add_190_195_groupi_n_5366 ,csa_tree_add_190_195_groupi_n_3761 ,csa_tree_add_190_195_groupi_n_1689);
  xnor csa_tree_add_190_195_groupi_g43864(csa_tree_add_190_195_groupi_n_5365 ,csa_tree_add_190_195_groupi_n_4066 ,csa_tree_add_190_195_groupi_n_1899);
  xnor csa_tree_add_190_195_groupi_g43865(csa_tree_add_190_195_groupi_n_5364 ,csa_tree_add_190_195_groupi_n_3975 ,csa_tree_add_190_195_groupi_n_1024);
  xnor csa_tree_add_190_195_groupi_g43866(csa_tree_add_190_195_groupi_n_5362 ,csa_tree_add_190_195_groupi_n_4062 ,csa_tree_add_190_195_groupi_n_2040);
  xnor csa_tree_add_190_195_groupi_g43867(csa_tree_add_190_195_groupi_n_5360 ,csa_tree_add_190_195_groupi_n_3805 ,csa_tree_add_190_195_groupi_n_1173);
  xnor csa_tree_add_190_195_groupi_g43868(csa_tree_add_190_195_groupi_n_5358 ,csa_tree_add_190_195_groupi_n_3739 ,csa_tree_add_190_195_groupi_n_1967);
  xnor csa_tree_add_190_195_groupi_g43869(csa_tree_add_190_195_groupi_n_5356 ,csa_tree_add_190_195_groupi_n_3950 ,csa_tree_add_190_195_groupi_n_2041);
  xnor csa_tree_add_190_195_groupi_g43870(csa_tree_add_190_195_groupi_n_5355 ,csa_tree_add_190_195_groupi_n_3983 ,csa_tree_add_190_195_groupi_n_1972);
  xnor csa_tree_add_190_195_groupi_g43871(csa_tree_add_190_195_groupi_n_5353 ,csa_tree_add_190_195_groupi_n_3775 ,csa_tree_add_190_195_groupi_n_1759);
  xnor csa_tree_add_190_195_groupi_g43872(csa_tree_add_190_195_groupi_n_5352 ,csa_tree_add_190_195_groupi_n_3919 ,csa_tree_add_190_195_groupi_n_1867);
  xnor csa_tree_add_190_195_groupi_g43873(csa_tree_add_190_195_groupi_n_5351 ,csa_tree_add_190_195_groupi_n_3957 ,csa_tree_add_190_195_groupi_n_1795);
  xnor csa_tree_add_190_195_groupi_g43874(csa_tree_add_190_195_groupi_n_5350 ,csa_tree_add_190_195_groupi_n_4047 ,csa_tree_add_190_195_groupi_n_1574);
  xnor csa_tree_add_190_195_groupi_g43875(csa_tree_add_190_195_groupi_n_5349 ,csa_tree_add_190_195_groupi_n_4079 ,csa_tree_add_190_195_groupi_n_2001);
  xnor csa_tree_add_190_195_groupi_g43876(csa_tree_add_190_195_groupi_n_5348 ,csa_tree_add_190_195_groupi_n_3967 ,csa_tree_add_190_195_groupi_n_1230);
  xnor csa_tree_add_190_195_groupi_g43877(csa_tree_add_190_195_groupi_n_5347 ,csa_tree_add_190_195_groupi_n_4131 ,csa_tree_add_190_195_groupi_n_1990);
  xnor csa_tree_add_190_195_groupi_g43878(csa_tree_add_190_195_groupi_n_5345 ,csa_tree_add_190_195_groupi_n_3847 ,csa_tree_add_190_195_groupi_n_1185);
  xnor csa_tree_add_190_195_groupi_g43879(csa_tree_add_190_195_groupi_n_5344 ,csa_tree_add_190_195_groupi_n_4063 ,csa_tree_add_190_195_groupi_n_1658);
  xnor csa_tree_add_190_195_groupi_g43880(csa_tree_add_190_195_groupi_n_5342 ,csa_tree_add_190_195_groupi_n_4019 ,csa_tree_add_190_195_groupi_n_1676);
  xnor csa_tree_add_190_195_groupi_g43881(csa_tree_add_190_195_groupi_n_5340 ,csa_tree_add_190_195_groupi_n_3734 ,csa_tree_add_190_195_groupi_n_1931);
  xnor csa_tree_add_190_195_groupi_g43882(csa_tree_add_190_195_groupi_n_5338 ,csa_tree_add_190_195_groupi_n_3922 ,csa_tree_add_190_195_groupi_n_2082);
  xnor csa_tree_add_190_195_groupi_g43883(csa_tree_add_190_195_groupi_n_5336 ,csa_tree_add_190_195_groupi_n_3737 ,csa_tree_add_190_195_groupi_n_2049);
  xnor csa_tree_add_190_195_groupi_g43884(csa_tree_add_190_195_groupi_n_5335 ,csa_tree_add_190_195_groupi_n_4086 ,csa_tree_add_190_195_groupi_n_1901);
  xnor csa_tree_add_190_195_groupi_g43885(csa_tree_add_190_195_groupi_n_5333 ,csa_tree_add_190_195_groupi_n_3810 ,csa_tree_add_190_195_groupi_n_1785);
  xnor csa_tree_add_190_195_groupi_g43886(csa_tree_add_190_195_groupi_n_5331 ,csa_tree_add_190_195_groupi_n_3833 ,csa_tree_add_190_195_groupi_n_1761);
  xnor csa_tree_add_190_195_groupi_g43887(csa_tree_add_190_195_groupi_n_5329 ,csa_tree_add_190_195_groupi_n_4107 ,csa_tree_add_190_195_groupi_n_1810);
  xnor csa_tree_add_190_195_groupi_g43888(csa_tree_add_190_195_groupi_n_5328 ,csa_tree_add_190_195_groupi_n_44 ,csa_tree_add_190_195_groupi_n_1948);
  xnor csa_tree_add_190_195_groupi_g43889(csa_tree_add_190_195_groupi_n_5326 ,csa_tree_add_190_195_groupi_n_3839 ,csa_tree_add_190_195_groupi_n_1973);
  xnor csa_tree_add_190_195_groupi_g43890(csa_tree_add_190_195_groupi_n_5325 ,csa_tree_add_190_195_groupi_n_3894 ,csa_tree_add_190_195_groupi_n_1873);
  xnor csa_tree_add_190_195_groupi_g43891(csa_tree_add_190_195_groupi_n_5323 ,csa_tree_add_190_195_groupi_n_3992 ,csa_tree_add_190_195_groupi_n_1932);
  xnor csa_tree_add_190_195_groupi_g43892(csa_tree_add_190_195_groupi_n_5322 ,csa_tree_add_190_195_groupi_n_4042 ,csa_tree_add_190_195_groupi_n_2118);
  xnor csa_tree_add_190_195_groupi_g43893(csa_tree_add_190_195_groupi_n_5321 ,csa_tree_add_190_195_groupi_n_3997 ,csa_tree_add_190_195_groupi_n_2000);
  xnor csa_tree_add_190_195_groupi_g43894(csa_tree_add_190_195_groupi_n_5320 ,csa_tree_add_190_195_groupi_n_4121 ,csa_tree_add_190_195_groupi_n_1992);
  xnor csa_tree_add_190_195_groupi_g43895(csa_tree_add_190_195_groupi_n_5318 ,csa_tree_add_190_195_groupi_n_3749 ,csa_tree_add_190_195_groupi_n_2053);
  xnor csa_tree_add_190_195_groupi_g43896(csa_tree_add_190_195_groupi_n_5315 ,csa_tree_add_190_195_groupi_n_4037 ,csa_tree_add_190_195_groupi_n_1767);
  xnor csa_tree_add_190_195_groupi_g43897(csa_tree_add_190_195_groupi_n_5313 ,csa_tree_add_190_195_groupi_n_4083 ,in58[0]);
  xnor csa_tree_add_190_195_groupi_g43898(csa_tree_add_190_195_groupi_n_5312 ,csa_tree_add_190_195_groupi_n_3990 ,csa_tree_add_190_195_groupi_n_1700);
  xnor csa_tree_add_190_195_groupi_g43899(csa_tree_add_190_195_groupi_n_5311 ,csa_tree_add_190_195_groupi_n_82 ,csa_tree_add_190_195_groupi_n_1677);
  xnor csa_tree_add_190_195_groupi_g43900(csa_tree_add_190_195_groupi_n_5310 ,csa_tree_add_190_195_groupi_n_3865 ,in55[9]);
  xnor csa_tree_add_190_195_groupi_g43902(csa_tree_add_190_195_groupi_n_5306 ,csa_tree_add_190_195_groupi_n_4055 ,csa_tree_add_190_195_groupi_n_2674);
  xnor csa_tree_add_190_195_groupi_g43904(csa_tree_add_190_195_groupi_n_5304 ,csa_tree_add_190_195_groupi_n_4125 ,csa_tree_add_190_195_groupi_n_1941);
  xnor csa_tree_add_190_195_groupi_g43905(csa_tree_add_190_195_groupi_n_5302 ,csa_tree_add_190_195_groupi_n_3746 ,csa_tree_add_190_195_groupi_n_1677);
  xnor csa_tree_add_190_195_groupi_g43906(csa_tree_add_190_195_groupi_n_5301 ,csa_tree_add_190_195_groupi_n_3759 ,csa_tree_add_190_195_groupi_n_1718);
  xnor csa_tree_add_190_195_groupi_g43907(csa_tree_add_190_195_groupi_n_5299 ,csa_tree_add_190_195_groupi_n_3822 ,csa_tree_add_190_195_groupi_n_1701);
  xnor csa_tree_add_190_195_groupi_g43908(csa_tree_add_190_195_groupi_n_5298 ,csa_tree_add_190_195_groupi_n_3796 ,csa_tree_add_190_195_groupi_n_2213);
  xnor csa_tree_add_190_195_groupi_g43909(csa_tree_add_190_195_groupi_n_5297 ,csa_tree_add_190_195_groupi_n_3826 ,in55[11]);
  xnor csa_tree_add_190_195_groupi_g43910(csa_tree_add_190_195_groupi_n_5296 ,csa_tree_add_190_195_groupi_n_3 ,csa_tree_add_190_195_groupi_n_1883);
  xnor csa_tree_add_190_195_groupi_g43911(csa_tree_add_190_195_groupi_n_5294 ,csa_tree_add_190_195_groupi_n_4085 ,csa_tree_add_190_195_groupi_n_1698);
  xnor csa_tree_add_190_195_groupi_g43912(csa_tree_add_190_195_groupi_n_5292 ,csa_tree_add_190_195_groupi_n_3852 ,in59[0]);
  xnor csa_tree_add_190_195_groupi_g43913(csa_tree_add_190_195_groupi_n_5291 ,csa_tree_add_190_195_groupi_n_4032 ,csa_tree_add_190_195_groupi_n_2211);
  xnor csa_tree_add_190_195_groupi_g43915(csa_tree_add_190_195_groupi_n_5289 ,csa_tree_add_190_195_groupi_n_4023 ,csa_tree_add_190_195_groupi_n_1766);
  xnor csa_tree_add_190_195_groupi_g43916(csa_tree_add_190_195_groupi_n_5287 ,csa_tree_add_190_195_groupi_n_3858 ,csa_tree_add_190_195_groupi_n_1842);
  xnor csa_tree_add_190_195_groupi_g43917(csa_tree_add_190_195_groupi_n_5286 ,csa_tree_add_190_195_groupi_n_3736 ,csa_tree_add_190_195_groupi_n_1936);
  xnor csa_tree_add_190_195_groupi_g43918(csa_tree_add_190_195_groupi_n_5285 ,csa_tree_add_190_195_groupi_n_3928 ,csa_tree_add_190_195_groupi_n_1696);
  xnor csa_tree_add_190_195_groupi_g43919(csa_tree_add_190_195_groupi_n_5283 ,csa_tree_add_190_195_groupi_n_3208 ,csa_tree_add_190_195_groupi_n_3841);
  xnor csa_tree_add_190_195_groupi_g43920(csa_tree_add_190_195_groupi_n_5282 ,csa_tree_add_190_195_groupi_n_4132 ,csa_tree_add_190_195_groupi_n_488);
  xnor csa_tree_add_190_195_groupi_g43921(csa_tree_add_190_195_groupi_n_5281 ,csa_tree_add_190_195_groupi_n_3994 ,csa_tree_add_190_195_groupi_n_1661);
  xnor csa_tree_add_190_195_groupi_g43922(csa_tree_add_190_195_groupi_n_5280 ,csa_tree_add_190_195_groupi_n_3962 ,csa_tree_add_190_195_groupi_n_1830);
  xnor csa_tree_add_190_195_groupi_g43923(csa_tree_add_190_195_groupi_n_5278 ,csa_tree_add_190_195_groupi_n_3831 ,in57[13]);
  xnor csa_tree_add_190_195_groupi_g43924(csa_tree_add_190_195_groupi_n_5277 ,csa_tree_add_190_195_groupi_n_4057 ,csa_tree_add_190_195_groupi_n_1742);
  xnor csa_tree_add_190_195_groupi_g43925(csa_tree_add_190_195_groupi_n_5275 ,csa_tree_add_190_195_groupi_n_3988 ,in60[7]);
  xnor csa_tree_add_190_195_groupi_g43926(csa_tree_add_190_195_groupi_n_5274 ,csa_tree_add_190_195_groupi_n_3732 ,csa_tree_add_190_195_groupi_n_1745);
  xnor csa_tree_add_190_195_groupi_g43927(csa_tree_add_190_195_groupi_n_5272 ,csa_tree_add_190_195_groupi_n_4108 ,csa_tree_add_190_195_groupi_n_1652);
  xnor csa_tree_add_190_195_groupi_g43928(csa_tree_add_190_195_groupi_n_5270 ,csa_tree_add_190_195_groupi_n_3814 ,csa_tree_add_190_195_groupi_n_1749);
  xnor csa_tree_add_190_195_groupi_g43929(csa_tree_add_190_195_groupi_n_5269 ,csa_tree_add_190_195_groupi_n_4082 ,csa_tree_add_190_195_groupi_n_1603);
  xnor csa_tree_add_190_195_groupi_g43930(csa_tree_add_190_195_groupi_n_5268 ,csa_tree_add_190_195_groupi_n_3955 ,csa_tree_add_190_195_groupi_n_1894);
  xnor csa_tree_add_190_195_groupi_g43931(csa_tree_add_190_195_groupi_n_5266 ,csa_tree_add_190_195_groupi_n_3993 ,csa_tree_add_190_195_groupi_n_1050);
  xnor csa_tree_add_190_195_groupi_g43932(csa_tree_add_190_195_groupi_n_5265 ,csa_tree_add_190_195_groupi_n_4017 ,csa_tree_add_190_195_groupi_n_2000);
  xnor csa_tree_add_190_195_groupi_g43933(csa_tree_add_190_195_groupi_n_5263 ,csa_tree_add_190_195_groupi_n_3836 ,in57[10]);
  xnor csa_tree_add_190_195_groupi_g43934(csa_tree_add_190_195_groupi_n_5262 ,csa_tree_add_190_195_groupi_n_3901 ,csa_tree_add_190_195_groupi_n_1871);
  xnor csa_tree_add_190_195_groupi_g43935(csa_tree_add_190_195_groupi_n_5260 ,csa_tree_add_190_195_groupi_n_4070 ,csa_tree_add_190_195_groupi_n_1711);
  xnor csa_tree_add_190_195_groupi_g43936(csa_tree_add_190_195_groupi_n_5259 ,csa_tree_add_190_195_groupi_n_4068 ,csa_tree_add_190_195_groupi_n_1168);
  xnor csa_tree_add_190_195_groupi_g43937(csa_tree_add_190_195_groupi_n_5258 ,csa_tree_add_190_195_groupi_n_3959 ,csa_tree_add_190_195_groupi_n_1015);
  xnor csa_tree_add_190_195_groupi_g43938(csa_tree_add_190_195_groupi_n_5257 ,csa_tree_add_190_195_groupi_n_3902 ,csa_tree_add_190_195_groupi_n_1186);
  xnor csa_tree_add_190_195_groupi_g43939(csa_tree_add_190_195_groupi_n_5256 ,csa_tree_add_190_195_groupi_n_4008 ,csa_tree_add_190_195_groupi_n_990);
  xnor csa_tree_add_190_195_groupi_g43940(csa_tree_add_190_195_groupi_n_5255 ,csa_tree_add_190_195_groupi_n_4095 ,csa_tree_add_190_195_groupi_n_963);
  xnor csa_tree_add_190_195_groupi_g43941(csa_tree_add_190_195_groupi_n_5253 ,csa_tree_add_190_195_groupi_n_4029 ,csa_tree_add_190_195_groupi_n_1598);
  xnor csa_tree_add_190_195_groupi_g43942(csa_tree_add_190_195_groupi_n_5252 ,csa_tree_add_190_195_groupi_n_4112 ,csa_tree_add_190_195_groupi_n_1886);
  xnor csa_tree_add_190_195_groupi_g43944(csa_tree_add_190_195_groupi_n_5250 ,csa_tree_add_190_195_groupi_n_3890 ,csa_tree_add_190_195_groupi_n_1896);
  xnor csa_tree_add_190_195_groupi_g43945(csa_tree_add_190_195_groupi_n_5248 ,csa_tree_add_190_195_groupi_n_3939 ,csa_tree_add_190_195_groupi_n_1626);
  xnor csa_tree_add_190_195_groupi_g43946(csa_tree_add_190_195_groupi_n_5245 ,csa_tree_add_190_195_groupi_n_3766 ,csa_tree_add_190_195_groupi_n_1922);
  xnor csa_tree_add_190_195_groupi_g43947(csa_tree_add_190_195_groupi_n_5244 ,csa_tree_add_190_195_groupi_n_3995 ,csa_tree_add_190_195_groupi_n_1893);
  xnor csa_tree_add_190_195_groupi_g43948(csa_tree_add_190_195_groupi_n_5243 ,csa_tree_add_190_195_groupi_n_4022 ,csa_tree_add_190_195_groupi_n_1997);
  xnor csa_tree_add_190_195_groupi_g43949(csa_tree_add_190_195_groupi_n_5242 ,csa_tree_add_190_195_groupi_n_4025 ,csa_tree_add_190_195_groupi_n_1935);
  xnor csa_tree_add_190_195_groupi_g43950(csa_tree_add_190_195_groupi_n_5241 ,csa_tree_add_190_195_groupi_n_3900 ,csa_tree_add_190_195_groupi_n_2213);
  xnor csa_tree_add_190_195_groupi_g43951(csa_tree_add_190_195_groupi_n_5240 ,csa_tree_add_190_195_groupi_n_4072 ,csa_tree_add_190_195_groupi_n_1711);
  xnor csa_tree_add_190_195_groupi_g43952(csa_tree_add_190_195_groupi_n_5239 ,csa_tree_add_190_195_groupi_n_4103 ,csa_tree_add_190_195_groupi_n_1942);
  xnor csa_tree_add_190_195_groupi_g43953(csa_tree_add_190_195_groupi_n_5238 ,csa_tree_add_190_195_groupi_n_3752 ,csa_tree_add_190_195_groupi_n_2063);
  xnor csa_tree_add_190_195_groupi_g43954(csa_tree_add_190_195_groupi_n_5236 ,csa_tree_add_190_195_groupi_n_3817 ,csa_tree_add_190_195_groupi_n_1899);
  xnor csa_tree_add_190_195_groupi_g43955(csa_tree_add_190_195_groupi_n_5234 ,csa_tree_add_190_195_groupi_n_4132 ,csa_tree_add_190_195_groupi_n_1390);
  xnor csa_tree_add_190_195_groupi_g43956(csa_tree_add_190_195_groupi_n_5233 ,csa_tree_add_190_195_groupi_n_3968 ,csa_tree_add_190_195_groupi_n_1887);
  xnor csa_tree_add_190_195_groupi_g43957(csa_tree_add_190_195_groupi_n_5232 ,csa_tree_add_190_195_groupi_n_3879 ,csa_tree_add_190_195_groupi_n_1774);
  xnor csa_tree_add_190_195_groupi_g43958(csa_tree_add_190_195_groupi_n_5230 ,csa_tree_add_190_195_groupi_n_4074 ,csa_tree_add_190_195_groupi_n_1891);
  xnor csa_tree_add_190_195_groupi_g43959(csa_tree_add_190_195_groupi_n_5228 ,csa_tree_add_190_195_groupi_n_3859 ,csa_tree_add_190_195_groupi_n_1765);
  xnor csa_tree_add_190_195_groupi_g43960(csa_tree_add_190_195_groupi_n_5227 ,csa_tree_add_190_195_groupi_n_3945 ,csa_tree_add_190_195_groupi_n_1890);
  xnor csa_tree_add_190_195_groupi_g43961(csa_tree_add_190_195_groupi_n_5225 ,csa_tree_add_190_195_groupi_n_3906 ,csa_tree_add_190_195_groupi_n_1047);
  xnor csa_tree_add_190_195_groupi_g43962(csa_tree_add_190_195_groupi_n_5224 ,csa_tree_add_190_195_groupi_n_3778 ,csa_tree_add_190_195_groupi_n_1688);
  xnor csa_tree_add_190_195_groupi_g43963(csa_tree_add_190_195_groupi_n_5223 ,csa_tree_add_190_195_groupi_n_4128 ,csa_tree_add_190_195_groupi_n_2090);
  xnor csa_tree_add_190_195_groupi_g43965(csa_tree_add_190_195_groupi_n_5220 ,csa_tree_add_190_195_groupi_n_4065 ,csa_tree_add_190_195_groupi_n_2052);
  xnor csa_tree_add_190_195_groupi_g43966(csa_tree_add_190_195_groupi_n_5218 ,csa_tree_add_190_195_groupi_n_3964 ,csa_tree_add_190_195_groupi_n_1830);
  xnor csa_tree_add_190_195_groupi_g43967(csa_tree_add_190_195_groupi_n_5217 ,csa_tree_add_190_195_groupi_n_3935 ,csa_tree_add_190_195_groupi_n_506);
  xnor csa_tree_add_190_195_groupi_g43968(csa_tree_add_190_195_groupi_n_5216 ,csa_tree_add_190_195_groupi_n_3954 ,csa_tree_add_190_195_groupi_n_2054);
  xnor csa_tree_add_190_195_groupi_g43969(csa_tree_add_190_195_groupi_n_5214 ,csa_tree_add_190_195_groupi_n_4061 ,csa_tree_add_190_195_groupi_n_1122);
  xnor csa_tree_add_190_195_groupi_g43970(csa_tree_add_190_195_groupi_n_5212 ,csa_tree_add_190_195_groupi_n_3874 ,in60[2]);
  xnor csa_tree_add_190_195_groupi_g43971(csa_tree_add_190_195_groupi_n_5210 ,csa_tree_add_190_195_groupi_n_4001 ,csa_tree_add_190_195_groupi_n_1987);
  xnor csa_tree_add_190_195_groupi_g43972(csa_tree_add_190_195_groupi_n_5209 ,csa_tree_add_190_195_groupi_n_3892 ,csa_tree_add_190_195_groupi_n_2090);
  xnor csa_tree_add_190_195_groupi_g43973(csa_tree_add_190_195_groupi_n_5207 ,csa_tree_add_190_195_groupi_n_3986 ,csa_tree_add_190_195_groupi_n_1911);
  xnor csa_tree_add_190_195_groupi_g43974(csa_tree_add_190_195_groupi_n_5206 ,csa_tree_add_190_195_groupi_n_3827 ,in55[10]);
  xnor csa_tree_add_190_195_groupi_g43975(csa_tree_add_190_195_groupi_n_5205 ,csa_tree_add_190_195_groupi_n_3867 ,csa_tree_add_190_195_groupi_n_499);
  xnor csa_tree_add_190_195_groupi_g43976(csa_tree_add_190_195_groupi_n_5203 ,csa_tree_add_190_195_groupi_n_3862 ,in58[15]);
  xnor csa_tree_add_190_195_groupi_g43977(csa_tree_add_190_195_groupi_n_5202 ,csa_tree_add_190_195_groupi_n_4013 ,csa_tree_add_190_195_groupi_n_1293);
  xnor csa_tree_add_190_195_groupi_g43978(csa_tree_add_190_195_groupi_n_5201 ,csa_tree_add_190_195_groupi_n_3845 ,in55[12]);
  xnor csa_tree_add_190_195_groupi_g43979(csa_tree_add_190_195_groupi_n_5200 ,csa_tree_add_190_195_groupi_n_3940 ,csa_tree_add_190_195_groupi_n_1901);
  xnor csa_tree_add_190_195_groupi_g43980(csa_tree_add_190_195_groupi_n_5199 ,csa_tree_add_190_195_groupi_n_4092 ,csa_tree_add_190_195_groupi_n_987);
  xnor csa_tree_add_190_195_groupi_g43981(csa_tree_add_190_195_groupi_n_5198 ,csa_tree_add_190_195_groupi_n_3893 ,csa_tree_add_190_195_groupi_n_1585);
  xnor csa_tree_add_190_195_groupi_g43982(csa_tree_add_190_195_groupi_n_5196 ,csa_tree_add_190_195_groupi_n_3774 ,csa_tree_add_190_195_groupi_n_1581);
  xnor csa_tree_add_190_195_groupi_g43984(csa_tree_add_190_195_groupi_n_5193 ,csa_tree_add_190_195_groupi_n_3973 ,csa_tree_add_190_195_groupi_n_1603);
  xnor csa_tree_add_190_195_groupi_g43985(csa_tree_add_190_195_groupi_n_5191 ,csa_tree_add_190_195_groupi_n_3809 ,csa_tree_add_190_195_groupi_n_1688);
  xnor csa_tree_add_190_195_groupi_g43986(csa_tree_add_190_195_groupi_n_5189 ,csa_tree_add_190_195_groupi_n_4007 ,csa_tree_add_190_195_groupi_n_1779);
  xnor csa_tree_add_190_195_groupi_g43987(csa_tree_add_190_195_groupi_n_5187 ,csa_tree_add_190_195_groupi_n_3937 ,csa_tree_add_190_195_groupi_n_1853);
  xnor csa_tree_add_190_195_groupi_g43988(csa_tree_add_190_195_groupi_n_5185 ,csa_tree_add_190_195_groupi_n_3876 ,csa_tree_add_190_195_groupi_n_1617);
  xnor csa_tree_add_190_195_groupi_g43989(csa_tree_add_190_195_groupi_n_5183 ,csa_tree_add_190_195_groupi_n_4036 ,csa_tree_add_190_195_groupi_n_1755);
  xnor csa_tree_add_190_195_groupi_g43990(csa_tree_add_190_195_groupi_n_5181 ,csa_tree_add_190_195_groupi_n_3777 ,csa_tree_add_190_195_groupi_n_1668);
  not csa_tree_add_190_195_groupi_g43992(csa_tree_add_190_195_groupi_n_5171 ,csa_tree_add_190_195_groupi_n_5170);
  not csa_tree_add_190_195_groupi_g43993(csa_tree_add_190_195_groupi_n_5165 ,csa_tree_add_190_195_groupi_n_5164);
  not csa_tree_add_190_195_groupi_g43995(csa_tree_add_190_195_groupi_n_5158 ,csa_tree_add_190_195_groupi_n_5157);
  not csa_tree_add_190_195_groupi_g43997(csa_tree_add_190_195_groupi_n_5124 ,csa_tree_add_190_195_groupi_n_5123);
  not csa_tree_add_190_195_groupi_g43998(csa_tree_add_190_195_groupi_n_5111 ,csa_tree_add_190_195_groupi_n_5110);
  not csa_tree_add_190_195_groupi_g43999(csa_tree_add_190_195_groupi_n_5109 ,csa_tree_add_190_195_groupi_n_5108);
  not csa_tree_add_190_195_groupi_g44000(csa_tree_add_190_195_groupi_n_5095 ,csa_tree_add_190_195_groupi_n_5096);
  not csa_tree_add_190_195_groupi_g44001(csa_tree_add_190_195_groupi_n_5094 ,csa_tree_add_190_195_groupi_n_5093);
  not csa_tree_add_190_195_groupi_g44002(csa_tree_add_190_195_groupi_n_5091 ,csa_tree_add_190_195_groupi_n_5092);
  not csa_tree_add_190_195_groupi_g44003(csa_tree_add_190_195_groupi_n_5089 ,csa_tree_add_190_195_groupi_n_5088);
  not csa_tree_add_190_195_groupi_g44004(csa_tree_add_190_195_groupi_n_5086 ,csa_tree_add_190_195_groupi_n_5085);
  not csa_tree_add_190_195_groupi_g44005(csa_tree_add_190_195_groupi_n_5083 ,csa_tree_add_190_195_groupi_n_5084);
  not csa_tree_add_190_195_groupi_g44006(csa_tree_add_190_195_groupi_n_5081 ,csa_tree_add_190_195_groupi_n_5082);
  not csa_tree_add_190_195_groupi_g44007(csa_tree_add_190_195_groupi_n_5078 ,csa_tree_add_190_195_groupi_n_5079);
  not csa_tree_add_190_195_groupi_g44008(csa_tree_add_190_195_groupi_n_5077 ,csa_tree_add_190_195_groupi_n_5076);
  not csa_tree_add_190_195_groupi_g44009(csa_tree_add_190_195_groupi_n_5074 ,csa_tree_add_190_195_groupi_n_5075);
  not csa_tree_add_190_195_groupi_g44010(csa_tree_add_190_195_groupi_n_5073 ,csa_tree_add_190_195_groupi_n_5072);
  not csa_tree_add_190_195_groupi_g44011(csa_tree_add_190_195_groupi_n_5070 ,csa_tree_add_190_195_groupi_n_5071);
  not csa_tree_add_190_195_groupi_g44012(csa_tree_add_190_195_groupi_n_5068 ,csa_tree_add_190_195_groupi_n_5069);
  not csa_tree_add_190_195_groupi_g44013(csa_tree_add_190_195_groupi_n_5066 ,csa_tree_add_190_195_groupi_n_5067);
  not csa_tree_add_190_195_groupi_g44014(csa_tree_add_190_195_groupi_n_5063 ,csa_tree_add_190_195_groupi_n_5064);
  not csa_tree_add_190_195_groupi_g44015(csa_tree_add_190_195_groupi_n_5061 ,csa_tree_add_190_195_groupi_n_5062);
  not csa_tree_add_190_195_groupi_g44016(csa_tree_add_190_195_groupi_n_5059 ,csa_tree_add_190_195_groupi_n_5060);
  not csa_tree_add_190_195_groupi_g44017(csa_tree_add_190_195_groupi_n_5057 ,csa_tree_add_190_195_groupi_n_5058);
  not csa_tree_add_190_195_groupi_g44018(csa_tree_add_190_195_groupi_n_5054 ,csa_tree_add_190_195_groupi_n_5055);
  not csa_tree_add_190_195_groupi_g44019(csa_tree_add_190_195_groupi_n_5052 ,csa_tree_add_190_195_groupi_n_5053);
  not csa_tree_add_190_195_groupi_g44020(csa_tree_add_190_195_groupi_n_5050 ,csa_tree_add_190_195_groupi_n_5051);
  not csa_tree_add_190_195_groupi_g44021(csa_tree_add_190_195_groupi_n_5048 ,csa_tree_add_190_195_groupi_n_5049);
  not csa_tree_add_190_195_groupi_g44022(csa_tree_add_190_195_groupi_n_5046 ,csa_tree_add_190_195_groupi_n_5047);
  not csa_tree_add_190_195_groupi_g44023(csa_tree_add_190_195_groupi_n_5044 ,csa_tree_add_190_195_groupi_n_5045);
  not csa_tree_add_190_195_groupi_g44024(csa_tree_add_190_195_groupi_n_5042 ,csa_tree_add_190_195_groupi_n_5043);
  not csa_tree_add_190_195_groupi_g44025(csa_tree_add_190_195_groupi_n_5040 ,csa_tree_add_190_195_groupi_n_5041);
  not csa_tree_add_190_195_groupi_g44026(csa_tree_add_190_195_groupi_n_5038 ,csa_tree_add_190_195_groupi_n_5037);
  not csa_tree_add_190_195_groupi_g44027(csa_tree_add_190_195_groupi_n_5035 ,csa_tree_add_190_195_groupi_n_5036);
  not csa_tree_add_190_195_groupi_g44028(csa_tree_add_190_195_groupi_n_5033 ,csa_tree_add_190_195_groupi_n_5034);
  not csa_tree_add_190_195_groupi_g44029(csa_tree_add_190_195_groupi_n_5030 ,csa_tree_add_190_195_groupi_n_5031);
  not csa_tree_add_190_195_groupi_g44030(csa_tree_add_190_195_groupi_n_5028 ,csa_tree_add_190_195_groupi_n_5029);
  not csa_tree_add_190_195_groupi_g44031(csa_tree_add_190_195_groupi_n_5026 ,csa_tree_add_190_195_groupi_n_5027);
  not csa_tree_add_190_195_groupi_g44032(csa_tree_add_190_195_groupi_n_5023 ,csa_tree_add_190_195_groupi_n_5024);
  not csa_tree_add_190_195_groupi_g44033(csa_tree_add_190_195_groupi_n_5021 ,csa_tree_add_190_195_groupi_n_5022);
  not csa_tree_add_190_195_groupi_g44034(csa_tree_add_190_195_groupi_n_5019 ,csa_tree_add_190_195_groupi_n_5020);
  not csa_tree_add_190_195_groupi_g44035(csa_tree_add_190_195_groupi_n_5015 ,csa_tree_add_190_195_groupi_n_5016);
  not csa_tree_add_190_195_groupi_g44036(csa_tree_add_190_195_groupi_n_5013 ,csa_tree_add_190_195_groupi_n_5014);
  not csa_tree_add_190_195_groupi_g44037(csa_tree_add_190_195_groupi_n_5011 ,csa_tree_add_190_195_groupi_n_5010);
  not csa_tree_add_190_195_groupi_g44038(csa_tree_add_190_195_groupi_n_5008 ,csa_tree_add_190_195_groupi_n_5009);
  not csa_tree_add_190_195_groupi_g44039(csa_tree_add_190_195_groupi_n_5006 ,csa_tree_add_190_195_groupi_n_5007);
  not csa_tree_add_190_195_groupi_g44040(csa_tree_add_190_195_groupi_n_5001 ,csa_tree_add_190_195_groupi_n_5002);
  not csa_tree_add_190_195_groupi_g44041(csa_tree_add_190_195_groupi_n_5000 ,csa_tree_add_190_195_groupi_n_4999);
  not csa_tree_add_190_195_groupi_g44042(csa_tree_add_190_195_groupi_n_4997 ,csa_tree_add_190_195_groupi_n_4998);
  not csa_tree_add_190_195_groupi_g44043(csa_tree_add_190_195_groupi_n_4995 ,csa_tree_add_190_195_groupi_n_4996);
  not csa_tree_add_190_195_groupi_g44044(csa_tree_add_190_195_groupi_n_4993 ,csa_tree_add_190_195_groupi_n_4994);
  not csa_tree_add_190_195_groupi_g44045(csa_tree_add_190_195_groupi_n_4990 ,csa_tree_add_190_195_groupi_n_4991);
  not csa_tree_add_190_195_groupi_g44046(csa_tree_add_190_195_groupi_n_4989 ,csa_tree_add_190_195_groupi_n_4988);
  not csa_tree_add_190_195_groupi_g44047(csa_tree_add_190_195_groupi_n_4984 ,csa_tree_add_190_195_groupi_n_4985);
  not csa_tree_add_190_195_groupi_g44048(csa_tree_add_190_195_groupi_n_4982 ,csa_tree_add_190_195_groupi_n_4983);
  not csa_tree_add_190_195_groupi_g44049(csa_tree_add_190_195_groupi_n_4980 ,csa_tree_add_190_195_groupi_n_4981);
  not csa_tree_add_190_195_groupi_g44050(csa_tree_add_190_195_groupi_n_4976 ,csa_tree_add_190_195_groupi_n_4977);
  not csa_tree_add_190_195_groupi_g44051(csa_tree_add_190_195_groupi_n_4974 ,csa_tree_add_190_195_groupi_n_4975);
  not csa_tree_add_190_195_groupi_g44052(csa_tree_add_190_195_groupi_n_4972 ,csa_tree_add_190_195_groupi_n_4973);
  not csa_tree_add_190_195_groupi_g44053(csa_tree_add_190_195_groupi_n_4970 ,csa_tree_add_190_195_groupi_n_4971);
  not csa_tree_add_190_195_groupi_g44054(csa_tree_add_190_195_groupi_n_4968 ,csa_tree_add_190_195_groupi_n_4969);
  not csa_tree_add_190_195_groupi_g44055(csa_tree_add_190_195_groupi_n_4965 ,csa_tree_add_190_195_groupi_n_4966);
  not csa_tree_add_190_195_groupi_g44056(csa_tree_add_190_195_groupi_n_4964 ,csa_tree_add_190_195_groupi_n_4963);
  not csa_tree_add_190_195_groupi_g44057(csa_tree_add_190_195_groupi_n_4961 ,csa_tree_add_190_195_groupi_n_4962);
  not csa_tree_add_190_195_groupi_g44058(csa_tree_add_190_195_groupi_n_4959 ,csa_tree_add_190_195_groupi_n_4960);
  not csa_tree_add_190_195_groupi_g44059(csa_tree_add_190_195_groupi_n_4956 ,csa_tree_add_190_195_groupi_n_4957);
  not csa_tree_add_190_195_groupi_g44060(csa_tree_add_190_195_groupi_n_4953 ,csa_tree_add_190_195_groupi_n_4954);
  not csa_tree_add_190_195_groupi_g44061(csa_tree_add_190_195_groupi_n_4952 ,csa_tree_add_190_195_groupi_n_4951);
  not csa_tree_add_190_195_groupi_g44062(csa_tree_add_190_195_groupi_n_4949 ,csa_tree_add_190_195_groupi_n_4950);
  not csa_tree_add_190_195_groupi_g44063(csa_tree_add_190_195_groupi_n_4947 ,csa_tree_add_190_195_groupi_n_4948);
  not csa_tree_add_190_195_groupi_g44064(csa_tree_add_190_195_groupi_n_4945 ,csa_tree_add_190_195_groupi_n_4946);
  not csa_tree_add_190_195_groupi_g44065(csa_tree_add_190_195_groupi_n_4942 ,csa_tree_add_190_195_groupi_n_4943);
  not csa_tree_add_190_195_groupi_g44066(csa_tree_add_190_195_groupi_n_4940 ,csa_tree_add_190_195_groupi_n_4941);
  not csa_tree_add_190_195_groupi_g44067(csa_tree_add_190_195_groupi_n_4939 ,csa_tree_add_190_195_groupi_n_4938);
  not csa_tree_add_190_195_groupi_g44068(csa_tree_add_190_195_groupi_n_4936 ,csa_tree_add_190_195_groupi_n_4937);
  not csa_tree_add_190_195_groupi_g44069(csa_tree_add_190_195_groupi_n_4935 ,csa_tree_add_190_195_groupi_n_4934);
  not csa_tree_add_190_195_groupi_g44070(csa_tree_add_190_195_groupi_n_4932 ,csa_tree_add_190_195_groupi_n_4933);
  not csa_tree_add_190_195_groupi_g44071(csa_tree_add_190_195_groupi_n_4929 ,csa_tree_add_190_195_groupi_n_4930);
  not csa_tree_add_190_195_groupi_g44072(csa_tree_add_190_195_groupi_n_4927 ,csa_tree_add_190_195_groupi_n_4926);
  not csa_tree_add_190_195_groupi_g44073(csa_tree_add_190_195_groupi_n_4923 ,csa_tree_add_190_195_groupi_n_4924);
  not csa_tree_add_190_195_groupi_g44074(csa_tree_add_190_195_groupi_n_4921 ,csa_tree_add_190_195_groupi_n_4922);
  not csa_tree_add_190_195_groupi_g44075(csa_tree_add_190_195_groupi_n_4919 ,csa_tree_add_190_195_groupi_n_4920);
  not csa_tree_add_190_195_groupi_g44076(csa_tree_add_190_195_groupi_n_4914 ,csa_tree_add_190_195_groupi_n_4915);
  not csa_tree_add_190_195_groupi_g44077(csa_tree_add_190_195_groupi_n_4912 ,csa_tree_add_190_195_groupi_n_4913);
  not csa_tree_add_190_195_groupi_g44078(csa_tree_add_190_195_groupi_n_4910 ,csa_tree_add_190_195_groupi_n_4911);
  not csa_tree_add_190_195_groupi_g44079(csa_tree_add_190_195_groupi_n_4905 ,csa_tree_add_190_195_groupi_n_4906);
  not csa_tree_add_190_195_groupi_g44080(csa_tree_add_190_195_groupi_n_4902 ,csa_tree_add_190_195_groupi_n_4903);
  not csa_tree_add_190_195_groupi_g44081(csa_tree_add_190_195_groupi_n_4900 ,csa_tree_add_190_195_groupi_n_4901);
  not csa_tree_add_190_195_groupi_g44082(csa_tree_add_190_195_groupi_n_4895 ,csa_tree_add_190_195_groupi_n_4896);
  not csa_tree_add_190_195_groupi_g44083(csa_tree_add_190_195_groupi_n_4889 ,csa_tree_add_190_195_groupi_n_4890);
  not csa_tree_add_190_195_groupi_g44084(csa_tree_add_190_195_groupi_n_4884 ,csa_tree_add_190_195_groupi_n_4885);
  not csa_tree_add_190_195_groupi_g44085(csa_tree_add_190_195_groupi_n_4880 ,csa_tree_add_190_195_groupi_n_4879);
  and csa_tree_add_190_195_groupi_g44086(csa_tree_add_190_195_groupi_n_4878 ,csa_tree_add_190_195_groupi_n_720 ,csa_tree_add_190_195_groupi_n_4136);
  or csa_tree_add_190_195_groupi_g44087(csa_tree_add_190_195_groupi_n_4877 ,csa_tree_add_190_195_groupi_n_1537 ,csa_tree_add_190_195_groupi_n_4136);
  or csa_tree_add_190_195_groupi_g44088(csa_tree_add_190_195_groupi_n_4876 ,csa_tree_add_190_195_groupi_n_3471 ,csa_tree_add_190_195_groupi_n_4141);
  and csa_tree_add_190_195_groupi_g44089(csa_tree_add_190_195_groupi_n_4875 ,csa_tree_add_190_195_groupi_n_3338 ,csa_tree_add_190_195_groupi_n_4138);
  or csa_tree_add_190_195_groupi_g44090(csa_tree_add_190_195_groupi_n_4874 ,csa_tree_add_190_195_groupi_n_3687 ,csa_tree_add_190_195_groupi_n_4140);
  and csa_tree_add_190_195_groupi_g44091(csa_tree_add_190_195_groupi_n_4873 ,csa_tree_add_190_195_groupi_n_1846 ,csa_tree_add_190_195_groupi_n_4567);
  and csa_tree_add_190_195_groupi_g44092(csa_tree_add_190_195_groupi_n_5174 ,csa_tree_add_190_195_groupi_n_2982 ,csa_tree_add_190_195_groupi_n_4323);
  and csa_tree_add_190_195_groupi_g44093(csa_tree_add_190_195_groupi_n_5173 ,csa_tree_add_190_195_groupi_n_3001 ,csa_tree_add_190_195_groupi_n_4203);
  and csa_tree_add_190_195_groupi_g44094(csa_tree_add_190_195_groupi_n_5172 ,csa_tree_add_190_195_groupi_n_3506 ,csa_tree_add_190_195_groupi_n_4238);
  or csa_tree_add_190_195_groupi_g44095(csa_tree_add_190_195_groupi_n_5170 ,csa_tree_add_190_195_groupi_n_3548 ,csa_tree_add_190_195_groupi_n_4241);
  and csa_tree_add_190_195_groupi_g44096(csa_tree_add_190_195_groupi_n_5169 ,csa_tree_add_190_195_groupi_n_3082 ,csa_tree_add_190_195_groupi_n_4515);
  or csa_tree_add_190_195_groupi_g44097(csa_tree_add_190_195_groupi_n_5168 ,csa_tree_add_190_195_groupi_n_3099 ,csa_tree_add_190_195_groupi_n_4499);
  or csa_tree_add_190_195_groupi_g44098(csa_tree_add_190_195_groupi_n_5167 ,csa_tree_add_190_195_groupi_n_2795 ,csa_tree_add_190_195_groupi_n_4557);
  and csa_tree_add_190_195_groupi_g44099(csa_tree_add_190_195_groupi_n_5166 ,csa_tree_add_190_195_groupi_n_3485 ,csa_tree_add_190_195_groupi_n_4467);
  or csa_tree_add_190_195_groupi_g44100(csa_tree_add_190_195_groupi_n_5164 ,csa_tree_add_190_195_groupi_n_2960 ,csa_tree_add_190_195_groupi_n_4245);
  and csa_tree_add_190_195_groupi_g44101(csa_tree_add_190_195_groupi_n_5163 ,csa_tree_add_190_195_groupi_n_3599 ,csa_tree_add_190_195_groupi_n_4309);
  and csa_tree_add_190_195_groupi_g44102(csa_tree_add_190_195_groupi_n_5162 ,csa_tree_add_190_195_groupi_n_3685 ,csa_tree_add_190_195_groupi_n_4164);
  and csa_tree_add_190_195_groupi_g44103(csa_tree_add_190_195_groupi_n_5161 ,csa_tree_add_190_195_groupi_n_2748 ,csa_tree_add_190_195_groupi_n_4433);
  or csa_tree_add_190_195_groupi_g44104(csa_tree_add_190_195_groupi_n_5160 ,csa_tree_add_190_195_groupi_n_3141 ,csa_tree_add_190_195_groupi_n_4502);
  and csa_tree_add_190_195_groupi_g44105(csa_tree_add_190_195_groupi_n_5159 ,csa_tree_add_190_195_groupi_n_3670 ,csa_tree_add_190_195_groupi_n_4267);
  or csa_tree_add_190_195_groupi_g44106(csa_tree_add_190_195_groupi_n_5157 ,csa_tree_add_190_195_groupi_n_3092 ,csa_tree_add_190_195_groupi_n_4505);
  and csa_tree_add_190_195_groupi_g44107(csa_tree_add_190_195_groupi_n_5156 ,csa_tree_add_190_195_groupi_n_2768 ,csa_tree_add_190_195_groupi_n_4306);
  and csa_tree_add_190_195_groupi_g44108(csa_tree_add_190_195_groupi_n_5155 ,csa_tree_add_190_195_groupi_n_3540 ,csa_tree_add_190_195_groupi_n_4160);
  and csa_tree_add_190_195_groupi_g44109(csa_tree_add_190_195_groupi_n_5154 ,csa_tree_add_190_195_groupi_n_3019 ,csa_tree_add_190_195_groupi_n_4320);
  and csa_tree_add_190_195_groupi_g44110(csa_tree_add_190_195_groupi_n_5153 ,csa_tree_add_190_195_groupi_n_3672 ,csa_tree_add_190_195_groupi_n_4282);
  or csa_tree_add_190_195_groupi_g44111(csa_tree_add_190_195_groupi_n_5152 ,csa_tree_add_190_195_groupi_n_3065 ,csa_tree_add_190_195_groupi_n_4277);
  and csa_tree_add_190_195_groupi_g44112(csa_tree_add_190_195_groupi_n_5151 ,csa_tree_add_190_195_groupi_n_3047 ,csa_tree_add_190_195_groupi_n_4247);
  and csa_tree_add_190_195_groupi_g44113(csa_tree_add_190_195_groupi_n_5150 ,csa_tree_add_190_195_groupi_n_3139 ,csa_tree_add_190_195_groupi_n_4234);
  and csa_tree_add_190_195_groupi_g44114(csa_tree_add_190_195_groupi_n_5149 ,csa_tree_add_190_195_groupi_n_3443 ,csa_tree_add_190_195_groupi_n_4343);
  and csa_tree_add_190_195_groupi_g44115(csa_tree_add_190_195_groupi_n_5148 ,csa_tree_add_190_195_groupi_n_3237 ,csa_tree_add_190_195_groupi_n_4202);
  and csa_tree_add_190_195_groupi_g44116(csa_tree_add_190_195_groupi_n_5147 ,csa_tree_add_190_195_groupi_n_2888 ,csa_tree_add_190_195_groupi_n_4363);
  or csa_tree_add_190_195_groupi_g44117(csa_tree_add_190_195_groupi_n_5146 ,csa_tree_add_190_195_groupi_n_2908 ,csa_tree_add_190_195_groupi_n_4496);
  or csa_tree_add_190_195_groupi_g44118(csa_tree_add_190_195_groupi_n_5145 ,csa_tree_add_190_195_groupi_n_3278 ,csa_tree_add_190_195_groupi_n_4272);
  and csa_tree_add_190_195_groupi_g44119(csa_tree_add_190_195_groupi_n_5144 ,csa_tree_add_190_195_groupi_n_3612 ,csa_tree_add_190_195_groupi_n_4326);
  and csa_tree_add_190_195_groupi_g44120(csa_tree_add_190_195_groupi_n_5143 ,csa_tree_add_190_195_groupi_n_3285 ,csa_tree_add_190_195_groupi_n_4337);
  and csa_tree_add_190_195_groupi_g44121(csa_tree_add_190_195_groupi_n_5142 ,csa_tree_add_190_195_groupi_n_2882 ,csa_tree_add_190_195_groupi_n_4316);
  and csa_tree_add_190_195_groupi_g44122(csa_tree_add_190_195_groupi_n_5141 ,csa_tree_add_190_195_groupi_n_2969 ,csa_tree_add_190_195_groupi_n_4477);
  and csa_tree_add_190_195_groupi_g44123(csa_tree_add_190_195_groupi_n_5140 ,csa_tree_add_190_195_groupi_n_3722 ,csa_tree_add_190_195_groupi_n_4352);
  and csa_tree_add_190_195_groupi_g44124(csa_tree_add_190_195_groupi_n_5139 ,csa_tree_add_190_195_groupi_n_3113 ,csa_tree_add_190_195_groupi_n_4218);
  and csa_tree_add_190_195_groupi_g44125(csa_tree_add_190_195_groupi_n_5138 ,csa_tree_add_190_195_groupi_n_3229 ,csa_tree_add_190_195_groupi_n_4541);
  or csa_tree_add_190_195_groupi_g44126(csa_tree_add_190_195_groupi_n_5137 ,csa_tree_add_190_195_groupi_n_2863 ,csa_tree_add_190_195_groupi_n_4447);
  and csa_tree_add_190_195_groupi_g44127(csa_tree_add_190_195_groupi_n_5136 ,csa_tree_add_190_195_groupi_n_3677 ,csa_tree_add_190_195_groupi_n_4553);
  and csa_tree_add_190_195_groupi_g44128(csa_tree_add_190_195_groupi_n_5135 ,csa_tree_add_190_195_groupi_n_2905 ,csa_tree_add_190_195_groupi_n_4332);
  or csa_tree_add_190_195_groupi_g44129(csa_tree_add_190_195_groupi_n_5134 ,csa_tree_add_190_195_groupi_n_3155 ,csa_tree_add_190_195_groupi_n_4298);
  or csa_tree_add_190_195_groupi_g44130(csa_tree_add_190_195_groupi_n_5133 ,csa_tree_add_190_195_groupi_n_3233 ,csa_tree_add_190_195_groupi_n_4531);
  and csa_tree_add_190_195_groupi_g44131(csa_tree_add_190_195_groupi_n_5132 ,csa_tree_add_190_195_groupi_n_3169 ,csa_tree_add_190_195_groupi_n_4315);
  and csa_tree_add_190_195_groupi_g44132(csa_tree_add_190_195_groupi_n_5131 ,csa_tree_add_190_195_groupi_n_2993 ,csa_tree_add_190_195_groupi_n_4176);
  and csa_tree_add_190_195_groupi_g44133(csa_tree_add_190_195_groupi_n_5130 ,csa_tree_add_190_195_groupi_n_3585 ,csa_tree_add_190_195_groupi_n_4372);
  and csa_tree_add_190_195_groupi_g44134(csa_tree_add_190_195_groupi_n_5129 ,csa_tree_add_190_195_groupi_n_2782 ,csa_tree_add_190_195_groupi_n_4222);
  and csa_tree_add_190_195_groupi_g44135(csa_tree_add_190_195_groupi_n_5128 ,csa_tree_add_190_195_groupi_n_2994 ,csa_tree_add_190_195_groupi_n_4550);
  or csa_tree_add_190_195_groupi_g44136(csa_tree_add_190_195_groupi_n_5127 ,csa_tree_add_190_195_groupi_n_2988 ,csa_tree_add_190_195_groupi_n_4305);
  or csa_tree_add_190_195_groupi_g44137(csa_tree_add_190_195_groupi_n_5126 ,csa_tree_add_190_195_groupi_n_2784 ,csa_tree_add_190_195_groupi_n_4500);
  and csa_tree_add_190_195_groupi_g44138(csa_tree_add_190_195_groupi_n_5125 ,csa_tree_add_190_195_groupi_n_3231 ,csa_tree_add_190_195_groupi_n_4464);
  or csa_tree_add_190_195_groupi_g44139(csa_tree_add_190_195_groupi_n_5123 ,csa_tree_add_190_195_groupi_n_2816 ,csa_tree_add_190_195_groupi_n_4430);
  and csa_tree_add_190_195_groupi_g44140(csa_tree_add_190_195_groupi_n_5122 ,csa_tree_add_190_195_groupi_n_3194 ,csa_tree_add_190_195_groupi_n_4253);
  or csa_tree_add_190_195_groupi_g44141(csa_tree_add_190_195_groupi_n_5121 ,csa_tree_add_190_195_groupi_n_2950 ,csa_tree_add_190_195_groupi_n_4549);
  and csa_tree_add_190_195_groupi_g44142(csa_tree_add_190_195_groupi_n_5120 ,csa_tree_add_190_195_groupi_n_2989 ,csa_tree_add_190_195_groupi_n_4458);
  and csa_tree_add_190_195_groupi_g44143(csa_tree_add_190_195_groupi_n_5119 ,csa_tree_add_190_195_groupi_n_3727 ,csa_tree_add_190_195_groupi_n_4504);
  or csa_tree_add_190_195_groupi_g44144(csa_tree_add_190_195_groupi_n_5118 ,csa_tree_add_190_195_groupi_n_2978 ,csa_tree_add_190_195_groupi_n_4520);
  or csa_tree_add_190_195_groupi_g44145(csa_tree_add_190_195_groupi_n_5117 ,csa_tree_add_190_195_groupi_n_2750 ,csa_tree_add_190_195_groupi_n_4527);
  and csa_tree_add_190_195_groupi_g44146(csa_tree_add_190_195_groupi_n_5116 ,csa_tree_add_190_195_groupi_n_2973 ,csa_tree_add_190_195_groupi_n_4193);
  and csa_tree_add_190_195_groupi_g44147(csa_tree_add_190_195_groupi_n_5115 ,csa_tree_add_190_195_groupi_n_3455 ,csa_tree_add_190_195_groupi_n_4280);
  and csa_tree_add_190_195_groupi_g44148(csa_tree_add_190_195_groupi_n_5114 ,csa_tree_add_190_195_groupi_n_3546 ,csa_tree_add_190_195_groupi_n_4281);
  and csa_tree_add_190_195_groupi_g44149(csa_tree_add_190_195_groupi_n_5113 ,csa_tree_add_190_195_groupi_n_3450 ,csa_tree_add_190_195_groupi_n_4210);
  and csa_tree_add_190_195_groupi_g44150(csa_tree_add_190_195_groupi_n_5112 ,csa_tree_add_190_195_groupi_n_3429 ,csa_tree_add_190_195_groupi_n_4167);
  or csa_tree_add_190_195_groupi_g44151(csa_tree_add_190_195_groupi_n_5110 ,csa_tree_add_190_195_groupi_n_2926 ,csa_tree_add_190_195_groupi_n_4461);
  or csa_tree_add_190_195_groupi_g44152(csa_tree_add_190_195_groupi_n_5108 ,csa_tree_add_190_195_groupi_n_3176 ,csa_tree_add_190_195_groupi_n_4285);
  and csa_tree_add_190_195_groupi_g44153(csa_tree_add_190_195_groupi_n_5107 ,csa_tree_add_190_195_groupi_n_3588 ,csa_tree_add_190_195_groupi_n_4219);
  and csa_tree_add_190_195_groupi_g44154(csa_tree_add_190_195_groupi_n_5106 ,csa_tree_add_190_195_groupi_n_3404 ,csa_tree_add_190_195_groupi_n_4448);
  and csa_tree_add_190_195_groupi_g44155(csa_tree_add_190_195_groupi_n_5105 ,csa_tree_add_190_195_groupi_n_3125 ,csa_tree_add_190_195_groupi_n_4333);
  or csa_tree_add_190_195_groupi_g44156(csa_tree_add_190_195_groupi_n_5104 ,csa_tree_add_190_195_groupi_n_3190 ,csa_tree_add_190_195_groupi_n_4422);
  or csa_tree_add_190_195_groupi_g44157(csa_tree_add_190_195_groupi_n_5103 ,csa_tree_add_190_195_groupi_n_3478 ,csa_tree_add_190_195_groupi_n_4264);
  or csa_tree_add_190_195_groupi_g44158(csa_tree_add_190_195_groupi_n_5102 ,csa_tree_add_190_195_groupi_n_3503 ,csa_tree_add_190_195_groupi_n_4493);
  and csa_tree_add_190_195_groupi_g44159(csa_tree_add_190_195_groupi_n_5101 ,csa_tree_add_190_195_groupi_n_2790 ,csa_tree_add_190_195_groupi_n_4379);
  or csa_tree_add_190_195_groupi_g44160(csa_tree_add_190_195_groupi_n_5100 ,csa_tree_add_190_195_groupi_n_3532 ,csa_tree_add_190_195_groupi_n_4412);
  and csa_tree_add_190_195_groupi_g44161(csa_tree_add_190_195_groupi_n_5099 ,csa_tree_add_190_195_groupi_n_3167 ,csa_tree_add_190_195_groupi_n_4457);
  and csa_tree_add_190_195_groupi_g44162(csa_tree_add_190_195_groupi_n_5098 ,csa_tree_add_190_195_groupi_n_2913 ,csa_tree_add_190_195_groupi_n_4423);
  or csa_tree_add_190_195_groupi_g44163(csa_tree_add_190_195_groupi_n_5097 ,csa_tree_add_190_195_groupi_n_3230 ,csa_tree_add_190_195_groupi_n_4440);
  and csa_tree_add_190_195_groupi_g44164(csa_tree_add_190_195_groupi_n_5096 ,csa_tree_add_190_195_groupi_n_2907 ,csa_tree_add_190_195_groupi_n_4237);
  or csa_tree_add_190_195_groupi_g44165(csa_tree_add_190_195_groupi_n_5093 ,csa_tree_add_190_195_groupi_n_3498 ,csa_tree_add_190_195_groupi_n_4252);
  and csa_tree_add_190_195_groupi_g44166(csa_tree_add_190_195_groupi_n_5092 ,csa_tree_add_190_195_groupi_n_2900 ,csa_tree_add_190_195_groupi_n_4556);
  and csa_tree_add_190_195_groupi_g44167(csa_tree_add_190_195_groupi_n_5090 ,csa_tree_add_190_195_groupi_n_2738 ,csa_tree_add_190_195_groupi_n_4174);
  or csa_tree_add_190_195_groupi_g44168(csa_tree_add_190_195_groupi_n_5088 ,csa_tree_add_190_195_groupi_n_2771 ,csa_tree_add_190_195_groupi_n_4246);
  or csa_tree_add_190_195_groupi_g44169(csa_tree_add_190_195_groupi_n_5087 ,csa_tree_add_190_195_groupi_n_3581 ,csa_tree_add_190_195_groupi_n_4294);
  and csa_tree_add_190_195_groupi_g44170(csa_tree_add_190_195_groupi_n_5085 ,csa_tree_add_190_195_groupi_n_3256 ,csa_tree_add_190_195_groupi_n_4150);
  or csa_tree_add_190_195_groupi_g44171(csa_tree_add_190_195_groupi_n_5084 ,csa_tree_add_190_195_groupi_n_3067 ,csa_tree_add_190_195_groupi_n_4552);
  or csa_tree_add_190_195_groupi_g44172(csa_tree_add_190_195_groupi_n_5082 ,csa_tree_add_190_195_groupi_n_3709 ,csa_tree_add_190_195_groupi_n_4300);
  or csa_tree_add_190_195_groupi_g44173(csa_tree_add_190_195_groupi_n_5080 ,csa_tree_add_190_195_groupi_n_2824 ,csa_tree_add_190_195_groupi_n_4335);
  and csa_tree_add_190_195_groupi_g44174(csa_tree_add_190_195_groupi_n_5079 ,csa_tree_add_190_195_groupi_n_3363 ,csa_tree_add_190_195_groupi_n_4184);
  and csa_tree_add_190_195_groupi_g44175(csa_tree_add_190_195_groupi_n_5076 ,csa_tree_add_190_195_groupi_n_2927 ,csa_tree_add_190_195_groupi_n_4293);
  and csa_tree_add_190_195_groupi_g44176(csa_tree_add_190_195_groupi_n_5075 ,csa_tree_add_190_195_groupi_n_3323 ,csa_tree_add_190_195_groupi_n_4400);
  or csa_tree_add_190_195_groupi_g44177(csa_tree_add_190_195_groupi_n_5072 ,csa_tree_add_190_195_groupi_n_2813 ,csa_tree_add_190_195_groupi_n_4491);
  and csa_tree_add_190_195_groupi_g44178(csa_tree_add_190_195_groupi_n_5071 ,csa_tree_add_190_195_groupi_n_3308 ,csa_tree_add_190_195_groupi_n_4397);
  or csa_tree_add_190_195_groupi_g44179(csa_tree_add_190_195_groupi_n_5069 ,csa_tree_add_190_195_groupi_n_3528 ,csa_tree_add_190_195_groupi_n_4414);
  or csa_tree_add_190_195_groupi_g44180(csa_tree_add_190_195_groupi_n_5067 ,csa_tree_add_190_195_groupi_n_2968 ,csa_tree_add_190_195_groupi_n_4366);
  or csa_tree_add_190_195_groupi_g44181(csa_tree_add_190_195_groupi_n_5065 ,csa_tree_add_190_195_groupi_n_3122 ,csa_tree_add_190_195_groupi_n_4425);
  or csa_tree_add_190_195_groupi_g44182(csa_tree_add_190_195_groupi_n_5064 ,csa_tree_add_190_195_groupi_n_3287 ,csa_tree_add_190_195_groupi_n_4248);
  or csa_tree_add_190_195_groupi_g44183(csa_tree_add_190_195_groupi_n_5062 ,csa_tree_add_190_195_groupi_n_3559 ,csa_tree_add_190_195_groupi_n_4374);
  and csa_tree_add_190_195_groupi_g44184(csa_tree_add_190_195_groupi_n_5060 ,csa_tree_add_190_195_groupi_n_3587 ,csa_tree_add_190_195_groupi_n_4373);
  and csa_tree_add_190_195_groupi_g44185(csa_tree_add_190_195_groupi_n_5058 ,csa_tree_add_190_195_groupi_n_2914 ,csa_tree_add_190_195_groupi_n_4276);
  or csa_tree_add_190_195_groupi_g44186(csa_tree_add_190_195_groupi_n_5056 ,csa_tree_add_190_195_groupi_n_3276 ,csa_tree_add_190_195_groupi_n_4274);
  and csa_tree_add_190_195_groupi_g44187(csa_tree_add_190_195_groupi_n_5055 ,csa_tree_add_190_195_groupi_n_3479 ,csa_tree_add_190_195_groupi_n_4360);
  or csa_tree_add_190_195_groupi_g44188(csa_tree_add_190_195_groupi_n_5053 ,csa_tree_add_190_195_groupi_n_3000 ,csa_tree_add_190_195_groupi_n_4523);
  and csa_tree_add_190_195_groupi_g44189(csa_tree_add_190_195_groupi_n_5051 ,csa_tree_add_190_195_groupi_n_2948 ,csa_tree_add_190_195_groupi_n_4304);
  or csa_tree_add_190_195_groupi_g44190(csa_tree_add_190_195_groupi_n_5049 ,csa_tree_add_190_195_groupi_n_3290 ,csa_tree_add_190_195_groupi_n_4286);
  and csa_tree_add_190_195_groupi_g44191(csa_tree_add_190_195_groupi_n_5047 ,csa_tree_add_190_195_groupi_n_3610 ,csa_tree_add_190_195_groupi_n_4152);
  or csa_tree_add_190_195_groupi_g44192(csa_tree_add_190_195_groupi_n_5045 ,csa_tree_add_190_195_groupi_n_3302 ,csa_tree_add_190_195_groupi_n_4348);
  and csa_tree_add_190_195_groupi_g44193(csa_tree_add_190_195_groupi_n_5043 ,csa_tree_add_190_195_groupi_n_3441 ,csa_tree_add_190_195_groupi_n_4344);
  or csa_tree_add_190_195_groupi_g44194(csa_tree_add_190_195_groupi_n_5041 ,csa_tree_add_190_195_groupi_n_3192 ,csa_tree_add_190_195_groupi_n_4497);
  or csa_tree_add_190_195_groupi_g44195(csa_tree_add_190_195_groupi_n_5039 ,csa_tree_add_190_195_groupi_n_2792 ,csa_tree_add_190_195_groupi_n_4460);
  or csa_tree_add_190_195_groupi_g44196(csa_tree_add_190_195_groupi_n_5037 ,csa_tree_add_190_195_groupi_n_3569 ,csa_tree_add_190_195_groupi_n_4215);
  or csa_tree_add_190_195_groupi_g44197(csa_tree_add_190_195_groupi_n_5036 ,csa_tree_add_190_195_groupi_n_2835 ,csa_tree_add_190_195_groupi_n_4528);
  and csa_tree_add_190_195_groupi_g44198(csa_tree_add_190_195_groupi_n_5034 ,csa_tree_add_190_195_groupi_n_2929 ,csa_tree_add_190_195_groupi_n_4327);
  and csa_tree_add_190_195_groupi_g44199(csa_tree_add_190_195_groupi_n_5032 ,csa_tree_add_190_195_groupi_n_3440 ,csa_tree_add_190_195_groupi_n_4205);
  or csa_tree_add_190_195_groupi_g44200(csa_tree_add_190_195_groupi_n_5031 ,csa_tree_add_190_195_groupi_n_3578 ,csa_tree_add_190_195_groupi_n_4473);
  and csa_tree_add_190_195_groupi_g44201(csa_tree_add_190_195_groupi_n_5029 ,csa_tree_add_190_195_groupi_n_3409 ,csa_tree_add_190_195_groupi_n_4445);
  and csa_tree_add_190_195_groupi_g44202(csa_tree_add_190_195_groupi_n_5027 ,csa_tree_add_190_195_groupi_n_3463 ,csa_tree_add_190_195_groupi_n_4472);
  or csa_tree_add_190_195_groupi_g44203(csa_tree_add_190_195_groupi_n_5025 ,csa_tree_add_190_195_groupi_n_3166 ,csa_tree_add_190_195_groupi_n_4480);
  or csa_tree_add_190_195_groupi_g44204(csa_tree_add_190_195_groupi_n_5024 ,csa_tree_add_190_195_groupi_n_3448 ,csa_tree_add_190_195_groupi_n_4279);
  or csa_tree_add_190_195_groupi_g44205(csa_tree_add_190_195_groupi_n_5022 ,csa_tree_add_190_195_groupi_n_3277 ,csa_tree_add_190_195_groupi_n_4231);
  and csa_tree_add_190_195_groupi_g44206(csa_tree_add_190_195_groupi_n_5020 ,csa_tree_add_190_195_groupi_n_3519 ,csa_tree_add_190_195_groupi_n_4406);
  or csa_tree_add_190_195_groupi_g44207(csa_tree_add_190_195_groupi_n_5018 ,csa_tree_add_190_195_groupi_n_3590 ,csa_tree_add_190_195_groupi_n_4410);
  or csa_tree_add_190_195_groupi_g44208(csa_tree_add_190_195_groupi_n_5017 ,csa_tree_add_190_195_groupi_n_3013 ,csa_tree_add_190_195_groupi_n_4367);
  or csa_tree_add_190_195_groupi_g44209(csa_tree_add_190_195_groupi_n_5016 ,csa_tree_add_190_195_groupi_n_3095 ,csa_tree_add_190_195_groupi_n_4485);
  or csa_tree_add_190_195_groupi_g44210(csa_tree_add_190_195_groupi_n_5014 ,csa_tree_add_190_195_groupi_n_3138 ,csa_tree_add_190_195_groupi_n_4488);
  and csa_tree_add_190_195_groupi_g44211(csa_tree_add_190_195_groupi_n_5012 ,csa_tree_add_190_195_groupi_n_3012 ,csa_tree_add_190_195_groupi_n_4289);
  and csa_tree_add_190_195_groupi_g44212(csa_tree_add_190_195_groupi_n_5010 ,csa_tree_add_190_195_groupi_n_3241 ,csa_tree_add_190_195_groupi_n_4308);
  or csa_tree_add_190_195_groupi_g44213(csa_tree_add_190_195_groupi_n_5009 ,csa_tree_add_190_195_groupi_n_3052 ,csa_tree_add_190_195_groupi_n_4474);
  or csa_tree_add_190_195_groupi_g44214(csa_tree_add_190_195_groupi_n_5007 ,csa_tree_add_190_195_groupi_n_2815 ,csa_tree_add_190_195_groupi_n_4519);
  or csa_tree_add_190_195_groupi_g44215(csa_tree_add_190_195_groupi_n_5005 ,csa_tree_add_190_195_groupi_n_3116 ,csa_tree_add_190_195_groupi_n_4435);
  or csa_tree_add_190_195_groupi_g44216(csa_tree_add_190_195_groupi_n_5004 ,csa_tree_add_190_195_groupi_n_3543 ,csa_tree_add_190_195_groupi_n_4384);
  or csa_tree_add_190_195_groupi_g44217(csa_tree_add_190_195_groupi_n_5003 ,csa_tree_add_190_195_groupi_n_2776 ,csa_tree_add_190_195_groupi_n_4243);
  and csa_tree_add_190_195_groupi_g44218(csa_tree_add_190_195_groupi_n_5002 ,csa_tree_add_190_195_groupi_n_3195 ,csa_tree_add_190_195_groupi_n_4510);
  or csa_tree_add_190_195_groupi_g44219(csa_tree_add_190_195_groupi_n_4999 ,csa_tree_add_190_195_groupi_n_3031 ,csa_tree_add_190_195_groupi_n_4487);
  or csa_tree_add_190_195_groupi_g44220(csa_tree_add_190_195_groupi_n_4998 ,csa_tree_add_190_195_groupi_n_3331 ,csa_tree_add_190_195_groupi_n_4266);
  or csa_tree_add_190_195_groupi_g44221(csa_tree_add_190_195_groupi_n_4996 ,csa_tree_add_190_195_groupi_n_3613 ,csa_tree_add_190_195_groupi_n_4538);
  or csa_tree_add_190_195_groupi_g44222(csa_tree_add_190_195_groupi_n_4994 ,csa_tree_add_190_195_groupi_n_3185 ,csa_tree_add_190_195_groupi_n_4513);
  and csa_tree_add_190_195_groupi_g44223(csa_tree_add_190_195_groupi_n_4992 ,csa_tree_add_190_195_groupi_n_3247 ,csa_tree_add_190_195_groupi_n_4221);
  or csa_tree_add_190_195_groupi_g44224(csa_tree_add_190_195_groupi_n_4991 ,csa_tree_add_190_195_groupi_n_3483 ,csa_tree_add_190_195_groupi_n_4559);
  or csa_tree_add_190_195_groupi_g44225(csa_tree_add_190_195_groupi_n_4988 ,csa_tree_add_190_195_groupi_n_3456 ,csa_tree_add_190_195_groupi_n_4361);
  and csa_tree_add_190_195_groupi_g44226(csa_tree_add_190_195_groupi_n_4987 ,csa_tree_add_190_195_groupi_n_2895 ,csa_tree_add_190_195_groupi_n_4498);
  or csa_tree_add_190_195_groupi_g44227(csa_tree_add_190_195_groupi_n_4986 ,csa_tree_add_190_195_groupi_n_3412 ,csa_tree_add_190_195_groupi_n_4295);
  and csa_tree_add_190_195_groupi_g44228(csa_tree_add_190_195_groupi_n_4985 ,csa_tree_add_190_195_groupi_n_3079 ,csa_tree_add_190_195_groupi_n_4534);
  or csa_tree_add_190_195_groupi_g44229(csa_tree_add_190_195_groupi_n_4983 ,csa_tree_add_190_195_groupi_n_3390 ,csa_tree_add_190_195_groupi_n_4273);
  or csa_tree_add_190_195_groupi_g44230(csa_tree_add_190_195_groupi_n_4981 ,csa_tree_add_190_195_groupi_n_2919 ,csa_tree_add_190_195_groupi_n_4530);
  or csa_tree_add_190_195_groupi_g44231(csa_tree_add_190_195_groupi_n_4979 ,csa_tree_add_190_195_groupi_n_3539 ,csa_tree_add_190_195_groupi_n_4232);
  and csa_tree_add_190_195_groupi_g44232(csa_tree_add_190_195_groupi_n_4978 ,csa_tree_add_190_195_groupi_n_3351 ,csa_tree_add_190_195_groupi_n_4399);
  or csa_tree_add_190_195_groupi_g44233(csa_tree_add_190_195_groupi_n_4977 ,csa_tree_add_190_195_groupi_n_3630 ,csa_tree_add_190_195_groupi_n_4470);
  or csa_tree_add_190_195_groupi_g44234(csa_tree_add_190_195_groupi_n_4975 ,csa_tree_add_190_195_groupi_n_2858 ,csa_tree_add_190_195_groupi_n_4334);
  or csa_tree_add_190_195_groupi_g44235(csa_tree_add_190_195_groupi_n_4973 ,csa_tree_add_190_195_groupi_n_3481 ,csa_tree_add_190_195_groupi_n_4346);
  and csa_tree_add_190_195_groupi_g44236(csa_tree_add_190_195_groupi_n_4971 ,csa_tree_add_190_195_groupi_n_3586 ,csa_tree_add_190_195_groupi_n_4371);
  or csa_tree_add_190_195_groupi_g44237(csa_tree_add_190_195_groupi_n_4969 ,csa_tree_add_190_195_groupi_n_3090 ,csa_tree_add_190_195_groupi_n_4429);
  and csa_tree_add_190_195_groupi_g44238(csa_tree_add_190_195_groupi_n_4967 ,csa_tree_add_190_195_groupi_n_3558 ,csa_tree_add_190_195_groupi_n_4413);
  or csa_tree_add_190_195_groupi_g44239(csa_tree_add_190_195_groupi_n_4966 ,csa_tree_add_190_195_groupi_n_3571 ,csa_tree_add_190_195_groupi_n_4269);
  and csa_tree_add_190_195_groupi_g44240(csa_tree_add_190_195_groupi_n_4963 ,csa_tree_add_190_195_groupi_n_2794 ,csa_tree_add_190_195_groupi_n_4196);
  and csa_tree_add_190_195_groupi_g44241(csa_tree_add_190_195_groupi_n_4962 ,csa_tree_add_190_195_groupi_n_3327 ,csa_tree_add_190_195_groupi_n_4405);
  or csa_tree_add_190_195_groupi_g44242(csa_tree_add_190_195_groupi_n_4960 ,csa_tree_add_190_195_groupi_n_3652 ,csa_tree_add_190_195_groupi_n_4451);
  and csa_tree_add_190_195_groupi_g44243(csa_tree_add_190_195_groupi_n_4958 ,csa_tree_add_190_195_groupi_n_3621 ,csa_tree_add_190_195_groupi_n_4476);
  or csa_tree_add_190_195_groupi_g44244(csa_tree_add_190_195_groupi_n_4957 ,csa_tree_add_190_195_groupi_n_3361 ,csa_tree_add_190_195_groupi_n_4303);
  or csa_tree_add_190_195_groupi_g44245(csa_tree_add_190_195_groupi_n_4955 ,csa_tree_add_190_195_groupi_n_3303 ,csa_tree_add_190_195_groupi_n_4339);
  or csa_tree_add_190_195_groupi_g44246(csa_tree_add_190_195_groupi_n_4954 ,csa_tree_add_190_195_groupi_n_2755 ,csa_tree_add_190_195_groupi_n_4546);
  or csa_tree_add_190_195_groupi_g44247(csa_tree_add_190_195_groupi_n_4951 ,csa_tree_add_190_195_groupi_n_3006 ,csa_tree_add_190_195_groupi_n_4301);
  or csa_tree_add_190_195_groupi_g44248(csa_tree_add_190_195_groupi_n_4950 ,csa_tree_add_190_195_groupi_n_2979 ,csa_tree_add_190_195_groupi_n_4486);
  or csa_tree_add_190_195_groupi_g44249(csa_tree_add_190_195_groupi_n_4948 ,csa_tree_add_190_195_groupi_n_3305 ,csa_tree_add_190_195_groupi_n_4325);
  or csa_tree_add_190_195_groupi_g44250(csa_tree_add_190_195_groupi_n_4946 ,csa_tree_add_190_195_groupi_n_2812 ,csa_tree_add_190_195_groupi_n_4554);
  or csa_tree_add_190_195_groupi_g44251(csa_tree_add_190_195_groupi_n_4944 ,csa_tree_add_190_195_groupi_n_2845 ,csa_tree_add_190_195_groupi_n_4437);
  and csa_tree_add_190_195_groupi_g44252(csa_tree_add_190_195_groupi_n_4943 ,csa_tree_add_190_195_groupi_n_3322 ,csa_tree_add_190_195_groupi_n_4389);
  or csa_tree_add_190_195_groupi_g44253(csa_tree_add_190_195_groupi_n_4941 ,csa_tree_add_190_195_groupi_n_2820 ,csa_tree_add_190_195_groupi_n_4438);
  and csa_tree_add_190_195_groupi_g44254(csa_tree_add_190_195_groupi_n_4938 ,csa_tree_add_190_195_groupi_n_2999 ,csa_tree_add_190_195_groupi_n_4242);
  or csa_tree_add_190_195_groupi_g44255(csa_tree_add_190_195_groupi_n_4937 ,csa_tree_add_190_195_groupi_n_2998 ,csa_tree_add_190_195_groupi_n_4482);
  or csa_tree_add_190_195_groupi_g44256(csa_tree_add_190_195_groupi_n_4934 ,csa_tree_add_190_195_groupi_n_2866 ,csa_tree_add_190_195_groupi_n_4200);
  and csa_tree_add_190_195_groupi_g44257(csa_tree_add_190_195_groupi_n_4933 ,csa_tree_add_190_195_groupi_n_3666 ,csa_tree_add_190_195_groupi_n_4317);
  and csa_tree_add_190_195_groupi_g44258(csa_tree_add_190_195_groupi_n_4931 ,csa_tree_add_190_195_groupi_n_3023 ,csa_tree_add_190_195_groupi_n_4494);
  or csa_tree_add_190_195_groupi_g44259(csa_tree_add_190_195_groupi_n_4930 ,csa_tree_add_190_195_groupi_n_3366 ,csa_tree_add_190_195_groupi_n_4209);
  and csa_tree_add_190_195_groupi_g44260(csa_tree_add_190_195_groupi_n_4928 ,csa_tree_add_190_195_groupi_n_3597 ,csa_tree_add_190_195_groupi_n_4415);
  and csa_tree_add_190_195_groupi_g44261(csa_tree_add_190_195_groupi_n_4926 ,csa_tree_add_190_195_groupi_n_3711 ,csa_tree_add_190_195_groupi_n_4385);
  and csa_tree_add_190_195_groupi_g44262(csa_tree_add_190_195_groupi_n_4925 ,csa_tree_add_190_195_groupi_n_3426 ,csa_tree_add_190_195_groupi_n_4341);
  or csa_tree_add_190_195_groupi_g44263(csa_tree_add_190_195_groupi_n_4924 ,csa_tree_add_190_195_groupi_n_3461 ,csa_tree_add_190_195_groupi_n_4358);
  and csa_tree_add_190_195_groupi_g44264(csa_tree_add_190_195_groupi_n_4922 ,csa_tree_add_190_195_groupi_n_3165 ,csa_tree_add_190_195_groupi_n_4249);
  or csa_tree_add_190_195_groupi_g44265(csa_tree_add_190_195_groupi_n_4920 ,csa_tree_add_190_195_groupi_n_3118 ,csa_tree_add_190_195_groupi_n_4524);
  or csa_tree_add_190_195_groupi_g44266(csa_tree_add_190_195_groupi_n_4918 ,csa_tree_add_190_195_groupi_n_2744 ,csa_tree_add_190_195_groupi_n_4465);
  and csa_tree_add_190_195_groupi_g44267(csa_tree_add_190_195_groupi_n_4917 ,csa_tree_add_190_195_groupi_n_3360 ,csa_tree_add_190_195_groupi_n_4403);
  or csa_tree_add_190_195_groupi_g44268(csa_tree_add_190_195_groupi_n_4916 ,csa_tree_add_190_195_groupi_n_3209 ,csa_tree_add_190_195_groupi_n_4466);
  or csa_tree_add_190_195_groupi_g44269(csa_tree_add_190_195_groupi_n_4915 ,csa_tree_add_190_195_groupi_n_3457 ,csa_tree_add_190_195_groupi_n_4391);
  or csa_tree_add_190_195_groupi_g44270(csa_tree_add_190_195_groupi_n_4913 ,csa_tree_add_190_195_groupi_n_3294 ,csa_tree_add_190_195_groupi_n_4227);
  and csa_tree_add_190_195_groupi_g44271(csa_tree_add_190_195_groupi_n_4911 ,csa_tree_add_190_195_groupi_n_3312 ,csa_tree_add_190_195_groupi_n_4387);
  or csa_tree_add_190_195_groupi_g44272(csa_tree_add_190_195_groupi_n_4909 ,csa_tree_add_190_195_groupi_n_3089 ,csa_tree_add_190_195_groupi_n_4181);
  and csa_tree_add_190_195_groupi_g44273(csa_tree_add_190_195_groupi_n_4908 ,csa_tree_add_190_195_groupi_n_3514 ,csa_tree_add_190_195_groupi_n_4478);
  and csa_tree_add_190_195_groupi_g44274(csa_tree_add_190_195_groupi_n_4907 ,csa_tree_add_190_195_groupi_n_3374 ,csa_tree_add_190_195_groupi_n_4362);
  and csa_tree_add_190_195_groupi_g44275(csa_tree_add_190_195_groupi_n_4906 ,csa_tree_add_190_195_groupi_n_3093 ,csa_tree_add_190_195_groupi_n_4168);
  and csa_tree_add_190_195_groupi_g44276(csa_tree_add_190_195_groupi_n_4904 ,csa_tree_add_190_195_groupi_n_3191 ,csa_tree_add_190_195_groupi_n_4220);
  or csa_tree_add_190_195_groupi_g44277(csa_tree_add_190_195_groupi_n_4903 ,csa_tree_add_190_195_groupi_n_2869 ,csa_tree_add_190_195_groupi_n_4368);
  or csa_tree_add_190_195_groupi_g44278(csa_tree_add_190_195_groupi_n_4901 ,csa_tree_add_190_195_groupi_n_3644 ,csa_tree_add_190_195_groupi_n_4452);
  or csa_tree_add_190_195_groupi_g44279(csa_tree_add_190_195_groupi_n_4899 ,csa_tree_add_190_195_groupi_n_2876 ,csa_tree_add_190_195_groupi_n_4544);
  and csa_tree_add_190_195_groupi_g44280(csa_tree_add_190_195_groupi_n_4898 ,csa_tree_add_190_195_groupi_n_3719 ,csa_tree_add_190_195_groupi_n_4431);
  or csa_tree_add_190_195_groupi_g44281(csa_tree_add_190_195_groupi_n_4897 ,csa_tree_add_190_195_groupi_n_3580 ,csa_tree_add_190_195_groupi_n_4383);
  and csa_tree_add_190_195_groupi_g44282(csa_tree_add_190_195_groupi_n_4896 ,csa_tree_add_190_195_groupi_n_3270 ,csa_tree_add_190_195_groupi_n_4302);
  or csa_tree_add_190_195_groupi_g44283(csa_tree_add_190_195_groupi_n_4894 ,csa_tree_add_190_195_groupi_n_3026 ,csa_tree_add_190_195_groupi_n_4310);
  and csa_tree_add_190_195_groupi_g44284(csa_tree_add_190_195_groupi_n_4893 ,csa_tree_add_190_195_groupi_n_3689 ,csa_tree_add_190_195_groupi_n_4537);
  or csa_tree_add_190_195_groupi_g44285(csa_tree_add_190_195_groupi_n_4892 ,csa_tree_add_190_195_groupi_n_3377 ,csa_tree_add_190_195_groupi_n_4312);
  or csa_tree_add_190_195_groupi_g44286(csa_tree_add_190_195_groupi_n_4891 ,csa_tree_add_190_195_groupi_n_3310 ,csa_tree_add_190_195_groupi_n_4250);
  or csa_tree_add_190_195_groupi_g44287(csa_tree_add_190_195_groupi_n_4890 ,csa_tree_add_190_195_groupi_n_3357 ,csa_tree_add_190_195_groupi_n_4380);
  or csa_tree_add_190_195_groupi_g44288(csa_tree_add_190_195_groupi_n_4888 ,csa_tree_add_190_195_groupi_n_3510 ,csa_tree_add_190_195_groupi_n_4178);
  and csa_tree_add_190_195_groupi_g44289(csa_tree_add_190_195_groupi_n_4887 ,csa_tree_add_190_195_groupi_n_3210 ,csa_tree_add_190_195_groupi_n_4330);
  and csa_tree_add_190_195_groupi_g44290(csa_tree_add_190_195_groupi_n_4886 ,csa_tree_add_190_195_groupi_n_2740 ,csa_tree_add_190_195_groupi_n_4177);
  and csa_tree_add_190_195_groupi_g44291(csa_tree_add_190_195_groupi_n_4885 ,csa_tree_add_190_195_groupi_n_3145 ,csa_tree_add_190_195_groupi_n_4259);
  or csa_tree_add_190_195_groupi_g44292(csa_tree_add_190_195_groupi_n_4883 ,csa_tree_add_190_195_groupi_n_3142 ,csa_tree_add_190_195_groupi_n_4314);
  or csa_tree_add_190_195_groupi_g44293(csa_tree_add_190_195_groupi_n_4882 ,csa_tree_add_190_195_groupi_n_3253 ,csa_tree_add_190_195_groupi_n_4347);
  or csa_tree_add_190_195_groupi_g44294(csa_tree_add_190_195_groupi_n_4881 ,csa_tree_add_190_195_groupi_n_3663 ,csa_tree_add_190_195_groupi_n_4357);
  or csa_tree_add_190_195_groupi_g44295(csa_tree_add_190_195_groupi_n_4879 ,csa_tree_add_190_195_groupi_n_3157 ,csa_tree_add_190_195_groupi_n_4481);
  not csa_tree_add_190_195_groupi_g44296(csa_tree_add_190_195_groupi_n_4868 ,csa_tree_add_190_195_groupi_n_4867);
  not csa_tree_add_190_195_groupi_g44297(csa_tree_add_190_195_groupi_n_4864 ,csa_tree_add_190_195_groupi_n_4863);
  not csa_tree_add_190_195_groupi_g44298(csa_tree_add_190_195_groupi_n_4859 ,csa_tree_add_190_195_groupi_n_4858);
  not csa_tree_add_190_195_groupi_g44299(csa_tree_add_190_195_groupi_n_4854 ,csa_tree_add_190_195_groupi_n_4853);
  not csa_tree_add_190_195_groupi_g44300(csa_tree_add_190_195_groupi_n_4835 ,csa_tree_add_190_195_groupi_n_4834);
  not csa_tree_add_190_195_groupi_g44302(csa_tree_add_190_195_groupi_n_4823 ,csa_tree_add_190_195_groupi_n_4822);
  not csa_tree_add_190_195_groupi_g44303(csa_tree_add_190_195_groupi_n_4819 ,csa_tree_add_190_195_groupi_n_4818);
  not csa_tree_add_190_195_groupi_g44305(csa_tree_add_190_195_groupi_n_4810 ,csa_tree_add_190_195_groupi_n_4809);
  not csa_tree_add_190_195_groupi_g44306(csa_tree_add_190_195_groupi_n_4795 ,csa_tree_add_190_195_groupi_n_4796);
  not csa_tree_add_190_195_groupi_g44307(csa_tree_add_190_195_groupi_n_4792 ,csa_tree_add_190_195_groupi_n_4793);
  not csa_tree_add_190_195_groupi_g44308(csa_tree_add_190_195_groupi_n_4790 ,csa_tree_add_190_195_groupi_n_4791);
  not csa_tree_add_190_195_groupi_g44309(csa_tree_add_190_195_groupi_n_4788 ,csa_tree_add_190_195_groupi_n_4789);
  not csa_tree_add_190_195_groupi_g44310(csa_tree_add_190_195_groupi_n_4786 ,csa_tree_add_190_195_groupi_n_4785);
  not csa_tree_add_190_195_groupi_g44311(csa_tree_add_190_195_groupi_n_4784 ,csa_tree_add_190_195_groupi_n_4783);
  not csa_tree_add_190_195_groupi_g44312(csa_tree_add_190_195_groupi_n_4779 ,csa_tree_add_190_195_groupi_n_4780);
  not csa_tree_add_190_195_groupi_g44313(csa_tree_add_190_195_groupi_n_4778 ,csa_tree_add_190_195_groupi_n_4777);
  not csa_tree_add_190_195_groupi_g44314(csa_tree_add_190_195_groupi_n_4774 ,csa_tree_add_190_195_groupi_n_4775);
  not csa_tree_add_190_195_groupi_g44315(csa_tree_add_190_195_groupi_n_4772 ,csa_tree_add_190_195_groupi_n_4773);
  not csa_tree_add_190_195_groupi_g44316(csa_tree_add_190_195_groupi_n_4770 ,csa_tree_add_190_195_groupi_n_4771);
  not csa_tree_add_190_195_groupi_g44317(csa_tree_add_190_195_groupi_n_4768 ,csa_tree_add_190_195_groupi_n_4769);
  not csa_tree_add_190_195_groupi_g44318(csa_tree_add_190_195_groupi_n_4766 ,csa_tree_add_190_195_groupi_n_4767);
  not csa_tree_add_190_195_groupi_g44319(csa_tree_add_190_195_groupi_n_4764 ,csa_tree_add_190_195_groupi_n_4765);
  not csa_tree_add_190_195_groupi_g44320(csa_tree_add_190_195_groupi_n_4762 ,csa_tree_add_190_195_groupi_n_4763);
  not csa_tree_add_190_195_groupi_g44321(csa_tree_add_190_195_groupi_n_4761 ,csa_tree_add_190_195_groupi_n_4760);
  not csa_tree_add_190_195_groupi_g44322(csa_tree_add_190_195_groupi_n_4754 ,csa_tree_add_190_195_groupi_n_4755);
  not csa_tree_add_190_195_groupi_g44323(csa_tree_add_190_195_groupi_n_4750 ,csa_tree_add_190_195_groupi_n_4749);
  not csa_tree_add_190_195_groupi_g44324(csa_tree_add_190_195_groupi_n_4747 ,csa_tree_add_190_195_groupi_n_4748);
  not csa_tree_add_190_195_groupi_g44325(csa_tree_add_190_195_groupi_n_4746 ,csa_tree_add_190_195_groupi_n_4745);
  not csa_tree_add_190_195_groupi_g44326(csa_tree_add_190_195_groupi_n_4742 ,csa_tree_add_190_195_groupi_n_4743);
  not csa_tree_add_190_195_groupi_g44327(csa_tree_add_190_195_groupi_n_4740 ,csa_tree_add_190_195_groupi_n_4741);
  not csa_tree_add_190_195_groupi_g44328(csa_tree_add_190_195_groupi_n_4738 ,csa_tree_add_190_195_groupi_n_4737);
  not csa_tree_add_190_195_groupi_g44329(csa_tree_add_190_195_groupi_n_4735 ,csa_tree_add_190_195_groupi_n_4736);
  not csa_tree_add_190_195_groupi_g44330(csa_tree_add_190_195_groupi_n_4733 ,csa_tree_add_190_195_groupi_n_4734);
  not csa_tree_add_190_195_groupi_g44331(csa_tree_add_190_195_groupi_n_4730 ,csa_tree_add_190_195_groupi_n_4731);
  not csa_tree_add_190_195_groupi_g44332(csa_tree_add_190_195_groupi_n_4727 ,csa_tree_add_190_195_groupi_n_4728);
  not csa_tree_add_190_195_groupi_g44333(csa_tree_add_190_195_groupi_n_4725 ,csa_tree_add_190_195_groupi_n_4726);
  not csa_tree_add_190_195_groupi_g44334(csa_tree_add_190_195_groupi_n_4723 ,csa_tree_add_190_195_groupi_n_4724);
  not csa_tree_add_190_195_groupi_g44335(csa_tree_add_190_195_groupi_n_4722 ,csa_tree_add_190_195_groupi_n_4721);
  not csa_tree_add_190_195_groupi_g44336(csa_tree_add_190_195_groupi_n_4719 ,csa_tree_add_190_195_groupi_n_4720);
  not csa_tree_add_190_195_groupi_g44337(csa_tree_add_190_195_groupi_n_4717 ,csa_tree_add_190_195_groupi_n_4718);
  not csa_tree_add_190_195_groupi_g44338(csa_tree_add_190_195_groupi_n_4713 ,csa_tree_add_190_195_groupi_n_4714);
  not csa_tree_add_190_195_groupi_g44339(csa_tree_add_190_195_groupi_n_4711 ,csa_tree_add_190_195_groupi_n_4712);
  not csa_tree_add_190_195_groupi_g44340(csa_tree_add_190_195_groupi_n_4709 ,csa_tree_add_190_195_groupi_n_4710);
  not csa_tree_add_190_195_groupi_g44341(csa_tree_add_190_195_groupi_n_4708 ,csa_tree_add_190_195_groupi_n_4707);
  not csa_tree_add_190_195_groupi_g44342(csa_tree_add_190_195_groupi_n_4703 ,csa_tree_add_190_195_groupi_n_4704);
  not csa_tree_add_190_195_groupi_g44343(csa_tree_add_190_195_groupi_n_4702 ,csa_tree_add_190_195_groupi_n_4701);
  not csa_tree_add_190_195_groupi_g44344(csa_tree_add_190_195_groupi_n_4698 ,csa_tree_add_190_195_groupi_n_4699);
  not csa_tree_add_190_195_groupi_g44345(csa_tree_add_190_195_groupi_n_4695 ,csa_tree_add_190_195_groupi_n_4696);
  not csa_tree_add_190_195_groupi_g44346(csa_tree_add_190_195_groupi_n_4692 ,csa_tree_add_190_195_groupi_n_4693);
  not csa_tree_add_190_195_groupi_g44347(csa_tree_add_190_195_groupi_n_4687 ,csa_tree_add_190_195_groupi_n_4688);
  not csa_tree_add_190_195_groupi_g44348(csa_tree_add_190_195_groupi_n_4684 ,csa_tree_add_190_195_groupi_n_4685);
  not csa_tree_add_190_195_groupi_g44349(csa_tree_add_190_195_groupi_n_4681 ,csa_tree_add_190_195_groupi_n_4680);
  not csa_tree_add_190_195_groupi_g44350(csa_tree_add_190_195_groupi_n_4679 ,csa_tree_add_190_195_groupi_n_4678);
  not csa_tree_add_190_195_groupi_g44351(csa_tree_add_190_195_groupi_n_4674 ,csa_tree_add_190_195_groupi_n_4675);
  not csa_tree_add_190_195_groupi_g44352(csa_tree_add_190_195_groupi_n_4673 ,csa_tree_add_190_195_groupi_n_4672);
  not csa_tree_add_190_195_groupi_g44353(csa_tree_add_190_195_groupi_n_4667 ,csa_tree_add_190_195_groupi_n_4666);
  not csa_tree_add_190_195_groupi_g44354(csa_tree_add_190_195_groupi_n_4663 ,csa_tree_add_190_195_groupi_n_4664);
  not csa_tree_add_190_195_groupi_g44355(csa_tree_add_190_195_groupi_n_4662 ,csa_tree_add_190_195_groupi_n_4661);
  not csa_tree_add_190_195_groupi_g44356(csa_tree_add_190_195_groupi_n_4658 ,csa_tree_add_190_195_groupi_n_4659);
  not csa_tree_add_190_195_groupi_g44357(csa_tree_add_190_195_groupi_n_4657 ,csa_tree_add_190_195_groupi_n_4656);
  not csa_tree_add_190_195_groupi_g44358(csa_tree_add_190_195_groupi_n_4654 ,csa_tree_add_190_195_groupi_n_4655);
  not csa_tree_add_190_195_groupi_g44359(csa_tree_add_190_195_groupi_n_4652 ,csa_tree_add_190_195_groupi_n_4653);
  not csa_tree_add_190_195_groupi_g44360(csa_tree_add_190_195_groupi_n_4651 ,csa_tree_add_190_195_groupi_n_4650);
  not csa_tree_add_190_195_groupi_g44361(csa_tree_add_190_195_groupi_n_4648 ,csa_tree_add_190_195_groupi_n_4649);
  not csa_tree_add_190_195_groupi_g44362(csa_tree_add_190_195_groupi_n_4646 ,csa_tree_add_190_195_groupi_n_4645);
  not csa_tree_add_190_195_groupi_g44363(csa_tree_add_190_195_groupi_n_4641 ,csa_tree_add_190_195_groupi_n_4642);
  not csa_tree_add_190_195_groupi_g44364(csa_tree_add_190_195_groupi_n_4639 ,csa_tree_add_190_195_groupi_n_4640);
  not csa_tree_add_190_195_groupi_g44365(csa_tree_add_190_195_groupi_n_4637 ,csa_tree_add_190_195_groupi_n_4638);
  not csa_tree_add_190_195_groupi_g44366(csa_tree_add_190_195_groupi_n_4636 ,csa_tree_add_190_195_groupi_n_4635);
  not csa_tree_add_190_195_groupi_g44367(csa_tree_add_190_195_groupi_n_4634 ,csa_tree_add_190_195_groupi_n_4633);
  not csa_tree_add_190_195_groupi_g44368(csa_tree_add_190_195_groupi_n_4631 ,csa_tree_add_190_195_groupi_n_4632);
  not csa_tree_add_190_195_groupi_g44369(csa_tree_add_190_195_groupi_n_4629 ,csa_tree_add_190_195_groupi_n_4630);
  not csa_tree_add_190_195_groupi_g44370(csa_tree_add_190_195_groupi_n_4626 ,csa_tree_add_190_195_groupi_n_4627);
  not csa_tree_add_190_195_groupi_g44371(csa_tree_add_190_195_groupi_n_4624 ,csa_tree_add_190_195_groupi_n_4625);
  not csa_tree_add_190_195_groupi_g44372(csa_tree_add_190_195_groupi_n_4622 ,csa_tree_add_190_195_groupi_n_4623);
  not csa_tree_add_190_195_groupi_g44373(csa_tree_add_190_195_groupi_n_4620 ,csa_tree_add_190_195_groupi_n_4621);
  not csa_tree_add_190_195_groupi_g44374(csa_tree_add_190_195_groupi_n_4614 ,csa_tree_add_190_195_groupi_n_4615);
  not csa_tree_add_190_195_groupi_g44375(csa_tree_add_190_195_groupi_n_4610 ,csa_tree_add_190_195_groupi_n_4611);
  not csa_tree_add_190_195_groupi_g44376(csa_tree_add_190_195_groupi_n_4608 ,csa_tree_add_190_195_groupi_n_4609);
  not csa_tree_add_190_195_groupi_g44377(csa_tree_add_190_195_groupi_n_4607 ,csa_tree_add_190_195_groupi_n_4606);
  not csa_tree_add_190_195_groupi_g44378(csa_tree_add_190_195_groupi_n_4605 ,csa_tree_add_190_195_groupi_n_4604);
  not csa_tree_add_190_195_groupi_g44379(csa_tree_add_190_195_groupi_n_4602 ,csa_tree_add_190_195_groupi_n_4603);
  not csa_tree_add_190_195_groupi_g44380(csa_tree_add_190_195_groupi_n_4601 ,csa_tree_add_190_195_groupi_n_4600);
  not csa_tree_add_190_195_groupi_g44381(csa_tree_add_190_195_groupi_n_4598 ,csa_tree_add_190_195_groupi_n_4599);
  not csa_tree_add_190_195_groupi_g44382(csa_tree_add_190_195_groupi_n_4596 ,csa_tree_add_190_195_groupi_n_4597);
  not csa_tree_add_190_195_groupi_g44383(csa_tree_add_190_195_groupi_n_4594 ,csa_tree_add_190_195_groupi_n_4595);
  not csa_tree_add_190_195_groupi_g44384(csa_tree_add_190_195_groupi_n_4592 ,csa_tree_add_190_195_groupi_n_4593);
  not csa_tree_add_190_195_groupi_g44385(csa_tree_add_190_195_groupi_n_4589 ,csa_tree_add_190_195_groupi_n_4590);
  not csa_tree_add_190_195_groupi_g44386(csa_tree_add_190_195_groupi_n_4587 ,csa_tree_add_190_195_groupi_n_4588);
  not csa_tree_add_190_195_groupi_g44387(csa_tree_add_190_195_groupi_n_4585 ,csa_tree_add_190_195_groupi_n_4586);
  not csa_tree_add_190_195_groupi_g44388(csa_tree_add_190_195_groupi_n_4584 ,csa_tree_add_190_195_groupi_n_4583);
  not csa_tree_add_190_195_groupi_g44389(csa_tree_add_190_195_groupi_n_4581 ,csa_tree_add_190_195_groupi_n_4582);
  or csa_tree_add_190_195_groupi_g44390(csa_tree_add_190_195_groupi_n_4580 ,csa_tree_add_190_195_groupi_n_1846 ,csa_tree_add_190_195_groupi_n_4567);
  and csa_tree_add_190_195_groupi_g44391(csa_tree_add_190_195_groupi_n_4579 ,csa_tree_add_190_195_groupi_n_2955 ,csa_tree_add_190_195_groupi_n_4139);
  or csa_tree_add_190_195_groupi_g44392(csa_tree_add_190_195_groupi_n_4578 ,csa_tree_add_190_195_groupi_n_1499 ,csa_tree_add_190_195_groupi_n_4118);
  and csa_tree_add_190_195_groupi_g44393(csa_tree_add_190_195_groupi_n_4577 ,csa_tree_add_190_195_groupi_n_3488 ,csa_tree_add_190_195_groupi_n_4142);
  and csa_tree_add_190_195_groupi_g44394(csa_tree_add_190_195_groupi_n_4576 ,csa_tree_add_190_195_groupi_n_1498 ,csa_tree_add_190_195_groupi_n_4118);
  xnor csa_tree_add_190_195_groupi_g44395(csa_tree_add_190_195_groupi_n_4575 ,csa_tree_add_190_195_groupi_n_3205 ,in56[6]);
  xnor csa_tree_add_190_195_groupi_g44396(csa_tree_add_190_195_groupi_n_4574 ,csa_tree_add_190_195_groupi_n_3207 ,in56[8]);
  xnor csa_tree_add_190_195_groupi_g44397(csa_tree_add_190_195_groupi_n_4573 ,csa_tree_add_190_195_groupi_n_3206 ,in55[15]);
  xnor csa_tree_add_190_195_groupi_g44398(csa_tree_add_190_195_groupi_n_4572 ,csa_tree_add_190_195_groupi_n_3704 ,csa_tree_add_190_195_groupi_n_1995);
  xnor csa_tree_add_190_195_groupi_g44399(csa_tree_add_190_195_groupi_n_4571 ,csa_tree_add_190_195_groupi_n_3701 ,csa_tree_add_190_195_groupi_n_2209);
  or csa_tree_add_190_195_groupi_g44400(csa_tree_add_190_195_groupi_n_4872 ,csa_tree_add_190_195_groupi_n_3077 ,csa_tree_add_190_195_groupi_n_4186);
  and csa_tree_add_190_195_groupi_g44401(csa_tree_add_190_195_groupi_n_4871 ,csa_tree_add_190_195_groupi_n_2779 ,csa_tree_add_190_195_groupi_n_4532);
  or csa_tree_add_190_195_groupi_g44402(csa_tree_add_190_195_groupi_n_4870 ,csa_tree_add_190_195_groupi_n_3468 ,csa_tree_add_190_195_groupi_n_4359);
  or csa_tree_add_190_195_groupi_g44403(csa_tree_add_190_195_groupi_n_4869 ,csa_tree_add_190_195_groupi_n_3639 ,csa_tree_add_190_195_groupi_n_4468);
  or csa_tree_add_190_195_groupi_g44404(csa_tree_add_190_195_groupi_n_4867 ,csa_tree_add_190_195_groupi_n_3563 ,csa_tree_add_190_195_groupi_n_4382);
  and csa_tree_add_190_195_groupi_g44405(csa_tree_add_190_195_groupi_n_4866 ,csa_tree_add_190_195_groupi_n_2871 ,csa_tree_add_190_195_groupi_n_4170);
  or csa_tree_add_190_195_groupi_g44406(csa_tree_add_190_195_groupi_n_4865 ,csa_tree_add_190_195_groupi_n_3709 ,csa_tree_add_190_195_groupi_n_4236);
  or csa_tree_add_190_195_groupi_g44407(csa_tree_add_190_195_groupi_n_4863 ,csa_tree_add_190_195_groupi_n_3710 ,csa_tree_add_190_195_groupi_n_4503);
  and csa_tree_add_190_195_groupi_g44408(csa_tree_add_190_195_groupi_n_4862 ,csa_tree_add_190_195_groupi_n_3127 ,csa_tree_add_190_195_groupi_n_4275);
  or csa_tree_add_190_195_groupi_g44409(csa_tree_add_190_195_groupi_n_4861 ,csa_tree_add_190_195_groupi_n_2737 ,csa_tree_add_190_195_groupi_n_4509);
  or csa_tree_add_190_195_groupi_g44410(csa_tree_add_190_195_groupi_n_4860 ,csa_tree_add_190_195_groupi_n_3549 ,csa_tree_add_190_195_groupi_n_4407);
  or csa_tree_add_190_195_groupi_g44411(csa_tree_add_190_195_groupi_n_4858 ,csa_tree_add_190_195_groupi_n_3538 ,csa_tree_add_190_195_groupi_n_4287);
  and csa_tree_add_190_195_groupi_g44412(csa_tree_add_190_195_groupi_n_4857 ,csa_tree_add_190_195_groupi_n_3499 ,csa_tree_add_190_195_groupi_n_4427);
  or csa_tree_add_190_195_groupi_g44413(csa_tree_add_190_195_groupi_n_4856 ,csa_tree_add_190_195_groupi_n_3119 ,csa_tree_add_190_195_groupi_n_4535);
  or csa_tree_add_190_195_groupi_g44414(csa_tree_add_190_195_groupi_n_4855 ,csa_tree_add_190_195_groupi_n_3420 ,csa_tree_add_190_195_groupi_n_4345);
  or csa_tree_add_190_195_groupi_g44415(csa_tree_add_190_195_groupi_n_4853 ,csa_tree_add_190_195_groupi_n_3324 ,csa_tree_add_190_195_groupi_n_4208);
  and csa_tree_add_190_195_groupi_g44416(csa_tree_add_190_195_groupi_n_4852 ,csa_tree_add_190_195_groupi_n_3215 ,csa_tree_add_190_195_groupi_n_4173);
  or csa_tree_add_190_195_groupi_g44417(csa_tree_add_190_195_groupi_n_4851 ,csa_tree_add_190_195_groupi_n_2928 ,csa_tree_add_190_195_groupi_n_4555);
  and csa_tree_add_190_195_groupi_g44418(csa_tree_add_190_195_groupi_n_4850 ,csa_tree_add_190_195_groupi_n_3042 ,csa_tree_add_190_195_groupi_n_4508);
  or csa_tree_add_190_195_groupi_g44419(csa_tree_add_190_195_groupi_n_4849 ,csa_tree_add_190_195_groupi_n_3209 ,csa_tree_add_190_195_groupi_n_4446);
  or csa_tree_add_190_195_groupi_g44420(csa_tree_add_190_195_groupi_n_4848 ,csa_tree_add_190_195_groupi_n_3051 ,csa_tree_add_190_195_groupi_n_4506);
  and csa_tree_add_190_195_groupi_g44421(csa_tree_add_190_195_groupi_n_4847 ,csa_tree_add_190_195_groupi_n_3250 ,csa_tree_add_190_195_groupi_n_4365);
  or csa_tree_add_190_195_groupi_g44422(csa_tree_add_190_195_groupi_n_4846 ,csa_tree_add_190_195_groupi_n_3306 ,csa_tree_add_190_195_groupi_n_4353);
  and csa_tree_add_190_195_groupi_g44423(csa_tree_add_190_195_groupi_n_4845 ,csa_tree_add_190_195_groupi_n_3568 ,csa_tree_add_190_195_groupi_n_4381);
  and csa_tree_add_190_195_groupi_g44424(csa_tree_add_190_195_groupi_n_4844 ,csa_tree_add_190_195_groupi_n_2890 ,csa_tree_add_190_195_groupi_n_4419);
  and csa_tree_add_190_195_groupi_g44425(csa_tree_add_190_195_groupi_n_4843 ,csa_tree_add_190_195_groupi_n_3708 ,csa_tree_add_190_195_groupi_n_4442);
  or csa_tree_add_190_195_groupi_g44426(csa_tree_add_190_195_groupi_n_4842 ,csa_tree_add_190_195_groupi_n_3088 ,csa_tree_add_190_195_groupi_n_4418);
  and csa_tree_add_190_195_groupi_g44427(csa_tree_add_190_195_groupi_n_4841 ,csa_tree_add_190_195_groupi_n_3564 ,csa_tree_add_190_195_groupi_n_4411);
  and csa_tree_add_190_195_groupi_g44428(csa_tree_add_190_195_groupi_n_4840 ,csa_tree_add_190_195_groupi_n_3396 ,csa_tree_add_190_195_groupi_n_4398);
  and csa_tree_add_190_195_groupi_g44429(csa_tree_add_190_195_groupi_n_4839 ,csa_tree_add_190_195_groupi_n_2951 ,csa_tree_add_190_195_groupi_n_4495);
  and csa_tree_add_190_195_groupi_g44430(csa_tree_add_190_195_groupi_n_4838 ,csa_tree_add_190_195_groupi_n_3271 ,csa_tree_add_190_195_groupi_n_4179);
  and csa_tree_add_190_195_groupi_g44431(csa_tree_add_190_195_groupi_n_4837 ,csa_tree_add_190_195_groupi_n_3059 ,csa_tree_add_190_195_groupi_n_4270);
  or csa_tree_add_190_195_groupi_g44432(csa_tree_add_190_195_groupi_n_4836 ,csa_tree_add_190_195_groupi_n_3321 ,csa_tree_add_190_195_groupi_n_4201);
  or csa_tree_add_190_195_groupi_g44434(csa_tree_add_190_195_groupi_n_4833 ,csa_tree_add_190_195_groupi_n_3216 ,csa_tree_add_190_195_groupi_n_4336);
  and csa_tree_add_190_195_groupi_g44435(csa_tree_add_190_195_groupi_n_4832 ,csa_tree_add_190_195_groupi_n_2935 ,csa_tree_add_190_195_groupi_n_4211);
  and csa_tree_add_190_195_groupi_g44436(csa_tree_add_190_195_groupi_n_4831 ,csa_tree_add_190_195_groupi_n_2893 ,csa_tree_add_190_195_groupi_n_4175);
  and csa_tree_add_190_195_groupi_g44437(csa_tree_add_190_195_groupi_n_4830 ,csa_tree_add_190_195_groupi_n_3283 ,csa_tree_add_190_195_groupi_n_4459);
  or csa_tree_add_190_195_groupi_g44438(csa_tree_add_190_195_groupi_n_4829 ,csa_tree_add_190_195_groupi_n_3071 ,csa_tree_add_190_195_groupi_n_4151);
  and csa_tree_add_190_195_groupi_g44439(csa_tree_add_190_195_groupi_n_4828 ,csa_tree_add_190_195_groupi_n_2823 ,csa_tree_add_190_195_groupi_n_4518);
  or csa_tree_add_190_195_groupi_g44440(csa_tree_add_190_195_groupi_n_4827 ,csa_tree_add_190_195_groupi_n_3177 ,csa_tree_add_190_195_groupi_n_4182);
  or csa_tree_add_190_195_groupi_g44441(csa_tree_add_190_195_groupi_n_4826 ,csa_tree_add_190_195_groupi_n_3624 ,csa_tree_add_190_195_groupi_n_4355);
  and csa_tree_add_190_195_groupi_g44442(csa_tree_add_190_195_groupi_n_4825 ,csa_tree_add_190_195_groupi_n_2917 ,csa_tree_add_190_195_groupi_n_4420);
  and csa_tree_add_190_195_groupi_g44443(csa_tree_add_190_195_groupi_n_4824 ,csa_tree_add_190_195_groupi_n_3527 ,csa_tree_add_190_195_groupi_n_4213);
  or csa_tree_add_190_195_groupi_g44444(csa_tree_add_190_195_groupi_n_4822 ,csa_tree_add_190_195_groupi_n_3245 ,csa_tree_add_190_195_groupi_n_4311);
  or csa_tree_add_190_195_groupi_g44445(csa_tree_add_190_195_groupi_n_4821 ,csa_tree_add_190_195_groupi_n_3718 ,csa_tree_add_190_195_groupi_n_4290);
  or csa_tree_add_190_195_groupi_g44446(csa_tree_add_190_195_groupi_n_4820 ,csa_tree_add_190_195_groupi_n_3584 ,csa_tree_add_190_195_groupi_n_4229);
  or csa_tree_add_190_195_groupi_g44447(csa_tree_add_190_195_groupi_n_4818 ,csa_tree_add_190_195_groupi_n_3295 ,csa_tree_add_190_195_groupi_n_4225);
  and csa_tree_add_190_195_groupi_g44448(csa_tree_add_190_195_groupi_n_4817 ,csa_tree_add_190_195_groupi_n_3501 ,csa_tree_add_190_195_groupi_n_4525);
  and csa_tree_add_190_195_groupi_g44449(csa_tree_add_190_195_groupi_n_4816 ,csa_tree_add_190_195_groupi_n_3526 ,csa_tree_add_190_195_groupi_n_4199);
  or csa_tree_add_190_195_groupi_g44450(csa_tree_add_190_195_groupi_n_4815 ,csa_tree_add_190_195_groupi_n_2938 ,csa_tree_add_190_195_groupi_n_4543);
  and csa_tree_add_190_195_groupi_g44451(csa_tree_add_190_195_groupi_n_4814 ,csa_tree_add_190_195_groupi_n_2881 ,csa_tree_add_190_195_groupi_n_4318);
  and csa_tree_add_190_195_groupi_g44452(csa_tree_add_190_195_groupi_n_4813 ,csa_tree_add_190_195_groupi_n_3288 ,csa_tree_add_190_195_groupi_n_4370);
  or csa_tree_add_190_195_groupi_g44453(csa_tree_add_190_195_groupi_n_4812 ,csa_tree_add_190_195_groupi_n_3617 ,csa_tree_add_190_195_groupi_n_4329);
  or csa_tree_add_190_195_groupi_g44454(csa_tree_add_190_195_groupi_n_4811 ,csa_tree_add_190_195_groupi_n_3080 ,csa_tree_add_190_195_groupi_n_4536);
  or csa_tree_add_190_195_groupi_g44455(csa_tree_add_190_195_groupi_n_4809 ,csa_tree_add_190_195_groupi_n_3316 ,csa_tree_add_190_195_groupi_n_4375);
  and csa_tree_add_190_195_groupi_g44456(csa_tree_add_190_195_groupi_n_4808 ,csa_tree_add_190_195_groupi_n_3197 ,csa_tree_add_190_195_groupi_n_4484);
  and csa_tree_add_190_195_groupi_g44457(csa_tree_add_190_195_groupi_n_4807 ,csa_tree_add_190_195_groupi_n_3325 ,csa_tree_add_190_195_groupi_n_4402);
  and csa_tree_add_190_195_groupi_g44458(csa_tree_add_190_195_groupi_n_4806 ,csa_tree_add_190_195_groupi_n_3315 ,csa_tree_add_190_195_groupi_n_4155);
  and csa_tree_add_190_195_groupi_g44459(csa_tree_add_190_195_groupi_n_4805 ,csa_tree_add_190_195_groupi_n_3260 ,csa_tree_add_190_195_groupi_n_4492);
  or csa_tree_add_190_195_groupi_g44460(csa_tree_add_190_195_groupi_n_4804 ,csa_tree_add_190_195_groupi_n_3126 ,csa_tree_add_190_195_groupi_n_4434);
  or csa_tree_add_190_195_groupi_g44461(csa_tree_add_190_195_groupi_n_4803 ,csa_tree_add_190_195_groupi_n_3117 ,csa_tree_add_190_195_groupi_n_4443);
  and csa_tree_add_190_195_groupi_g44462(csa_tree_add_190_195_groupi_n_4802 ,csa_tree_add_190_195_groupi_n_3534 ,csa_tree_add_190_195_groupi_n_4257);
  and csa_tree_add_190_195_groupi_g44463(csa_tree_add_190_195_groupi_n_4801 ,csa_tree_add_190_195_groupi_n_3679 ,csa_tree_add_190_195_groupi_n_4149);
  or csa_tree_add_190_195_groupi_g44464(csa_tree_add_190_195_groupi_n_4800 ,csa_tree_add_190_195_groupi_n_3469 ,csa_tree_add_190_195_groupi_n_4268);
  or csa_tree_add_190_195_groupi_g44465(csa_tree_add_190_195_groupi_n_4799 ,csa_tree_add_190_195_groupi_n_3600 ,csa_tree_add_190_195_groupi_n_4185);
  and csa_tree_add_190_195_groupi_g44466(csa_tree_add_190_195_groupi_n_4798 ,csa_tree_add_190_195_groupi_n_3474 ,csa_tree_add_190_195_groupi_n_4299);
  or csa_tree_add_190_195_groupi_g44467(csa_tree_add_190_195_groupi_n_4797 ,csa_tree_add_190_195_groupi_n_3058 ,csa_tree_add_190_195_groupi_n_4426);
  and csa_tree_add_190_195_groupi_g44468(csa_tree_add_190_195_groupi_n_4796 ,csa_tree_add_190_195_groupi_n_3401 ,csa_tree_add_190_195_groupi_n_4342);
  or csa_tree_add_190_195_groupi_g44469(csa_tree_add_190_195_groupi_n_4794 ,csa_tree_add_190_195_groupi_n_3173 ,csa_tree_add_190_195_groupi_n_4558);
  or csa_tree_add_190_195_groupi_g44470(csa_tree_add_190_195_groupi_n_4793 ,csa_tree_add_190_195_groupi_n_3379 ,csa_tree_add_190_195_groupi_n_4216);
  and csa_tree_add_190_195_groupi_g44471(csa_tree_add_190_195_groupi_n_4791 ,csa_tree_add_190_195_groupi_n_3131 ,csa_tree_add_190_195_groupi_n_4501);
  and csa_tree_add_190_195_groupi_g44472(csa_tree_add_190_195_groupi_n_4789 ,csa_tree_add_190_195_groupi_n_3337 ,csa_tree_add_190_195_groupi_n_4263);
  and csa_tree_add_190_195_groupi_g44473(csa_tree_add_190_195_groupi_n_4787 ,csa_tree_add_190_195_groupi_n_3494 ,csa_tree_add_190_195_groupi_n_4297);
  and csa_tree_add_190_195_groupi_g44474(csa_tree_add_190_195_groupi_n_4785 ,csa_tree_add_190_195_groupi_n_3066 ,csa_tree_add_190_195_groupi_n_4251);
  or csa_tree_add_190_195_groupi_g44475(csa_tree_add_190_195_groupi_n_4783 ,csa_tree_add_190_195_groupi_n_3193 ,csa_tree_add_190_195_groupi_n_4529);
  and csa_tree_add_190_195_groupi_g44476(csa_tree_add_190_195_groupi_n_4782 ,csa_tree_add_190_195_groupi_n_2765 ,csa_tree_add_190_195_groupi_n_4261);
  or csa_tree_add_190_195_groupi_g44477(csa_tree_add_190_195_groupi_n_4781 ,csa_tree_add_190_195_groupi_n_2850 ,csa_tree_add_190_195_groupi_n_4183);
  or csa_tree_add_190_195_groupi_g44478(csa_tree_add_190_195_groupi_n_4780 ,csa_tree_add_190_195_groupi_n_3002 ,csa_tree_add_190_195_groupi_n_4436);
  and csa_tree_add_190_195_groupi_g44479(csa_tree_add_190_195_groupi_n_4777 ,csa_tree_add_190_195_groupi_n_3213 ,csa_tree_add_190_195_groupi_n_4165);
  or csa_tree_add_190_195_groupi_g44480(csa_tree_add_190_195_groupi_n_4776 ,csa_tree_add_190_195_groupi_n_2904 ,csa_tree_add_190_195_groupi_n_4511);
  or csa_tree_add_190_195_groupi_g44481(csa_tree_add_190_195_groupi_n_4775 ,csa_tree_add_190_195_groupi_n_3178 ,csa_tree_add_190_195_groupi_n_4490);
  and csa_tree_add_190_195_groupi_g44482(csa_tree_add_190_195_groupi_n_4773 ,csa_tree_add_190_195_groupi_n_3275 ,csa_tree_add_190_195_groupi_n_4313);
  or csa_tree_add_190_195_groupi_g44483(csa_tree_add_190_195_groupi_n_4771 ,csa_tree_add_190_195_groupi_n_3400 ,csa_tree_add_190_195_groupi_n_4224);
  and csa_tree_add_190_195_groupi_g44484(csa_tree_add_190_195_groupi_n_4769 ,csa_tree_add_190_195_groupi_n_2842 ,csa_tree_add_190_195_groupi_n_4207);
  or csa_tree_add_190_195_groupi_g44485(csa_tree_add_190_195_groupi_n_4767 ,csa_tree_add_190_195_groupi_n_3034 ,csa_tree_add_190_195_groupi_n_4439);
  or csa_tree_add_190_195_groupi_g44486(csa_tree_add_190_195_groupi_n_4765 ,csa_tree_add_190_195_groupi_n_2943 ,csa_tree_add_190_195_groupi_n_4507);
  or csa_tree_add_190_195_groupi_g44487(csa_tree_add_190_195_groupi_n_4763 ,csa_tree_add_190_195_groupi_n_2934 ,csa_tree_add_190_195_groupi_n_4475);
  and csa_tree_add_190_195_groupi_g44488(csa_tree_add_190_195_groupi_n_4760 ,csa_tree_add_190_195_groupi_n_2963 ,csa_tree_add_190_195_groupi_n_4328);
  and csa_tree_add_190_195_groupi_g44489(csa_tree_add_190_195_groupi_n_4759 ,csa_tree_add_190_195_groupi_n_2791 ,csa_tree_add_190_195_groupi_n_4321);
  and csa_tree_add_190_195_groupi_g44490(csa_tree_add_190_195_groupi_n_4758 ,csa_tree_add_190_195_groupi_n_3460 ,csa_tree_add_190_195_groupi_n_4454);
  or csa_tree_add_190_195_groupi_g44491(csa_tree_add_190_195_groupi_n_4757 ,csa_tree_add_190_195_groupi_n_3365 ,csa_tree_add_190_195_groupi_n_4194);
  and csa_tree_add_190_195_groupi_g44492(csa_tree_add_190_195_groupi_n_4756 ,csa_tree_add_190_195_groupi_n_2758 ,csa_tree_add_190_195_groupi_n_4456);
  or csa_tree_add_190_195_groupi_g44493(csa_tree_add_190_195_groupi_n_4755 ,csa_tree_add_190_195_groupi_n_2774 ,csa_tree_add_190_195_groupi_n_4522);
  or csa_tree_add_190_195_groupi_g44494(csa_tree_add_190_195_groupi_n_4753 ,csa_tree_add_190_195_groupi_n_3508 ,csa_tree_add_190_195_groupi_n_4517);
  and csa_tree_add_190_195_groupi_g44495(csa_tree_add_190_195_groupi_n_4752 ,csa_tree_add_190_195_groupi_n_3495 ,csa_tree_add_190_195_groupi_n_4424);
  or csa_tree_add_190_195_groupi_g44496(csa_tree_add_190_195_groupi_n_4751 ,csa_tree_add_190_195_groupi_n_2997 ,csa_tree_add_190_195_groupi_n_4547);
  and csa_tree_add_190_195_groupi_g44497(csa_tree_add_190_195_groupi_n_4749 ,csa_tree_add_190_195_groupi_n_3004 ,csa_tree_add_190_195_groupi_n_4154);
  or csa_tree_add_190_195_groupi_g44498(csa_tree_add_190_195_groupi_n_4748 ,csa_tree_add_190_195_groupi_n_3262 ,csa_tree_add_190_195_groupi_n_4291);
  and csa_tree_add_190_195_groupi_g44499(csa_tree_add_190_195_groupi_n_4745 ,csa_tree_add_190_195_groupi_n_2747 ,csa_tree_add_190_195_groupi_n_4331);
  or csa_tree_add_190_195_groupi_g44500(csa_tree_add_190_195_groupi_n_4744 ,csa_tree_add_190_195_groupi_n_3329 ,csa_tree_add_190_195_groupi_n_4230);
  and csa_tree_add_190_195_groupi_g44501(csa_tree_add_190_195_groupi_n_4743 ,csa_tree_add_190_195_groupi_n_3130 ,csa_tree_add_190_195_groupi_n_4441);
  or csa_tree_add_190_195_groupi_g44502(csa_tree_add_190_195_groupi_n_4741 ,csa_tree_add_190_195_groupi_n_3728 ,csa_tree_add_190_195_groupi_n_4378);
  and csa_tree_add_190_195_groupi_g44503(csa_tree_add_190_195_groupi_n_4739 ,csa_tree_add_190_195_groupi_n_3168 ,csa_tree_add_190_195_groupi_n_4278);
  or csa_tree_add_190_195_groupi_g44504(csa_tree_add_190_195_groupi_n_4737 ,csa_tree_add_190_195_groupi_n_3243 ,csa_tree_add_190_195_groupi_n_4262);
  and csa_tree_add_190_195_groupi_g44505(csa_tree_add_190_195_groupi_n_4736 ,csa_tree_add_190_195_groupi_n_2769 ,csa_tree_add_190_195_groupi_n_4489);
  or csa_tree_add_190_195_groupi_g44506(csa_tree_add_190_195_groupi_n_4734 ,csa_tree_add_190_195_groupi_n_3472 ,csa_tree_add_190_195_groupi_n_4390);
  or csa_tree_add_190_195_groupi_g44507(csa_tree_add_190_195_groupi_n_4732 ,csa_tree_add_190_195_groupi_n_2849 ,csa_tree_add_190_195_groupi_n_4516);
  or csa_tree_add_190_195_groupi_g44508(csa_tree_add_190_195_groupi_n_4731 ,csa_tree_add_190_195_groupi_n_3320 ,csa_tree_add_190_195_groupi_n_4223);
  or csa_tree_add_190_195_groupi_g44509(csa_tree_add_190_195_groupi_n_4729 ,csa_tree_add_190_195_groupi_n_3660 ,csa_tree_add_190_195_groupi_n_4449);
  or csa_tree_add_190_195_groupi_g44510(csa_tree_add_190_195_groupi_n_4728 ,csa_tree_add_190_195_groupi_n_3642 ,csa_tree_add_190_195_groupi_n_4469);
  and csa_tree_add_190_195_groupi_g44511(csa_tree_add_190_195_groupi_n_4726 ,csa_tree_add_190_195_groupi_n_3388 ,csa_tree_add_190_195_groupi_n_4388);
  or csa_tree_add_190_195_groupi_g44512(csa_tree_add_190_195_groupi_n_4724 ,csa_tree_add_190_195_groupi_n_3598 ,csa_tree_add_190_195_groupi_n_4255);
  or csa_tree_add_190_195_groupi_g44513(csa_tree_add_190_195_groupi_n_4721 ,csa_tree_add_190_195_groupi_n_3724 ,csa_tree_add_190_195_groupi_n_4169);
  or csa_tree_add_190_195_groupi_g44514(csa_tree_add_190_195_groupi_n_4720 ,csa_tree_add_190_195_groupi_n_3184 ,csa_tree_add_190_195_groupi_n_4514);
  or csa_tree_add_190_195_groupi_g44515(csa_tree_add_190_195_groupi_n_4718 ,csa_tree_add_190_195_groupi_n_3713 ,csa_tree_add_190_195_groupi_n_4217);
  or csa_tree_add_190_195_groupi_g44516(csa_tree_add_190_195_groupi_n_4716 ,csa_tree_add_190_195_groupi_n_2886 ,csa_tree_add_190_195_groupi_n_4539);
  or csa_tree_add_190_195_groupi_g44517(csa_tree_add_190_195_groupi_n_4715 ,csa_tree_add_190_195_groupi_n_3128 ,csa_tree_add_190_195_groupi_n_4455);
  and csa_tree_add_190_195_groupi_g44518(csa_tree_add_190_195_groupi_n_4714 ,csa_tree_add_190_195_groupi_n_2991 ,csa_tree_add_190_195_groupi_n_4521);
  or csa_tree_add_190_195_groupi_g44519(csa_tree_add_190_195_groupi_n_4712 ,csa_tree_add_190_195_groupi_n_3313 ,csa_tree_add_190_195_groupi_n_4187);
  or csa_tree_add_190_195_groupi_g44520(csa_tree_add_190_195_groupi_n_4710 ,csa_tree_add_190_195_groupi_n_3286 ,csa_tree_add_190_195_groupi_n_4338);
  and csa_tree_add_190_195_groupi_g44521(csa_tree_add_190_195_groupi_n_4707 ,csa_tree_add_190_195_groupi_n_2761 ,csa_tree_add_190_195_groupi_n_4319);
  or csa_tree_add_190_195_groupi_g44522(csa_tree_add_190_195_groupi_n_4706 ,csa_tree_add_190_195_groupi_n_3418 ,csa_tree_add_190_195_groupi_n_4198);
  and csa_tree_add_190_195_groupi_g44523(csa_tree_add_190_195_groupi_n_4705 ,csa_tree_add_190_195_groupi_n_3725 ,csa_tree_add_190_195_groupi_n_4428);
  and csa_tree_add_190_195_groupi_g44524(csa_tree_add_190_195_groupi_n_4704 ,csa_tree_add_190_195_groupi_n_3199 ,csa_tree_add_190_195_groupi_n_4239);
  and csa_tree_add_190_195_groupi_g44525(csa_tree_add_190_195_groupi_n_4701 ,csa_tree_add_190_195_groupi_n_2865 ,csa_tree_add_190_195_groupi_n_4258);
  or csa_tree_add_190_195_groupi_g44526(csa_tree_add_190_195_groupi_n_4700 ,csa_tree_add_190_195_groupi_n_2752 ,csa_tree_add_190_195_groupi_n_4364);
  or csa_tree_add_190_195_groupi_g44527(csa_tree_add_190_195_groupi_n_4699 ,csa_tree_add_190_195_groupi_n_3423 ,csa_tree_add_190_195_groupi_n_4197);
  or csa_tree_add_190_195_groupi_g44528(csa_tree_add_190_195_groupi_n_4697 ,csa_tree_add_190_195_groupi_n_3234 ,csa_tree_add_190_195_groupi_n_4180);
  or csa_tree_add_190_195_groupi_g44529(csa_tree_add_190_195_groupi_n_4696 ,csa_tree_add_190_195_groupi_n_2800 ,csa_tree_add_190_195_groupi_n_4421);
  and csa_tree_add_190_195_groupi_g44530(csa_tree_add_190_195_groupi_n_4694 ,csa_tree_add_190_195_groupi_n_2825 ,csa_tree_add_190_195_groupi_n_4235);
  or csa_tree_add_190_195_groupi_g44531(csa_tree_add_190_195_groupi_n_4693 ,csa_tree_add_190_195_groupi_n_3622 ,csa_tree_add_190_195_groupi_n_4540);
  or csa_tree_add_190_195_groupi_g44532(csa_tree_add_190_195_groupi_n_4691 ,csa_tree_add_190_195_groupi_n_2841 ,csa_tree_add_190_195_groupi_n_4416);
  and csa_tree_add_190_195_groupi_g44533(csa_tree_add_190_195_groupi_n_4690 ,csa_tree_add_190_195_groupi_n_3708 ,csa_tree_add_190_195_groupi_n_4192);
  or csa_tree_add_190_195_groupi_g44534(csa_tree_add_190_195_groupi_n_4689 ,csa_tree_add_190_195_groupi_n_3609 ,csa_tree_add_190_195_groupi_n_4188);
  and csa_tree_add_190_195_groupi_g44535(csa_tree_add_190_195_groupi_n_4688 ,csa_tree_add_190_195_groupi_n_3583 ,csa_tree_add_190_195_groupi_n_4256);
  or csa_tree_add_190_195_groupi_g44536(csa_tree_add_190_195_groupi_n_4686 ,csa_tree_add_190_195_groupi_n_3048 ,csa_tree_add_190_195_groupi_n_4548);
  and csa_tree_add_190_195_groupi_g44537(csa_tree_add_190_195_groupi_n_4685 ,csa_tree_add_190_195_groupi_n_3529 ,csa_tree_add_190_195_groupi_n_4386);
  or csa_tree_add_190_195_groupi_g44538(csa_tree_add_190_195_groupi_n_4683 ,csa_tree_add_190_195_groupi_n_3530 ,csa_tree_add_190_195_groupi_n_4233);
  or csa_tree_add_190_195_groupi_g44539(csa_tree_add_190_195_groupi_n_4682 ,csa_tree_add_190_195_groupi_n_3415 ,csa_tree_add_190_195_groupi_n_4189);
  and csa_tree_add_190_195_groupi_g44540(csa_tree_add_190_195_groupi_n_4680 ,csa_tree_add_190_195_groupi_n_2981 ,csa_tree_add_190_195_groupi_n_4228);
  and csa_tree_add_190_195_groupi_g44541(csa_tree_add_190_195_groupi_n_4678 ,csa_tree_add_190_195_groupi_n_2786 ,csa_tree_add_190_195_groupi_n_4191);
  and csa_tree_add_190_195_groupi_g44542(csa_tree_add_190_195_groupi_n_4677 ,csa_tree_add_190_195_groupi_n_2830 ,csa_tree_add_190_195_groupi_n_4172);
  or csa_tree_add_190_195_groupi_g44543(csa_tree_add_190_195_groupi_n_4676 ,csa_tree_add_190_195_groupi_n_3405 ,csa_tree_add_190_195_groupi_n_4148);
  or csa_tree_add_190_195_groupi_g44544(csa_tree_add_190_195_groupi_n_4675 ,csa_tree_add_190_195_groupi_n_3371 ,csa_tree_add_190_195_groupi_n_4396);
  and csa_tree_add_190_195_groupi_g44545(csa_tree_add_190_195_groupi_n_4672 ,csa_tree_add_190_195_groupi_n_2821 ,csa_tree_add_190_195_groupi_n_4204);
  or csa_tree_add_190_195_groupi_g44546(csa_tree_add_190_195_groupi_n_4671 ,csa_tree_add_190_195_groupi_n_3172 ,csa_tree_add_190_195_groupi_n_4432);
  or csa_tree_add_190_195_groupi_g44547(csa_tree_add_190_195_groupi_n_4670 ,csa_tree_add_190_195_groupi_n_3257 ,csa_tree_add_190_195_groupi_n_4162);
  or csa_tree_add_190_195_groupi_g44548(csa_tree_add_190_195_groupi_n_4669 ,csa_tree_add_190_195_groupi_n_2887 ,csa_tree_add_190_195_groupi_n_4349);
  or csa_tree_add_190_195_groupi_g44549(csa_tree_add_190_195_groupi_n_4668 ,csa_tree_add_190_195_groupi_n_2797 ,csa_tree_add_190_195_groupi_n_4533);
  or csa_tree_add_190_195_groupi_g44550(csa_tree_add_190_195_groupi_n_4666 ,csa_tree_add_190_195_groupi_n_2880 ,csa_tree_add_190_195_groupi_n_4284);
  or csa_tree_add_190_195_groupi_g44551(csa_tree_add_190_195_groupi_n_4665 ,csa_tree_add_190_195_groupi_n_3710 ,csa_tree_add_190_195_groupi_n_4350);
  or csa_tree_add_190_195_groupi_g44552(csa_tree_add_190_195_groupi_n_4664 ,csa_tree_add_190_195_groupi_n_2915 ,csa_tree_add_190_195_groupi_n_4542);
  or csa_tree_add_190_195_groupi_g44553(csa_tree_add_190_195_groupi_n_4661 ,csa_tree_add_190_195_groupi_n_3347 ,csa_tree_add_190_195_groupi_n_4214);
  and csa_tree_add_190_195_groupi_g44554(csa_tree_add_190_195_groupi_n_4660 ,csa_tree_add_190_195_groupi_n_3350 ,csa_tree_add_190_195_groupi_n_4404);
  or csa_tree_add_190_195_groupi_g44555(csa_tree_add_190_195_groupi_n_4659 ,csa_tree_add_190_195_groupi_n_2843 ,csa_tree_add_190_195_groupi_n_4417);
  and csa_tree_add_190_195_groupi_g44556(csa_tree_add_190_195_groupi_n_4656 ,csa_tree_add_190_195_groupi_n_3537 ,csa_tree_add_190_195_groupi_n_4296);
  or csa_tree_add_190_195_groupi_g44557(csa_tree_add_190_195_groupi_n_4655 ,csa_tree_add_190_195_groupi_n_2949 ,csa_tree_add_190_195_groupi_n_4526);
  or csa_tree_add_190_195_groupi_g44558(csa_tree_add_190_195_groupi_n_4653 ,csa_tree_add_190_195_groupi_n_3606 ,csa_tree_add_190_195_groupi_n_4409);
  or csa_tree_add_190_195_groupi_g44559(csa_tree_add_190_195_groupi_n_4650 ,csa_tree_add_190_195_groupi_n_3513 ,csa_tree_add_190_195_groupi_n_4206);
  or csa_tree_add_190_195_groupi_g44560(csa_tree_add_190_195_groupi_n_4649 ,csa_tree_add_190_195_groupi_n_3096 ,csa_tree_add_190_195_groupi_n_4462);
  or csa_tree_add_190_195_groupi_g44561(csa_tree_add_190_195_groupi_n_4647 ,csa_tree_add_190_195_groupi_n_2906 ,csa_tree_add_190_195_groupi_n_4161);
  and csa_tree_add_190_195_groupi_g44562(csa_tree_add_190_195_groupi_n_4645 ,csa_tree_add_190_195_groupi_n_2909 ,csa_tree_add_190_195_groupi_n_4190);
  or csa_tree_add_190_195_groupi_g44563(csa_tree_add_190_195_groupi_n_4644 ,csa_tree_add_190_195_groupi_n_3554 ,csa_tree_add_190_195_groupi_n_4408);
  or csa_tree_add_190_195_groupi_g44564(csa_tree_add_190_195_groupi_n_4643 ,csa_tree_add_190_195_groupi_n_3164 ,csa_tree_add_190_195_groupi_n_4377);
  or csa_tree_add_190_195_groupi_g44565(csa_tree_add_190_195_groupi_n_4642 ,csa_tree_add_190_195_groupi_n_3248 ,csa_tree_add_190_195_groupi_n_4369);
  or csa_tree_add_190_195_groupi_g44566(csa_tree_add_190_195_groupi_n_4640 ,csa_tree_add_190_195_groupi_n_3411 ,csa_tree_add_190_195_groupi_n_4288);
  and csa_tree_add_190_195_groupi_g44567(csa_tree_add_190_195_groupi_n_4638 ,csa_tree_add_190_195_groupi_n_3140 ,csa_tree_add_190_195_groupi_n_4158);
  and csa_tree_add_190_195_groupi_g44568(csa_tree_add_190_195_groupi_n_4635 ,csa_tree_add_190_195_groupi_n_3035 ,csa_tree_add_190_195_groupi_n_4157);
  or csa_tree_add_190_195_groupi_g44569(csa_tree_add_190_195_groupi_n_4633 ,csa_tree_add_190_195_groupi_n_3439 ,csa_tree_add_190_195_groupi_n_4156);
  or csa_tree_add_190_195_groupi_g44570(csa_tree_add_190_195_groupi_n_4632 ,csa_tree_add_190_195_groupi_n_3497 ,csa_tree_add_190_195_groupi_n_4551);
  or csa_tree_add_190_195_groupi_g44571(csa_tree_add_190_195_groupi_n_4630 ,csa_tree_add_190_195_groupi_n_2940 ,csa_tree_add_190_195_groupi_n_4512);
  and csa_tree_add_190_195_groupi_g44572(csa_tree_add_190_195_groupi_n_4628 ,csa_tree_add_190_195_groupi_n_3636 ,csa_tree_add_190_195_groupi_n_4159);
  and csa_tree_add_190_195_groupi_g44573(csa_tree_add_190_195_groupi_n_4627 ,csa_tree_add_190_195_groupi_n_2811 ,csa_tree_add_190_195_groupi_n_4254);
  and csa_tree_add_190_195_groupi_g44574(csa_tree_add_190_195_groupi_n_4625 ,csa_tree_add_190_195_groupi_n_2801 ,csa_tree_add_190_195_groupi_n_4545);
  or csa_tree_add_190_195_groupi_g44575(csa_tree_add_190_195_groupi_n_4623 ,csa_tree_add_190_195_groupi_n_3226 ,csa_tree_add_190_195_groupi_n_4483);
  or csa_tree_add_190_195_groupi_g44576(csa_tree_add_190_195_groupi_n_4621 ,csa_tree_add_190_195_groupi_n_3631 ,csa_tree_add_190_195_groupi_n_4283);
  or csa_tree_add_190_195_groupi_g44577(csa_tree_add_190_195_groupi_n_4619 ,csa_tree_add_190_195_groupi_n_3311 ,csa_tree_add_190_195_groupi_n_4153);
  or csa_tree_add_190_195_groupi_g44578(csa_tree_add_190_195_groupi_n_4618 ,csa_tree_add_190_195_groupi_n_3682 ,csa_tree_add_190_195_groupi_n_4166);
  and csa_tree_add_190_195_groupi_g44579(csa_tree_add_190_195_groupi_n_4617 ,csa_tree_add_190_195_groupi_n_3722 ,csa_tree_add_190_195_groupi_n_4351);
  or csa_tree_add_190_195_groupi_g44580(csa_tree_add_190_195_groupi_n_4616 ,csa_tree_add_190_195_groupi_n_3110 ,csa_tree_add_190_195_groupi_n_4226);
  or csa_tree_add_190_195_groupi_g44581(csa_tree_add_190_195_groupi_n_4615 ,csa_tree_add_190_195_groupi_n_3198 ,csa_tree_add_190_195_groupi_n_4444);
  and csa_tree_add_190_195_groupi_g44582(csa_tree_add_190_195_groupi_n_4613 ,csa_tree_add_190_195_groupi_n_3556 ,csa_tree_add_190_195_groupi_n_4212);
  and csa_tree_add_190_195_groupi_g44583(csa_tree_add_190_195_groupi_n_4612 ,csa_tree_add_190_195_groupi_n_2852 ,csa_tree_add_190_195_groupi_n_4265);
  or csa_tree_add_190_195_groupi_g44584(csa_tree_add_190_195_groupi_n_4611 ,csa_tree_add_190_195_groupi_n_3435 ,csa_tree_add_190_195_groupi_n_4376);
  or csa_tree_add_190_195_groupi_g44585(csa_tree_add_190_195_groupi_n_4609 ,csa_tree_add_190_195_groupi_n_3656 ,csa_tree_add_190_195_groupi_n_4450);
  or csa_tree_add_190_195_groupi_g44586(csa_tree_add_190_195_groupi_n_4606 ,csa_tree_add_190_195_groupi_n_2805 ,csa_tree_add_190_195_groupi_n_4292);
  or csa_tree_add_190_195_groupi_g44587(csa_tree_add_190_195_groupi_n_4604 ,csa_tree_add_190_195_groupi_n_2987 ,csa_tree_add_190_195_groupi_n_4147);
  or csa_tree_add_190_195_groupi_g44588(csa_tree_add_190_195_groupi_n_4603 ,csa_tree_add_190_195_groupi_n_3632 ,csa_tree_add_190_195_groupi_n_4453);
  or csa_tree_add_190_195_groupi_g44589(csa_tree_add_190_195_groupi_n_4600 ,csa_tree_add_190_195_groupi_n_3103 ,csa_tree_add_190_195_groupi_n_4146);
  and csa_tree_add_190_195_groupi_g44590(csa_tree_add_190_195_groupi_n_4599 ,csa_tree_add_190_195_groupi_n_3267 ,csa_tree_add_190_195_groupi_n_4340);
  or csa_tree_add_190_195_groupi_g44591(csa_tree_add_190_195_groupi_n_4597 ,csa_tree_add_190_195_groupi_n_3566 ,csa_tree_add_190_195_groupi_n_4307);
  or csa_tree_add_190_195_groupi_g44592(csa_tree_add_190_195_groupi_n_4595 ,csa_tree_add_190_195_groupi_n_3333 ,csa_tree_add_190_195_groupi_n_4163);
  or csa_tree_add_190_195_groupi_g44593(csa_tree_add_190_195_groupi_n_4593 ,csa_tree_add_190_195_groupi_n_3649 ,csa_tree_add_190_195_groupi_n_4471);
  or csa_tree_add_190_195_groupi_g44594(csa_tree_add_190_195_groupi_n_4591 ,csa_tree_add_190_195_groupi_n_3542 ,csa_tree_add_190_195_groupi_n_4271);
  and csa_tree_add_190_195_groupi_g44595(csa_tree_add_190_195_groupi_n_4590 ,csa_tree_add_190_195_groupi_n_3674 ,csa_tree_add_190_195_groupi_n_4479);
  and csa_tree_add_190_195_groupi_g44596(csa_tree_add_190_195_groupi_n_4588 ,csa_tree_add_190_195_groupi_n_3354 ,csa_tree_add_190_195_groupi_n_4401);
  or csa_tree_add_190_195_groupi_g44597(csa_tree_add_190_195_groupi_n_4586 ,csa_tree_add_190_195_groupi_n_62 ,csa_tree_add_190_195_groupi_n_4260);
  and csa_tree_add_190_195_groupi_g44598(csa_tree_add_190_195_groupi_n_4583 ,csa_tree_add_190_195_groupi_n_3009 ,csa_tree_add_190_195_groupi_n_4240);
  or csa_tree_add_190_195_groupi_g44599(csa_tree_add_190_195_groupi_n_4582 ,csa_tree_add_190_195_groupi_n_2829 ,csa_tree_add_190_195_groupi_n_4463);
  not csa_tree_add_190_195_groupi_g44600(csa_tree_add_190_195_groupi_n_4564 ,csa_tree_add_190_195_groupi_n_4565);
  not csa_tree_add_190_195_groupi_g44601(csa_tree_add_190_195_groupi_n_4562 ,csa_tree_add_190_195_groupi_n_4563);
  not csa_tree_add_190_195_groupi_g44602(csa_tree_add_190_195_groupi_n_4560 ,csa_tree_add_190_195_groupi_n_4561);
  and csa_tree_add_190_195_groupi_g44603(csa_tree_add_190_195_groupi_n_4559 ,csa_tree_add_190_195_groupi_n_1997 ,csa_tree_add_190_195_groupi_n_3462);
  and csa_tree_add_190_195_groupi_g44604(csa_tree_add_190_195_groupi_n_4558 ,csa_tree_add_190_195_groupi_n_1764 ,csa_tree_add_190_195_groupi_n_2874);
  and csa_tree_add_190_195_groupi_g44605(csa_tree_add_190_195_groupi_n_4557 ,csa_tree_add_190_195_groupi_n_1585 ,csa_tree_add_190_195_groupi_n_2826);
  or csa_tree_add_190_195_groupi_g44606(csa_tree_add_190_195_groupi_n_4556 ,csa_tree_add_190_195_groupi_n_1873 ,csa_tree_add_190_195_groupi_n_3188);
  and csa_tree_add_190_195_groupi_g44607(csa_tree_add_190_195_groupi_n_4555 ,in61[12] ,csa_tree_add_190_195_groupi_n_3069);
  and csa_tree_add_190_195_groupi_g44608(csa_tree_add_190_195_groupi_n_4554 ,csa_tree_add_190_195_groupi_n_1686 ,csa_tree_add_190_195_groupi_n_3242);
  or csa_tree_add_190_195_groupi_g44609(csa_tree_add_190_195_groupi_n_4553 ,csa_tree_add_190_195_groupi_n_1671 ,csa_tree_add_190_195_groupi_n_2809);
  and csa_tree_add_190_195_groupi_g44610(csa_tree_add_190_195_groupi_n_4552 ,csa_tree_add_190_195_groupi_n_2002 ,csa_tree_add_190_195_groupi_n_2739);
  and csa_tree_add_190_195_groupi_g44611(csa_tree_add_190_195_groupi_n_4551 ,csa_tree_add_190_195_groupi_n_1602 ,csa_tree_add_190_195_groupi_n_3509);
  or csa_tree_add_190_195_groupi_g44612(csa_tree_add_190_195_groupi_n_4550 ,csa_tree_add_190_195_groupi_n_2714 ,csa_tree_add_190_195_groupi_n_2911);
  and csa_tree_add_190_195_groupi_g44613(csa_tree_add_190_195_groupi_n_4549 ,in59[3] ,csa_tree_add_190_195_groupi_n_2772);
  and csa_tree_add_190_195_groupi_g44614(csa_tree_add_190_195_groupi_n_4548 ,csa_tree_add_190_195_groupi_n_1709 ,csa_tree_add_190_195_groupi_n_2933);
  and csa_tree_add_190_195_groupi_g44615(csa_tree_add_190_195_groupi_n_4547 ,csa_tree_add_190_195_groupi_n_1601 ,csa_tree_add_190_195_groupi_n_3124);
  and csa_tree_add_190_195_groupi_g44616(csa_tree_add_190_195_groupi_n_4546 ,csa_tree_add_190_195_groupi_n_1894 ,csa_tree_add_190_195_groupi_n_2734);
  or csa_tree_add_190_195_groupi_g44617(csa_tree_add_190_195_groupi_n_4545 ,csa_tree_add_190_195_groupi_n_1580 ,csa_tree_add_190_195_groupi_n_2749);
  and csa_tree_add_190_195_groupi_g44618(csa_tree_add_190_195_groupi_n_4544 ,csa_tree_add_190_195_groupi_n_1861 ,csa_tree_add_190_195_groupi_n_2877);
  and csa_tree_add_190_195_groupi_g44619(csa_tree_add_190_195_groupi_n_4543 ,in59[8] ,csa_tree_add_190_195_groupi_n_3102);
  and csa_tree_add_190_195_groupi_g44620(csa_tree_add_190_195_groupi_n_4542 ,csa_tree_add_190_195_groupi_n_1640 ,csa_tree_add_190_195_groupi_n_2857);
  or csa_tree_add_190_195_groupi_g44621(csa_tree_add_190_195_groupi_n_4541 ,csa_tree_add_190_195_groupi_n_1842 ,csa_tree_add_190_195_groupi_n_2931);
  and csa_tree_add_190_195_groupi_g44622(csa_tree_add_190_195_groupi_n_4540 ,csa_tree_add_190_195_groupi_n_1608 ,csa_tree_add_190_195_groupi_n_3620);
  and csa_tree_add_190_195_groupi_g44623(csa_tree_add_190_195_groupi_n_4539 ,csa_tree_add_190_195_groupi_n_1898 ,csa_tree_add_190_195_groupi_n_3097);
  and csa_tree_add_190_195_groupi_g44624(csa_tree_add_190_195_groupi_n_4538 ,csa_tree_add_190_195_groupi_n_1837 ,csa_tree_add_190_195_groupi_n_2947);
  or csa_tree_add_190_195_groupi_g44625(csa_tree_add_190_195_groupi_n_4537 ,csa_tree_add_190_195_groupi_n_2005 ,csa_tree_add_190_195_groupi_n_3105);
  and csa_tree_add_190_195_groupi_g44626(csa_tree_add_190_195_groupi_n_4536 ,csa_tree_add_190_195_groupi_n_1754 ,csa_tree_add_190_195_groupi_n_3114);
  and csa_tree_add_190_195_groupi_g44627(csa_tree_add_190_195_groupi_n_4535 ,csa_tree_add_190_195_groupi_n_1612 ,csa_tree_add_190_195_groupi_n_2840);
  or csa_tree_add_190_195_groupi_g44628(csa_tree_add_190_195_groupi_n_4534 ,csa_tree_add_190_195_groupi_n_1701 ,csa_tree_add_190_195_groupi_n_3240);
  and csa_tree_add_190_195_groupi_g44629(csa_tree_add_190_195_groupi_n_4533 ,csa_tree_add_190_195_groupi_n_1916 ,csa_tree_add_190_195_groupi_n_2892);
  or csa_tree_add_190_195_groupi_g44630(csa_tree_add_190_195_groupi_n_4532 ,csa_tree_add_190_195_groupi_n_2544 ,csa_tree_add_190_195_groupi_n_2746);
  and csa_tree_add_190_195_groupi_g44631(csa_tree_add_190_195_groupi_n_4531 ,csa_tree_add_190_195_groupi_n_1709 ,csa_tree_add_190_195_groupi_n_3022);
  and csa_tree_add_190_195_groupi_g44632(csa_tree_add_190_195_groupi_n_4530 ,in58[3] ,csa_tree_add_190_195_groupi_n_2777);
  and csa_tree_add_190_195_groupi_g44633(csa_tree_add_190_195_groupi_n_4529 ,csa_tree_add_190_195_groupi_n_2004 ,csa_tree_add_190_195_groupi_n_2961);
  and csa_tree_add_190_195_groupi_g44634(csa_tree_add_190_195_groupi_n_4528 ,csa_tree_add_190_195_groupi_n_1759 ,csa_tree_add_190_195_groupi_n_2996);
  and csa_tree_add_190_195_groupi_g44635(csa_tree_add_190_195_groupi_n_4527 ,csa_tree_add_190_195_groupi_n_1756 ,csa_tree_add_190_195_groupi_n_2966);
  and csa_tree_add_190_195_groupi_g44636(csa_tree_add_190_195_groupi_n_4526 ,csa_tree_add_190_195_groupi_n_1852 ,csa_tree_add_190_195_groupi_n_2983);
  or csa_tree_add_190_195_groupi_g44637(csa_tree_add_190_195_groupi_n_4525 ,csa_tree_add_190_195_groupi_n_1900 ,csa_tree_add_190_195_groupi_n_3505);
  and csa_tree_add_190_195_groupi_g44638(csa_tree_add_190_195_groupi_n_4524 ,csa_tree_add_190_195_groupi_n_1690 ,csa_tree_add_190_195_groupi_n_2793);
  and csa_tree_add_190_195_groupi_g44639(csa_tree_add_190_195_groupi_n_4523 ,csa_tree_add_190_195_groupi_n_1696 ,csa_tree_add_190_195_groupi_n_3619);
  and csa_tree_add_190_195_groupi_g44640(csa_tree_add_190_195_groupi_n_4522 ,csa_tree_add_190_195_groupi_n_1896 ,csa_tree_add_190_195_groupi_n_2847);
  or csa_tree_add_190_195_groupi_g44641(csa_tree_add_190_195_groupi_n_4521 ,csa_tree_add_190_195_groupi_n_1899 ,csa_tree_add_190_195_groupi_n_2802);
  and csa_tree_add_190_195_groupi_g44642(csa_tree_add_190_195_groupi_n_4520 ,in58[2] ,csa_tree_add_190_195_groupi_n_2885);
  and csa_tree_add_190_195_groupi_g44643(csa_tree_add_190_195_groupi_n_4519 ,csa_tree_add_190_195_groupi_n_1646 ,csa_tree_add_190_195_groupi_n_3087);
  or csa_tree_add_190_195_groupi_g44644(csa_tree_add_190_195_groupi_n_4518 ,csa_tree_add_190_195_groupi_n_1747 ,csa_tree_add_190_195_groupi_n_2920);
  and csa_tree_add_190_195_groupi_g44645(csa_tree_add_190_195_groupi_n_4517 ,csa_tree_add_190_195_groupi_n_1653 ,csa_tree_add_190_195_groupi_n_3493);
  and csa_tree_add_190_195_groupi_g44646(csa_tree_add_190_195_groupi_n_4516 ,csa_tree_add_190_195_groupi_n_1749 ,csa_tree_add_190_195_groupi_n_3043);
  or csa_tree_add_190_195_groupi_g44647(csa_tree_add_190_195_groupi_n_4515 ,csa_tree_add_190_195_groupi_n_1842 ,csa_tree_add_190_195_groupi_n_2985);
  and csa_tree_add_190_195_groupi_g44648(csa_tree_add_190_195_groupi_n_4514 ,csa_tree_add_190_195_groupi_n_1647 ,csa_tree_add_190_195_groupi_n_2846);
  and csa_tree_add_190_195_groupi_g44649(csa_tree_add_190_195_groupi_n_4513 ,csa_tree_add_190_195_groupi_n_1589 ,csa_tree_add_190_195_groupi_n_2796);
  and csa_tree_add_190_195_groupi_g44650(csa_tree_add_190_195_groupi_n_4512 ,in59[6] ,csa_tree_add_190_195_groupi_n_2875);
  and csa_tree_add_190_195_groupi_g44651(csa_tree_add_190_195_groupi_n_4511 ,csa_tree_add_190_195_groupi_n_1752 ,csa_tree_add_190_195_groupi_n_3246);
  or csa_tree_add_190_195_groupi_g44652(csa_tree_add_190_195_groupi_n_4510 ,csa_tree_add_190_195_groupi_n_1710 ,csa_tree_add_190_195_groupi_n_2868);
  and csa_tree_add_190_195_groupi_g44653(csa_tree_add_190_195_groupi_n_4509 ,csa_tree_add_190_195_groupi_n_1611 ,csa_tree_add_190_195_groupi_n_3084);
  or csa_tree_add_190_195_groupi_g44654(csa_tree_add_190_195_groupi_n_4508 ,csa_tree_add_190_195_groupi_n_2695 ,csa_tree_add_190_195_groupi_n_2804);
  and csa_tree_add_190_195_groupi_g44655(csa_tree_add_190_195_groupi_n_4507 ,csa_tree_add_190_195_groupi_n_1851 ,csa_tree_add_190_195_groupi_n_3039);
  and csa_tree_add_190_195_groupi_g44656(csa_tree_add_190_195_groupi_n_4506 ,in58[4] ,csa_tree_add_190_195_groupi_n_2898);
  and csa_tree_add_190_195_groupi_g44657(csa_tree_add_190_195_groupi_n_4505 ,csa_tree_add_190_195_groupi_n_1765 ,csa_tree_add_190_195_groupi_n_2783);
  or csa_tree_add_190_195_groupi_g44658(csa_tree_add_190_195_groupi_n_4504 ,csa_tree_add_190_195_groupi_n_2538 ,csa_tree_add_190_195_groupi_n_3225);
  and csa_tree_add_190_195_groupi_g44659(csa_tree_add_190_195_groupi_n_4503 ,csa_tree_add_190_195_groupi_n_1756 ,csa_tree_add_190_195_groupi_n_3223);
  and csa_tree_add_190_195_groupi_g44660(csa_tree_add_190_195_groupi_n_4502 ,csa_tree_add_190_195_groupi_n_1621 ,csa_tree_add_190_195_groupi_n_2745);
  or csa_tree_add_190_195_groupi_g44661(csa_tree_add_190_195_groupi_n_4501 ,csa_tree_add_190_195_groupi_n_1762 ,csa_tree_add_190_195_groupi_n_3008);
  and csa_tree_add_190_195_groupi_g44662(csa_tree_add_190_195_groupi_n_4500 ,in59[11] ,csa_tree_add_190_195_groupi_n_2884);
  and csa_tree_add_190_195_groupi_g44663(csa_tree_add_190_195_groupi_n_4499 ,csa_tree_add_190_195_groupi_n_1752 ,csa_tree_add_190_195_groupi_n_2848);
  or csa_tree_add_190_195_groupi_g44664(csa_tree_add_190_195_groupi_n_4498 ,csa_tree_add_190_195_groupi_n_2388 ,csa_tree_add_190_195_groupi_n_2944);
  and csa_tree_add_190_195_groupi_g44665(csa_tree_add_190_195_groupi_n_4497 ,csa_tree_add_190_195_groupi_n_1895 ,csa_tree_add_190_195_groupi_n_3033);
  and csa_tree_add_190_195_groupi_g44666(csa_tree_add_190_195_groupi_n_4496 ,in59[14] ,csa_tree_add_190_195_groupi_n_3484);
  or csa_tree_add_190_195_groupi_g44667(csa_tree_add_190_195_groupi_n_4495 ,csa_tree_add_190_195_groupi_n_1623 ,csa_tree_add_190_195_groupi_n_2957);
  or csa_tree_add_190_195_groupi_g44668(csa_tree_add_190_195_groupi_n_4494 ,csa_tree_add_190_195_groupi_n_1689 ,csa_tree_add_190_195_groupi_n_2976);
  and csa_tree_add_190_195_groupi_g44669(csa_tree_add_190_195_groupi_n_4493 ,csa_tree_add_190_195_groupi_n_1698 ,csa_tree_add_190_195_groupi_n_3504);
  or csa_tree_add_190_195_groupi_g44670(csa_tree_add_190_195_groupi_n_4492 ,csa_tree_add_190_195_groupi_n_2730 ,csa_tree_add_190_195_groupi_n_2799);
  and csa_tree_add_190_195_groupi_g44671(csa_tree_add_190_195_groupi_n_4491 ,csa_tree_add_190_195_groupi_n_1649 ,csa_tree_add_190_195_groupi_n_2856);
  and csa_tree_add_190_195_groupi_g44672(csa_tree_add_190_195_groupi_n_4490 ,csa_tree_add_190_195_groupi_n_1697 ,csa_tree_add_190_195_groupi_n_3134);
  or csa_tree_add_190_195_groupi_g44673(csa_tree_add_190_195_groupi_n_4489 ,csa_tree_add_190_195_groupi_n_1746 ,csa_tree_add_190_195_groupi_n_3653);
  and csa_tree_add_190_195_groupi_g44674(csa_tree_add_190_195_groupi_n_4488 ,csa_tree_add_190_195_groupi_n_1630 ,csa_tree_add_190_195_groupi_n_3162);
  and csa_tree_add_190_195_groupi_g44675(csa_tree_add_190_195_groupi_n_4487 ,csa_tree_add_190_195_groupi_n_1896 ,csa_tree_add_190_195_groupi_n_3101);
  and csa_tree_add_190_195_groupi_g44676(csa_tree_add_190_195_groupi_n_4486 ,csa_tree_add_190_195_groupi_n_1943 ,csa_tree_add_190_195_groupi_n_3137);
  and csa_tree_add_190_195_groupi_g44677(csa_tree_add_190_195_groupi_n_4485 ,csa_tree_add_190_195_groupi_n_1871 ,csa_tree_add_190_195_groupi_n_2860);
  or csa_tree_add_190_195_groupi_g44678(csa_tree_add_190_195_groupi_n_4484 ,csa_tree_add_190_195_groupi_n_2565 ,csa_tree_add_190_195_groupi_n_2867);
  and csa_tree_add_190_195_groupi_g44679(csa_tree_add_190_195_groupi_n_4483 ,csa_tree_add_190_195_groupi_n_1692 ,csa_tree_add_190_195_groupi_n_3212);
  and csa_tree_add_190_195_groupi_g44680(csa_tree_add_190_195_groupi_n_4482 ,csa_tree_add_190_195_groupi_n_1854 ,csa_tree_add_190_195_groupi_n_3158);
  and csa_tree_add_190_195_groupi_g44681(csa_tree_add_190_195_groupi_n_4481 ,csa_tree_add_190_195_groupi_n_1710 ,csa_tree_add_190_195_groupi_n_2956);
  and csa_tree_add_190_195_groupi_g44682(csa_tree_add_190_195_groupi_n_4480 ,csa_tree_add_190_195_groupi_n_1859 ,csa_tree_add_190_195_groupi_n_3261);
  or csa_tree_add_190_195_groupi_g44683(csa_tree_add_190_195_groupi_n_4479 ,csa_tree_add_190_195_groupi_n_1608 ,csa_tree_add_190_195_groupi_n_3675);
  or csa_tree_add_190_195_groupi_g44684(csa_tree_add_190_195_groupi_n_4478 ,csa_tree_add_190_195_groupi_n_1972 ,csa_tree_add_190_195_groupi_n_3490);
  or csa_tree_add_190_195_groupi_g44685(csa_tree_add_190_195_groupi_n_4477 ,csa_tree_add_190_195_groupi_n_1825 ,csa_tree_add_190_195_groupi_n_3030);
  or csa_tree_add_190_195_groupi_g44686(csa_tree_add_190_195_groupi_n_4476 ,csa_tree_add_190_195_groupi_n_1990 ,csa_tree_add_190_195_groupi_n_3255);
  nor csa_tree_add_190_195_groupi_g44687(csa_tree_add_190_195_groupi_n_4475 ,csa_tree_add_190_195_groupi_n_2678 ,csa_tree_add_190_195_groupi_n_2836);
  nor csa_tree_add_190_195_groupi_g44688(csa_tree_add_190_195_groupi_n_4474 ,csa_tree_add_190_195_groupi_n_2515 ,csa_tree_add_190_195_groupi_n_3146);
  and csa_tree_add_190_195_groupi_g44689(csa_tree_add_190_195_groupi_n_4473 ,csa_tree_add_190_195_groupi_n_1899 ,csa_tree_add_190_195_groupi_n_3604);
  or csa_tree_add_190_195_groupi_g44690(csa_tree_add_190_195_groupi_n_4472 ,csa_tree_add_190_195_groupi_n_1543 ,csa_tree_add_190_195_groupi_n_3480);
  and csa_tree_add_190_195_groupi_g44691(csa_tree_add_190_195_groupi_n_4471 ,csa_tree_add_190_195_groupi_n_1776 ,csa_tree_add_190_195_groupi_n_3648);
  and csa_tree_add_190_195_groupi_g44692(csa_tree_add_190_195_groupi_n_4470 ,csa_tree_add_190_195_groupi_n_1662 ,csa_tree_add_190_195_groupi_n_3635);
  and csa_tree_add_190_195_groupi_g44693(csa_tree_add_190_195_groupi_n_4469 ,csa_tree_add_190_195_groupi_n_1852 ,csa_tree_add_190_195_groupi_n_3662);
  and csa_tree_add_190_195_groupi_g44694(csa_tree_add_190_195_groupi_n_4468 ,csa_tree_add_190_195_groupi_n_1618 ,csa_tree_add_190_195_groupi_n_3628);
  or csa_tree_add_190_195_groupi_g44695(csa_tree_add_190_195_groupi_n_4467 ,csa_tree_add_190_195_groupi_n_1964 ,csa_tree_add_190_195_groupi_n_3486);
  nor csa_tree_add_190_195_groupi_g44696(csa_tree_add_190_195_groupi_n_4466 ,csa_tree_add_190_195_groupi_n_2666 ,csa_tree_add_190_195_groupi_n_3217);
  nor csa_tree_add_190_195_groupi_g44697(csa_tree_add_190_195_groupi_n_4465 ,csa_tree_add_190_195_groupi_n_2668 ,csa_tree_add_190_195_groupi_n_3015);
  or csa_tree_add_190_195_groupi_g44698(csa_tree_add_190_195_groupi_n_4464 ,csa_tree_add_190_195_groupi_n_2672 ,csa_tree_add_190_195_groupi_n_3196);
  nor csa_tree_add_190_195_groupi_g44699(csa_tree_add_190_195_groupi_n_4463 ,csa_tree_add_190_195_groupi_n_2344 ,csa_tree_add_190_195_groupi_n_3063);
  nor csa_tree_add_190_195_groupi_g44700(csa_tree_add_190_195_groupi_n_4462 ,csa_tree_add_190_195_groupi_n_2675 ,csa_tree_add_190_195_groupi_n_3018);
  nor csa_tree_add_190_195_groupi_g44701(csa_tree_add_190_195_groupi_n_4461 ,csa_tree_add_190_195_groupi_n_2665 ,csa_tree_add_190_195_groupi_n_3144);
  nor csa_tree_add_190_195_groupi_g44702(csa_tree_add_190_195_groupi_n_4460 ,csa_tree_add_190_195_groupi_n_2667 ,csa_tree_add_190_195_groupi_n_2995);
  or csa_tree_add_190_195_groupi_g44703(csa_tree_add_190_195_groupi_n_4459 ,csa_tree_add_190_195_groupi_n_2157 ,csa_tree_add_190_195_groupi_n_3014);
  or csa_tree_add_190_195_groupi_g44704(csa_tree_add_190_195_groupi_n_4458 ,csa_tree_add_190_195_groupi_n_2669 ,csa_tree_add_190_195_groupi_n_51);
  or csa_tree_add_190_195_groupi_g44705(csa_tree_add_190_195_groupi_n_4457 ,csa_tree_add_190_195_groupi_n_2661 ,csa_tree_add_190_195_groupi_n_3111);
  or csa_tree_add_190_195_groupi_g44706(csa_tree_add_190_195_groupi_n_4456 ,csa_tree_add_190_195_groupi_n_2662 ,csa_tree_add_190_195_groupi_n_2859);
  nor csa_tree_add_190_195_groupi_g44707(csa_tree_add_190_195_groupi_n_4455 ,csa_tree_add_190_195_groupi_n_2673 ,csa_tree_add_190_195_groupi_n_2851);
  or csa_tree_add_190_195_groupi_g44708(csa_tree_add_190_195_groupi_n_4454 ,csa_tree_add_190_195_groupi_n_1851 ,csa_tree_add_190_195_groupi_n_3476);
  and csa_tree_add_190_195_groupi_g44709(csa_tree_add_190_195_groupi_n_4453 ,csa_tree_add_190_195_groupi_n_1627 ,csa_tree_add_190_195_groupi_n_3650);
  and csa_tree_add_190_195_groupi_g44710(csa_tree_add_190_195_groupi_n_4452 ,csa_tree_add_190_195_groupi_n_2001 ,csa_tree_add_190_195_groupi_n_3640);
  and csa_tree_add_190_195_groupi_g44711(csa_tree_add_190_195_groupi_n_4451 ,csa_tree_add_190_195_groupi_n_1697 ,csa_tree_add_190_195_groupi_n_3661);
  and csa_tree_add_190_195_groupi_g44712(csa_tree_add_190_195_groupi_n_4450 ,csa_tree_add_190_195_groupi_n_1853 ,csa_tree_add_190_195_groupi_n_3657);
  and csa_tree_add_190_195_groupi_g44713(csa_tree_add_190_195_groupi_n_4449 ,csa_tree_add_190_195_groupi_n_1742 ,csa_tree_add_190_195_groupi_n_3658);
  or csa_tree_add_190_195_groupi_g44714(csa_tree_add_190_195_groupi_n_4448 ,csa_tree_add_190_195_groupi_n_1998 ,csa_tree_add_190_195_groupi_n_3413);
  nor csa_tree_add_190_195_groupi_g44715(csa_tree_add_190_195_groupi_n_4447 ,csa_tree_add_190_195_groupi_n_2634 ,csa_tree_add_190_195_groupi_n_3057);
  nor csa_tree_add_190_195_groupi_g44716(csa_tree_add_190_195_groupi_n_4446 ,csa_tree_add_190_195_groupi_n_1535 ,csa_tree_add_190_195_groupi_n_3217);
  or csa_tree_add_190_195_groupi_g44717(csa_tree_add_190_195_groupi_n_4445 ,csa_tree_add_190_195_groupi_n_2042 ,csa_tree_add_190_195_groupi_n_3447);
  nor csa_tree_add_190_195_groupi_g44718(csa_tree_add_190_195_groupi_n_4444 ,csa_tree_add_190_195_groupi_n_2640 ,csa_tree_add_190_195_groupi_n_2743);
  nor csa_tree_add_190_195_groupi_g44719(csa_tree_add_190_195_groupi_n_4443 ,csa_tree_add_190_195_groupi_n_2485 ,csa_tree_add_190_195_groupi_n_2822);
  or csa_tree_add_190_195_groupi_g44720(csa_tree_add_190_195_groupi_n_4442 ,csa_tree_add_190_195_groupi_n_882 ,csa_tree_add_190_195_groupi_n_3726);
  or csa_tree_add_190_195_groupi_g44721(csa_tree_add_190_195_groupi_n_4441 ,csa_tree_add_190_195_groupi_n_1974 ,csa_tree_add_190_195_groupi_n_2828);
  nor csa_tree_add_190_195_groupi_g44722(csa_tree_add_190_195_groupi_n_4440 ,csa_tree_add_190_195_groupi_n_2650 ,csa_tree_add_190_195_groupi_n_2910);
  nor csa_tree_add_190_195_groupi_g44723(csa_tree_add_190_195_groupi_n_4439 ,csa_tree_add_190_195_groupi_n_1566 ,csa_tree_add_190_195_groupi_n_2990);
  nor csa_tree_add_190_195_groupi_g44724(csa_tree_add_190_195_groupi_n_4438 ,csa_tree_add_190_195_groupi_n_2488 ,csa_tree_add_190_195_groupi_n_3032);
  nor csa_tree_add_190_195_groupi_g44725(csa_tree_add_190_195_groupi_n_4437 ,csa_tree_add_190_195_groupi_n_2647 ,csa_tree_add_190_195_groupi_n_3239);
  nor csa_tree_add_190_195_groupi_g44726(csa_tree_add_190_195_groupi_n_4436 ,csa_tree_add_190_195_groupi_n_2492 ,csa_tree_add_190_195_groupi_n_3028);
  nor csa_tree_add_190_195_groupi_g44727(csa_tree_add_190_195_groupi_n_4435 ,csa_tree_add_190_195_groupi_n_2653 ,csa_tree_add_190_195_groupi_n_3053);
  nor csa_tree_add_190_195_groupi_g44728(csa_tree_add_190_195_groupi_n_4434 ,csa_tree_add_190_195_groupi_n_2643 ,csa_tree_add_190_195_groupi_n_2912);
  or csa_tree_add_190_195_groupi_g44729(csa_tree_add_190_195_groupi_n_4433 ,csa_tree_add_190_195_groupi_n_2646 ,csa_tree_add_190_195_groupi_n_3076);
  nor csa_tree_add_190_195_groupi_g44730(csa_tree_add_190_195_groupi_n_4432 ,csa_tree_add_190_195_groupi_n_2645 ,csa_tree_add_190_195_groupi_n_2967);
  or csa_tree_add_190_195_groupi_g44731(csa_tree_add_190_195_groupi_n_4431 ,csa_tree_add_190_195_groupi_n_2118 ,csa_tree_add_190_195_groupi_n_3717);
  nor csa_tree_add_190_195_groupi_g44732(csa_tree_add_190_195_groupi_n_4430 ,csa_tree_add_190_195_groupi_n_2652 ,csa_tree_add_190_195_groupi_n_2903);
  nor csa_tree_add_190_195_groupi_g44733(csa_tree_add_190_195_groupi_n_4429 ,csa_tree_add_190_195_groupi_n_2639 ,csa_tree_add_190_195_groupi_n_3236);
  or csa_tree_add_190_195_groupi_g44734(csa_tree_add_190_195_groupi_n_4428 ,csa_tree_add_190_195_groupi_n_1775 ,csa_tree_add_190_195_groupi_n_3707);
  or csa_tree_add_190_195_groupi_g44735(csa_tree_add_190_195_groupi_n_4427 ,csa_tree_add_190_195_groupi_n_2216 ,csa_tree_add_190_195_groupi_n_3500);
  nor csa_tree_add_190_195_groupi_g44736(csa_tree_add_190_195_groupi_n_4426 ,csa_tree_add_190_195_groupi_n_2659 ,csa_tree_add_190_195_groupi_n_3668);
  nor csa_tree_add_190_195_groupi_g44737(csa_tree_add_190_195_groupi_n_4425 ,csa_tree_add_190_195_groupi_n_2656 ,csa_tree_add_190_195_groupi_n_2959);
  or csa_tree_add_190_195_groupi_g44738(csa_tree_add_190_195_groupi_n_4424 ,csa_tree_add_190_195_groupi_n_982 ,csa_tree_add_190_195_groupi_n_3491);
  or csa_tree_add_190_195_groupi_g44739(csa_tree_add_190_195_groupi_n_4423 ,csa_tree_add_190_195_groupi_n_1353 ,csa_tree_add_190_195_groupi_n_2759);
  nor csa_tree_add_190_195_groupi_g44740(csa_tree_add_190_195_groupi_n_4422 ,csa_tree_add_190_195_groupi_n_2483 ,csa_tree_add_190_195_groupi_n_3133);
  nor csa_tree_add_190_195_groupi_g44741(csa_tree_add_190_195_groupi_n_4421 ,csa_tree_add_190_195_groupi_n_2493 ,csa_tree_add_190_195_groupi_n_2763);
  or csa_tree_add_190_195_groupi_g44742(csa_tree_add_190_195_groupi_n_4420 ,csa_tree_add_190_195_groupi_n_1174 ,csa_tree_add_190_195_groupi_n_2964);
  or csa_tree_add_190_195_groupi_g44743(csa_tree_add_190_195_groupi_n_4419 ,csa_tree_add_190_195_groupi_n_2657 ,csa_tree_add_190_195_groupi_n_3003);
  nor csa_tree_add_190_195_groupi_g44744(csa_tree_add_190_195_groupi_n_4418 ,csa_tree_add_190_195_groupi_n_2649 ,csa_tree_add_190_195_groupi_n_3676);
  nor csa_tree_add_190_195_groupi_g44745(csa_tree_add_190_195_groupi_n_4417 ,csa_tree_add_190_195_groupi_n_2494 ,csa_tree_add_190_195_groupi_n_3098);
  nor csa_tree_add_190_195_groupi_g44746(csa_tree_add_190_195_groupi_n_4416 ,csa_tree_add_190_195_groupi_n_2495 ,csa_tree_add_190_195_groupi_n_2831);
  or csa_tree_add_190_195_groupi_g44747(csa_tree_add_190_195_groupi_n_4415 ,in56[1] ,csa_tree_add_190_195_groupi_n_3602);
  and csa_tree_add_190_195_groupi_g44748(csa_tree_add_190_195_groupi_n_4414 ,csa_tree_add_190_195_groupi_n_1626 ,csa_tree_add_190_195_groupi_n_3596);
  or csa_tree_add_190_195_groupi_g44749(csa_tree_add_190_195_groupi_n_4413 ,csa_tree_add_190_195_groupi_n_1819 ,csa_tree_add_190_195_groupi_n_3603);
  and csa_tree_add_190_195_groupi_g44750(csa_tree_add_190_195_groupi_n_4412 ,csa_tree_add_190_195_groupi_n_1705 ,csa_tree_add_190_195_groupi_n_3572);
  or csa_tree_add_190_195_groupi_g44751(csa_tree_add_190_195_groupi_n_4411 ,csa_tree_add_190_195_groupi_n_1834 ,csa_tree_add_190_195_groupi_n_3573);
  and csa_tree_add_190_195_groupi_g44752(csa_tree_add_190_195_groupi_n_4410 ,csa_tree_add_190_195_groupi_n_1900 ,csa_tree_add_190_195_groupi_n_3605);
  and csa_tree_add_190_195_groupi_g44753(csa_tree_add_190_195_groupi_n_4409 ,csa_tree_add_190_195_groupi_n_1887 ,csa_tree_add_190_195_groupi_n_3524);
  and csa_tree_add_190_195_groupi_g44754(csa_tree_add_190_195_groupi_n_4408 ,csa_tree_add_190_195_groupi_n_1661 ,csa_tree_add_190_195_groupi_n_3579);
  and csa_tree_add_190_195_groupi_g44755(csa_tree_add_190_195_groupi_n_4407 ,csa_tree_add_190_195_groupi_n_1894 ,csa_tree_add_190_195_groupi_n_3560);
  or csa_tree_add_190_195_groupi_g44756(csa_tree_add_190_195_groupi_n_4406 ,csa_tree_add_190_195_groupi_n_2215 ,csa_tree_add_190_195_groupi_n_3595);
  or csa_tree_add_190_195_groupi_g44757(csa_tree_add_190_195_groupi_n_4405 ,csa_tree_add_190_195_groupi_n_1659 ,csa_tree_add_190_195_groupi_n_3383);
  or csa_tree_add_190_195_groupi_g44758(csa_tree_add_190_195_groupi_n_4404 ,csa_tree_add_190_195_groupi_n_1892 ,csa_tree_add_190_195_groupi_n_3330);
  or csa_tree_add_190_195_groupi_g44759(csa_tree_add_190_195_groupi_n_4403 ,csa_tree_add_190_195_groupi_n_2058 ,csa_tree_add_190_195_groupi_n_3346);
  or csa_tree_add_190_195_groupi_g44760(csa_tree_add_190_195_groupi_n_4402 ,csa_tree_add_190_195_groupi_n_1987 ,csa_tree_add_190_195_groupi_n_3397);
  or csa_tree_add_190_195_groupi_g44761(csa_tree_add_190_195_groupi_n_4401 ,csa_tree_add_190_195_groupi_n_760 ,csa_tree_add_190_195_groupi_n_3317);
  or csa_tree_add_190_195_groupi_g44762(csa_tree_add_190_195_groupi_n_4400 ,csa_tree_add_190_195_groupi_n_1009 ,csa_tree_add_190_195_groupi_n_3335);
  or csa_tree_add_190_195_groupi_g44763(csa_tree_add_190_195_groupi_n_4399 ,csa_tree_add_190_195_groupi_n_1994 ,csa_tree_add_190_195_groupi_n_3382);
  or csa_tree_add_190_195_groupi_g44764(csa_tree_add_190_195_groupi_n_4398 ,csa_tree_add_190_195_groupi_n_1767 ,csa_tree_add_190_195_groupi_n_3344);
  or csa_tree_add_190_195_groupi_g44765(csa_tree_add_190_195_groupi_n_4397 ,csa_tree_add_190_195_groupi_n_1993 ,csa_tree_add_190_195_groupi_n_3348);
  and csa_tree_add_190_195_groupi_g44766(csa_tree_add_190_195_groupi_n_4396 ,csa_tree_add_190_195_groupi_n_1643 ,csa_tree_add_190_195_groupi_n_3370);
  and csa_tree_add_190_195_groupi_g44767(csa_tree_add_190_195_groupi_n_4395 ,csa_tree_add_190_195_groupi_n_2473 ,csa_tree_add_190_195_groupi_n_1348);
  or csa_tree_add_190_195_groupi_g44768(csa_tree_add_190_195_groupi_n_4394 ,csa_tree_add_190_195_groupi_n_1528 ,csa_tree_add_190_195_groupi_n_3201);
  or csa_tree_add_190_195_groupi_g44769(csa_tree_add_190_195_groupi_n_4393 ,csa_tree_add_190_195_groupi_n_1988 ,csa_tree_add_190_195_groupi_n_3200);
  nor csa_tree_add_190_195_groupi_g44770(csa_tree_add_190_195_groupi_n_4392 ,csa_tree_add_190_195_groupi_n_2460 ,csa_tree_add_190_195_groupi_n_1329);
  and csa_tree_add_190_195_groupi_g44771(csa_tree_add_190_195_groupi_n_4391 ,csa_tree_add_190_195_groupi_n_2087 ,csa_tree_add_190_195_groupi_n_3482);
  and csa_tree_add_190_195_groupi_g44772(csa_tree_add_190_195_groupi_n_4390 ,csa_tree_add_190_195_groupi_n_1942 ,csa_tree_add_190_195_groupi_n_3464);
  or csa_tree_add_190_195_groupi_g44773(csa_tree_add_190_195_groupi_n_4389 ,csa_tree_add_190_195_groupi_n_1905 ,csa_tree_add_190_195_groupi_n_3341);
  or csa_tree_add_190_195_groupi_g44774(csa_tree_add_190_195_groupi_n_4388 ,csa_tree_add_190_195_groupi_n_2006 ,csa_tree_add_190_195_groupi_n_3352);
  or csa_tree_add_190_195_groupi_g44775(csa_tree_add_190_195_groupi_n_4387 ,csa_tree_add_190_195_groupi_n_1856 ,csa_tree_add_190_195_groupi_n_3384);
  or csa_tree_add_190_195_groupi_g44776(csa_tree_add_190_195_groupi_n_4386 ,csa_tree_add_190_195_groupi_n_2119 ,csa_tree_add_190_195_groupi_n_3555);
  or csa_tree_add_190_195_groupi_g44777(csa_tree_add_190_195_groupi_n_4385 ,csa_tree_add_190_195_groupi_n_2713 ,csa_tree_add_190_195_groupi_n_3714);
  and csa_tree_add_190_195_groupi_g44778(csa_tree_add_190_195_groupi_n_4384 ,csa_tree_add_190_195_groupi_n_1767 ,csa_tree_add_190_195_groupi_n_3520);
  and csa_tree_add_190_195_groupi_g44779(csa_tree_add_190_195_groupi_n_4383 ,csa_tree_add_190_195_groupi_n_1650 ,csa_tree_add_190_195_groupi_n_3608);
  and csa_tree_add_190_195_groupi_g44780(csa_tree_add_190_195_groupi_n_4382 ,in61[0] ,csa_tree_add_190_195_groupi_n_3553);
  or csa_tree_add_190_195_groupi_g44781(csa_tree_add_190_195_groupi_n_4381 ,csa_tree_add_190_195_groupi_n_1822 ,csa_tree_add_190_195_groupi_n_3577);
  and csa_tree_add_190_195_groupi_g44782(csa_tree_add_190_195_groupi_n_4380 ,csa_tree_add_190_195_groupi_n_2058 ,csa_tree_add_190_195_groupi_n_3373);
  or csa_tree_add_190_195_groupi_g44783(csa_tree_add_190_195_groupi_n_4379 ,csa_tree_add_190_195_groupi_n_1462 ,csa_tree_add_190_195_groupi_n_2879);
  nor csa_tree_add_190_195_groupi_g44784(csa_tree_add_190_195_groupi_n_4378 ,csa_tree_add_190_195_groupi_n_2601 ,csa_tree_add_190_195_groupi_n_3225);
  nor csa_tree_add_190_195_groupi_g44785(csa_tree_add_190_195_groupi_n_4377 ,csa_tree_add_190_195_groupi_n_2601 ,csa_tree_add_190_195_groupi_n_3060);
  and csa_tree_add_190_195_groupi_g44786(csa_tree_add_190_195_groupi_n_4376 ,csa_tree_add_190_195_groupi_n_1008 ,csa_tree_add_190_195_groupi_n_3434);
  and csa_tree_add_190_195_groupi_g44787(csa_tree_add_190_195_groupi_n_4375 ,csa_tree_add_190_195_groupi_n_1901 ,csa_tree_add_190_195_groupi_n_3332);
  and csa_tree_add_190_195_groupi_g44788(csa_tree_add_190_195_groupi_n_4374 ,csa_tree_add_190_195_groupi_n_1696 ,csa_tree_add_190_195_groupi_n_3552);
  or csa_tree_add_190_195_groupi_g44789(csa_tree_add_190_195_groupi_n_4373 ,csa_tree_add_190_195_groupi_n_1753 ,csa_tree_add_190_195_groupi_n_3589);
  or csa_tree_add_190_195_groupi_g44790(csa_tree_add_190_195_groupi_n_4372 ,csa_tree_add_190_195_groupi_n_1910 ,csa_tree_add_190_195_groupi_n_3592);
  or csa_tree_add_190_195_groupi_g44791(csa_tree_add_190_195_groupi_n_4371 ,csa_tree_add_190_195_groupi_n_1814 ,csa_tree_add_190_195_groupi_n_3547);
  or csa_tree_add_190_195_groupi_g44792(csa_tree_add_190_195_groupi_n_4370 ,csa_tree_add_190_195_groupi_n_1743 ,csa_tree_add_190_195_groupi_n_3281);
  nor csa_tree_add_190_195_groupi_g44793(csa_tree_add_190_195_groupi_n_4369 ,csa_tree_add_190_195_groupi_n_3163 ,csa_tree_add_190_195_groupi_n_2594);
  nor csa_tree_add_190_195_groupi_g44794(csa_tree_add_190_195_groupi_n_4368 ,csa_tree_add_190_195_groupi_n_2984 ,csa_tree_add_190_195_groupi_n_2432);
  nor csa_tree_add_190_195_groupi_g44795(csa_tree_add_190_195_groupi_n_4367 ,csa_tree_add_190_195_groupi_n_1469 ,csa_tree_add_190_195_groupi_n_3046);
  nor csa_tree_add_190_195_groupi_g44796(csa_tree_add_190_195_groupi_n_4366 ,csa_tree_add_190_195_groupi_n_1523 ,csa_tree_add_190_195_groupi_n_3149);
  or csa_tree_add_190_195_groupi_g44797(csa_tree_add_190_195_groupi_n_4365 ,csa_tree_add_190_195_groupi_n_1519 ,csa_tree_add_190_195_groupi_n_2896);
  nor csa_tree_add_190_195_groupi_g44798(csa_tree_add_190_195_groupi_n_4364 ,csa_tree_add_190_195_groupi_n_2429 ,csa_tree_add_190_195_groupi_n_3040);
  or csa_tree_add_190_195_groupi_g44799(csa_tree_add_190_195_groupi_n_4363 ,csa_tree_add_190_195_groupi_n_1533 ,csa_tree_add_190_195_groupi_n_2861);
  or csa_tree_add_190_195_groupi_g44800(csa_tree_add_190_195_groupi_n_4362 ,csa_tree_add_190_195_groupi_n_1675 ,csa_tree_add_190_195_groupi_n_3392);
  and csa_tree_add_190_195_groupi_g44801(csa_tree_add_190_195_groupi_n_4361 ,csa_tree_add_190_195_groupi_n_1591 ,csa_tree_add_190_195_groupi_n_3473);
  or csa_tree_add_190_195_groupi_g44802(csa_tree_add_190_195_groupi_n_4360 ,csa_tree_add_190_195_groupi_n_969 ,csa_tree_add_190_195_groupi_n_3475);
  and csa_tree_add_190_195_groupi_g44803(csa_tree_add_190_195_groupi_n_4359 ,csa_tree_add_190_195_groupi_n_1990 ,csa_tree_add_190_195_groupi_n_3466);
  and csa_tree_add_190_195_groupi_g44804(csa_tree_add_190_195_groupi_n_4358 ,csa_tree_add_190_195_groupi_n_1833 ,csa_tree_add_190_195_groupi_n_3454);
  and csa_tree_add_190_195_groupi_g44805(csa_tree_add_190_195_groupi_n_4357 ,csa_tree_add_190_195_groupi_n_1603 ,csa_tree_add_190_195_groupi_n_3623);
  nor csa_tree_add_190_195_groupi_g44806(csa_tree_add_190_195_groupi_n_4356 ,csa_tree_add_190_195_groupi_n_2450 ,csa_tree_add_190_195_groupi_n_3701);
  and csa_tree_add_190_195_groupi_g44807(csa_tree_add_190_195_groupi_n_4355 ,csa_tree_add_190_195_groupi_n_1910 ,csa_tree_add_190_195_groupi_n_3626);
  or csa_tree_add_190_195_groupi_g44808(csa_tree_add_190_195_groupi_n_4354 ,csa_tree_add_190_195_groupi_n_2209 ,csa_tree_add_190_195_groupi_n_3700);
  and csa_tree_add_190_195_groupi_g44809(csa_tree_add_190_195_groupi_n_4353 ,in59[13] ,csa_tree_add_190_195_groupi_n_3304);
  or csa_tree_add_190_195_groupi_g44810(csa_tree_add_190_195_groupi_n_4352 ,csa_tree_add_190_195_groupi_n_1701 ,csa_tree_add_190_195_groupi_n_3723);
  or csa_tree_add_190_195_groupi_g44811(csa_tree_add_190_195_groupi_n_4351 ,csa_tree_add_190_195_groupi_n_951 ,csa_tree_add_190_195_groupi_n_3723);
  nor csa_tree_add_190_195_groupi_g44812(csa_tree_add_190_195_groupi_n_4350 ,csa_tree_add_190_195_groupi_n_1562 ,csa_tree_add_190_195_groupi_n_3224);
  nor csa_tree_add_190_195_groupi_g44813(csa_tree_add_190_195_groupi_n_4349 ,csa_tree_add_190_195_groupi_n_2585 ,csa_tree_add_190_195_groupi_n_3143);
  and csa_tree_add_190_195_groupi_g44814(csa_tree_add_190_195_groupi_n_4348 ,in61[10] ,csa_tree_add_190_195_groupi_n_3299);
  and csa_tree_add_190_195_groupi_g44815(csa_tree_add_190_195_groupi_n_4347 ,csa_tree_add_190_195_groupi_n_1600 ,csa_tree_add_190_195_groupi_n_2742);
  and csa_tree_add_190_195_groupi_g44816(csa_tree_add_190_195_groupi_n_4346 ,csa_tree_add_190_195_groupi_n_1693 ,csa_tree_add_190_195_groupi_n_3467);
  and csa_tree_add_190_195_groupi_g44817(csa_tree_add_190_195_groupi_n_4345 ,csa_tree_add_190_195_groupi_n_1779 ,csa_tree_add_190_195_groupi_n_3432);
  or csa_tree_add_190_195_groupi_g44818(csa_tree_add_190_195_groupi_n_4344 ,csa_tree_add_190_195_groupi_n_2052 ,csa_tree_add_190_195_groupi_n_3442);
  or csa_tree_add_190_195_groupi_g44819(csa_tree_add_190_195_groupi_n_4343 ,csa_tree_add_190_195_groupi_n_2391 ,csa_tree_add_190_195_groupi_n_3449);
  or csa_tree_add_190_195_groupi_g44820(csa_tree_add_190_195_groupi_n_4342 ,csa_tree_add_190_195_groupi_n_1949 ,csa_tree_add_190_195_groupi_n_3431);
  or csa_tree_add_190_195_groupi_g44821(csa_tree_add_190_195_groupi_n_4341 ,csa_tree_add_190_195_groupi_n_1005 ,csa_tree_add_190_195_groupi_n_3438);
  or csa_tree_add_190_195_groupi_g44822(csa_tree_add_190_195_groupi_n_4340 ,csa_tree_add_190_195_groupi_n_1689 ,csa_tree_add_190_195_groupi_n_3264);
  and csa_tree_add_190_195_groupi_g44823(csa_tree_add_190_195_groupi_n_4339 ,in60[7] ,csa_tree_add_190_195_groupi_n_3301);
  and csa_tree_add_190_195_groupi_g44824(csa_tree_add_190_195_groupi_n_4338 ,in61[6] ,csa_tree_add_190_195_groupi_n_3293);
  or csa_tree_add_190_195_groupi_g44825(csa_tree_add_190_195_groupi_n_4337 ,csa_tree_add_190_195_groupi_n_2569 ,csa_tree_add_190_195_groupi_n_3280);
  nor csa_tree_add_190_195_groupi_g44826(csa_tree_add_190_195_groupi_n_4336 ,csa_tree_add_190_195_groupi_n_1541 ,csa_tree_add_190_195_groupi_n_3218);
  nor csa_tree_add_190_195_groupi_g44827(csa_tree_add_190_195_groupi_n_4335 ,csa_tree_add_190_195_groupi_n_1546 ,csa_tree_add_190_195_groupi_n_2889);
  nor csa_tree_add_190_195_groupi_g44828(csa_tree_add_190_195_groupi_n_4334 ,csa_tree_add_190_195_groupi_n_1539 ,csa_tree_add_190_195_groupi_n_2932);
  or csa_tree_add_190_195_groupi_g44829(csa_tree_add_190_195_groupi_n_4333 ,csa_tree_add_190_195_groupi_n_1672 ,csa_tree_add_190_195_groupi_n_3258);
  or csa_tree_add_190_195_groupi_g44830(csa_tree_add_190_195_groupi_n_4332 ,in57[7] ,csa_tree_add_190_195_groupi_n_3182);
  or csa_tree_add_190_195_groupi_g44831(csa_tree_add_190_195_groupi_n_4331 ,csa_tree_add_190_195_groupi_n_2542 ,csa_tree_add_190_195_groupi_n_2780);
  or csa_tree_add_190_195_groupi_g44832(csa_tree_add_190_195_groupi_n_4330 ,csa_tree_add_190_195_groupi_n_1156 ,csa_tree_add_190_195_groupi_n_3222);
  and csa_tree_add_190_195_groupi_g44833(csa_tree_add_190_195_groupi_n_4329 ,csa_tree_add_190_195_groupi_n_1753 ,csa_tree_add_190_195_groupi_n_3615);
  or csa_tree_add_190_195_groupi_g44834(csa_tree_add_190_195_groupi_n_4328 ,csa_tree_add_190_195_groupi_n_1902 ,csa_tree_add_190_195_groupi_n_2808);
  or csa_tree_add_190_195_groupi_g44835(csa_tree_add_190_195_groupi_n_4327 ,csa_tree_add_190_195_groupi_n_2059 ,csa_tree_add_190_195_groupi_n_2736);
  or csa_tree_add_190_195_groupi_g44836(csa_tree_add_190_195_groupi_n_4326 ,csa_tree_add_190_195_groupi_n_2117 ,csa_tree_add_190_195_groupi_n_3068);
  and csa_tree_add_190_195_groupi_g44837(csa_tree_add_190_195_groupi_n_4325 ,in61[9] ,csa_tree_add_190_195_groupi_n_3307);
  and csa_tree_add_190_195_groupi_g44838(csa_tree_add_190_195_groupi_n_4324 ,csa_tree_add_190_195_groupi_n_3696 ,csa_tree_add_190_195_groupi_n_3697);
  or csa_tree_add_190_195_groupi_g44839(csa_tree_add_190_195_groupi_n_4323 ,csa_tree_add_190_195_groupi_n_1002 ,csa_tree_add_190_195_groupi_n_3121);
  or csa_tree_add_190_195_groupi_g44840(csa_tree_add_190_195_groupi_n_4322 ,csa_tree_add_190_195_groupi_n_3697 ,csa_tree_add_190_195_groupi_n_3696);
  or csa_tree_add_190_195_groupi_g44841(csa_tree_add_190_195_groupi_n_4321 ,csa_tree_add_190_195_groupi_n_2541 ,csa_tree_add_190_195_groupi_n_3489);
  or csa_tree_add_190_195_groupi_g44842(csa_tree_add_190_195_groupi_n_4320 ,in57[3] ,csa_tree_add_190_195_groupi_n_3238);
  or csa_tree_add_190_195_groupi_g44843(csa_tree_add_190_195_groupi_n_4319 ,csa_tree_add_190_195_groupi_n_1699 ,csa_tree_add_190_195_groupi_n_2883);
  or csa_tree_add_190_195_groupi_g44844(csa_tree_add_190_195_groupi_n_4318 ,csa_tree_add_190_195_groupi_n_2356 ,csa_tree_add_190_195_groupi_n_3183);
  or csa_tree_add_190_195_groupi_g44845(csa_tree_add_190_195_groupi_n_4317 ,csa_tree_add_190_195_groupi_n_1816 ,csa_tree_add_190_195_groupi_n_3641);
  or csa_tree_add_190_195_groupi_g44846(csa_tree_add_190_195_groupi_n_4316 ,csa_tree_add_190_195_groupi_n_2570 ,csa_tree_add_190_195_groupi_n_3050);
  or csa_tree_add_190_195_groupi_g44847(csa_tree_add_190_195_groupi_n_4315 ,csa_tree_add_190_195_groupi_n_3594 ,csa_tree_add_190_195_groupi_n_3703);
  nor csa_tree_add_190_195_groupi_g44848(csa_tree_add_190_195_groupi_n_4314 ,csa_tree_add_190_195_groupi_n_3235 ,csa_tree_add_190_195_groupi_n_966);
  or csa_tree_add_190_195_groupi_g44849(csa_tree_add_190_195_groupi_n_4313 ,csa_tree_add_190_195_groupi_n_919 ,csa_tree_add_190_195_groupi_n_3274);
  and csa_tree_add_190_195_groupi_g44850(csa_tree_add_190_195_groupi_n_4312 ,csa_tree_add_190_195_groupi_n_1692 ,csa_tree_add_190_195_groupi_n_3336);
  nor csa_tree_add_190_195_groupi_g44851(csa_tree_add_190_195_groupi_n_4311 ,csa_tree_add_190_195_groupi_n_1902 ,csa_tree_add_190_195_groupi_n_3062);
  nor csa_tree_add_190_195_groupi_g44852(csa_tree_add_190_195_groupi_n_4310 ,csa_tree_add_190_195_groupi_n_3232 ,csa_tree_add_190_195_groupi_n_784);
  or csa_tree_add_190_195_groupi_g44853(csa_tree_add_190_195_groupi_n_4309 ,csa_tree_add_190_195_groupi_n_2710 ,csa_tree_add_190_195_groupi_n_3576);
  or csa_tree_add_190_195_groupi_g44854(csa_tree_add_190_195_groupi_n_4308 ,in57[2] ,csa_tree_add_190_195_groupi_n_2810);
  and csa_tree_add_190_195_groupi_g44855(csa_tree_add_190_195_groupi_n_4307 ,csa_tree_add_190_195_groupi_n_1632 ,csa_tree_add_190_195_groupi_n_3582);
  or csa_tree_add_190_195_groupi_g44856(csa_tree_add_190_195_groupi_n_4306 ,csa_tree_add_190_195_groupi_n_2008 ,csa_tree_add_190_195_groupi_n_3154);
  and csa_tree_add_190_195_groupi_g44857(csa_tree_add_190_195_groupi_n_4305 ,csa_tree_add_190_195_groupi_n_1578 ,csa_tree_add_190_195_groupi_n_3085);
  or csa_tree_add_190_195_groupi_g44858(csa_tree_add_190_195_groupi_n_4304 ,csa_tree_add_190_195_groupi_n_2674 ,csa_tree_add_190_195_groupi_n_3010);
  and csa_tree_add_190_195_groupi_g44859(csa_tree_add_190_195_groupi_n_4303 ,csa_tree_add_190_195_groupi_n_1641 ,csa_tree_add_190_195_groupi_n_3314);
  or csa_tree_add_190_195_groupi_g44860(csa_tree_add_190_195_groupi_n_4302 ,in56[14] ,csa_tree_add_190_195_groupi_n_3269);
  nor csa_tree_add_190_195_groupi_g44861(csa_tree_add_190_195_groupi_n_4301 ,csa_tree_add_190_195_groupi_n_67 ,csa_tree_add_190_195_groupi_n_1815);
  and csa_tree_add_190_195_groupi_g44862(csa_tree_add_190_195_groupi_n_4300 ,csa_tree_add_190_195_groupi_n_2050 ,csa_tree_add_190_195_groupi_n_3729);
  or csa_tree_add_190_195_groupi_g44863(csa_tree_add_190_195_groupi_n_4299 ,csa_tree_add_190_195_groupi_n_2390 ,csa_tree_add_190_195_groupi_n_3459);
  nor csa_tree_add_190_195_groupi_g44864(csa_tree_add_190_195_groupi_n_4298 ,csa_tree_add_190_195_groupi_n_3159 ,csa_tree_add_190_195_groupi_n_2082);
  or csa_tree_add_190_195_groupi_g44865(csa_tree_add_190_195_groupi_n_4297 ,csa_tree_add_190_195_groupi_n_2547 ,csa_tree_add_190_195_groupi_n_3511);
  or csa_tree_add_190_195_groupi_g44866(csa_tree_add_190_195_groupi_n_4296 ,csa_tree_add_190_195_groupi_n_2545 ,csa_tree_add_190_195_groupi_n_3249);
  and csa_tree_add_190_195_groupi_g44867(csa_tree_add_190_195_groupi_n_4295 ,csa_tree_add_190_195_groupi_n_1972 ,csa_tree_add_190_195_groupi_n_3445);
  and csa_tree_add_190_195_groupi_g44868(csa_tree_add_190_195_groupi_n_4294 ,csa_tree_add_190_195_groupi_n_1811 ,csa_tree_add_190_195_groupi_n_3574);
  or csa_tree_add_190_195_groupi_g44869(csa_tree_add_190_195_groupi_n_4293 ,csa_tree_add_190_195_groupi_n_1872 ,csa_tree_add_190_195_groupi_n_3029);
  nor csa_tree_add_190_195_groupi_g44870(csa_tree_add_190_195_groupi_n_4292 ,csa_tree_add_190_195_groupi_n_2965 ,csa_tree_add_190_195_groupi_n_1948);
  and csa_tree_add_190_195_groupi_g44871(csa_tree_add_190_195_groupi_n_4291 ,csa_tree_add_190_195_groupi_n_2059 ,csa_tree_add_190_195_groupi_n_3263);
  and csa_tree_add_190_195_groupi_g44872(csa_tree_add_190_195_groupi_n_4290 ,csa_tree_add_190_195_groupi_n_223 ,csa_tree_add_190_195_groupi_n_3716);
  or csa_tree_add_190_195_groupi_g44873(csa_tree_add_190_195_groupi_n_4289 ,csa_tree_add_190_195_groupi_n_918 ,csa_tree_add_190_195_groupi_n_3106);
  and csa_tree_add_190_195_groupi_g44874(csa_tree_add_190_195_groupi_n_4288 ,csa_tree_add_190_195_groupi_n_749 ,csa_tree_add_190_195_groupi_n_3428);
  and csa_tree_add_190_195_groupi_g44875(csa_tree_add_190_195_groupi_n_4287 ,csa_tree_add_190_195_groupi_n_1821 ,csa_tree_add_190_195_groupi_n_3591);
  and csa_tree_add_190_195_groupi_g44876(csa_tree_add_190_195_groupi_n_4286 ,csa_tree_add_190_195_groupi_n_1764 ,csa_tree_add_190_195_groupi_n_3291);
  nor csa_tree_add_190_195_groupi_g44877(csa_tree_add_190_195_groupi_n_4285 ,csa_tree_add_190_195_groupi_n_1774 ,csa_tree_add_190_195_groupi_n_3112);
  nor csa_tree_add_190_195_groupi_g44878(csa_tree_add_190_195_groupi_n_4284 ,csa_tree_add_190_195_groupi_n_2902 ,csa_tree_add_190_195_groupi_n_2212);
  and csa_tree_add_190_195_groupi_g44879(csa_tree_add_190_195_groupi_n_4283 ,csa_tree_add_190_195_groupi_n_1766 ,csa_tree_add_190_195_groupi_n_3638);
  or csa_tree_add_190_195_groupi_g44880(csa_tree_add_190_195_groupi_n_4282 ,in56[2] ,csa_tree_add_190_195_groupi_n_3673);
  or csa_tree_add_190_195_groupi_g44881(csa_tree_add_190_195_groupi_n_4281 ,csa_tree_add_190_195_groupi_n_2722 ,csa_tree_add_190_195_groupi_n_3607);
  or csa_tree_add_190_195_groupi_g44882(csa_tree_add_190_195_groupi_n_4280 ,csa_tree_add_190_195_groupi_n_2548 ,csa_tree_add_190_195_groupi_n_3470);
  and csa_tree_add_190_195_groupi_g44883(csa_tree_add_190_195_groupi_n_4279 ,csa_tree_add_190_195_groupi_n_2000 ,csa_tree_add_190_195_groupi_n_3417);
  or csa_tree_add_190_195_groupi_g44884(csa_tree_add_190_195_groupi_n_4278 ,in56[13] ,csa_tree_add_190_195_groupi_n_2952);
  nor csa_tree_add_190_195_groupi_g44885(csa_tree_add_190_195_groupi_n_4277 ,csa_tree_add_190_195_groupi_n_2862 ,csa_tree_add_190_195_groupi_n_756);
  or csa_tree_add_190_195_groupi_g44886(csa_tree_add_190_195_groupi_n_4276 ,csa_tree_add_190_195_groupi_n_2549 ,csa_tree_add_190_195_groupi_n_2923);
  or csa_tree_add_190_195_groupi_g44887(csa_tree_add_190_195_groupi_n_4275 ,csa_tree_add_190_195_groupi_n_1038 ,csa_tree_add_190_195_groupi_n_2901);
  and csa_tree_add_190_195_groupi_g44888(csa_tree_add_190_195_groupi_n_4274 ,csa_tree_add_190_195_groupi_n_922 ,csa_tree_add_190_195_groupi_n_3273);
  and csa_tree_add_190_195_groupi_g44889(csa_tree_add_190_195_groupi_n_4273 ,csa_tree_add_190_195_groupi_n_1813 ,csa_tree_add_190_195_groupi_n_3355);
  and csa_tree_add_190_195_groupi_g44890(csa_tree_add_190_195_groupi_n_4272 ,in60[5] ,csa_tree_add_190_195_groupi_n_3296);
  and csa_tree_add_190_195_groupi_g44891(csa_tree_add_190_195_groupi_n_4271 ,csa_tree_add_190_195_groupi_n_1757 ,csa_tree_add_190_195_groupi_n_3523);
  or csa_tree_add_190_195_groupi_g44892(csa_tree_add_190_195_groupi_n_4270 ,csa_tree_add_190_195_groupi_n_1995 ,csa_tree_add_190_195_groupi_n_2975);
  and csa_tree_add_190_195_groupi_g44893(csa_tree_add_190_195_groupi_n_4269 ,csa_tree_add_190_195_groupi_n_2053 ,csa_tree_add_190_195_groupi_n_3545);
  and csa_tree_add_190_195_groupi_g44894(csa_tree_add_190_195_groupi_n_4268 ,csa_tree_add_190_195_groupi_n_1932 ,csa_tree_add_190_195_groupi_n_3477);
  or csa_tree_add_190_195_groupi_g44895(csa_tree_add_190_195_groupi_n_4267 ,in57[1] ,csa_tree_add_190_195_groupi_n_3671);
  and csa_tree_add_190_195_groupi_g44896(csa_tree_add_190_195_groupi_n_4266 ,csa_tree_add_190_195_groupi_n_1080 ,csa_tree_add_190_195_groupi_n_3362);
  or csa_tree_add_190_195_groupi_g44897(csa_tree_add_190_195_groupi_n_4265 ,csa_tree_add_190_195_groupi_n_2545 ,csa_tree_add_190_195_groupi_n_3156);
  and csa_tree_add_190_195_groupi_g44898(csa_tree_add_190_195_groupi_n_4264 ,csa_tree_add_190_195_groupi_n_1588 ,csa_tree_add_190_195_groupi_n_3465);
  or csa_tree_add_190_195_groupi_g44899(csa_tree_add_190_195_groupi_n_4263 ,csa_tree_add_190_195_groupi_n_1658 ,csa_tree_add_190_195_groupi_n_3391);
  nor csa_tree_add_190_195_groupi_g44900(csa_tree_add_190_195_groupi_n_4262 ,csa_tree_add_190_195_groupi_n_3254 ,csa_tree_add_190_195_groupi_n_1606);
  or csa_tree_add_190_195_groupi_g44901(csa_tree_add_190_195_groupi_n_4261 ,csa_tree_add_190_195_groupi_n_1670 ,csa_tree_add_190_195_groupi_n_3129);
  and csa_tree_add_190_195_groupi_g44902(csa_tree_add_190_195_groupi_n_4260 ,csa_tree_add_190_195_groupi_n_1998 ,csa_tree_add_190_195_groupi_n_2922);
  or csa_tree_add_190_195_groupi_g44903(csa_tree_add_190_195_groupi_n_4259 ,csa_tree_add_190_195_groupi_n_2663 ,csa_tree_add_190_195_groupi_n_2925);
  or csa_tree_add_190_195_groupi_g44904(csa_tree_add_190_195_groupi_n_4258 ,in56[5] ,csa_tree_add_190_195_groupi_n_3086);
  or csa_tree_add_190_195_groupi_g44905(csa_tree_add_190_195_groupi_n_4257 ,csa_tree_add_190_195_groupi_n_1920 ,csa_tree_add_190_195_groupi_n_3565);
  or csa_tree_add_190_195_groupi_g44906(csa_tree_add_190_195_groupi_n_4256 ,csa_tree_add_190_195_groupi_n_1898 ,csa_tree_add_190_195_groupi_n_3531);
  and csa_tree_add_190_195_groupi_g44907(csa_tree_add_190_195_groupi_n_4255 ,csa_tree_add_190_195_groupi_n_1575 ,csa_tree_add_190_195_groupi_n_3570);
  or csa_tree_add_190_195_groupi_g44908(csa_tree_add_190_195_groupi_n_4254 ,csa_tree_add_190_195_groupi_n_2358 ,csa_tree_add_190_195_groupi_n_3187);
  or csa_tree_add_190_195_groupi_g44909(csa_tree_add_190_195_groupi_n_4253 ,csa_tree_add_190_195_groupi_n_1924 ,csa_tree_add_190_195_groupi_n_3135);
  and csa_tree_add_190_195_groupi_g44910(csa_tree_add_190_195_groupi_n_4252 ,csa_tree_add_190_195_groupi_n_2003 ,csa_tree_add_190_195_groupi_n_3502);
  or csa_tree_add_190_195_groupi_g44911(csa_tree_add_190_195_groupi_n_4251 ,csa_tree_add_190_195_groupi_n_2549 ,csa_tree_add_190_195_groupi_n_2864);
  and csa_tree_add_190_195_groupi_g44912(csa_tree_add_190_195_groupi_n_4250 ,csa_tree_add_190_195_groupi_n_1693 ,csa_tree_add_190_195_groupi_n_3380);
  or csa_tree_add_190_195_groupi_g44913(csa_tree_add_190_195_groupi_n_4249 ,csa_tree_add_190_195_groupi_n_2546 ,csa_tree_add_190_195_groupi_n_2962);
  and csa_tree_add_190_195_groupi_g44914(csa_tree_add_190_195_groupi_n_4248 ,in61[8] ,csa_tree_add_190_195_groupi_n_3284);
  or csa_tree_add_190_195_groupi_g44915(csa_tree_add_190_195_groupi_n_4247 ,csa_tree_add_190_195_groupi_n_3704 ,csa_tree_add_190_195_groupi_n_2814);
  nor csa_tree_add_190_195_groupi_g44916(csa_tree_add_190_195_groupi_n_4246 ,csa_tree_add_190_195_groupi_n_2958 ,csa_tree_add_190_195_groupi_n_1989);
  nor csa_tree_add_190_195_groupi_g44917(csa_tree_add_190_195_groupi_n_4245 ,csa_tree_add_190_195_groupi_n_2970 ,csa_tree_add_190_195_groupi_n_844);
  or csa_tree_add_190_195_groupi_g44918(csa_tree_add_190_195_groupi_n_4244 ,csa_tree_add_190_195_groupi_n_2089 ,csa_tree_add_190_195_groupi_n_3694);
  nor csa_tree_add_190_195_groupi_g44919(csa_tree_add_190_195_groupi_n_4243 ,in57[4] ,csa_tree_add_190_195_groupi_n_2873);
  or csa_tree_add_190_195_groupi_g44920(csa_tree_add_190_195_groupi_n_4242 ,csa_tree_add_190_195_groupi_n_2116 ,csa_tree_add_190_195_groupi_n_2980);
  and csa_tree_add_190_195_groupi_g44921(csa_tree_add_190_195_groupi_n_4241 ,csa_tree_add_190_195_groupi_n_1765 ,csa_tree_add_190_195_groupi_n_3557);
  or csa_tree_add_190_195_groupi_g44922(csa_tree_add_190_195_groupi_n_4240 ,csa_tree_add_190_195_groupi_n_2511 ,csa_tree_add_190_195_groupi_n_2918);
  or csa_tree_add_190_195_groupi_g44923(csa_tree_add_190_195_groupi_n_4239 ,csa_tree_add_190_195_groupi_n_1827 ,csa_tree_add_190_195_groupi_n_3175);
  or csa_tree_add_190_195_groupi_g44924(csa_tree_add_190_195_groupi_n_4238 ,csa_tree_add_190_195_groupi_n_3205 ,csa_tree_add_190_195_groupi_n_3515);
  or csa_tree_add_190_195_groupi_g44925(csa_tree_add_190_195_groupi_n_4237 ,csa_tree_add_190_195_groupi_n_2381 ,csa_tree_add_190_195_groupi_n_3083);
  and csa_tree_add_190_195_groupi_g44926(csa_tree_add_190_195_groupi_n_4236 ,csa_tree_add_190_195_groupi_n_524 ,csa_tree_add_190_195_groupi_n_3729);
  or csa_tree_add_190_195_groupi_g44927(csa_tree_add_190_195_groupi_n_4235 ,csa_tree_add_190_195_groupi_n_1759 ,csa_tree_add_190_195_groupi_n_2839);
  or csa_tree_add_190_195_groupi_g44928(csa_tree_add_190_195_groupi_n_4234 ,in57[5] ,csa_tree_add_190_195_groupi_n_2971);
  and csa_tree_add_190_195_groupi_g44929(csa_tree_add_190_195_groupi_n_4233 ,csa_tree_add_190_195_groupi_n_1895 ,csa_tree_add_190_195_groupi_n_3593);
  nor csa_tree_add_190_195_groupi_g44930(csa_tree_add_190_195_groupi_n_4232 ,csa_tree_add_190_195_groupi_n_2056 ,csa_tree_add_190_195_groupi_n_3533);
  and csa_tree_add_190_195_groupi_g44931(csa_tree_add_190_195_groupi_n_4231 ,csa_tree_add_190_195_groupi_n_1644 ,csa_tree_add_190_195_groupi_n_3272);
  and csa_tree_add_190_195_groupi_g44932(csa_tree_add_190_195_groupi_n_4230 ,csa_tree_add_190_195_groupi_n_1870 ,csa_tree_add_190_195_groupi_n_3319);
  and csa_tree_add_190_195_groupi_g44933(csa_tree_add_190_195_groupi_n_4229 ,csa_tree_add_190_195_groupi_n_1777 ,csa_tree_add_190_195_groupi_n_3561);
  or csa_tree_add_190_195_groupi_g44934(csa_tree_add_190_195_groupi_n_4228 ,csa_tree_add_190_195_groupi_n_1617 ,csa_tree_add_190_195_groupi_n_3298);
  and csa_tree_add_190_195_groupi_g44935(csa_tree_add_190_195_groupi_n_4227 ,in61[11] ,csa_tree_add_190_195_groupi_n_3289);
  nor csa_tree_add_190_195_groupi_g44936(csa_tree_add_190_195_groupi_n_4226 ,csa_tree_add_190_195_groupi_n_68 ,csa_tree_add_190_195_groupi_n_1915);
  and csa_tree_add_190_195_groupi_g44937(csa_tree_add_190_195_groupi_n_4225 ,in59[4] ,csa_tree_add_190_195_groupi_n_3292);
  and csa_tree_add_190_195_groupi_g44938(csa_tree_add_190_195_groupi_n_4224 ,csa_tree_add_190_195_groupi_n_2156 ,csa_tree_add_190_195_groupi_n_3398);
  and csa_tree_add_190_195_groupi_g44939(csa_tree_add_190_195_groupi_n_4223 ,csa_tree_add_190_195_groupi_n_1635 ,csa_tree_add_190_195_groupi_n_3326);
  or csa_tree_add_190_195_groupi_g44940(csa_tree_add_190_195_groupi_n_4222 ,csa_tree_add_190_195_groupi_n_906 ,csa_tree_add_190_195_groupi_n_2832);
  or csa_tree_add_190_195_groupi_g44941(csa_tree_add_190_195_groupi_n_4221 ,csa_tree_add_190_195_groupi_n_2543 ,csa_tree_add_190_195_groupi_n_3036);
  or csa_tree_add_190_195_groupi_g44942(csa_tree_add_190_195_groupi_n_4220 ,csa_tree_add_190_195_groupi_n_1888 ,csa_tree_add_190_195_groupi_n_3041);
  or csa_tree_add_190_195_groupi_g44943(csa_tree_add_190_195_groupi_n_4219 ,in57[9] ,csa_tree_add_190_195_groupi_n_2741);
  or csa_tree_add_190_195_groupi_g44944(csa_tree_add_190_195_groupi_n_4218 ,in57[11] ,csa_tree_add_190_195_groupi_n_2924);
  and csa_tree_add_190_195_groupi_g44945(csa_tree_add_190_195_groupi_n_4217 ,csa_tree_add_190_195_groupi_n_1755 ,csa_tree_add_190_195_groupi_n_3721);
  and csa_tree_add_190_195_groupi_g44946(csa_tree_add_190_195_groupi_n_4216 ,csa_tree_add_190_195_groupi_n_1853 ,csa_tree_add_190_195_groupi_n_3342);
  and csa_tree_add_190_195_groupi_g44947(csa_tree_add_190_195_groupi_n_4215 ,csa_tree_add_190_195_groupi_n_1755 ,csa_tree_add_190_195_groupi_n_3544);
  and csa_tree_add_190_195_groupi_g44948(csa_tree_add_190_195_groupi_n_4214 ,csa_tree_add_190_195_groupi_n_1987 ,csa_tree_add_190_195_groupi_n_3393);
  or csa_tree_add_190_195_groupi_g44949(csa_tree_add_190_195_groupi_n_4213 ,csa_tree_add_190_195_groupi_n_2711 ,csa_tree_add_190_195_groupi_n_3518);
  or csa_tree_add_190_195_groupi_g44950(csa_tree_add_190_195_groupi_n_4212 ,csa_tree_add_190_195_groupi_n_1699 ,csa_tree_add_190_195_groupi_n_3536);
  or csa_tree_add_190_195_groupi_g44951(csa_tree_add_190_195_groupi_n_4211 ,in58[15] ,csa_tree_add_190_195_groupi_n_3297);
  or csa_tree_add_190_195_groupi_g44952(csa_tree_add_190_195_groupi_n_4210 ,csa_tree_add_190_195_groupi_n_1655 ,csa_tree_add_190_195_groupi_n_3421);
  and csa_tree_add_190_195_groupi_g44953(csa_tree_add_190_195_groupi_n_4209 ,csa_tree_add_190_195_groupi_n_1633 ,csa_tree_add_190_195_groupi_n_3395);
  and csa_tree_add_190_195_groupi_g44954(csa_tree_add_190_195_groupi_n_4208 ,csa_tree_add_190_195_groupi_n_1605 ,csa_tree_add_190_195_groupi_n_3394);
  or csa_tree_add_190_195_groupi_g44955(csa_tree_add_190_195_groupi_n_4207 ,csa_tree_add_190_195_groupi_n_2514 ,csa_tree_add_190_195_groupi_n_3150);
  and csa_tree_add_190_195_groupi_g44956(csa_tree_add_190_195_groupi_n_4206 ,csa_tree_add_190_195_groupi_n_1891 ,csa_tree_add_190_195_groupi_n_3512);
  or csa_tree_add_190_195_groupi_g44957(csa_tree_add_190_195_groupi_n_4205 ,csa_tree_add_190_195_groupi_n_945 ,csa_tree_add_190_195_groupi_n_3406);
  or csa_tree_add_190_195_groupi_g44958(csa_tree_add_190_195_groupi_n_4204 ,csa_tree_add_190_195_groupi_n_2717 ,csa_tree_add_190_195_groupi_n_3115);
  or csa_tree_add_190_195_groupi_g44959(csa_tree_add_190_195_groupi_n_4203 ,csa_tree_add_190_195_groupi_n_1963 ,csa_tree_add_190_195_groupi_n_2788);
  or csa_tree_add_190_195_groupi_g44960(csa_tree_add_190_195_groupi_n_4202 ,in57[13] ,csa_tree_add_190_195_groupi_n_3551);
  and csa_tree_add_190_195_groupi_g44961(csa_tree_add_190_195_groupi_n_4201 ,csa_tree_add_190_195_groupi_n_1810 ,csa_tree_add_190_195_groupi_n_3386);
  nor csa_tree_add_190_195_groupi_g44962(csa_tree_add_190_195_groupi_n_4200 ,csa_tree_add_190_195_groupi_n_1867 ,csa_tree_add_190_195_groupi_n_3045);
  or csa_tree_add_190_195_groupi_g44963(csa_tree_add_190_195_groupi_n_4199 ,csa_tree_add_190_195_groupi_n_2664 ,csa_tree_add_190_195_groupi_n_3525);
  and csa_tree_add_190_195_groupi_g44964(csa_tree_add_190_195_groupi_n_4198 ,csa_tree_add_190_195_groupi_n_1577 ,csa_tree_add_190_195_groupi_n_3444);
  and csa_tree_add_190_195_groupi_g44965(csa_tree_add_190_195_groupi_n_4197 ,csa_tree_add_190_195_groupi_n_1592 ,csa_tree_add_190_195_groupi_n_3399);
  or csa_tree_add_190_195_groupi_g44966(csa_tree_add_190_195_groupi_n_4196 ,csa_tree_add_190_195_groupi_n_1949 ,csa_tree_add_190_195_groupi_n_2941);
  and csa_tree_add_190_195_groupi_g44967(csa_tree_add_190_195_groupi_n_4195 ,csa_tree_add_190_195_groupi_n_2089 ,csa_tree_add_190_195_groupi_n_3694);
  and csa_tree_add_190_195_groupi_g44968(csa_tree_add_190_195_groupi_n_4194 ,csa_tree_add_190_195_groupi_n_1744 ,csa_tree_add_190_195_groupi_n_3328);
  or csa_tree_add_190_195_groupi_g44969(csa_tree_add_190_195_groupi_n_4193 ,csa_tree_add_190_195_groupi_n_921 ,csa_tree_add_190_195_groupi_n_2833);
  or csa_tree_add_190_195_groupi_g44970(csa_tree_add_190_195_groupi_n_4192 ,csa_tree_add_190_195_groupi_n_2378 ,csa_tree_add_190_195_groupi_n_3726);
  or csa_tree_add_190_195_groupi_g44971(csa_tree_add_190_195_groupi_n_4191 ,csa_tree_add_190_195_groupi_n_1704 ,csa_tree_add_190_195_groupi_n_3054);
  or csa_tree_add_190_195_groupi_g44972(csa_tree_add_190_195_groupi_n_4190 ,csa_tree_add_190_195_groupi_n_2507 ,csa_tree_add_190_195_groupi_n_2798);
  and csa_tree_add_190_195_groupi_g44973(csa_tree_add_190_195_groupi_n_4189 ,csa_tree_add_190_195_groupi_n_2116 ,csa_tree_add_190_195_groupi_n_3446);
  and csa_tree_add_190_195_groupi_g44974(csa_tree_add_190_195_groupi_n_4188 ,csa_tree_add_190_195_groupi_n_1574 ,csa_tree_add_190_195_groupi_n_3521);
  and csa_tree_add_190_195_groupi_g44975(csa_tree_add_190_195_groupi_n_4187 ,csa_tree_add_190_195_groupi_n_1673 ,csa_tree_add_190_195_groupi_n_3340);
  nor csa_tree_add_190_195_groupi_g44976(csa_tree_add_190_195_groupi_n_4186 ,csa_tree_add_190_195_groupi_n_2992 ,csa_tree_add_190_195_groupi_n_1068);
  nor csa_tree_add_190_195_groupi_g44977(csa_tree_add_190_195_groupi_n_4185 ,csa_tree_add_190_195_groupi_n_3522 ,csa_tree_add_190_195_groupi_n_3705);
  or csa_tree_add_190_195_groupi_g44978(csa_tree_add_190_195_groupi_n_4184 ,csa_tree_add_190_195_groupi_n_1856 ,csa_tree_add_190_195_groupi_n_3389);
  nor csa_tree_add_190_195_groupi_g44979(csa_tree_add_190_195_groupi_n_4183 ,csa_tree_add_190_195_groupi_n_1624 ,csa_tree_add_190_195_groupi_n_3541);
  nor csa_tree_add_190_195_groupi_g44980(csa_tree_add_190_195_groupi_n_4182 ,in57[8] ,csa_tree_add_190_195_groupi_n_2767);
  and csa_tree_add_190_195_groupi_g44981(csa_tree_add_190_195_groupi_n_4181 ,in59[0] ,csa_tree_add_190_195_groupi_n_2806);
  and csa_tree_add_190_195_groupi_g44982(csa_tree_add_190_195_groupi_n_4180 ,csa_tree_add_190_195_groupi_n_1629 ,csa_tree_add_190_195_groupi_n_3174);
  or csa_tree_add_190_195_groupi_g44983(csa_tree_add_190_195_groupi_n_4179 ,csa_tree_add_190_195_groupi_n_3206 ,csa_tree_add_190_195_groupi_n_3268);
  and csa_tree_add_190_195_groupi_g44984(csa_tree_add_190_195_groupi_n_4178 ,csa_tree_add_190_195_groupi_n_1817 ,csa_tree_add_190_195_groupi_n_3496);
  or csa_tree_add_190_195_groupi_g44985(csa_tree_add_190_195_groupi_n_4177 ,csa_tree_add_190_195_groupi_n_864 ,csa_tree_add_190_195_groupi_n_3148);
  or csa_tree_add_190_195_groupi_g44986(csa_tree_add_190_195_groupi_n_4176 ,csa_tree_add_190_195_groupi_n_2546 ,csa_tree_add_190_195_groupi_n_2818);
  or csa_tree_add_190_195_groupi_g44987(csa_tree_add_190_195_groupi_n_4175 ,in56[4] ,csa_tree_add_190_195_groupi_n_2954);
  or csa_tree_add_190_195_groupi_g44988(csa_tree_add_190_195_groupi_n_4174 ,csa_tree_add_190_195_groupi_n_2513 ,csa_tree_add_190_195_groupi_n_3005);
  or csa_tree_add_190_195_groupi_g44989(csa_tree_add_190_195_groupi_n_4173 ,csa_tree_add_190_195_groupi_n_1846 ,csa_tree_add_190_195_groupi_n_3218);
  or csa_tree_add_190_195_groupi_g44990(csa_tree_add_190_195_groupi_n_4172 ,csa_tree_add_190_195_groupi_n_2064 ,csa_tree_add_190_195_groupi_n_3244);
  nor csa_tree_add_190_195_groupi_g44991(csa_tree_add_190_195_groupi_n_4171 ,csa_tree_add_190_195_groupi_n_3136 ,csa_tree_add_190_195_groupi_n_3208);
  or csa_tree_add_190_195_groupi_g44992(csa_tree_add_190_195_groupi_n_4170 ,in57[6] ,csa_tree_add_190_195_groupi_n_2953);
  and csa_tree_add_190_195_groupi_g44993(csa_tree_add_190_195_groupi_n_4169 ,csa_tree_add_190_195_groupi_n_1963 ,csa_tree_add_190_195_groupi_n_3706);
  or csa_tree_add_190_195_groupi_g44994(csa_tree_add_190_195_groupi_n_4168 ,csa_tree_add_190_195_groupi_n_1119 ,csa_tree_add_190_195_groupi_n_3073);
  or csa_tree_add_190_195_groupi_g44995(csa_tree_add_190_195_groupi_n_4167 ,csa_tree_add_190_195_groupi_n_1017 ,csa_tree_add_190_195_groupi_n_3419);
  and csa_tree_add_190_195_groupi_g44996(csa_tree_add_190_195_groupi_n_4166 ,csa_tree_add_190_195_groupi_n_1686 ,csa_tree_add_190_195_groupi_n_3681);
  or csa_tree_add_190_195_groupi_g44997(csa_tree_add_190_195_groupi_n_4165 ,csa_tree_add_190_195_groupi_n_1911 ,csa_tree_add_190_195_groupi_n_3219);
  or csa_tree_add_190_195_groupi_g44998(csa_tree_add_190_195_groupi_n_4164 ,in57[0] ,csa_tree_add_190_195_groupi_n_3688);
  and csa_tree_add_190_195_groupi_g44999(csa_tree_add_190_195_groupi_n_4163 ,csa_tree_add_190_195_groupi_n_1949 ,csa_tree_add_190_195_groupi_n_3334);
  and csa_tree_add_190_195_groupi_g45000(csa_tree_add_190_195_groupi_n_4162 ,csa_tree_add_190_195_groupi_n_1703 ,csa_tree_add_190_195_groupi_n_2762);
  nor csa_tree_add_190_195_groupi_g45001(csa_tree_add_190_195_groupi_n_4161 ,csa_tree_add_190_195_groupi_n_3108 ,csa_tree_add_190_195_groupi_n_1844);
  or csa_tree_add_190_195_groupi_g45002(csa_tree_add_190_195_groupi_n_4160 ,in56[12] ,csa_tree_add_190_195_groupi_n_3104);
  or csa_tree_add_190_195_groupi_g45003(csa_tree_add_190_195_groupi_n_4159 ,csa_tree_add_190_195_groupi_n_1897 ,csa_tree_add_190_195_groupi_n_3664);
  or csa_tree_add_190_195_groupi_g45004(csa_tree_add_190_195_groupi_n_4158 ,csa_tree_add_190_195_groupi_n_2357 ,csa_tree_add_190_195_groupi_n_2773);
  or csa_tree_add_190_195_groupi_g45005(csa_tree_add_190_195_groupi_n_4157 ,csa_tree_add_190_195_groupi_n_1762 ,csa_tree_add_190_195_groupi_n_2807);
  and csa_tree_add_190_195_groupi_g45006(csa_tree_add_190_195_groupi_n_4156 ,csa_tree_add_190_195_groupi_n_2056 ,csa_tree_add_190_195_groupi_n_3453);
  or csa_tree_add_190_195_groupi_g45007(csa_tree_add_190_195_groupi_n_4155 ,csa_tree_add_190_195_groupi_n_1997 ,csa_tree_add_190_195_groupi_n_3381);
  or csa_tree_add_190_195_groupi_g45008(csa_tree_add_190_195_groupi_n_4154 ,csa_tree_add_190_195_groupi_n_1656 ,csa_tree_add_190_195_groupi_n_2760);
  and csa_tree_add_190_195_groupi_g45009(csa_tree_add_190_195_groupi_n_4153 ,csa_tree_add_190_195_groupi_n_1652 ,csa_tree_add_190_195_groupi_n_3387);
  or csa_tree_add_190_195_groupi_g45010(csa_tree_add_190_195_groupi_n_4152 ,csa_tree_add_190_195_groupi_n_2678 ,csa_tree_add_190_195_groupi_n_3016);
  nor csa_tree_add_190_195_groupi_g45011(csa_tree_add_190_195_groupi_n_4151 ,in57[10] ,csa_tree_add_190_195_groupi_n_3123);
  or csa_tree_add_190_195_groupi_g45012(csa_tree_add_190_195_groupi_n_4150 ,csa_tree_add_190_195_groupi_n_2566 ,csa_tree_add_190_195_groupi_n_2785);
  or csa_tree_add_190_195_groupi_g45013(csa_tree_add_190_195_groupi_n_4149 ,csa_tree_add_190_195_groupi_n_3207 ,csa_tree_add_190_195_groupi_n_3678);
  and csa_tree_add_190_195_groupi_g45014(csa_tree_add_190_195_groupi_n_4148 ,csa_tree_add_190_195_groupi_n_1594 ,csa_tree_add_190_195_groupi_n_3433);
  nor csa_tree_add_190_195_groupi_g45015(csa_tree_add_190_195_groupi_n_4147 ,csa_tree_add_190_195_groupi_n_3075 ,csa_tree_add_190_195_groupi_n_2087);
  nor csa_tree_add_190_195_groupi_g45016(csa_tree_add_190_195_groupi_n_4146 ,csa_tree_add_190_195_groupi_n_3078 ,csa_tree_add_190_195_groupi_n_2039);
  or csa_tree_add_190_195_groupi_g45017(csa_tree_add_190_195_groupi_n_4145 ,csa_tree_add_190_195_groupi_n_3720 ,csa_tree_add_190_195_groupi_n_3713);
  nor csa_tree_add_190_195_groupi_g45018(csa_tree_add_190_195_groupi_n_4144 ,csa_tree_add_190_195_groupi_n_3226 ,csa_tree_add_190_195_groupi_n_3211);
  and csa_tree_add_190_195_groupi_g45019(csa_tree_add_190_195_groupi_n_4143 ,csa_tree_add_190_195_groupi_n_3210 ,csa_tree_add_190_195_groupi_n_3221);
  or csa_tree_add_190_195_groupi_g45020(csa_tree_add_190_195_groupi_n_4570 ,csa_tree_add_190_195_groupi_n_2764 ,csa_tree_add_190_195_groupi_n_1354);
  and csa_tree_add_190_195_groupi_g45021(csa_tree_add_190_195_groupi_n_4569 ,csa_tree_add_190_195_groupi_n_3056 ,csa_tree_add_190_195_groupi_n_3204);
  xnor csa_tree_add_190_195_groupi_g45022(csa_tree_add_190_195_groupi_n_4568 ,csa_tree_add_190_195_groupi_n_1916 ,csa_tree_add_190_195_groupi_n_1842);
  or csa_tree_add_190_195_groupi_g45023(csa_tree_add_190_195_groupi_n_4567 ,csa_tree_add_190_195_groupi_n_3151 ,csa_tree_add_190_195_groupi_n_1348);
  and csa_tree_add_190_195_groupi_g45024(csa_tree_add_190_195_groupi_n_4566 ,csa_tree_add_190_195_groupi_n_3614 ,csa_tree_add_190_195_groupi_n_1314);
  and csa_tree_add_190_195_groupi_g45025(csa_tree_add_190_195_groupi_n_4565 ,csa_tree_add_190_195_groupi_n_3695 ,csa_tree_add_190_195_groupi_n_3669);
  and csa_tree_add_190_195_groupi_g45026(csa_tree_add_190_195_groupi_n_4563 ,csa_tree_add_190_195_groupi_n_3683 ,csa_tree_add_190_195_groupi_n_3692);
  or csa_tree_add_190_195_groupi_g45027(csa_tree_add_190_195_groupi_n_4561 ,csa_tree_add_190_195_groupi_n_3011 ,csa_tree_add_190_195_groupi_n_1329);
  not csa_tree_add_190_195_groupi_g45028(csa_tree_add_190_195_groupi_n_4133 ,csa_tree_add_190_195_groupi_n_4134);
  not csa_tree_add_190_195_groupi_g45029(csa_tree_add_190_195_groupi_n_4126 ,csa_tree_add_190_195_groupi_n_4127);
  not csa_tree_add_190_195_groupi_g45030(csa_tree_add_190_195_groupi_n_4116 ,csa_tree_add_190_195_groupi_n_4117);
  not csa_tree_add_190_195_groupi_g45031(csa_tree_add_190_195_groupi_n_4115 ,csa_tree_add_190_195_groupi_n_4114);
  xnor csa_tree_add_190_195_groupi_g45032(csa_tree_add_190_195_groupi_n_4113 ,csa_tree_add_190_195_groupi_n_742 ,csa_tree_add_190_195_groupi_n_970);
  xnor csa_tree_add_190_195_groupi_g45033(csa_tree_add_190_195_groupi_n_4112 ,in55[2] ,in55[0]);
  xnor csa_tree_add_190_195_groupi_g45034(csa_tree_add_190_195_groupi_n_4111 ,csa_tree_add_190_195_groupi_n_564 ,csa_tree_add_190_195_groupi_n_2117);
  xnor csa_tree_add_190_195_groupi_g45035(csa_tree_add_190_195_groupi_n_4110 ,csa_tree_add_190_195_groupi_n_538 ,csa_tree_add_190_195_groupi_n_1998);
  xnor csa_tree_add_190_195_groupi_g45036(csa_tree_add_190_195_groupi_n_4109 ,csa_tree_add_190_195_groupi_n_362 ,csa_tree_add_190_195_groupi_n_1900);
  xnor csa_tree_add_190_195_groupi_g45037(csa_tree_add_190_195_groupi_n_4108 ,csa_tree_add_190_195_groupi_n_411 ,csa_tree_add_190_195_groupi_n_1165);
  xnor csa_tree_add_190_195_groupi_g45038(csa_tree_add_190_195_groupi_n_4107 ,csa_tree_add_190_195_groupi_n_1030 ,in55[1]);
  xnor csa_tree_add_190_195_groupi_g45039(csa_tree_add_190_195_groupi_n_4106 ,csa_tree_add_190_195_groupi_n_973 ,csa_tree_add_190_195_groupi_n_1005);
  xnor csa_tree_add_190_195_groupi_g45040(csa_tree_add_190_195_groupi_n_4105 ,csa_tree_add_190_195_groupi_n_1824 ,csa_tree_add_190_195_groupi_n_1819);
  xnor csa_tree_add_190_195_groupi_g45041(csa_tree_add_190_195_groupi_n_4104 ,csa_tree_add_190_195_groupi_n_865 ,csa_tree_add_190_195_groupi_n_1578);
  xnor csa_tree_add_190_195_groupi_g45042(csa_tree_add_190_195_groupi_n_4103 ,csa_tree_add_190_195_groupi_n_1904 ,csa_tree_add_190_195_groupi_n_1963);
  xnor csa_tree_add_190_195_groupi_g45043(csa_tree_add_190_195_groupi_n_4102 ,csa_tree_add_190_195_groupi_n_266 ,csa_tree_add_190_195_groupi_n_1840);
  xnor csa_tree_add_190_195_groupi_g45044(csa_tree_add_190_195_groupi_n_4101 ,csa_tree_add_190_195_groupi_n_610 ,csa_tree_add_190_195_groupi_n_1653);
  xnor csa_tree_add_190_195_groupi_g45045(csa_tree_add_190_195_groupi_n_4100 ,csa_tree_add_190_195_groupi_n_1921 ,csa_tree_add_190_195_groupi_n_1641);
  xnor csa_tree_add_190_195_groupi_g45046(csa_tree_add_190_195_groupi_n_4099 ,csa_tree_add_190_195_groupi_n_1970 ,csa_tree_add_190_195_groupi_n_1758);
  xnor csa_tree_add_190_195_groupi_g45047(csa_tree_add_190_195_groupi_n_4098 ,csa_tree_add_190_195_groupi_n_1974 ,csa_tree_add_190_195_groupi_n_1868);
  xnor csa_tree_add_190_195_groupi_g45048(csa_tree_add_190_195_groupi_n_4097 ,csa_tree_add_190_195_groupi_n_2051 ,csa_tree_add_190_195_groupi_n_1972);
  xnor csa_tree_add_190_195_groupi_g45049(csa_tree_add_190_195_groupi_n_4096 ,csa_tree_add_190_195_groupi_n_1877 ,csa_tree_add_190_195_groupi_n_1618);
  xnor csa_tree_add_190_195_groupi_g45050(csa_tree_add_190_195_groupi_n_4095 ,csa_tree_add_190_195_groupi_n_1973 ,csa_tree_add_190_195_groupi_n_1762);
  xnor csa_tree_add_190_195_groupi_g45051(csa_tree_add_190_195_groupi_n_4094 ,csa_tree_add_190_195_groupi_n_1060 ,csa_tree_add_190_195_groupi_n_1679);
  xnor csa_tree_add_190_195_groupi_g45052(csa_tree_add_190_195_groupi_n_4093 ,csa_tree_add_190_195_groupi_n_1960 ,csa_tree_add_190_195_groupi_n_1694);
  xnor csa_tree_add_190_195_groupi_g45053(csa_tree_add_190_195_groupi_n_4092 ,csa_tree_add_190_195_groupi_n_1845 ,csa_tree_add_190_195_groupi_n_1671);
  xnor csa_tree_add_190_195_groupi_g45054(csa_tree_add_190_195_groupi_n_4091 ,csa_tree_add_190_195_groupi_n_2084 ,csa_tree_add_190_195_groupi_n_2003);
  xnor csa_tree_add_190_195_groupi_g45055(csa_tree_add_190_195_groupi_n_4090 ,in55[14] ,in55[10]);
  xnor csa_tree_add_190_195_groupi_g45056(csa_tree_add_190_195_groupi_n_4089 ,csa_tree_add_190_195_groupi_n_2057 ,csa_tree_add_190_195_groupi_n_1869);
  xnor csa_tree_add_190_195_groupi_g45057(csa_tree_add_190_195_groupi_n_4088 ,in60[13] ,in56[13]);
  xnor csa_tree_add_190_195_groupi_g45058(csa_tree_add_190_195_groupi_n_4087 ,csa_tree_add_190_195_groupi_n_386 ,csa_tree_add_190_195_groupi_n_1960);
  xnor csa_tree_add_190_195_groupi_g45059(csa_tree_add_190_195_groupi_n_4086 ,csa_tree_add_190_195_groupi_n_1255 ,csa_tree_add_190_195_groupi_n_1027);
  xnor csa_tree_add_190_195_groupi_g45060(csa_tree_add_190_195_groupi_n_4085 ,csa_tree_add_190_195_groupi_n_230 ,csa_tree_add_190_195_groupi_n_1822);
  xnor csa_tree_add_190_195_groupi_g45061(csa_tree_add_190_195_groupi_n_4084 ,csa_tree_add_190_195_groupi_n_1923 ,csa_tree_add_190_195_groupi_n_1922);
  xnor csa_tree_add_190_195_groupi_g45062(csa_tree_add_190_195_groupi_n_4083 ,in56[0] ,in57[0]);
  xnor csa_tree_add_190_195_groupi_g45063(csa_tree_add_190_195_groupi_n_4082 ,csa_tree_add_190_195_groupi_n_1604 ,csa_tree_add_190_195_groupi_n_1605);
  xnor csa_tree_add_190_195_groupi_g45064(csa_tree_add_190_195_groupi_n_4081 ,in58[7] ,in56[7]);
  xnor csa_tree_add_190_195_groupi_g45065(csa_tree_add_190_195_groupi_n_4080 ,csa_tree_add_190_195_groupi_n_2062 ,csa_tree_add_190_195_groupi_n_999);
  xnor csa_tree_add_190_195_groupi_g45066(csa_tree_add_190_195_groupi_n_4079 ,csa_tree_add_190_195_groupi_n_2086 ,csa_tree_add_190_195_groupi_n_2003);
  xnor csa_tree_add_190_195_groupi_g45067(csa_tree_add_190_195_groupi_n_4078 ,in61[2] ,in57[2]);
  xnor csa_tree_add_190_195_groupi_g45068(csa_tree_add_190_195_groupi_n_4077 ,csa_tree_add_190_195_groupi_n_405 ,csa_tree_add_190_195_groupi_n_1146);
  xnor csa_tree_add_190_195_groupi_g45069(csa_tree_add_190_195_groupi_n_4076 ,csa_tree_add_190_195_groupi_n_852 ,csa_tree_add_190_195_groupi_n_1713);
  xnor csa_tree_add_190_195_groupi_g45070(csa_tree_add_190_195_groupi_n_4075 ,csa_tree_add_190_195_groupi_n_1847 ,csa_tree_add_190_195_groupi_n_1586);
  xnor csa_tree_add_190_195_groupi_g45071(csa_tree_add_190_195_groupi_n_4074 ,csa_tree_add_190_195_groupi_n_375 ,csa_tree_add_190_195_groupi_n_1890);
  xnor csa_tree_add_190_195_groupi_g45072(csa_tree_add_190_195_groupi_n_4073 ,csa_tree_add_190_195_groupi_n_222 ,csa_tree_add_190_195_groupi_n_1897);
  xnor csa_tree_add_190_195_groupi_g45073(csa_tree_add_190_195_groupi_n_4072 ,csa_tree_add_190_195_groupi_n_1820 ,csa_tree_add_190_195_groupi_n_1697);
  xnor csa_tree_add_190_195_groupi_g45074(csa_tree_add_190_195_groupi_n_4071 ,csa_tree_add_190_195_groupi_n_2005 ,csa_tree_add_190_195_groupi_n_2004);
  xnor csa_tree_add_190_195_groupi_g45075(csa_tree_add_190_195_groupi_n_4070 ,csa_tree_add_190_195_groupi_n_2061 ,csa_tree_add_190_195_groupi_n_1835);
  xnor csa_tree_add_190_195_groupi_g45076(csa_tree_add_190_195_groupi_n_4069 ,csa_tree_add_190_195_groupi_n_2007 ,csa_tree_add_190_195_groupi_n_1902);
  xnor csa_tree_add_190_195_groupi_g45077(csa_tree_add_190_195_groupi_n_4068 ,csa_tree_add_190_195_groupi_n_1892 ,csa_tree_add_190_195_groupi_n_1766);
  xnor csa_tree_add_190_195_groupi_g45078(csa_tree_add_190_195_groupi_n_4067 ,csa_tree_add_190_195_groupi_n_332 ,csa_tree_add_190_195_groupi_n_2063);
  xnor csa_tree_add_190_195_groupi_g45079(csa_tree_add_190_195_groupi_n_4066 ,csa_tree_add_190_195_groupi_n_2090 ,csa_tree_add_190_195_groupi_n_1991);
  xnor csa_tree_add_190_195_groupi_g45080(csa_tree_add_190_195_groupi_n_4065 ,csa_tree_add_190_195_groupi_n_2055 ,csa_tree_add_190_195_groupi_n_2053);
  xnor csa_tree_add_190_195_groupi_g45082(csa_tree_add_190_195_groupi_n_4064 ,csa_tree_add_190_195_groupi_n_1014 ,csa_tree_add_190_195_groupi_n_1678);
  xnor csa_tree_add_190_195_groupi_g45083(csa_tree_add_190_195_groupi_n_4063 ,csa_tree_add_190_195_groupi_n_574 ,csa_tree_add_190_195_groupi_n_1914);
  xnor csa_tree_add_190_195_groupi_g45084(csa_tree_add_190_195_groupi_n_4062 ,csa_tree_add_190_195_groupi_n_2158 ,csa_tree_add_190_195_groupi_n_1744);
  xnor csa_tree_add_190_195_groupi_g45085(csa_tree_add_190_195_groupi_n_4061 ,csa_tree_add_190_195_groupi_n_199 ,csa_tree_add_190_195_groupi_n_1623);
  xnor csa_tree_add_190_195_groupi_g45086(csa_tree_add_190_195_groupi_n_4060 ,csa_tree_add_190_195_groupi_n_1962 ,csa_tree_add_190_195_groupi_n_1856);
  xnor csa_tree_add_190_195_groupi_g45087(csa_tree_add_190_195_groupi_n_4059 ,csa_tree_add_190_195_groupi_n_384 ,csa_tree_add_190_195_groupi_n_2060);
  xnor csa_tree_add_190_195_groupi_g45088(csa_tree_add_190_195_groupi_n_4058 ,csa_tree_add_190_195_groupi_n_1844 ,csa_tree_add_190_195_groupi_n_2008);
  xnor csa_tree_add_190_195_groupi_g45089(csa_tree_add_190_195_groupi_n_4057 ,csa_tree_add_190_195_groupi_n_985 ,csa_tree_add_190_195_groupi_n_1743);
  xnor csa_tree_add_190_195_groupi_g45090(csa_tree_add_190_195_groupi_n_4056 ,csa_tree_add_190_195_groupi_n_1706 ,csa_tree_add_190_195_groupi_n_922);
  xnor csa_tree_add_190_195_groupi_g45091(csa_tree_add_190_195_groupi_n_4055 ,csa_tree_add_190_195_groupi_n_317 ,csa_tree_add_190_195_groupi_n_1815);
  xnor csa_tree_add_190_195_groupi_g45092(csa_tree_add_190_195_groupi_n_4054 ,csa_tree_add_190_195_groupi_n_2063 ,csa_tree_add_190_195_groupi_n_1989);
  xnor csa_tree_add_190_195_groupi_g45093(csa_tree_add_190_195_groupi_n_4053 ,in59[15] ,in56[15]);
  xnor csa_tree_add_190_195_groupi_g45094(csa_tree_add_190_195_groupi_n_4052 ,csa_tree_add_190_195_groupi_n_491 ,csa_tree_add_190_195_groupi_n_1269);
  xnor csa_tree_add_190_195_groupi_g45095(csa_tree_add_190_195_groupi_n_4051 ,csa_tree_add_190_195_groupi_n_2054 ,csa_tree_add_190_195_groupi_n_1036);
  xnor csa_tree_add_190_195_groupi_g45096(csa_tree_add_190_195_groupi_n_4050 ,in60[4] ,in57[4]);
  xnor csa_tree_add_190_195_groupi_g45097(csa_tree_add_190_195_groupi_n_4049 ,csa_tree_add_190_195_groupi_n_1029 ,csa_tree_add_190_195_groupi_n_919);
  xnor csa_tree_add_190_195_groupi_g45098(csa_tree_add_190_195_groupi_n_4048 ,csa_tree_add_190_195_groupi_n_970 ,csa_tree_add_190_195_groupi_n_1592);
  xnor csa_tree_add_190_195_groupi_g45099(csa_tree_add_190_195_groupi_n_4047 ,csa_tree_add_190_195_groupi_n_1607 ,csa_tree_add_190_195_groupi_n_1950);
  xnor csa_tree_add_190_195_groupi_g45100(csa_tree_add_190_195_groupi_n_4046 ,csa_tree_add_190_195_groupi_n_1976 ,csa_tree_add_190_195_groupi_n_1693);
  xnor csa_tree_add_190_195_groupi_g45101(csa_tree_add_190_195_groupi_n_4045 ,csa_tree_add_190_195_groupi_n_2156 ,csa_tree_add_190_195_groupi_n_2082);
  xnor csa_tree_add_190_195_groupi_g45102(csa_tree_add_190_195_groupi_n_4044 ,csa_tree_add_190_195_groupi_n_2050 ,csa_tree_add_190_195_groupi_n_1977);
  xnor csa_tree_add_190_195_groupi_g45103(csa_tree_add_190_195_groupi_n_4043 ,csa_tree_add_190_195_groupi_n_1869 ,csa_tree_add_190_195_groupi_n_2058);
  xnor csa_tree_add_190_195_groupi_g45104(csa_tree_add_190_195_groupi_n_4042 ,csa_tree_add_190_195_groupi_n_616 ,csa_tree_add_190_195_groupi_n_1119);
  xnor csa_tree_add_190_195_groupi_g45105(csa_tree_add_190_195_groupi_n_4041 ,csa_tree_add_190_195_groupi_n_2040 ,csa_tree_add_190_195_groupi_n_1924);
  xnor csa_tree_add_190_195_groupi_g45106(csa_tree_add_190_195_groupi_n_4040 ,csa_tree_add_190_195_groupi_n_486 ,csa_tree_add_190_195_groupi_n_2060);
  xnor csa_tree_add_190_195_groupi_g45107(csa_tree_add_190_195_groupi_n_4039 ,csa_tree_add_190_195_groupi_n_508 ,csa_tree_add_190_195_groupi_n_973);
  xnor csa_tree_add_190_195_groupi_g45108(csa_tree_add_190_195_groupi_n_4038 ,csa_tree_add_190_195_groupi_n_1095 ,csa_tree_add_190_195_groupi_n_1872);
  xnor csa_tree_add_190_195_groupi_g45109(csa_tree_add_190_195_groupi_n_4037 ,csa_tree_add_190_195_groupi_n_1836 ,csa_tree_add_190_195_groupi_n_1935);
  xnor csa_tree_add_190_195_groupi_g45111(csa_tree_add_190_195_groupi_n_4036 ,csa_tree_add_190_195_groupi_n_1928 ,csa_tree_add_190_195_groupi_n_1850);
  xnor csa_tree_add_190_195_groupi_g45112(csa_tree_add_190_195_groupi_n_4035 ,csa_tree_add_190_195_groupi_n_2055 ,csa_tree_add_190_195_groupi_n_1757);
  xnor csa_tree_add_190_195_groupi_g45113(csa_tree_add_190_195_groupi_n_4034 ,csa_tree_add_190_195_groupi_n_2082 ,csa_tree_add_190_195_groupi_n_1630);
  xnor csa_tree_add_190_195_groupi_g45114(csa_tree_add_190_195_groupi_n_4033 ,csa_tree_add_190_195_groupi_n_1780 ,csa_tree_add_190_195_groupi_n_1777);
  xnor csa_tree_add_190_195_groupi_g45115(csa_tree_add_190_195_groupi_n_4032 ,csa_tree_add_190_195_groupi_n_2214 ,csa_tree_add_190_195_groupi_n_1949);
  xnor csa_tree_add_190_195_groupi_g45116(csa_tree_add_190_195_groupi_n_4031 ,csa_tree_add_190_195_groupi_n_423 ,csa_tree_add_190_195_groupi_n_1606);
  xnor csa_tree_add_190_195_groupi_g45117(csa_tree_add_190_195_groupi_n_4030 ,csa_tree_add_190_195_groupi_n_305 ,csa_tree_add_190_195_groupi_n_1003);
  xnor csa_tree_add_190_195_groupi_g45118(csa_tree_add_190_195_groupi_n_4029 ,csa_tree_add_190_195_groupi_n_1674 ,csa_tree_add_190_195_groupi_n_760);
  xnor csa_tree_add_190_195_groupi_g45119(csa_tree_add_190_195_groupi_n_4028 ,csa_tree_add_190_195_groupi_n_1975 ,csa_tree_add_190_195_groupi_n_1692);
  xnor csa_tree_add_190_195_groupi_g45120(csa_tree_add_190_195_groupi_n_4027 ,csa_tree_add_190_195_groupi_n_609 ,csa_tree_add_190_195_groupi_n_1902);
  xnor csa_tree_add_190_195_groupi_g45121(csa_tree_add_190_195_groupi_n_4026 ,in58[14] ,in59[14]);
  xnor csa_tree_add_190_195_groupi_g45123(csa_tree_add_190_195_groupi_n_4025 ,csa_tree_add_190_195_groupi_n_366 ,csa_tree_add_190_195_groupi_n_1888);
  xnor csa_tree_add_190_195_groupi_g45124(csa_tree_add_190_195_groupi_n_4024 ,csa_tree_add_190_195_groupi_n_1020 ,csa_tree_add_190_195_groupi_n_1703);
  xnor csa_tree_add_190_195_groupi_g45125(csa_tree_add_190_195_groupi_n_4023 ,csa_tree_add_190_195_groupi_n_202 ,csa_tree_add_190_195_groupi_n_1838);
  xnor csa_tree_add_190_195_groupi_g45126(csa_tree_add_190_195_groupi_n_4022 ,csa_tree_add_190_195_groupi_n_1995 ,csa_tree_add_190_195_groupi_n_1998);
  xnor csa_tree_add_190_195_groupi_g45127(csa_tree_add_190_195_groupi_n_4021 ,csa_tree_add_190_195_groupi_n_1996 ,csa_tree_add_190_195_groupi_n_1995);
  xnor csa_tree_add_190_195_groupi_g45128(csa_tree_add_190_195_groupi_n_4020 ,in55[4] ,in55[2]);
  xnor csa_tree_add_190_195_groupi_g45129(csa_tree_add_190_195_groupi_n_4019 ,csa_tree_add_190_195_groupi_n_334 ,csa_tree_add_190_195_groupi_n_1583);
  xnor csa_tree_add_190_195_groupi_g45130(csa_tree_add_190_195_groupi_n_4018 ,csa_tree_add_190_195_groupi_n_1021 ,csa_tree_add_190_195_groupi_n_1707);
  xnor csa_tree_add_190_195_groupi_g45131(csa_tree_add_190_195_groupi_n_4017 ,csa_tree_add_190_195_groupi_n_1116 ,csa_tree_add_190_195_groupi_n_1852);
  xnor csa_tree_add_190_195_groupi_g45132(csa_tree_add_190_195_groupi_n_4016 ,csa_tree_add_190_195_groupi_n_1924 ,csa_tree_add_190_195_groupi_n_1656);
  xnor csa_tree_add_190_195_groupi_g45133(csa_tree_add_190_195_groupi_n_4015 ,in55[7] ,in55[5]);
  xnor csa_tree_add_190_195_groupi_g45134(csa_tree_add_190_195_groupi_n_4014 ,csa_tree_add_190_195_groupi_n_1931 ,csa_tree_add_190_195_groupi_n_889);
  xnor csa_tree_add_190_195_groupi_g45135(csa_tree_add_190_195_groupi_n_4013 ,csa_tree_add_190_195_groupi_n_876 ,csa_tree_add_190_195_groupi_n_1720);
  xnor csa_tree_add_190_195_groupi_g45136(csa_tree_add_190_195_groupi_n_4012 ,csa_tree_add_190_195_groupi_n_877 ,csa_tree_add_190_195_groupi_n_862);
  xnor csa_tree_add_190_195_groupi_g45137(csa_tree_add_190_195_groupi_n_4011 ,csa_tree_add_190_195_groupi_n_347 ,csa_tree_add_190_195_groupi_n_2049);
  xnor csa_tree_add_190_195_groupi_g45138(csa_tree_add_190_195_groupi_n_4010 ,csa_tree_add_190_195_groupi_n_957 ,csa_tree_add_190_195_groupi_n_796);
  xnor csa_tree_add_190_195_groupi_g45139(csa_tree_add_190_195_groupi_n_4009 ,csa_tree_add_190_195_groupi_n_230 ,csa_tree_add_190_195_groupi_n_1069);
  xnor csa_tree_add_190_195_groupi_g45140(csa_tree_add_190_195_groupi_n_4008 ,csa_tree_add_190_195_groupi_n_1923 ,csa_tree_add_190_195_groupi_n_1635);
  xnor csa_tree_add_190_195_groupi_g45141(csa_tree_add_190_195_groupi_n_4007 ,csa_tree_add_190_195_groupi_n_1975 ,csa_tree_add_190_195_groupi_n_1776);
  xnor csa_tree_add_190_195_groupi_g45142(csa_tree_add_190_195_groupi_n_4006 ,csa_tree_add_190_195_groupi_n_355 ,csa_tree_add_190_195_groupi_n_1220);
  xnor csa_tree_add_190_195_groupi_g45143(csa_tree_add_190_195_groupi_n_4005 ,csa_tree_add_190_195_groupi_n_370 ,csa_tree_add_190_195_groupi_n_1149);
  xnor csa_tree_add_190_195_groupi_g45144(csa_tree_add_190_195_groupi_n_4004 ,csa_tree_add_190_195_groupi_n_751 ,csa_tree_add_190_195_groupi_n_1591);
  xnor csa_tree_add_190_195_groupi_g45145(csa_tree_add_190_195_groupi_n_4003 ,csa_tree_add_190_195_groupi_n_1942 ,csa_tree_add_190_195_groupi_n_1852);
  xnor csa_tree_add_190_195_groupi_g45146(csa_tree_add_190_195_groupi_n_4002 ,csa_tree_add_190_195_groupi_n_2118 ,csa_tree_add_190_195_groupi_n_1855);
  xnor csa_tree_add_190_195_groupi_g45147(csa_tree_add_190_195_groupi_n_4001 ,csa_tree_add_190_195_groupi_n_384 ,csa_tree_add_190_195_groupi_n_2061);
  xnor csa_tree_add_190_195_groupi_g45148(csa_tree_add_190_195_groupi_n_4000 ,csa_tree_add_190_195_groupi_n_1023 ,csa_tree_add_190_195_groupi_n_1860);
  xnor csa_tree_add_190_195_groupi_g45149(csa_tree_add_190_195_groupi_n_3999 ,csa_tree_add_190_195_groupi_n_1674 ,csa_tree_add_190_195_groupi_n_810);
  xnor csa_tree_add_190_195_groupi_g45150(csa_tree_add_190_195_groupi_n_3998 ,csa_tree_add_190_195_groupi_n_526 ,csa_tree_add_190_195_groupi_n_2058);
  xnor csa_tree_add_190_195_groupi_g45151(csa_tree_add_190_195_groupi_n_3997 ,csa_tree_add_190_195_groupi_n_2152 ,csa_tree_add_190_195_groupi_n_2039);
  xnor csa_tree_add_190_195_groupi_g45152(csa_tree_add_190_195_groupi_n_3996 ,in55[2] ,in57[5]);
  xnor csa_tree_add_190_195_groupi_g45153(csa_tree_add_190_195_groupi_n_3995 ,csa_tree_add_190_195_groupi_n_1936 ,csa_tree_add_190_195_groupi_n_1989);
  xnor csa_tree_add_190_195_groupi_g45154(csa_tree_add_190_195_groupi_n_3994 ,csa_tree_add_190_195_groupi_n_993 ,csa_tree_add_190_195_groupi_n_1851);
  xnor csa_tree_add_190_195_groupi_g45155(csa_tree_add_190_195_groupi_n_3993 ,csa_tree_add_190_195_groupi_n_1921 ,csa_tree_add_190_195_groupi_n_2039);
  xnor csa_tree_add_190_195_groupi_g45156(csa_tree_add_190_195_groupi_n_3992 ,csa_tree_add_190_195_groupi_n_475 ,csa_tree_add_190_195_groupi_n_1989);
  xnor csa_tree_add_190_195_groupi_g45157(csa_tree_add_190_195_groupi_n_3991 ,in55[4] ,in57[7]);
  xnor csa_tree_add_190_195_groupi_g45158(csa_tree_add_190_195_groupi_n_3990 ,csa_tree_add_190_195_groupi_n_1823 ,csa_tree_add_190_195_groupi_n_1910);
  xnor csa_tree_add_190_195_groupi_g45159(csa_tree_add_190_195_groupi_n_3989 ,in58[12] ,in59[12]);
  xnor csa_tree_add_190_195_groupi_g45160(csa_tree_add_190_195_groupi_n_3988 ,in55[8] ,in55[3]);
  xnor csa_tree_add_190_195_groupi_g45161(csa_tree_add_190_195_groupi_n_3987 ,csa_tree_add_190_195_groupi_n_1823 ,csa_tree_add_190_195_groupi_n_1821);
  xnor csa_tree_add_190_195_groupi_g45162(csa_tree_add_190_195_groupi_n_3986 ,csa_tree_add_190_195_groupi_n_951 ,csa_tree_add_190_195_groupi_n_1826);
  xnor csa_tree_add_190_195_groupi_g45163(csa_tree_add_190_195_groupi_n_3985 ,in58[5] ,in56[5]);
  xnor csa_tree_add_190_195_groupi_g45164(csa_tree_add_190_195_groupi_n_3984 ,in55[15] ,in55[11]);
  xnor csa_tree_add_190_195_groupi_g45165(csa_tree_add_190_195_groupi_n_3983 ,csa_tree_add_190_195_groupi_n_1113 ,csa_tree_add_190_195_groupi_n_1691);
  xnor csa_tree_add_190_195_groupi_g45166(csa_tree_add_190_195_groupi_n_3982 ,csa_tree_add_190_195_groupi_n_2213 ,csa_tree_add_190_195_groupi_n_2089);
  xnor csa_tree_add_190_195_groupi_g45167(csa_tree_add_190_195_groupi_n_3981 ,csa_tree_add_190_195_groupi_n_2214 ,csa_tree_add_190_195_groupi_n_1655);
  xnor csa_tree_add_190_195_groupi_g45168(csa_tree_add_190_195_groupi_n_3980 ,csa_tree_add_190_195_groupi_n_897 ,csa_tree_add_190_195_groupi_n_2212);
  xnor csa_tree_add_190_195_groupi_g45169(csa_tree_add_190_195_groupi_n_3979 ,csa_tree_add_190_195_groupi_n_1906 ,csa_tree_add_190_195_groupi_n_2116);
  xnor csa_tree_add_190_195_groupi_g45170(csa_tree_add_190_195_groupi_n_3978 ,csa_tree_add_190_195_groupi_n_502 ,csa_tree_add_190_195_groupi_n_1767);
  xnor csa_tree_add_190_195_groupi_g45171(csa_tree_add_190_195_groupi_n_3977 ,csa_tree_add_190_195_groupi_n_1826 ,csa_tree_add_190_195_groupi_n_1701);
  xnor csa_tree_add_190_195_groupi_g45172(csa_tree_add_190_195_groupi_n_3976 ,csa_tree_add_190_195_groupi_n_1283 ,csa_tree_add_190_195_groupi_n_1644);
  xnor csa_tree_add_190_195_groupi_g45173(csa_tree_add_190_195_groupi_n_3975 ,csa_tree_add_190_195_groupi_n_1951 ,csa_tree_add_190_195_groupi_n_1895);
  xnor csa_tree_add_190_195_groupi_g45174(csa_tree_add_190_195_groupi_n_3974 ,csa_tree_add_190_195_groupi_n_1877 ,in59[1]);
  xnor csa_tree_add_190_195_groupi_g45175(csa_tree_add_190_195_groupi_n_3973 ,csa_tree_add_190_195_groupi_n_283 ,csa_tree_add_190_195_groupi_n_1602);
  xnor csa_tree_add_190_195_groupi_g45176(csa_tree_add_190_195_groupi_n_3972 ,csa_tree_add_190_195_groupi_n_216 ,csa_tree_add_190_195_groupi_n_1949);
  xnor csa_tree_add_190_195_groupi_g45177(csa_tree_add_190_195_groupi_n_3971 ,csa_tree_add_190_195_groupi_n_293 ,csa_tree_add_190_195_groupi_n_1815);
  xnor csa_tree_add_190_195_groupi_g45178(csa_tree_add_190_195_groupi_n_3970 ,csa_tree_add_190_195_groupi_n_1971 ,csa_tree_add_190_195_groupi_n_1817);
  xnor csa_tree_add_190_195_groupi_g45179(csa_tree_add_190_195_groupi_n_3969 ,csa_tree_add_190_195_groupi_n_533 ,csa_tree_add_190_195_groupi_n_2216);
  xnor csa_tree_add_190_195_groupi_g45180(csa_tree_add_190_195_groupi_n_3968 ,csa_tree_add_190_195_groupi_n_1988 ,csa_tree_add_190_195_groupi_n_1933);
  xnor csa_tree_add_190_195_groupi_g45181(csa_tree_add_190_195_groupi_n_3967 ,csa_tree_add_190_195_groupi_n_907 ,csa_tree_add_190_195_groupi_n_1672);
  xnor csa_tree_add_190_195_groupi_g45182(csa_tree_add_190_195_groupi_n_3966 ,csa_tree_add_190_195_groupi_n_1909 ,csa_tree_add_190_195_groupi_n_1696);
  xnor csa_tree_add_190_195_groupi_g45183(csa_tree_add_190_195_groupi_n_3965 ,csa_tree_add_190_195_groupi_n_862 ,csa_tree_add_190_195_groupi_n_1580);
  xnor csa_tree_add_190_195_groupi_g45184(csa_tree_add_190_195_groupi_n_3964 ,csa_tree_add_190_195_groupi_n_1843 ,csa_tree_add_190_195_groupi_n_1650);
  xnor csa_tree_add_190_195_groupi_g45185(csa_tree_add_190_195_groupi_n_3963 ,csa_tree_add_190_195_groupi_n_843 ,csa_tree_add_190_195_groupi_n_1586);
  xnor csa_tree_add_190_195_groupi_g45186(csa_tree_add_190_195_groupi_n_3962 ,csa_tree_add_190_195_groupi_n_1863 ,csa_tree_add_190_195_groupi_n_1633);
  xnor csa_tree_add_190_195_groupi_g45187(csa_tree_add_190_195_groupi_n_3961 ,csa_tree_add_190_195_groupi_n_1991 ,csa_tree_add_190_195_groupi_n_1699);
  xnor csa_tree_add_190_195_groupi_g45188(csa_tree_add_190_195_groupi_n_3960 ,csa_tree_add_190_195_groupi_n_1708 ,csa_tree_add_190_195_groupi_n_1937);
  xnor csa_tree_add_190_195_groupi_g45189(csa_tree_add_190_195_groupi_n_3959 ,csa_tree_add_190_195_groupi_n_912 ,csa_tree_add_190_195_groupi_n_1637);
  xnor csa_tree_add_190_195_groupi_g45190(csa_tree_add_190_195_groupi_n_3958 ,csa_tree_add_190_195_groupi_n_858 ,csa_tree_add_190_195_groupi_n_794);
  xnor csa_tree_add_190_195_groupi_g45191(csa_tree_add_190_195_groupi_n_3957 ,csa_tree_add_190_195_groupi_n_477 ,csa_tree_add_190_195_groupi_n_967);
  xnor csa_tree_add_190_195_groupi_g45192(csa_tree_add_190_195_groupi_n_3956 ,csa_tree_add_190_195_groupi_n_855 ,csa_tree_add_190_195_groupi_n_1602);
  xnor csa_tree_add_190_195_groupi_g45193(csa_tree_add_190_195_groupi_n_3955 ,csa_tree_add_190_195_groupi_n_2154 ,csa_tree_add_190_195_groupi_n_2087);
  xnor csa_tree_add_190_195_groupi_g45194(csa_tree_add_190_195_groupi_n_3954 ,csa_tree_add_190_195_groupi_n_1818 ,csa_tree_add_190_195_groupi_n_1757);
  xnor csa_tree_add_190_195_groupi_g45195(csa_tree_add_190_195_groupi_n_3953 ,csa_tree_add_190_195_groupi_n_996 ,csa_tree_add_190_195_groupi_n_1080);
  xnor csa_tree_add_190_195_groupi_g45196(csa_tree_add_190_195_groupi_n_3952 ,csa_tree_add_190_195_groupi_n_937 ,csa_tree_add_190_195_groupi_n_1779);
  xnor csa_tree_add_190_195_groupi_g45197(csa_tree_add_190_195_groupi_n_3951 ,csa_tree_add_190_195_groupi_n_903 ,csa_tree_add_190_195_groupi_n_927);
  xnor csa_tree_add_190_195_groupi_g45198(csa_tree_add_190_195_groupi_n_3950 ,csa_tree_add_190_195_groupi_n_1922 ,csa_tree_add_190_195_groupi_n_1632);
  xnor csa_tree_add_190_195_groupi_g45199(csa_tree_add_190_195_groupi_n_3949 ,in55[6] ,in55[1]);
  xnor csa_tree_add_190_195_groupi_g45200(csa_tree_add_190_195_groupi_n_3948 ,csa_tree_add_190_195_groupi_n_213 ,csa_tree_add_190_195_groupi_n_1905);
  xnor csa_tree_add_190_195_groupi_g45201(csa_tree_add_190_195_groupi_n_3947 ,csa_tree_add_190_195_groupi_n_350 ,csa_tree_add_190_195_groupi_n_883);
  xnor csa_tree_add_190_195_groupi_g45202(csa_tree_add_190_195_groupi_n_3946 ,csa_tree_add_190_195_groupi_n_261 ,csa_tree_add_190_195_groupi_n_1873);
  xnor csa_tree_add_190_195_groupi_g45203(csa_tree_add_190_195_groupi_n_3945 ,csa_tree_add_190_195_groupi_n_1978 ,csa_tree_add_190_195_groupi_n_1834);
  xnor csa_tree_add_190_195_groupi_g45204(csa_tree_add_190_195_groupi_n_3944 ,csa_tree_add_190_195_groupi_n_1864 ,csa_tree_add_190_195_groupi_n_2056);
  xnor csa_tree_add_190_195_groupi_g45205(csa_tree_add_190_195_groupi_n_3943 ,csa_tree_add_190_195_groupi_n_394 ,csa_tree_add_190_195_groupi_n_1994);
  xnor csa_tree_add_190_195_groupi_g45206(csa_tree_add_190_195_groupi_n_3942 ,csa_tree_add_190_195_groupi_n_1871 ,csa_tree_add_190_195_groupi_n_1816);
  xnor csa_tree_add_190_195_groupi_g45207(csa_tree_add_190_195_groupi_n_3941 ,csa_tree_add_190_195_groupi_n_328 ,csa_tree_add_190_195_groupi_n_940);
  xnor csa_tree_add_190_195_groupi_g45208(csa_tree_add_190_195_groupi_n_3940 ,csa_tree_add_190_195_groupi_n_2158 ,csa_tree_add_190_195_groupi_n_2155);
  xnor csa_tree_add_190_195_groupi_g45209(csa_tree_add_190_195_groupi_n_3939 ,csa_tree_add_190_195_groupi_n_1921 ,csa_tree_add_190_195_groupi_n_1841);
  xnor csa_tree_add_190_195_groupi_g45210(csa_tree_add_190_195_groupi_n_3938 ,csa_tree_add_190_195_groupi_n_1907 ,csa_tree_add_190_195_groupi_n_2059);
  xnor csa_tree_add_190_195_groupi_g45212(csa_tree_add_190_195_groupi_n_3937 ,csa_tree_add_190_195_groupi_n_601 ,csa_tree_add_190_195_groupi_n_1054);
  xnor csa_tree_add_190_195_groupi_g45213(csa_tree_add_190_195_groupi_n_3936 ,csa_tree_add_190_195_groupi_n_2216 ,csa_tree_add_190_195_groupi_n_1861);
  xnor csa_tree_add_190_195_groupi_g45215(csa_tree_add_190_195_groupi_n_3935 ,csa_tree_add_190_195_groupi_n_777 ,csa_tree_add_190_195_groupi_n_907);
  xnor csa_tree_add_190_195_groupi_g45216(csa_tree_add_190_195_groupi_n_3934 ,csa_tree_add_190_195_groupi_n_600 ,csa_tree_add_190_195_groupi_n_1111);
  xnor csa_tree_add_190_195_groupi_g45217(csa_tree_add_190_195_groupi_n_3933 ,csa_tree_add_190_195_groupi_n_550 ,csa_tree_add_190_195_groupi_n_1748);
  xnor csa_tree_add_190_195_groupi_g45218(csa_tree_add_190_195_groupi_n_3932 ,csa_tree_add_190_195_groupi_n_309 ,in55[0]);
  xnor csa_tree_add_190_195_groupi_g45219(csa_tree_add_190_195_groupi_n_3931 ,csa_tree_add_190_195_groupi_n_224 ,csa_tree_add_190_195_groupi_n_1164);
  xnor csa_tree_add_190_195_groupi_g45220(csa_tree_add_190_195_groupi_n_3930 ,csa_tree_add_190_195_groupi_n_417 ,csa_tree_add_190_195_groupi_n_1934);
  xnor csa_tree_add_190_195_groupi_g45221(csa_tree_add_190_195_groupi_n_3929 ,csa_tree_add_190_195_groupi_n_237 ,csa_tree_add_190_195_groupi_n_812);
  xnor csa_tree_add_190_195_groupi_g45222(csa_tree_add_190_195_groupi_n_3928 ,csa_tree_add_190_195_groupi_n_595 ,csa_tree_add_190_195_groupi_n_1821);
  xnor csa_tree_add_190_195_groupi_g45224(csa_tree_add_190_195_groupi_n_3927 ,csa_tree_add_190_195_groupi_n_224 ,csa_tree_add_190_195_groupi_n_1202);
  xnor csa_tree_add_190_195_groupi_g45225(csa_tree_add_190_195_groupi_n_3926 ,csa_tree_add_190_195_groupi_n_353 ,csa_tree_add_190_195_groupi_n_1098);
  xnor csa_tree_add_190_195_groupi_g45226(csa_tree_add_190_195_groupi_n_3925 ,csa_tree_add_190_195_groupi_n_273 ,csa_tree_add_190_195_groupi_n_1126);
  xnor csa_tree_add_190_195_groupi_g45227(csa_tree_add_190_195_groupi_n_3924 ,csa_tree_add_190_195_groupi_n_594 ,csa_tree_add_190_195_groupi_n_1820);
  xnor csa_tree_add_190_195_groupi_g45228(csa_tree_add_190_195_groupi_n_3923 ,csa_tree_add_190_195_groupi_n_594 ,csa_tree_add_190_195_groupi_n_1700);
  xnor csa_tree_add_190_195_groupi_g45229(csa_tree_add_190_195_groupi_n_3922 ,csa_tree_add_190_195_groupi_n_465 ,csa_tree_add_190_195_groupi_n_2212);
  xnor csa_tree_add_190_195_groupi_g45230(csa_tree_add_190_195_groupi_n_3921 ,csa_tree_add_190_195_groupi_n_470 ,csa_tree_add_190_195_groupi_n_1752);
  xnor csa_tree_add_190_195_groupi_g45231(csa_tree_add_190_195_groupi_n_3920 ,csa_tree_add_190_195_groupi_n_259 ,csa_tree_add_190_195_groupi_n_1930);
  xnor csa_tree_add_190_195_groupi_g45232(csa_tree_add_190_195_groupi_n_3919 ,csa_tree_add_190_195_groupi_n_579 ,csa_tree_add_190_195_groupi_n_1761);
  xnor csa_tree_add_190_195_groupi_g45233(csa_tree_add_190_195_groupi_n_3918 ,csa_tree_add_190_195_groupi_n_499 ,csa_tree_add_190_195_groupi_n_1870);
  xnor csa_tree_add_190_195_groupi_g45234(csa_tree_add_190_195_groupi_n_3917 ,csa_tree_add_190_195_groupi_n_240 ,csa_tree_add_190_195_groupi_n_1826);
  xnor csa_tree_add_190_195_groupi_g45235(csa_tree_add_190_195_groupi_n_3916 ,csa_tree_add_190_195_groupi_n_535 ,csa_tree_add_190_195_groupi_n_1932);
  xnor csa_tree_add_190_195_groupi_g45236(csa_tree_add_190_195_groupi_n_3915 ,csa_tree_add_190_195_groupi_n_342 ,csa_tree_add_190_195_groupi_n_2157);
  xnor csa_tree_add_190_195_groupi_g45237(csa_tree_add_190_195_groupi_n_3914 ,csa_tree_add_190_195_groupi_n_366 ,csa_tree_add_190_195_groupi_n_1708);
  xnor csa_tree_add_190_195_groupi_g45238(csa_tree_add_190_195_groupi_n_3913 ,csa_tree_add_190_195_groupi_n_1107 ,csa_tree_add_190_195_groupi_n_1682);
  xnor csa_tree_add_190_195_groupi_g45239(csa_tree_add_190_195_groupi_n_3912 ,csa_tree_add_190_195_groupi_n_330 ,csa_tree_add_190_195_groupi_n_2051);
  xnor csa_tree_add_190_195_groupi_g45240(csa_tree_add_190_195_groupi_n_3911 ,csa_tree_add_190_195_groupi_n_391 ,csa_tree_add_190_195_groupi_n_1764);
  xnor csa_tree_add_190_195_groupi_g45241(csa_tree_add_190_195_groupi_n_3910 ,csa_tree_add_190_195_groupi_n_247 ,csa_tree_add_190_195_groupi_n_1277);
  xnor csa_tree_add_190_195_groupi_g45243(csa_tree_add_190_195_groupi_n_3909 ,csa_tree_add_190_195_groupi_n_606 ,csa_tree_add_190_195_groupi_n_1896);
  xnor csa_tree_add_190_195_groupi_g45244(csa_tree_add_190_195_groupi_n_3908 ,csa_tree_add_190_195_groupi_n_552 ,csa_tree_add_190_195_groupi_n_1776);
  xnor csa_tree_add_190_195_groupi_g45245(csa_tree_add_190_195_groupi_n_3907 ,csa_tree_add_190_195_groupi_n_612 ,csa_tree_add_190_195_groupi_n_1894);
  xnor csa_tree_add_190_195_groupi_g45246(csa_tree_add_190_195_groupi_n_3906 ,csa_tree_add_190_195_groupi_n_301 ,csa_tree_add_190_195_groupi_n_1747);
  xnor csa_tree_add_190_195_groupi_g45247(csa_tree_add_190_195_groupi_n_3905 ,csa_tree_add_190_195_groupi_n_377 ,csa_tree_add_190_195_groupi_n_2059);
  xnor csa_tree_add_190_195_groupi_g45248(csa_tree_add_190_195_groupi_n_3904 ,csa_tree_add_190_195_groupi_n_283 ,csa_tree_add_190_195_groupi_n_1303);
  xnor csa_tree_add_190_195_groupi_g45249(csa_tree_add_190_195_groupi_n_3903 ,csa_tree_add_190_195_groupi_n_312 ,csa_tree_add_190_195_groupi_n_1964);
  xnor csa_tree_add_190_195_groupi_g45251(csa_tree_add_190_195_groupi_n_3902 ,csa_tree_add_190_195_groupi_n_446 ,csa_tree_add_190_195_groupi_n_1962);
  xnor csa_tree_add_190_195_groupi_g45252(csa_tree_add_190_195_groupi_n_3901 ,csa_tree_add_190_195_groupi_n_247 ,csa_tree_add_190_195_groupi_n_1969);
  xnor csa_tree_add_190_195_groupi_g45254(csa_tree_add_190_195_groupi_n_3900 ,csa_tree_add_190_195_groupi_n_613 ,csa_tree_add_190_195_groupi_n_2090);
  xnor csa_tree_add_190_195_groupi_g45255(csa_tree_add_190_195_groupi_n_3899 ,csa_tree_add_190_195_groupi_n_309 ,csa_tree_add_190_195_groupi_n_1621);
  xnor csa_tree_add_190_195_groupi_g45256(csa_tree_add_190_195_groupi_n_3898 ,csa_tree_add_190_195_groupi_n_401 ,csa_tree_add_190_195_groupi_n_2119);
  xnor csa_tree_add_190_195_groupi_g45257(csa_tree_add_190_195_groupi_n_3897 ,csa_tree_add_190_195_groupi_n_403 ,csa_tree_add_190_195_groupi_n_1275);
  xnor csa_tree_add_190_195_groupi_g45258(csa_tree_add_190_195_groupi_n_3896 ,csa_tree_add_190_195_groupi_n_544 ,csa_tree_add_190_195_groupi_n_996);
  xnor csa_tree_add_190_195_groupi_g45259(csa_tree_add_190_195_groupi_n_3895 ,csa_tree_add_190_195_groupi_n_449 ,csa_tree_add_190_195_groupi_n_625);
  xnor csa_tree_add_190_195_groupi_g45260(csa_tree_add_190_195_groupi_n_3894 ,csa_tree_add_190_195_groupi_n_312 ,csa_tree_add_190_195_groupi_n_1977);
  xnor csa_tree_add_190_195_groupi_g45261(csa_tree_add_190_195_groupi_n_3893 ,csa_tree_add_190_195_groupi_n_336 ,csa_tree_add_190_195_groupi_n_1877);
  xnor csa_tree_add_190_195_groupi_g45262(csa_tree_add_190_195_groupi_n_3892 ,csa_tree_add_190_195_groupi_n_618 ,csa_tree_add_190_195_groupi_n_2004);
  xnor csa_tree_add_190_195_groupi_g45263(csa_tree_add_190_195_groupi_n_3891 ,csa_tree_add_190_195_groupi_n_325 ,csa_tree_add_190_195_groupi_n_1612);
  xnor csa_tree_add_190_195_groupi_g45264(csa_tree_add_190_195_groupi_n_3890 ,csa_tree_add_190_195_groupi_n_603 ,csa_tree_add_190_195_groupi_n_1102);
  xnor csa_tree_add_190_195_groupi_g45265(csa_tree_add_190_195_groupi_n_3889 ,csa_tree_add_190_195_groupi_n_1222 ,csa_tree_add_190_195_groupi_n_1594);
  xnor csa_tree_add_190_195_groupi_g45266(csa_tree_add_190_195_groupi_n_3888 ,csa_tree_add_190_195_groupi_n_504 ,csa_tree_add_190_195_groupi_n_1836);
  xnor csa_tree_add_190_195_groupi_g45268(csa_tree_add_190_195_groupi_n_3887 ,csa_tree_add_190_195_groupi_n_266 ,csa_tree_add_190_195_groupi_n_1291);
  xnor csa_tree_add_190_195_groupi_g45269(csa_tree_add_190_195_groupi_n_3886 ,csa_tree_add_190_195_groupi_n_577 ,csa_tree_add_190_195_groupi_n_1113);
  xnor csa_tree_add_190_195_groupi_g45270(csa_tree_add_190_195_groupi_n_3885 ,csa_tree_add_190_195_groupi_n_615 ,csa_tree_add_190_195_groupi_n_1774);
  xnor csa_tree_add_190_195_groupi_g45271(csa_tree_add_190_195_groupi_n_3884 ,csa_tree_add_190_195_groupi_n_572 ,csa_tree_add_190_195_groupi_n_2086);
  xnor csa_tree_add_190_195_groupi_g45272(csa_tree_add_190_195_groupi_n_3883 ,csa_tree_add_190_195_groupi_n_566 ,csa_tree_add_190_195_groupi_n_1647);
  xnor csa_tree_add_190_195_groupi_g45273(csa_tree_add_190_195_groupi_n_3882 ,csa_tree_add_190_195_groupi_n_451 ,csa_tree_add_190_195_groupi_n_2088);
  xnor csa_tree_add_190_195_groupi_g45274(csa_tree_add_190_195_groupi_n_3881 ,csa_tree_add_190_195_groupi_n_493 ,csa_tree_add_190_195_groupi_n_1974);
  xnor csa_tree_add_190_195_groupi_g45275(csa_tree_add_190_195_groupi_n_3880 ,csa_tree_add_190_195_groupi_n_895 ,csa_tree_add_190_195_groupi_n_491);
  xnor csa_tree_add_190_195_groupi_g45276(csa_tree_add_190_195_groupi_n_3879 ,csa_tree_add_190_195_groupi_n_516 ,csa_tree_add_190_195_groupi_n_1906);
  xnor csa_tree_add_190_195_groupi_g45277(csa_tree_add_190_195_groupi_n_3878 ,csa_tree_add_190_195_groupi_n_340 ,csa_tree_add_190_195_groupi_n_1963);
  xnor csa_tree_add_190_195_groupi_g45278(csa_tree_add_190_195_groupi_n_3877 ,csa_tree_add_190_195_groupi_n_264 ,csa_tree_add_190_195_groupi_n_1637);
  xnor csa_tree_add_190_195_groupi_g45279(csa_tree_add_190_195_groupi_n_3876 ,csa_tree_add_190_195_groupi_n_436 ,in55[0]);
  xnor csa_tree_add_190_195_groupi_g45281(csa_tree_add_190_195_groupi_n_3875 ,csa_tree_add_190_195_groupi_n_334 ,csa_tree_add_190_195_groupi_n_997);
  xnor csa_tree_add_190_195_groupi_g45282(csa_tree_add_190_195_groupi_n_3874 ,csa_tree_add_190_195_groupi_n_519 ,in58[2]);
  xnor csa_tree_add_190_195_groupi_g45283(csa_tree_add_190_195_groupi_n_3873 ,csa_tree_add_190_195_groupi_n_598 ,csa_tree_add_190_195_groupi_n_1646);
  xnor csa_tree_add_190_195_groupi_g45284(csa_tree_add_190_195_groupi_n_3872 ,csa_tree_add_190_195_groupi_n_368 ,csa_tree_add_190_195_groupi_n_1259);
  xnor csa_tree_add_190_195_groupi_g45285(csa_tree_add_190_195_groupi_n_3871 ,csa_tree_add_190_195_groupi_n_248 ,csa_tree_add_190_195_groupi_n_1844);
  xnor csa_tree_add_190_195_groupi_g45286(csa_tree_add_190_195_groupi_n_3870 ,csa_tree_add_190_195_groupi_n_597 ,csa_tree_add_190_195_groupi_n_1649);
  xnor csa_tree_add_190_195_groupi_g45288(csa_tree_add_190_195_groupi_n_3869 ,csa_tree_add_190_195_groupi_n_291 ,csa_tree_add_190_195_groupi_n_1756);
  xnor csa_tree_add_190_195_groupi_g45289(csa_tree_add_190_195_groupi_n_3868 ,csa_tree_add_190_195_groupi_n_409 ,csa_tree_add_190_195_groupi_n_1692);
  xnor csa_tree_add_190_195_groupi_g45290(csa_tree_add_190_195_groupi_n_3867 ,csa_tree_add_190_195_groupi_n_409 ,csa_tree_add_190_195_groupi_n_1969);
  xnor csa_tree_add_190_195_groupi_g45291(csa_tree_add_190_195_groupi_n_3866 ,csa_tree_add_190_195_groupi_n_382 ,csa_tree_add_190_195_groupi_n_1183);
  xnor csa_tree_add_190_195_groupi_g45292(csa_tree_add_190_195_groupi_n_3865 ,in55[11] ,in61[8]);
  xnor csa_tree_add_190_195_groupi_g45294(csa_tree_add_190_195_groupi_n_3864 ,csa_tree_add_190_195_groupi_n_276 ,in58[3]);
  xnor csa_tree_add_190_195_groupi_g45295(csa_tree_add_190_195_groupi_n_3863 ,csa_tree_add_190_195_groupi_n_252 ,csa_tree_add_190_195_groupi_n_1934);
  xnor csa_tree_add_190_195_groupi_g45296(csa_tree_add_190_195_groupi_n_3862 ,in55[12] ,in55[11]);
  xnor csa_tree_add_190_195_groupi_g45297(csa_tree_add_190_195_groupi_n_3861 ,csa_tree_add_190_195_groupi_n_229 ,csa_tree_add_190_195_groupi_n_1601);
  xnor csa_tree_add_190_195_groupi_g45298(csa_tree_add_190_195_groupi_n_3860 ,in55[7] ,in59[10]);
  xnor csa_tree_add_190_195_groupi_g45299(csa_tree_add_190_195_groupi_n_3859 ,csa_tree_add_190_195_groupi_n_231 ,csa_tree_add_190_195_groupi_n_1889);
  xnor csa_tree_add_190_195_groupi_g45300(csa_tree_add_190_195_groupi_n_3858 ,csa_tree_add_190_195_groupi_n_405 ,csa_tree_add_190_195_groupi_n_2152);
  xnor csa_tree_add_190_195_groupi_g45301(csa_tree_add_190_195_groupi_n_3857 ,csa_tree_add_190_195_groupi_n_1092 ,csa_tree_add_190_195_groupi_n_1753);
  xnor csa_tree_add_190_195_groupi_g45302(csa_tree_add_190_195_groupi_n_3856 ,csa_tree_add_190_195_groupi_n_355 ,csa_tree_add_190_195_groupi_n_1030);
  xnor csa_tree_add_190_195_groupi_g45303(csa_tree_add_190_195_groupi_n_3855 ,csa_tree_add_190_195_groupi_n_1285 ,csa_tree_add_190_195_groupi_n_2212);
  xnor csa_tree_add_190_195_groupi_g45304(csa_tree_add_190_195_groupi_n_3854 ,csa_tree_add_190_195_groupi_n_461 ,csa_tree_add_190_195_groupi_n_2056);
  xnor csa_tree_add_190_195_groupi_g45305(csa_tree_add_190_195_groupi_n_3853 ,in55[0] ,in58[4]);
  xnor csa_tree_add_190_195_groupi_g45306(csa_tree_add_190_195_groupi_n_3852 ,csa_tree_add_190_195_groupi_n_276 ,csa_tree_add_190_195_groupi_n_1707);
  xnor csa_tree_add_190_195_groupi_g45308(csa_tree_add_190_195_groupi_n_3851 ,csa_tree_add_190_195_groupi_n_874 ,csa_tree_add_190_195_groupi_n_1920);
  xnor csa_tree_add_190_195_groupi_g45309(csa_tree_add_190_195_groupi_n_3850 ,csa_tree_add_190_195_groupi_n_231 ,csa_tree_add_190_195_groupi_n_1837);
  xnor csa_tree_add_190_195_groupi_g45310(csa_tree_add_190_195_groupi_n_3849 ,in55[2] ,in60[6]);
  xnor csa_tree_add_190_195_groupi_g45311(csa_tree_add_190_195_groupi_n_3848 ,in55[7] ,in60[11]);
  xnor csa_tree_add_190_195_groupi_g45312(csa_tree_add_190_195_groupi_n_3847 ,csa_tree_add_190_195_groupi_n_319 ,csa_tree_add_190_195_groupi_n_1764);
  xnor csa_tree_add_190_195_groupi_g45313(csa_tree_add_190_195_groupi_n_3846 ,csa_tree_add_190_195_groupi_n_1050 ,csa_tree_add_190_195_groupi_n_1092);
  xnor csa_tree_add_190_195_groupi_g45314(csa_tree_add_190_195_groupi_n_3845 ,in55[14] ,in61[11]);
  xnor csa_tree_add_190_195_groupi_g45315(csa_tree_add_190_195_groupi_n_3844 ,csa_tree_add_190_195_groupi_n_1468 ,csa_tree_add_190_195_groupi_n_1399);
  xnor csa_tree_add_190_195_groupi_g45316(csa_tree_add_190_195_groupi_n_3843 ,csa_tree_add_190_195_groupi_n_837 ,csa_tree_add_190_195_groupi_n_1743);
  xnor csa_tree_add_190_195_groupi_g45317(csa_tree_add_190_195_groupi_n_3842 ,in55[9] ,in61[6]);
  xnor csa_tree_add_190_195_groupi_g45318(csa_tree_add_190_195_groupi_n_3841 ,in55[14] ,in55[13]);
  xnor csa_tree_add_190_195_groupi_g45319(csa_tree_add_190_195_groupi_n_3840 ,in55[5] ,in60[9]);
  xnor csa_tree_add_190_195_groupi_g45320(csa_tree_add_190_195_groupi_n_3839 ,csa_tree_add_190_195_groupi_n_1044 ,csa_tree_add_190_195_groupi_n_1870);
  xnor csa_tree_add_190_195_groupi_g45321(csa_tree_add_190_195_groupi_n_3838 ,in55[6] ,in59[9]);
  xnor csa_tree_add_190_195_groupi_g45322(csa_tree_add_190_195_groupi_n_3837 ,csa_tree_add_190_195_groupi_n_1132 ,csa_tree_add_190_195_groupi_n_1140);
  xnor csa_tree_add_190_195_groupi_g45323(csa_tree_add_190_195_groupi_n_3836 ,in55[6] ,in60[10]);
  xnor csa_tree_add_190_195_groupi_g45324(csa_tree_add_190_195_groupi_n_3835 ,in55[5] ,in59[8]);
  xnor csa_tree_add_190_195_groupi_g45325(csa_tree_add_190_195_groupi_n_3834 ,in55[8] ,in59[11]);
  xnor csa_tree_add_190_195_groupi_g45326(csa_tree_add_190_195_groupi_n_3833 ,csa_tree_add_190_195_groupi_n_924 ,csa_tree_add_190_195_groupi_n_1818);
  xnor csa_tree_add_190_195_groupi_g45327(csa_tree_add_190_195_groupi_n_3832 ,csa_tree_add_190_195_groupi_n_1887 ,csa_tree_add_190_195_groupi_n_1709);
  xnor csa_tree_add_190_195_groupi_g45328(csa_tree_add_190_195_groupi_n_3831 ,in55[9] ,in61[13]);
  xnor csa_tree_add_190_195_groupi_g45329(csa_tree_add_190_195_groupi_n_3830 ,in55[8] ,in61[12]);
  xnor csa_tree_add_190_195_groupi_g45330(csa_tree_add_190_195_groupi_n_3829 ,in55[4] ,in60[8]);
  xnor csa_tree_add_190_195_groupi_g45331(csa_tree_add_190_195_groupi_n_3828 ,csa_tree_add_190_195_groupi_n_1044 ,csa_tree_add_190_195_groupi_n_2050);
  xnor csa_tree_add_190_195_groupi_g45332(csa_tree_add_190_195_groupi_n_3827 ,in55[12] ,in61[9]);
  xnor csa_tree_add_190_195_groupi_g45333(csa_tree_add_190_195_groupi_n_3826 ,in55[13] ,in61[10]);
  xnor csa_tree_add_190_195_groupi_g45334(csa_tree_add_190_195_groupi_n_3825 ,in55[3] ,in59[6]);
  xnor csa_tree_add_190_195_groupi_g45335(csa_tree_add_190_195_groupi_n_3824 ,csa_tree_add_190_195_groupi_n_2062 ,csa_tree_add_190_195_groupi_n_1999);
  xnor csa_tree_add_190_195_groupi_g45336(csa_tree_add_190_195_groupi_n_3823 ,csa_tree_add_190_195_groupi_n_1888 ,csa_tree_add_190_195_groupi_n_1833);
  xnor csa_tree_add_190_195_groupi_g45337(csa_tree_add_190_195_groupi_n_3822 ,csa_tree_add_190_195_groupi_n_870 ,csa_tree_add_190_195_groupi_n_1125);
  xnor csa_tree_add_190_195_groupi_g45338(csa_tree_add_190_195_groupi_n_3821 ,csa_tree_add_190_195_groupi_n_2435 ,csa_tree_add_190_195_groupi_n_1566);
  xnor csa_tree_add_190_195_groupi_g45339(csa_tree_add_190_195_groupi_n_3820 ,csa_tree_add_190_195_groupi_n_870 ,csa_tree_add_190_195_groupi_n_1695);
  xnor csa_tree_add_190_195_groupi_g45340(csa_tree_add_190_195_groupi_n_3819 ,csa_tree_add_190_195_groupi_n_207 ,csa_tree_add_190_195_groupi_n_1839);
  xnor csa_tree_add_190_195_groupi_g45341(csa_tree_add_190_195_groupi_n_3818 ,csa_tree_add_190_195_groupi_n_994 ,csa_tree_add_190_195_groupi_n_1813);
  xnor csa_tree_add_190_195_groupi_g45342(csa_tree_add_190_195_groupi_n_3817 ,csa_tree_add_190_195_groupi_n_2209 ,csa_tree_add_190_195_groupi_n_2215);
  xnor csa_tree_add_190_195_groupi_g45343(csa_tree_add_190_195_groupi_n_3816 ,csa_tree_add_190_195_groupi_n_930 ,csa_tree_add_190_195_groupi_n_1893);
  xnor csa_tree_add_190_195_groupi_g45344(csa_tree_add_190_195_groupi_n_3815 ,csa_tree_add_190_195_groupi_n_888 ,csa_tree_add_190_195_groupi_n_1206);
  xnor csa_tree_add_190_195_groupi_g45345(csa_tree_add_190_195_groupi_n_3814 ,csa_tree_add_190_195_groupi_n_194 ,csa_tree_add_190_195_groupi_n_2086);
  xnor csa_tree_add_190_195_groupi_g45346(csa_tree_add_190_195_groupi_n_3813 ,csa_tree_add_190_195_groupi_n_2083 ,csa_tree_add_190_195_groupi_n_1271);
  xnor csa_tree_add_190_195_groupi_g45347(csa_tree_add_190_195_groupi_n_3812 ,csa_tree_add_190_195_groupi_n_2211 ,csa_tree_add_190_195_groupi_n_2156);
  xnor csa_tree_add_190_195_groupi_g45348(csa_tree_add_190_195_groupi_n_3811 ,csa_tree_add_190_195_groupi_n_975 ,csa_tree_add_190_195_groupi_n_1987);
  xnor csa_tree_add_190_195_groupi_g45349(csa_tree_add_190_195_groupi_n_3810 ,csa_tree_add_190_195_groupi_n_954 ,csa_tree_add_190_195_groupi_n_775);
  xnor csa_tree_add_190_195_groupi_g45350(csa_tree_add_190_195_groupi_n_3809 ,csa_tree_add_190_195_groupi_n_1961 ,csa_tree_add_190_195_groupi_n_1945);
  xnor csa_tree_add_190_195_groupi_g45351(csa_tree_add_190_195_groupi_n_3808 ,csa_tree_add_190_195_groupi_n_955 ,csa_tree_add_190_195_groupi_n_856);
  xnor csa_tree_add_190_195_groupi_g45352(csa_tree_add_190_195_groupi_n_3807 ,csa_tree_add_190_195_groupi_n_975 ,csa_tree_add_190_195_groupi_n_1825);
  xnor csa_tree_add_190_195_groupi_g45353(csa_tree_add_190_195_groupi_n_3806 ,csa_tree_add_190_195_groupi_n_1976 ,csa_tree_add_190_195_groupi_n_1758);
  xnor csa_tree_add_190_195_groupi_g45354(csa_tree_add_190_195_groupi_n_3805 ,csa_tree_add_190_195_groupi_n_1138 ,csa_tree_add_190_195_groupi_n_1905);
  xnor csa_tree_add_190_195_groupi_g45355(csa_tree_add_190_195_groupi_n_3804 ,csa_tree_add_190_195_groupi_n_1212 ,csa_tree_add_190_195_groupi_n_2015);
  xnor csa_tree_add_190_195_groupi_g45356(csa_tree_add_190_195_groupi_n_3803 ,csa_tree_add_190_195_groupi_n_2062 ,csa_tree_add_190_195_groupi_n_2060);
  xnor csa_tree_add_190_195_groupi_g45357(csa_tree_add_190_195_groupi_n_3802 ,csa_tree_add_190_195_groupi_n_380 ,csa_tree_add_190_195_groupi_n_1690);
  xnor csa_tree_add_190_195_groupi_g45358(csa_tree_add_190_195_groupi_n_3801 ,csa_tree_add_190_195_groupi_n_254 ,csa_tree_add_190_195_groupi_n_1086);
  xnor csa_tree_add_190_195_groupi_g45359(csa_tree_add_190_195_groupi_n_3800 ,csa_tree_add_190_195_groupi_n_207 ,csa_tree_add_190_195_groupi_n_1898);
  xnor csa_tree_add_190_195_groupi_g45360(csa_tree_add_190_195_groupi_n_3799 ,csa_tree_add_190_195_groupi_n_1026 ,csa_tree_add_190_195_groupi_n_1863);
  xnor csa_tree_add_190_195_groupi_g45361(csa_tree_add_190_195_groupi_n_3798 ,csa_tree_add_190_195_groupi_n_1191 ,in56[2]);
  xnor csa_tree_add_190_195_groupi_g45362(csa_tree_add_190_195_groupi_n_3797 ,csa_tree_add_190_195_groupi_n_930 ,csa_tree_add_190_195_groupi_n_1834);
  xnor csa_tree_add_190_195_groupi_g45363(csa_tree_add_190_195_groupi_n_3796 ,csa_tree_add_190_195_groupi_n_2154 ,csa_tree_add_190_195_groupi_n_2005);
  xnor csa_tree_add_190_195_groupi_g45364(csa_tree_add_190_195_groupi_n_3795 ,csa_tree_add_190_195_groupi_n_199 ,csa_tree_add_190_195_groupi_n_1808);
  xnor csa_tree_add_190_195_groupi_g45365(csa_tree_add_190_195_groupi_n_3794 ,csa_tree_add_190_195_groupi_n_2157 ,csa_tree_add_190_195_groupi_n_850);
  xnor csa_tree_add_190_195_groupi_g45366(csa_tree_add_190_195_groupi_n_3793 ,csa_tree_add_190_195_groupi_n_216 ,csa_tree_add_190_195_groupi_n_1829);
  xnor csa_tree_add_190_195_groupi_g45367(csa_tree_add_190_195_groupi_n_3792 ,csa_tree_add_190_195_groupi_n_1011 ,csa_tree_add_190_195_groupi_n_1859);
  xnor csa_tree_add_190_195_groupi_g45368(csa_tree_add_190_195_groupi_n_3791 ,csa_tree_add_190_195_groupi_n_710 ,csa_tree_add_190_195_groupi_n_746);
  xnor csa_tree_add_190_195_groupi_g45369(csa_tree_add_190_195_groupi_n_3790 ,csa_tree_add_190_195_groupi_n_226 ,csa_tree_add_190_195_groupi_n_1843);
  xnor csa_tree_add_190_195_groupi_g45370(csa_tree_add_190_195_groupi_n_3789 ,csa_tree_add_190_195_groupi_n_915 ,csa_tree_add_190_195_groupi_n_1861);
  xnor csa_tree_add_190_195_groupi_g45371(csa_tree_add_190_195_groupi_n_3788 ,csa_tree_add_190_195_groupi_n_210 ,csa_tree_add_190_195_groupi_n_1640);
  xnor csa_tree_add_190_195_groupi_g45372(csa_tree_add_190_195_groupi_n_3787 ,csa_tree_add_190_195_groupi_n_909 ,csa_tree_add_190_195_groupi_n_1673);
  xnor csa_tree_add_190_195_groupi_g45373(csa_tree_add_190_195_groupi_n_3786 ,csa_tree_add_190_195_groupi_n_1086 ,csa_tree_add_190_195_groupi_n_1134);
  xnor csa_tree_add_190_195_groupi_g45374(csa_tree_add_190_195_groupi_n_3785 ,csa_tree_add_190_195_groupi_n_2057 ,csa_tree_add_190_195_groupi_n_1965);
  xnor csa_tree_add_190_195_groupi_g45376(csa_tree_add_190_195_groupi_n_3784 ,csa_tree_add_190_195_groupi_n_942 ,csa_tree_add_190_195_groupi_n_1152);
  xnor csa_tree_add_190_195_groupi_g45377(csa_tree_add_190_195_groupi_n_3783 ,csa_tree_add_190_195_groupi_n_859 ,csa_tree_add_190_195_groupi_n_1604);
  xnor csa_tree_add_190_195_groupi_g45378(csa_tree_add_190_195_groupi_n_3782 ,csa_tree_add_190_195_groupi_n_834 ,csa_tree_add_190_195_groupi_n_1828);
  xnor csa_tree_add_190_195_groupi_g45379(csa_tree_add_190_195_groupi_n_3781 ,csa_tree_add_190_195_groupi_n_819 ,in57[1]);
  xnor csa_tree_add_190_195_groupi_g45381(csa_tree_add_190_195_groupi_n_3780 ,csa_tree_add_190_195_groupi_n_2214 ,csa_tree_add_190_195_groupi_n_1744);
  xnor csa_tree_add_190_195_groupi_g45382(csa_tree_add_190_195_groupi_n_3779 ,csa_tree_add_190_195_groupi_n_816 ,csa_tree_add_190_195_groupi_n_1703);
  xnor csa_tree_add_190_195_groupi_g45383(csa_tree_add_190_195_groupi_n_3778 ,csa_tree_add_190_195_groupi_n_939 ,csa_tree_add_190_195_groupi_n_2116);
  xnor csa_tree_add_190_195_groupi_g45384(csa_tree_add_190_195_groupi_n_3777 ,csa_tree_add_190_195_groupi_n_2209 ,csa_tree_add_190_195_groupi_n_2157);
  xnor csa_tree_add_190_195_groupi_g45385(csa_tree_add_190_195_groupi_n_3776 ,csa_tree_add_190_195_groupi_n_2437 ,csa_tree_add_190_195_groupi_n_1434);
  xnor csa_tree_add_190_195_groupi_g45386(csa_tree_add_190_195_groupi_n_3775 ,csa_tree_add_190_195_groupi_n_1975 ,csa_tree_add_190_195_groupi_n_1182);
  xnor csa_tree_add_190_195_groupi_g45387(csa_tree_add_190_195_groupi_n_3774 ,csa_tree_add_190_195_groupi_n_1197 ,csa_tree_add_190_195_groupi_n_1675);
  xnor csa_tree_add_190_195_groupi_g45388(csa_tree_add_190_195_groupi_n_3773 ,csa_tree_add_190_195_groupi_n_2211 ,csa_tree_add_190_195_groupi_n_1832);
  xnor csa_tree_add_190_195_groupi_g45389(csa_tree_add_190_195_groupi_n_3772 ,csa_tree_add_190_195_groupi_n_894 ,csa_tree_add_190_195_groupi_n_1684);
  xnor csa_tree_add_190_195_groupi_g45390(csa_tree_add_190_195_groupi_n_3771 ,csa_tree_add_190_195_groupi_n_748 ,csa_tree_add_190_195_groupi_n_1607);
  xnor csa_tree_add_190_195_groupi_g45391(csa_tree_add_190_195_groupi_n_3770 ,csa_tree_add_190_195_groupi_n_834 ,csa_tree_add_190_195_groupi_n_1829);
  xnor csa_tree_add_190_195_groupi_g45392(csa_tree_add_190_195_groupi_n_3769 ,csa_tree_add_190_195_groupi_n_1110 ,csa_tree_add_190_195_groupi_n_1177);
  xnor csa_tree_add_190_195_groupi_g45393(csa_tree_add_190_195_groupi_n_3768 ,csa_tree_add_190_195_groupi_n_967 ,csa_tree_add_190_195_groupi_n_1597);
  xnor csa_tree_add_190_195_groupi_g45394(csa_tree_add_190_195_groupi_n_3767 ,csa_tree_add_190_195_groupi_n_1893 ,csa_tree_add_190_195_groupi_n_1835);
  xnor csa_tree_add_190_195_groupi_g45395(csa_tree_add_190_195_groupi_n_3766 ,csa_tree_add_190_195_groupi_n_1831 ,csa_tree_add_190_195_groupi_n_1949);
  xnor csa_tree_add_190_195_groupi_g45396(csa_tree_add_190_195_groupi_n_3765 ,csa_tree_add_190_195_groupi_n_1831 ,csa_tree_add_190_195_groupi_n_2042);
  xnor csa_tree_add_190_195_groupi_g45397(csa_tree_add_190_195_groupi_n_3764 ,csa_tree_add_190_195_groupi_n_1775 ,csa_tree_add_190_195_groupi_n_1609);
  xnor csa_tree_add_190_195_groupi_g45398(csa_tree_add_190_195_groupi_n_3763 ,csa_tree_add_190_195_groupi_n_882 ,csa_tree_add_190_195_groupi_n_1589);
  xnor csa_tree_add_190_195_groupi_g45399(csa_tree_add_190_195_groupi_n_3762 ,csa_tree_add_190_195_groupi_n_1915 ,csa_tree_add_190_195_groupi_n_1831);
  xnor csa_tree_add_190_195_groupi_g45400(csa_tree_add_190_195_groupi_n_3761 ,csa_tree_add_190_195_groupi_n_2116 ,csa_tree_add_190_195_groupi_n_1176);
  xnor csa_tree_add_190_195_groupi_g45401(csa_tree_add_190_195_groupi_n_3760 ,csa_tree_add_190_195_groupi_n_2051 ,csa_tree_add_190_195_groupi_n_1691);
  xnor csa_tree_add_190_195_groupi_g45402(csa_tree_add_190_195_groupi_n_3759 ,csa_tree_add_190_195_groupi_n_775 ,csa_tree_add_190_195_groupi_n_1008);
  xnor csa_tree_add_190_195_groupi_g45403(csa_tree_add_190_195_groupi_n_3758 ,csa_tree_add_190_195_groupi_n_2042 ,csa_tree_add_190_195_groupi_n_1860);
  xnor csa_tree_add_190_195_groupi_g45404(csa_tree_add_190_195_groupi_n_3757 ,csa_tree_add_190_195_groupi_n_1836 ,csa_tree_add_190_195_groupi_n_1990);
  xnor csa_tree_add_190_195_groupi_g45405(csa_tree_add_190_195_groupi_n_3756 ,csa_tree_add_190_195_groupi_n_1069 ,csa_tree_add_190_195_groupi_n_946);
  xnor csa_tree_add_190_195_groupi_g45406(csa_tree_add_190_195_groupi_n_3755 ,csa_tree_add_190_195_groupi_n_2216 ,csa_tree_add_190_195_groupi_n_1746);
  xnor csa_tree_add_190_195_groupi_g45407(csa_tree_add_190_195_groupi_n_3754 ,csa_tree_add_190_195_groupi_n_1035 ,csa_tree_add_190_195_groupi_n_1967);
  xnor csa_tree_add_190_195_groupi_g45408(csa_tree_add_190_195_groupi_n_3753 ,csa_tree_add_190_195_groupi_n_1924 ,csa_tree_add_190_195_groupi_n_1752);
  xnor csa_tree_add_190_195_groupi_g45409(csa_tree_add_190_195_groupi_n_3752 ,csa_tree_add_190_195_groupi_n_1993 ,csa_tree_add_190_195_groupi_n_1990);
  xnor csa_tree_add_190_195_groupi_g45410(csa_tree_add_190_195_groupi_n_3751 ,csa_tree_add_190_195_groupi_n_1809 ,csa_tree_add_190_195_groupi_n_1705);
  xnor csa_tree_add_190_195_groupi_g45411(csa_tree_add_190_195_groupi_n_3750 ,csa_tree_add_190_195_groupi_n_1832 ,csa_tree_add_190_195_groupi_n_1827);
  xnor csa_tree_add_190_195_groupi_g45412(csa_tree_add_190_195_groupi_n_3749 ,csa_tree_add_190_195_groupi_n_1964 ,csa_tree_add_190_195_groupi_n_1693);
  xnor csa_tree_add_190_195_groupi_g45413(csa_tree_add_190_195_groupi_n_3748 ,csa_tree_add_190_195_groupi_n_1997 ,csa_tree_add_190_195_groupi_n_1833);
  xnor csa_tree_add_190_195_groupi_g45414(csa_tree_add_190_195_groupi_n_3747 ,csa_tree_add_190_195_groupi_n_1908 ,in61[0]);
  xnor csa_tree_add_190_195_groupi_g45415(csa_tree_add_190_195_groupi_n_3746 ,csa_tree_add_190_195_groupi_n_2007 ,csa_tree_add_190_195_groupi_n_1575);
  xnor csa_tree_add_190_195_groupi_g45416(csa_tree_add_190_195_groupi_n_3745 ,csa_tree_add_190_195_groupi_n_1966 ,csa_tree_add_190_195_groupi_n_1760);
  xnor csa_tree_add_190_195_groupi_g45417(csa_tree_add_190_195_groupi_n_3744 ,csa_tree_add_190_195_groupi_n_1970 ,csa_tree_add_190_195_groupi_n_1966);
  xnor csa_tree_add_190_195_groupi_g45418(csa_tree_add_190_195_groupi_n_3743 ,csa_tree_add_190_195_groupi_n_1903 ,csa_tree_add_190_195_groupi_n_1895);
  xnor csa_tree_add_190_195_groupi_g45419(csa_tree_add_190_195_groupi_n_3742 ,csa_tree_add_190_195_groupi_n_1748 ,csa_tree_add_190_195_groupi_n_1900);
  xnor csa_tree_add_190_195_groupi_g45420(csa_tree_add_190_195_groupi_n_3741 ,csa_tree_add_190_195_groupi_n_1702 ,csa_tree_add_190_195_groupi_n_1620);
  xnor csa_tree_add_190_195_groupi_g45421(csa_tree_add_190_195_groupi_n_3740 ,csa_tree_add_190_195_groupi_n_1706 ,csa_tree_add_190_195_groupi_n_1705);
  xnor csa_tree_add_190_195_groupi_g45422(csa_tree_add_190_195_groupi_n_3739 ,csa_tree_add_190_195_groupi_n_1812 ,csa_tree_add_190_195_groupi_n_1811);
  xnor csa_tree_add_190_195_groupi_g45423(csa_tree_add_190_195_groupi_n_3738 ,csa_tree_add_190_195_groupi_n_2085 ,csa_tree_add_190_195_groupi_n_1753);
  xnor csa_tree_add_190_195_groupi_g45424(csa_tree_add_190_195_groupi_n_3737 ,csa_tree_add_190_195_groupi_n_1763 ,csa_tree_add_190_195_groupi_n_1762);
  xnor csa_tree_add_190_195_groupi_g45425(csa_tree_add_190_195_groupi_n_3736 ,csa_tree_add_190_195_groupi_n_1933 ,csa_tree_add_190_195_groupi_n_1765);
  xnor csa_tree_add_190_195_groupi_g45426(csa_tree_add_190_195_groupi_n_3735 ,csa_tree_add_190_195_groupi_n_1937 ,csa_tree_add_190_195_groupi_n_1992);
  xnor csa_tree_add_190_195_groupi_g45427(csa_tree_add_190_195_groupi_n_3734 ,csa_tree_add_190_195_groupi_n_1665 ,csa_tree_add_190_195_groupi_n_1662);
  xnor csa_tree_add_190_195_groupi_g45428(csa_tree_add_190_195_groupi_n_3733 ,csa_tree_add_190_195_groupi_n_1943 ,csa_tree_add_190_195_groupi_n_1853);
  xnor csa_tree_add_190_195_groupi_g45429(csa_tree_add_190_195_groupi_n_3732 ,csa_tree_add_190_195_groupi_n_1747 ,csa_tree_add_190_195_groupi_n_1627);
  xnor csa_tree_add_190_195_groupi_g45430(csa_tree_add_190_195_groupi_n_3731 ,csa_tree_add_190_195_groupi_n_1867 ,csa_tree_add_190_195_groupi_n_1759);
  xnor csa_tree_add_190_195_groupi_g45431(csa_tree_add_190_195_groupi_n_3730 ,csa_tree_add_190_195_groupi_n_1777 ,csa_tree_add_190_195_groupi_n_1686);
  xnor csa_tree_add_190_195_groupi_g45432(csa_tree_add_190_195_groupi_n_4142 ,in55[3] ,in55[1]);
  xnor csa_tree_add_190_195_groupi_g45433(csa_tree_add_190_195_groupi_n_4141 ,in55[8] ,in61[5]);
  xnor csa_tree_add_190_195_groupi_g45434(csa_tree_add_190_195_groupi_n_4140 ,in55[10] ,in61[7]);
  xnor csa_tree_add_190_195_groupi_g45435(csa_tree_add_190_195_groupi_n_4139 ,in55[5] ,in55[3]);
  xnor csa_tree_add_190_195_groupi_g45436(csa_tree_add_190_195_groupi_n_4138 ,in55[6] ,in55[4]);
  xnor csa_tree_add_190_195_groupi_g45437(csa_tree_add_190_195_groupi_n_4137 ,csa_tree_add_190_195_groupi_n_846 ,csa_tree_add_190_195_groupi_n_1667);
  xnor csa_tree_add_190_195_groupi_g45438(csa_tree_add_190_195_groupi_n_4136 ,in55[13] ,in55[12]);
  xnor csa_tree_add_190_195_groupi_g45439(csa_tree_add_190_195_groupi_n_4135 ,in60[15] ,in57[15]);
  xnor csa_tree_add_190_195_groupi_g45440(csa_tree_add_190_195_groupi_n_4134 ,in60[3] ,in56[3]);
  xnor csa_tree_add_190_195_groupi_g45441(csa_tree_add_190_195_groupi_n_4132 ,csa_tree_add_190_195_groupi_n_1845 ,csa_tree_add_190_195_groupi_n_1550);
  xnor csa_tree_add_190_195_groupi_g45442(csa_tree_add_190_195_groupi_n_4131 ,csa_tree_add_190_195_groupi_n_1999 ,csa_tree_add_190_195_groupi_n_2064);
  xnor csa_tree_add_190_195_groupi_g45443(csa_tree_add_190_195_groupi_n_4130 ,csa_tree_add_190_195_groupi_n_961 ,csa_tree_add_190_195_groupi_n_1855);
  xnor csa_tree_add_190_195_groupi_g45444(csa_tree_add_190_195_groupi_n_4129 ,csa_tree_add_190_195_groupi_n_1695 ,csa_tree_add_190_195_groupi_n_1819);
  xnor csa_tree_add_190_195_groupi_g45445(csa_tree_add_190_195_groupi_n_4128 ,csa_tree_add_190_195_groupi_n_2091 ,csa_tree_add_190_195_groupi_n_2087);
  xnor csa_tree_add_190_195_groupi_g45446(csa_tree_add_190_195_groupi_n_4127 ,in55[9] ,in57[12]);
  xnor csa_tree_add_190_195_groupi_g45447(csa_tree_add_190_195_groupi_n_4125 ,csa_tree_add_190_195_groupi_n_1687 ,csa_tree_add_190_195_groupi_n_1854);
  xnor csa_tree_add_190_195_groupi_g45449(csa_tree_add_190_195_groupi_n_4124 ,csa_tree_add_190_195_groupi_n_1929 ,csa_tree_add_190_195_groupi_n_1851);
  xnor csa_tree_add_190_195_groupi_g45450(csa_tree_add_190_195_groupi_n_4123 ,csa_tree_add_190_195_groupi_n_2155 ,csa_tree_add_190_195_groupi_n_1754);
  xnor csa_tree_add_190_195_groupi_g45451(csa_tree_add_190_195_groupi_n_4122 ,csa_tree_add_190_195_groupi_n_1907 ,csa_tree_add_190_195_groupi_n_1763);
  xnor csa_tree_add_190_195_groupi_g45452(csa_tree_add_190_195_groupi_n_4121 ,csa_tree_add_190_195_groupi_n_1909 ,csa_tree_add_190_195_groupi_n_1910);
  xnor csa_tree_add_190_195_groupi_g45453(csa_tree_add_190_195_groupi_n_4120 ,csa_tree_add_190_195_groupi_n_1128 ,csa_tree_add_190_195_groupi_n_1572);
  xnor csa_tree_add_190_195_groupi_g45454(csa_tree_add_190_195_groupi_n_4119 ,csa_tree_add_190_195_groupi_n_1778 ,csa_tree_add_190_195_groupi_n_1608);
  xnor csa_tree_add_190_195_groupi_g45455(csa_tree_add_190_195_groupi_n_4118 ,in55[15] ,in55[14]);
  xnor csa_tree_add_190_195_groupi_g45456(csa_tree_add_190_195_groupi_n_4117 ,in55[15] ,in55[13]);
  xnor csa_tree_add_190_195_groupi_g45457(csa_tree_add_190_195_groupi_n_4114 ,csa_tree_add_190_195_groupi_n_2695 ,csa_tree_add_190_195_groupi_n_1615);
  not csa_tree_add_190_195_groupi_g45458(csa_tree_add_190_195_groupi_n_3728 ,csa_tree_add_190_195_groupi_n_3727);
  not csa_tree_add_190_195_groupi_g45459(csa_tree_add_190_195_groupi_n_3725 ,csa_tree_add_190_195_groupi_n_3724);
  not csa_tree_add_190_195_groupi_g45460(csa_tree_add_190_195_groupi_n_3721 ,csa_tree_add_190_195_groupi_n_3720);
  not csa_tree_add_190_195_groupi_g45461(csa_tree_add_190_195_groupi_n_3719 ,csa_tree_add_190_195_groupi_n_3718);
  not csa_tree_add_190_195_groupi_g45462(csa_tree_add_190_195_groupi_n_3717 ,csa_tree_add_190_195_groupi_n_3716);
  not csa_tree_add_190_195_groupi_g45463(csa_tree_add_190_195_groupi_n_3715 ,csa_tree_add_190_195_groupi_n_3714);
  not csa_tree_add_190_195_groupi_g45464(csa_tree_add_190_195_groupi_n_3712 ,csa_tree_add_190_195_groupi_n_3711);
  not csa_tree_add_190_195_groupi_g45465(csa_tree_add_190_195_groupi_n_3707 ,csa_tree_add_190_195_groupi_n_3706);
  not csa_tree_add_190_195_groupi_g45466(csa_tree_add_190_195_groupi_n_3703 ,csa_tree_add_190_195_groupi_n_3702);
  not csa_tree_add_190_195_groupi_g45467(csa_tree_add_190_195_groupi_n_3700 ,csa_tree_add_190_195_groupi_n_3701);
  not csa_tree_add_190_195_groupi_g45468(csa_tree_add_190_195_groupi_n_3698 ,csa_tree_add_190_195_groupi_n_3699);
  not csa_tree_add_190_195_groupi_g45470(csa_tree_add_190_195_groupi_n_3692 ,csa_tree_add_190_195_groupi_n_3693);
  not csa_tree_add_190_195_groupi_g45471(csa_tree_add_190_195_groupi_n_3691 ,csa_tree_add_190_195_groupi_n_3690);
  or csa_tree_add_190_195_groupi_g45472(csa_tree_add_190_195_groupi_n_3689 ,csa_tree_add_190_195_groupi_n_2213 ,csa_tree_add_190_195_groupi_n_2154);
  nor csa_tree_add_190_195_groupi_g45473(csa_tree_add_190_195_groupi_n_3688 ,csa_tree_add_190_195_groupi_n_2555 ,in58[0]);
  nor csa_tree_add_190_195_groupi_g45474(csa_tree_add_190_195_groupi_n_3687 ,csa_tree_add_190_195_groupi_n_2729 ,in58[7]);
  and csa_tree_add_190_195_groupi_g45475(csa_tree_add_190_195_groupi_n_3686 ,csa_tree_add_190_195_groupi_n_2083 ,csa_tree_add_190_195_groupi_n_1101);
  or csa_tree_add_190_195_groupi_g45476(csa_tree_add_190_195_groupi_n_3685 ,csa_tree_add_190_195_groupi_n_2558 ,in56[0]);
  or csa_tree_add_190_195_groupi_g45477(csa_tree_add_190_195_groupi_n_3684 ,csa_tree_add_190_195_groupi_n_2560 ,in56[7]);
  or csa_tree_add_190_195_groupi_g45478(csa_tree_add_190_195_groupi_n_3683 ,csa_tree_add_190_195_groupi_n_2718 ,csa_tree_add_190_195_groupi_n_1698);
  nor csa_tree_add_190_195_groupi_g45479(csa_tree_add_190_195_groupi_n_3682 ,csa_tree_add_190_195_groupi_n_2550 ,csa_tree_add_190_195_groupi_n_1854);
  or csa_tree_add_190_195_groupi_g45480(csa_tree_add_190_195_groupi_n_3681 ,csa_tree_add_190_195_groupi_n_2392 ,csa_tree_add_190_195_groupi_n_1687);
  or csa_tree_add_190_195_groupi_g45481(csa_tree_add_190_195_groupi_n_3680 ,csa_tree_add_190_195_groupi_n_1418 ,csa_tree_add_190_195_groupi_n_2668);
  or csa_tree_add_190_195_groupi_g45482(csa_tree_add_190_195_groupi_n_3679 ,csa_tree_add_190_195_groupi_n_2506 ,in56[8]);
  and csa_tree_add_190_195_groupi_g45483(csa_tree_add_190_195_groupi_n_3678 ,in56[8] ,csa_tree_add_190_195_groupi_n_2506);
  or csa_tree_add_190_195_groupi_g45484(csa_tree_add_190_195_groupi_n_3677 ,csa_tree_add_190_195_groupi_n_259 ,csa_tree_add_190_195_groupi_n_1930);
  nor csa_tree_add_190_195_groupi_g45485(csa_tree_add_190_195_groupi_n_3676 ,csa_tree_add_190_195_groupi_n_538 ,csa_tree_add_190_195_groupi_n_1265);
  nor csa_tree_add_190_195_groupi_g45486(csa_tree_add_190_195_groupi_n_3675 ,csa_tree_add_190_195_groupi_n_2389 ,csa_tree_add_190_195_groupi_n_2119);
  or csa_tree_add_190_195_groupi_g45487(csa_tree_add_190_195_groupi_n_3674 ,csa_tree_add_190_195_groupi_n_2655 ,csa_tree_add_190_195_groupi_n_1778);
  nor csa_tree_add_190_195_groupi_g45488(csa_tree_add_190_195_groupi_n_3673 ,csa_tree_add_190_195_groupi_n_2477 ,in59[2]);
  or csa_tree_add_190_195_groupi_g45489(csa_tree_add_190_195_groupi_n_3672 ,csa_tree_add_190_195_groupi_n_2720 ,csa_tree_add_190_195_groupi_n_204);
  nor csa_tree_add_190_195_groupi_g45490(csa_tree_add_190_195_groupi_n_3671 ,csa_tree_add_190_195_groupi_n_2614 ,in61[1]);
  or csa_tree_add_190_195_groupi_g45491(csa_tree_add_190_195_groupi_n_3670 ,csa_tree_add_190_195_groupi_n_2559 ,csa_tree_add_190_195_groupi_n_198);
  or csa_tree_add_190_195_groupi_g45492(csa_tree_add_190_195_groupi_n_3669 ,csa_tree_add_190_195_groupi_n_1334 ,in57[14]);
  nor csa_tree_add_190_195_groupi_g45493(csa_tree_add_190_195_groupi_n_3668 ,csa_tree_add_190_195_groupi_n_619 ,csa_tree_add_190_195_groupi_n_302);
  nor csa_tree_add_190_195_groupi_g45494(csa_tree_add_190_195_groupi_n_3667 ,csa_tree_add_190_195_groupi_n_2350 ,csa_tree_add_190_195_groupi_n_2156);
  or csa_tree_add_190_195_groupi_g45495(csa_tree_add_190_195_groupi_n_3666 ,csa_tree_add_190_195_groupi_n_2380 ,csa_tree_add_190_195_groupi_n_1976);
  or csa_tree_add_190_195_groupi_g45496(csa_tree_add_190_195_groupi_n_3665 ,csa_tree_add_190_195_groupi_n_2379 ,csa_tree_add_190_195_groupi_n_2056);
  nor csa_tree_add_190_195_groupi_g45497(csa_tree_add_190_195_groupi_n_3664 ,csa_tree_add_190_195_groupi_n_2386 ,csa_tree_add_190_195_groupi_n_2004);
  nor csa_tree_add_190_195_groupi_g45498(csa_tree_add_190_195_groupi_n_3663 ,csa_tree_add_190_195_groupi_n_2348 ,csa_tree_add_190_195_groupi_n_1604);
  or csa_tree_add_190_195_groupi_g45499(csa_tree_add_190_195_groupi_n_3662 ,csa_tree_add_190_195_groupi_n_2467 ,csa_tree_add_190_195_groupi_n_2000);
  or csa_tree_add_190_195_groupi_g45500(csa_tree_add_190_195_groupi_n_3661 ,csa_tree_add_190_195_groupi_n_1466 ,csa_tree_add_190_195_groupi_n_1711);
  nor csa_tree_add_190_195_groupi_g45501(csa_tree_add_190_195_groupi_n_3660 ,csa_tree_add_190_195_groupi_n_2351 ,csa_tree_add_190_195_groupi_n_982);
  nor csa_tree_add_190_195_groupi_g45502(csa_tree_add_190_195_groupi_n_3659 ,csa_tree_add_190_195_groupi_n_2657 ,csa_tree_add_190_195_groupi_n_1602);
  or csa_tree_add_190_195_groupi_g45503(csa_tree_add_190_195_groupi_n_3658 ,csa_tree_add_190_195_groupi_n_2484 ,csa_tree_add_190_195_groupi_n_1743);
  or csa_tree_add_190_195_groupi_g45504(csa_tree_add_190_195_groupi_n_3657 ,csa_tree_add_190_195_groupi_n_661 ,csa_tree_add_190_195_groupi_n_1943);
  and csa_tree_add_190_195_groupi_g45505(csa_tree_add_190_195_groupi_n_3656 ,csa_tree_add_190_195_groupi_n_1943 ,csa_tree_add_190_195_groupi_n_2639);
  or csa_tree_add_190_195_groupi_g45506(csa_tree_add_190_195_groupi_n_3655 ,csa_tree_add_190_195_groupi_n_667 ,csa_tree_add_190_195_groupi_n_1872);
  nor csa_tree_add_190_195_groupi_g45507(csa_tree_add_190_195_groupi_n_3654 ,csa_tree_add_190_195_groupi_n_2544 ,csa_tree_add_190_195_groupi_n_1866);
  and csa_tree_add_190_195_groupi_g45508(csa_tree_add_190_195_groupi_n_3653 ,csa_tree_add_190_195_groupi_n_2216 ,csa_tree_add_190_195_groupi_n_1920);
  nor csa_tree_add_190_195_groupi_g45509(csa_tree_add_190_195_groupi_n_3652 ,csa_tree_add_190_195_groupi_n_2711 ,csa_tree_add_190_195_groupi_n_1820);
  and csa_tree_add_190_195_groupi_g45510(csa_tree_add_190_195_groupi_n_3651 ,csa_tree_add_190_195_groupi_n_1872 ,csa_tree_add_190_195_groupi_n_667);
  or csa_tree_add_190_195_groupi_g45511(csa_tree_add_190_195_groupi_n_3650 ,csa_tree_add_190_195_groupi_n_2647 ,csa_tree_add_190_195_groupi_n_1747);
  nor csa_tree_add_190_195_groupi_g45512(csa_tree_add_190_195_groupi_n_3649 ,csa_tree_add_190_195_groupi_n_2353 ,csa_tree_add_190_195_groupi_n_1975);
  or csa_tree_add_190_195_groupi_g45513(csa_tree_add_190_195_groupi_n_3648 ,csa_tree_add_190_195_groupi_n_2610 ,csa_tree_add_190_195_groupi_n_1779);
  or csa_tree_add_190_195_groupi_g45514(csa_tree_add_190_195_groupi_n_3647 ,csa_tree_add_190_195_groupi_n_2501 ,csa_tree_add_190_195_groupi_n_2002);
  or csa_tree_add_190_195_groupi_g45515(csa_tree_add_190_195_groupi_n_3646 ,csa_tree_add_190_195_groupi_n_2349 ,csa_tree_add_190_195_groupi_n_1868);
  and csa_tree_add_190_195_groupi_g45516(csa_tree_add_190_195_groupi_n_3645 ,csa_tree_add_190_195_groupi_n_219 ,csa_tree_add_190_195_groupi_n_2541);
  and csa_tree_add_190_195_groupi_g45517(csa_tree_add_190_195_groupi_n_3644 ,csa_tree_add_190_195_groupi_n_2003 ,csa_tree_add_190_195_groupi_n_2640);
  nor csa_tree_add_190_195_groupi_g45518(csa_tree_add_190_195_groupi_n_3643 ,csa_tree_add_190_195_groupi_n_2670 ,csa_tree_add_190_195_groupi_n_1816);
  nor csa_tree_add_190_195_groupi_g45519(csa_tree_add_190_195_groupi_n_3642 ,csa_tree_add_190_195_groupi_n_2376 ,csa_tree_add_190_195_groupi_n_1117);
  nor csa_tree_add_190_195_groupi_g45520(csa_tree_add_190_195_groupi_n_3641 ,csa_tree_add_190_195_groupi_n_2451 ,csa_tree_add_190_195_groupi_n_1871);
  or csa_tree_add_190_195_groupi_g45521(csa_tree_add_190_195_groupi_n_3640 ,csa_tree_add_190_195_groupi_n_2640 ,csa_tree_add_190_195_groupi_n_2003);
  nor csa_tree_add_190_195_groupi_g45522(csa_tree_add_190_195_groupi_n_3639 ,csa_tree_add_190_195_groupi_n_2384 ,csa_tree_add_190_195_groupi_n_1877);
  or csa_tree_add_190_195_groupi_g45523(csa_tree_add_190_195_groupi_n_3638 ,csa_tree_add_190_195_groupi_n_2383 ,csa_tree_add_190_195_groupi_n_931);
  nor csa_tree_add_190_195_groupi_g45524(csa_tree_add_190_195_groupi_n_3637 ,csa_tree_add_190_195_groupi_n_2385 ,csa_tree_add_190_195_groupi_n_2216);
  or csa_tree_add_190_195_groupi_g45525(csa_tree_add_190_195_groupi_n_3636 ,csa_tree_add_190_195_groupi_n_2375 ,csa_tree_add_190_195_groupi_n_2005);
  or csa_tree_add_190_195_groupi_g45526(csa_tree_add_190_195_groupi_n_3635 ,csa_tree_add_190_195_groupi_n_2478 ,csa_tree_add_190_195_groupi_n_1664);
  nor csa_tree_add_190_195_groupi_g45527(csa_tree_add_190_195_groupi_n_3634 ,csa_tree_add_190_195_groupi_n_2709 ,csa_tree_add_190_195_groupi_n_1813);
  or csa_tree_add_190_195_groupi_g45528(csa_tree_add_190_195_groupi_n_3633 ,csa_tree_add_190_195_groupi_n_2541 ,csa_tree_add_190_195_groupi_n_218);
  and csa_tree_add_190_195_groupi_g45529(csa_tree_add_190_195_groupi_n_3632 ,csa_tree_add_190_195_groupi_n_1747 ,csa_tree_add_190_195_groupi_n_1458);
  nor csa_tree_add_190_195_groupi_g45530(csa_tree_add_190_195_groupi_n_3631 ,csa_tree_add_190_195_groupi_n_2609 ,csa_tree_add_190_195_groupi_n_1892);
  nor csa_tree_add_190_195_groupi_g45531(csa_tree_add_190_195_groupi_n_3630 ,csa_tree_add_190_195_groupi_n_2713 ,csa_tree_add_190_195_groupi_n_1931);
  or csa_tree_add_190_195_groupi_g45532(csa_tree_add_190_195_groupi_n_3629 ,csa_tree_add_190_195_groupi_n_2683 ,csa_tree_add_190_195_groupi_n_1760);
  or csa_tree_add_190_195_groupi_g45533(csa_tree_add_190_195_groupi_n_3628 ,csa_tree_add_190_195_groupi_n_2630 ,csa_tree_add_190_195_groupi_n_1704);
  or csa_tree_add_190_195_groupi_g45534(csa_tree_add_190_195_groupi_n_3627 ,csa_tree_add_190_195_groupi_n_2352 ,csa_tree_add_190_195_groupi_n_856);
  or csa_tree_add_190_195_groupi_g45535(csa_tree_add_190_195_groupi_n_3626 ,csa_tree_add_190_195_groupi_n_2530 ,csa_tree_add_190_195_groupi_n_1700);
  or csa_tree_add_190_195_groupi_g45536(csa_tree_add_190_195_groupi_n_3625 ,csa_tree_add_190_195_groupi_n_2502 ,csa_tree_add_190_195_groupi_n_1861);
  nor csa_tree_add_190_195_groupi_g45537(csa_tree_add_190_195_groupi_n_3624 ,csa_tree_add_190_195_groupi_n_2714 ,csa_tree_add_190_195_groupi_n_1823);
  or csa_tree_add_190_195_groupi_g45538(csa_tree_add_190_195_groupi_n_3623 ,csa_tree_add_190_195_groupi_n_2536 ,csa_tree_add_190_195_groupi_n_1605);
  and csa_tree_add_190_195_groupi_g45539(csa_tree_add_190_195_groupi_n_3622 ,csa_tree_add_190_195_groupi_n_1778 ,csa_tree_add_190_195_groupi_n_683);
  or csa_tree_add_190_195_groupi_g45540(csa_tree_add_190_195_groupi_n_3621 ,csa_tree_add_190_195_groupi_n_1999 ,csa_tree_add_190_195_groupi_n_2064);
  or csa_tree_add_190_195_groupi_g45541(csa_tree_add_190_195_groupi_n_3620 ,csa_tree_add_190_195_groupi_n_683 ,csa_tree_add_190_195_groupi_n_1778);
  or csa_tree_add_190_195_groupi_g45542(csa_tree_add_190_195_groupi_n_3619 ,csa_tree_add_190_195_groupi_n_273 ,csa_tree_add_190_195_groupi_n_1821);
  or csa_tree_add_190_195_groupi_g45543(csa_tree_add_190_195_groupi_n_3618 ,csa_tree_add_190_195_groupi_n_2355 ,csa_tree_add_190_195_groupi_n_229);
  nor csa_tree_add_190_195_groupi_g45544(csa_tree_add_190_195_groupi_n_3617 ,csa_tree_add_190_195_groupi_n_721 ,csa_tree_add_190_195_groupi_n_2008);
  nor csa_tree_add_190_195_groupi_g45545(csa_tree_add_190_195_groupi_n_3616 ,csa_tree_add_190_195_groupi_n_1392 ,csa_tree_add_190_195_groupi_n_1672);
  or csa_tree_add_190_195_groupi_g45546(csa_tree_add_190_195_groupi_n_3615 ,csa_tree_add_190_195_groupi_n_2347 ,csa_tree_add_190_195_groupi_n_873);
  or csa_tree_add_190_195_groupi_g45547(csa_tree_add_190_195_groupi_n_3614 ,csa_tree_add_190_195_groupi_n_2733 ,csa_tree_add_190_195_groupi_n_233);
  and csa_tree_add_190_195_groupi_g45548(csa_tree_add_190_195_groupi_n_3613 ,csa_tree_add_190_195_groupi_n_332 ,csa_tree_add_190_195_groupi_n_250);
  or csa_tree_add_190_195_groupi_g45549(csa_tree_add_190_195_groupi_n_3612 ,csa_tree_add_190_195_groupi_n_1526 ,csa_tree_add_190_195_groupi_n_1426);
  or csa_tree_add_190_195_groupi_g45550(csa_tree_add_190_195_groupi_n_3611 ,csa_tree_add_190_195_groupi_n_1928 ,csa_tree_add_190_195_groupi_n_1931);
  or csa_tree_add_190_195_groupi_g45551(csa_tree_add_190_195_groupi_n_3610 ,csa_tree_add_190_195_groupi_n_396 ,csa_tree_add_190_195_groupi_n_1173);
  nor csa_tree_add_190_195_groupi_g45552(csa_tree_add_190_195_groupi_n_3609 ,csa_tree_add_190_195_groupi_n_2534 ,csa_tree_add_190_195_groupi_n_1950);
  or csa_tree_add_190_195_groupi_g45553(csa_tree_add_190_195_groupi_n_3608 ,csa_tree_add_190_195_groupi_n_2485 ,csa_tree_add_190_195_groupi_n_1830);
  nor csa_tree_add_190_195_groupi_g45554(csa_tree_add_190_195_groupi_n_3607 ,csa_tree_add_190_195_groupi_n_2685 ,csa_tree_add_190_195_groupi_n_1715);
  and csa_tree_add_190_195_groupi_g45555(csa_tree_add_190_195_groupi_n_3606 ,csa_tree_add_190_195_groupi_n_1933 ,csa_tree_add_190_195_groupi_n_2460);
  or csa_tree_add_190_195_groupi_g45556(csa_tree_add_190_195_groupi_n_3605 ,csa_tree_add_190_195_groupi_n_2624 ,csa_tree_add_190_195_groupi_n_1748);
  or csa_tree_add_190_195_groupi_g45557(csa_tree_add_190_195_groupi_n_3604 ,csa_tree_add_190_195_groupi_n_678 ,csa_tree_add_190_195_groupi_n_1991);
  nor csa_tree_add_190_195_groupi_g45558(csa_tree_add_190_195_groupi_n_3603 ,csa_tree_add_190_195_groupi_n_2706 ,csa_tree_add_190_195_groupi_n_1978);
  nor csa_tree_add_190_195_groupi_g45559(csa_tree_add_190_195_groupi_n_3602 ,csa_tree_add_190_195_groupi_n_2696 ,csa_tree_add_190_195_groupi_n_798);
  nor csa_tree_add_190_195_groupi_g45560(csa_tree_add_190_195_groupi_n_3601 ,csa_tree_add_190_195_groupi_n_2709 ,csa_tree_add_190_195_groupi_n_1974);
  nor csa_tree_add_190_195_groupi_g45561(csa_tree_add_190_195_groupi_n_3600 ,csa_tree_add_190_195_groupi_n_754 ,csa_tree_add_190_195_groupi_n_1937);
  or csa_tree_add_190_195_groupi_g45562(csa_tree_add_190_195_groupi_n_3599 ,csa_tree_add_190_195_groupi_n_2499 ,csa_tree_add_190_195_groupi_n_1674);
  nor csa_tree_add_190_195_groupi_g45563(csa_tree_add_190_195_groupi_n_3598 ,csa_tree_add_190_195_groupi_n_2529 ,csa_tree_add_190_195_groupi_n_1677);
  or csa_tree_add_190_195_groupi_g45564(csa_tree_add_190_195_groupi_n_3597 ,csa_tree_add_190_195_groupi_n_2472 ,csa_tree_add_190_195_groupi_n_1707);
  or csa_tree_add_190_195_groupi_g45565(csa_tree_add_190_195_groupi_n_3596 ,csa_tree_add_190_195_groupi_n_2626 ,csa_tree_add_190_195_groupi_n_1841);
  nor csa_tree_add_190_195_groupi_g45566(csa_tree_add_190_195_groupi_n_3595 ,csa_tree_add_190_195_groupi_n_2517 ,csa_tree_add_190_195_groupi_n_2213);
  and csa_tree_add_190_195_groupi_g45567(csa_tree_add_190_195_groupi_n_3594 ,csa_tree_add_190_195_groupi_n_1937 ,csa_tree_add_190_195_groupi_n_1992);
  or csa_tree_add_190_195_groupi_g45568(csa_tree_add_190_195_groupi_n_3593 ,csa_tree_add_190_195_groupi_n_2707 ,csa_tree_add_190_195_groupi_n_1023);
  nor csa_tree_add_190_195_groupi_g45569(csa_tree_add_190_195_groupi_n_3592 ,csa_tree_add_190_195_groupi_n_2684 ,csa_tree_add_190_195_groupi_n_1909);
  or csa_tree_add_190_195_groupi_g45570(csa_tree_add_190_195_groupi_n_3591 ,csa_tree_add_190_195_groupi_n_2530 ,csa_tree_add_190_195_groupi_n_1066);
  nor csa_tree_add_190_195_groupi_g45571(csa_tree_add_190_195_groupi_n_3590 ,csa_tree_add_190_195_groupi_n_2700 ,csa_tree_add_190_195_groupi_n_1923);
  and csa_tree_add_190_195_groupi_g45572(csa_tree_add_190_195_groupi_n_3589 ,csa_tree_add_190_195_groupi_n_2085 ,csa_tree_add_190_195_groupi_n_2662);
  or csa_tree_add_190_195_groupi_g45573(csa_tree_add_190_195_groupi_n_3588 ,csa_tree_add_190_195_groupi_n_2592 ,csa_tree_add_190_195_groupi_n_2727);
  or csa_tree_add_190_195_groupi_g45574(csa_tree_add_190_195_groupi_n_3587 ,csa_tree_add_190_195_groupi_n_2662 ,csa_tree_add_190_195_groupi_n_2085);
  or csa_tree_add_190_195_groupi_g45575(csa_tree_add_190_195_groupi_n_3586 ,csa_tree_add_190_195_groupi_n_2510 ,csa_tree_add_190_195_groupi_n_1869);
  or csa_tree_add_190_195_groupi_g45576(csa_tree_add_190_195_groupi_n_3585 ,csa_tree_add_190_195_groupi_n_2671 ,csa_tree_add_190_195_groupi_n_1992);
  nor csa_tree_add_190_195_groupi_g45577(csa_tree_add_190_195_groupi_n_3584 ,csa_tree_add_190_195_groupi_n_2496 ,csa_tree_add_190_195_groupi_n_1780);
  or csa_tree_add_190_195_groupi_g45578(csa_tree_add_190_195_groupi_n_3583 ,csa_tree_add_190_195_groupi_n_2531 ,csa_tree_add_190_195_groupi_n_912);
  or csa_tree_add_190_195_groupi_g45579(csa_tree_add_190_195_groupi_n_3582 ,csa_tree_add_190_195_groupi_n_2537 ,csa_tree_add_190_195_groupi_n_1830);
  nor csa_tree_add_190_195_groupi_g45580(csa_tree_add_190_195_groupi_n_3581 ,csa_tree_add_190_195_groupi_n_2527 ,csa_tree_add_190_195_groupi_n_1967);
  and csa_tree_add_190_195_groupi_g45581(csa_tree_add_190_195_groupi_n_3580 ,csa_tree_add_190_195_groupi_n_1830 ,csa_tree_add_190_195_groupi_n_2485);
  or csa_tree_add_190_195_groupi_g45582(csa_tree_add_190_195_groupi_n_3579 ,csa_tree_add_190_195_groupi_n_2446 ,csa_tree_add_190_195_groupi_n_1851);
  and csa_tree_add_190_195_groupi_g45583(csa_tree_add_190_195_groupi_n_3578 ,csa_tree_add_190_195_groupi_n_1991 ,csa_tree_add_190_195_groupi_n_678);
  nor csa_tree_add_190_195_groupi_g45584(csa_tree_add_190_195_groupi_n_3577 ,csa_tree_add_190_195_groupi_n_2538 ,csa_tree_add_190_195_groupi_n_1824);
  nor csa_tree_add_190_195_groupi_g45585(csa_tree_add_190_195_groupi_n_3576 ,csa_tree_add_190_195_groupi_n_2698 ,csa_tree_add_190_195_groupi_n_972);
  or csa_tree_add_190_195_groupi_g45586(csa_tree_add_190_195_groupi_n_3575 ,csa_tree_add_190_195_groupi_n_419 ,csa_tree_add_190_195_groupi_n_228);
  or csa_tree_add_190_195_groupi_g45587(csa_tree_add_190_195_groupi_n_3574 ,csa_tree_add_190_195_groupi_n_2691 ,csa_tree_add_190_195_groupi_n_1812);
  nor csa_tree_add_190_195_groupi_g45588(csa_tree_add_190_195_groupi_n_3573 ,csa_tree_add_190_195_groupi_n_2693 ,csa_tree_add_190_195_groupi_n_1978);
  or csa_tree_add_190_195_groupi_g45589(csa_tree_add_190_195_groupi_n_3572 ,csa_tree_add_190_195_groupi_n_1372 ,csa_tree_add_190_195_groupi_n_1706);
  nor csa_tree_add_190_195_groupi_g45590(csa_tree_add_190_195_groupi_n_3571 ,csa_tree_add_190_195_groupi_n_2623 ,csa_tree_add_190_195_groupi_n_1869);
  or csa_tree_add_190_195_groupi_g45591(csa_tree_add_190_195_groupi_n_3570 ,csa_tree_add_190_195_groupi_n_2685 ,csa_tree_add_190_195_groupi_n_2007);
  nor csa_tree_add_190_195_groupi_g45592(csa_tree_add_190_195_groupi_n_3569 ,csa_tree_add_190_195_groupi_n_2454 ,csa_tree_add_190_195_groupi_n_1850);
  or csa_tree_add_190_195_groupi_g45593(csa_tree_add_190_195_groupi_n_3568 ,csa_tree_add_190_195_groupi_n_1464 ,csa_tree_add_190_195_groupi_n_1819);
  nor csa_tree_add_190_195_groupi_g45594(csa_tree_add_190_195_groupi_n_3567 ,csa_tree_add_190_195_groupi_n_2533 ,csa_tree_add_190_195_groupi_n_1929);
  nor csa_tree_add_190_195_groupi_g45595(csa_tree_add_190_195_groupi_n_3566 ,csa_tree_add_190_195_groupi_n_2704 ,csa_tree_add_190_195_groupi_n_1863);
  nor csa_tree_add_190_195_groupi_g45596(csa_tree_add_190_195_groupi_n_3565 ,csa_tree_add_190_195_groupi_n_1537 ,csa_tree_add_190_195_groupi_n_1862);
  or csa_tree_add_190_195_groupi_g45597(csa_tree_add_190_195_groupi_n_3564 ,csa_tree_add_190_195_groupi_n_2468 ,csa_tree_add_190_195_groupi_n_1890);
  and csa_tree_add_190_195_groupi_g45598(csa_tree_add_190_195_groupi_n_3563 ,csa_tree_add_190_195_groupi_n_1908 ,csa_tree_add_190_195_groupi_n_2652);
  or csa_tree_add_190_195_groupi_g45599(csa_tree_add_190_195_groupi_n_3562 ,csa_tree_add_190_195_groupi_n_2509 ,csa_tree_add_190_195_groupi_n_1751);
  or csa_tree_add_190_195_groupi_g45600(csa_tree_add_190_195_groupi_n_3561 ,csa_tree_add_190_195_groupi_n_2524 ,csa_tree_add_190_195_groupi_n_2117);
  or csa_tree_add_190_195_groupi_g45601(csa_tree_add_190_195_groupi_n_3560 ,csa_tree_add_190_195_groupi_n_2471 ,csa_tree_add_190_195_groupi_n_2087);
  nor csa_tree_add_190_195_groupi_g45602(csa_tree_add_190_195_groupi_n_3559 ,csa_tree_add_190_195_groupi_n_2374 ,csa_tree_add_190_195_groupi_n_1909);
  or csa_tree_add_190_195_groupi_g45603(csa_tree_add_190_195_groupi_n_3558 ,csa_tree_add_190_195_groupi_n_2468 ,csa_tree_add_190_195_groupi_n_1695);
  or csa_tree_add_190_195_groupi_g45604(csa_tree_add_190_195_groupi_n_3557 ,csa_tree_add_190_195_groupi_n_2705 ,csa_tree_add_190_195_groupi_n_1933);
  or csa_tree_add_190_195_groupi_g45605(csa_tree_add_190_195_groupi_n_3556 ,csa_tree_add_190_195_groupi_n_2519 ,csa_tree_add_190_195_groupi_n_1909);
  nor csa_tree_add_190_195_groupi_g45606(csa_tree_add_190_195_groupi_n_3555 ,csa_tree_add_190_195_groupi_n_2522 ,csa_tree_add_190_195_groupi_n_2118);
  nor csa_tree_add_190_195_groupi_g45607(csa_tree_add_190_195_groupi_n_3554 ,csa_tree_add_190_195_groupi_n_2518 ,csa_tree_add_190_195_groupi_n_993);
  or csa_tree_add_190_195_groupi_g45608(csa_tree_add_190_195_groupi_n_3553 ,csa_tree_add_190_195_groupi_n_1464 ,csa_tree_add_190_195_groupi_n_1908);
  or csa_tree_add_190_195_groupi_g45609(csa_tree_add_190_195_groupi_n_3552 ,csa_tree_add_190_195_groupi_n_2671 ,csa_tree_add_190_195_groupi_n_1908);
  nor csa_tree_add_190_195_groupi_g45610(csa_tree_add_190_195_groupi_n_3551 ,in55[9] ,in61[13]);
  or csa_tree_add_190_195_groupi_g45611(csa_tree_add_190_195_groupi_n_3550 ,csa_tree_add_190_195_groupi_n_2083 ,csa_tree_add_190_195_groupi_n_221);
  nor csa_tree_add_190_195_groupi_g45612(csa_tree_add_190_195_groupi_n_3549 ,csa_tree_add_190_195_groupi_n_2701 ,csa_tree_add_190_195_groupi_n_2154);
  nor csa_tree_add_190_195_groupi_g45613(csa_tree_add_190_195_groupi_n_3548 ,csa_tree_add_190_195_groupi_n_2346 ,csa_tree_add_190_195_groupi_n_1936);
  nor csa_tree_add_190_195_groupi_g45614(csa_tree_add_190_195_groupi_n_3547 ,csa_tree_add_190_195_groupi_n_2694 ,csa_tree_add_190_195_groupi_n_2058);
  or csa_tree_add_190_195_groupi_g45615(csa_tree_add_190_195_groupi_n_3546 ,csa_tree_add_190_195_groupi_n_2505 ,csa_tree_add_190_195_groupi_n_1677);
  or csa_tree_add_190_195_groupi_g45616(csa_tree_add_190_195_groupi_n_3545 ,csa_tree_add_190_195_groupi_n_2694 ,csa_tree_add_190_195_groupi_n_2057);
  or csa_tree_add_190_195_groupi_g45617(csa_tree_add_190_195_groupi_n_3544 ,csa_tree_add_190_195_groupi_n_2681 ,csa_tree_add_190_195_groupi_n_1928);
  and csa_tree_add_190_195_groupi_g45618(csa_tree_add_190_195_groupi_n_3543 ,csa_tree_add_190_195_groupi_n_1935 ,csa_tree_add_190_195_groupi_n_2659);
  nor csa_tree_add_190_195_groupi_g45619(csa_tree_add_190_195_groupi_n_3542 ,csa_tree_add_190_195_groupi_n_2439 ,csa_tree_add_190_195_groupi_n_1818);
  nor csa_tree_add_190_195_groupi_g45620(csa_tree_add_190_195_groupi_n_3541 ,csa_tree_add_190_195_groupi_n_1199 ,csa_tree_add_190_195_groupi_n_1123);
  nand csa_tree_add_190_195_groupi_g45621(csa_tree_add_190_195_groupi_n_3540 ,in58[12] ,in59[12]);
  nor csa_tree_add_190_195_groupi_g45622(csa_tree_add_190_195_groupi_n_3539 ,csa_tree_add_190_195_groupi_n_461 ,csa_tree_add_190_195_groupi_n_2708);
  nor csa_tree_add_190_195_groupi_g45623(csa_tree_add_190_195_groupi_n_3538 ,csa_tree_add_190_195_groupi_n_2651 ,csa_tree_add_190_195_groupi_n_1823);
  or csa_tree_add_190_195_groupi_g45624(csa_tree_add_190_195_groupi_n_3537 ,csa_tree_add_190_195_groupi_n_1152 ,csa_tree_add_190_195_groupi_n_1075);
  nor csa_tree_add_190_195_groupi_g45625(csa_tree_add_190_195_groupi_n_3536 ,csa_tree_add_190_195_groupi_n_2671 ,csa_tree_add_190_195_groupi_n_1910);
  or csa_tree_add_190_195_groupi_g45626(csa_tree_add_190_195_groupi_n_3535 ,csa_tree_add_190_195_groupi_n_2635 ,csa_tree_add_190_195_groupi_n_1868);
  or csa_tree_add_190_195_groupi_g45627(csa_tree_add_190_195_groupi_n_3534 ,csa_tree_add_190_195_groupi_n_2680 ,csa_tree_add_190_195_groupi_n_1093);
  and csa_tree_add_190_195_groupi_g45628(csa_tree_add_190_195_groupi_n_3533 ,csa_tree_add_190_195_groupi_n_293 ,csa_tree_add_190_195_groupi_n_712);
  nor csa_tree_add_190_195_groupi_g45629(csa_tree_add_190_195_groupi_n_3532 ,csa_tree_add_190_195_groupi_n_2679 ,csa_tree_add_190_195_groupi_n_1880);
  nor csa_tree_add_190_195_groupi_g45630(csa_tree_add_190_195_groupi_n_3531 ,csa_tree_add_190_195_groupi_n_2452 ,csa_tree_add_190_195_groupi_n_1860);
  nor csa_tree_add_190_195_groupi_g45631(csa_tree_add_190_195_groupi_n_3530 ,csa_tree_add_190_195_groupi_n_2452 ,csa_tree_add_190_195_groupi_n_1951);
  or csa_tree_add_190_195_groupi_g45632(csa_tree_add_190_195_groupi_n_3529 ,csa_tree_add_190_195_groupi_n_2481 ,csa_tree_add_190_195_groupi_n_1855);
  nor csa_tree_add_190_195_groupi_g45633(csa_tree_add_190_195_groupi_n_3528 ,csa_tree_add_190_195_groupi_n_2689 ,csa_tree_add_190_195_groupi_n_1921);
  or csa_tree_add_190_195_groupi_g45634(csa_tree_add_190_195_groupi_n_3527 ,csa_tree_add_190_195_groupi_n_2615 ,csa_tree_add_190_195_groupi_n_1835);
  or csa_tree_add_190_195_groupi_g45635(csa_tree_add_190_195_groupi_n_3526 ,csa_tree_add_190_195_groupi_n_2488 ,csa_tree_add_190_195_groupi_n_1936);
  and csa_tree_add_190_195_groupi_g45636(csa_tree_add_190_195_groupi_n_3525 ,csa_tree_add_190_195_groupi_n_1936 ,csa_tree_add_190_195_groupi_n_1508);
  or csa_tree_add_190_195_groupi_g45637(csa_tree_add_190_195_groupi_n_3524 ,csa_tree_add_190_195_groupi_n_1503 ,csa_tree_add_190_195_groupi_n_1933);
  or csa_tree_add_190_195_groupi_g45638(csa_tree_add_190_195_groupi_n_3523 ,csa_tree_add_190_195_groupi_n_2528 ,csa_tree_add_190_195_groupi_n_2054);
  and csa_tree_add_190_195_groupi_g45639(csa_tree_add_190_195_groupi_n_3522 ,csa_tree_add_190_195_groupi_n_1937 ,csa_tree_add_190_195_groupi_n_754);
  or csa_tree_add_190_195_groupi_g45640(csa_tree_add_190_195_groupi_n_3521 ,csa_tree_add_190_195_groupi_n_2699 ,csa_tree_add_190_195_groupi_n_1607);
  or csa_tree_add_190_195_groupi_g45641(csa_tree_add_190_195_groupi_n_3520 ,csa_tree_add_190_195_groupi_n_1482 ,csa_tree_add_190_195_groupi_n_1935);
  or csa_tree_add_190_195_groupi_g45642(csa_tree_add_190_195_groupi_n_3519 ,csa_tree_add_190_195_groupi_n_2447 ,csa_tree_add_190_195_groupi_n_2089);
  nor csa_tree_add_190_195_groupi_g45643(csa_tree_add_190_195_groupi_n_3518 ,csa_tree_add_190_195_groupi_n_2687 ,csa_tree_add_190_195_groupi_n_2061);
  nor csa_tree_add_190_195_groupi_g45644(csa_tree_add_190_195_groupi_n_3517 ,csa_tree_add_190_195_groupi_n_1472 ,csa_tree_add_190_195_groupi_n_2015);
  and csa_tree_add_190_195_groupi_g45645(csa_tree_add_190_195_groupi_n_3516 ,csa_tree_add_190_195_groupi_n_2015 ,csa_tree_add_190_195_groupi_n_1472);
  and csa_tree_add_190_195_groupi_g45646(csa_tree_add_190_195_groupi_n_3515 ,in56[6] ,csa_tree_add_190_195_groupi_n_676);
  or csa_tree_add_190_195_groupi_g45647(csa_tree_add_190_195_groupi_n_3514 ,csa_tree_add_190_195_groupi_n_700 ,csa_tree_add_190_195_groupi_n_1873);
  nor csa_tree_add_190_195_groupi_g45648(csa_tree_add_190_195_groupi_n_3513 ,csa_tree_add_190_195_groupi_n_1506 ,csa_tree_add_190_195_groupi_n_1890);
  or csa_tree_add_190_195_groupi_g45649(csa_tree_add_190_195_groupi_n_3512 ,csa_tree_add_190_195_groupi_n_2693 ,csa_tree_add_190_195_groupi_n_510);
  and csa_tree_add_190_195_groupi_g45650(csa_tree_add_190_195_groupi_n_3511 ,csa_tree_add_190_195_groupi_n_1606 ,csa_tree_add_190_195_groupi_n_765);
  nor csa_tree_add_190_195_groupi_g45651(csa_tree_add_190_195_groupi_n_3510 ,csa_tree_add_190_195_groupi_n_1560 ,csa_tree_add_190_195_groupi_n_1815);
  or csa_tree_add_190_195_groupi_g45652(csa_tree_add_190_195_groupi_n_3509 ,csa_tree_add_190_195_groupi_n_829 ,csa_tree_add_190_195_groupi_n_1603);
  and csa_tree_add_190_195_groupi_g45653(csa_tree_add_190_195_groupi_n_3508 ,csa_tree_add_190_195_groupi_n_1841 ,csa_tree_add_190_195_groupi_n_2413);
  or csa_tree_add_190_195_groupi_g45654(csa_tree_add_190_195_groupi_n_3507 ,csa_tree_add_190_195_groupi_n_2703 ,csa_tree_add_190_195_groupi_n_432);
  or csa_tree_add_190_195_groupi_g45655(csa_tree_add_190_195_groupi_n_3506 ,csa_tree_add_190_195_groupi_n_739 ,in56[6]);
  and csa_tree_add_190_195_groupi_g45656(csa_tree_add_190_195_groupi_n_3505 ,csa_tree_add_190_195_groupi_n_2085 ,csa_tree_add_190_195_groupi_n_1490);
  or csa_tree_add_190_195_groupi_g45657(csa_tree_add_190_195_groupi_n_3504 ,csa_tree_add_190_195_groupi_n_729 ,csa_tree_add_190_195_groupi_n_1822);
  and csa_tree_add_190_195_groupi_g45658(csa_tree_add_190_195_groupi_n_3503 ,csa_tree_add_190_195_groupi_n_1822 ,csa_tree_add_190_195_groupi_n_1548);
  or csa_tree_add_190_195_groupi_g45659(csa_tree_add_190_195_groupi_n_3502 ,csa_tree_add_190_195_groupi_n_2520 ,csa_tree_add_190_195_groupi_n_624);
  or csa_tree_add_190_195_groupi_g45660(csa_tree_add_190_195_groupi_n_3501 ,csa_tree_add_190_195_groupi_n_1491 ,csa_tree_add_190_195_groupi_n_2085);
  and csa_tree_add_190_195_groupi_g45661(csa_tree_add_190_195_groupi_n_3500 ,csa_tree_add_190_195_groupi_n_1950 ,csa_tree_add_190_195_groupi_n_1477);
  or csa_tree_add_190_195_groupi_g45662(csa_tree_add_190_195_groupi_n_3499 ,csa_tree_add_190_195_groupi_n_1478 ,csa_tree_add_190_195_groupi_n_1950);
  nor csa_tree_add_190_195_groupi_g45663(csa_tree_add_190_195_groupi_n_3498 ,csa_tree_add_190_195_groupi_n_2412 ,csa_tree_add_190_195_groupi_n_2084);
  and csa_tree_add_190_195_groupi_g45664(csa_tree_add_190_195_groupi_n_3497 ,csa_tree_add_190_195_groupi_n_1603 ,csa_tree_add_190_195_groupi_n_828);
  or csa_tree_add_190_195_groupi_g45665(csa_tree_add_190_195_groupi_n_3496 ,csa_tree_add_190_195_groupi_n_2387 ,csa_tree_add_190_195_groupi_n_317);
  or csa_tree_add_190_195_groupi_g45666(csa_tree_add_190_195_groupi_n_3495 ,csa_tree_add_190_195_groupi_n_726 ,csa_tree_add_190_195_groupi_n_1840);
  or csa_tree_add_190_195_groupi_g45667(csa_tree_add_190_195_groupi_n_3494 ,csa_tree_add_190_195_groupi_n_828 ,csa_tree_add_190_195_groupi_n_1606);
  or csa_tree_add_190_195_groupi_g45668(csa_tree_add_190_195_groupi_n_3493 ,csa_tree_add_190_195_groupi_n_2413 ,csa_tree_add_190_195_groupi_n_1841);
  nor csa_tree_add_190_195_groupi_g45669(csa_tree_add_190_195_groupi_n_3492 ,csa_tree_add_190_195_groupi_n_1525 ,csa_tree_add_190_195_groupi_n_1941);
  and csa_tree_add_190_195_groupi_g45670(csa_tree_add_190_195_groupi_n_3491 ,csa_tree_add_190_195_groupi_n_1840 ,csa_tree_add_190_195_groupi_n_745);
  and csa_tree_add_190_195_groupi_g45671(csa_tree_add_190_195_groupi_n_3490 ,csa_tree_add_190_195_groupi_n_1873 ,csa_tree_add_190_195_groupi_n_700);
  and csa_tree_add_190_195_groupi_g45672(csa_tree_add_190_195_groupi_n_3489 ,csa_tree_add_190_195_groupi_n_1147 ,csa_tree_add_190_195_groupi_n_1017);
  or csa_tree_add_190_195_groupi_g45673(csa_tree_add_190_195_groupi_n_3488 ,csa_tree_add_190_195_groupi_n_2372 ,csa_tree_add_190_195_groupi_n_466);
  nor csa_tree_add_190_195_groupi_g45674(csa_tree_add_190_195_groupi_n_3487 ,csa_tree_add_190_195_groupi_n_1505 ,csa_tree_add_190_195_groupi_n_2064);
  and csa_tree_add_190_195_groupi_g45675(csa_tree_add_190_195_groupi_n_3486 ,csa_tree_add_190_195_groupi_n_2052 ,csa_tree_add_190_195_groupi_n_685);
  or csa_tree_add_190_195_groupi_g45676(csa_tree_add_190_195_groupi_n_3485 ,csa_tree_add_190_195_groupi_n_1562 ,csa_tree_add_190_195_groupi_n_2052);
  or csa_tree_add_190_195_groupi_g45677(csa_tree_add_190_195_groupi_n_3484 ,in61[14] ,in58[14]);
  nor csa_tree_add_190_195_groupi_g45678(csa_tree_add_190_195_groupi_n_3483 ,csa_tree_add_190_195_groupi_n_2343 ,csa_tree_add_190_195_groupi_n_1995);
  or csa_tree_add_190_195_groupi_g45679(csa_tree_add_190_195_groupi_n_3482 ,csa_tree_add_190_195_groupi_n_681 ,csa_tree_add_190_195_groupi_n_2091);
  nor csa_tree_add_190_195_groupi_g45680(csa_tree_add_190_195_groupi_n_3481 ,csa_tree_add_190_195_groupi_n_2669 ,csa_tree_add_190_195_groupi_n_2053);
  nor csa_tree_add_190_195_groupi_g45681(csa_tree_add_190_195_groupi_n_3480 ,csa_tree_add_190_195_groupi_n_529 ,csa_tree_add_190_195_groupi_n_2505);
  or csa_tree_add_190_195_groupi_g45682(csa_tree_add_190_195_groupi_n_3479 ,csa_tree_add_190_195_groupi_n_2475 ,csa_tree_add_190_195_groupi_n_784);
  nor csa_tree_add_190_195_groupi_g45683(csa_tree_add_190_195_groupi_n_3478 ,csa_tree_add_190_195_groupi_n_2490 ,csa_tree_add_190_195_groupi_n_1715);
  or csa_tree_add_190_195_groupi_g45684(csa_tree_add_190_195_groupi_n_3477 ,csa_tree_add_190_195_groupi_n_2664 ,csa_tree_add_190_195_groupi_n_464);
  and csa_tree_add_190_195_groupi_g45685(csa_tree_add_190_195_groupi_n_3476 ,csa_tree_add_190_195_groupi_n_1929 ,csa_tree_add_190_195_groupi_n_733);
  nor csa_tree_add_190_195_groupi_g45686(csa_tree_add_190_195_groupi_n_3475 ,csa_tree_add_190_195_groupi_n_2511 ,csa_tree_add_190_195_groupi_n_1791);
  or csa_tree_add_190_195_groupi_g45687(csa_tree_add_190_195_groupi_n_3474 ,csa_tree_add_190_195_groupi_n_2612 ,csa_tree_add_190_195_groupi_n_2155);
  or csa_tree_add_190_195_groupi_g45688(csa_tree_add_190_195_groupi_n_3473 ,csa_tree_add_190_195_groupi_n_2480 ,csa_tree_add_190_195_groupi_n_746);
  and csa_tree_add_190_195_groupi_g45689(csa_tree_add_190_195_groupi_n_3472 ,csa_tree_add_190_195_groupi_n_1963 ,csa_tree_add_190_195_groupi_n_672);
  nor csa_tree_add_190_195_groupi_g45690(csa_tree_add_190_195_groupi_n_3471 ,csa_tree_add_190_195_groupi_n_2665 ,csa_tree_add_190_195_groupi_n_1253);
  nor csa_tree_add_190_195_groupi_g45691(csa_tree_add_190_195_groupi_n_3470 ,csa_tree_add_190_195_groupi_n_326 ,csa_tree_add_190_195_groupi_n_2508);
  nor csa_tree_add_190_195_groupi_g45692(csa_tree_add_190_195_groupi_n_3469 ,csa_tree_add_190_195_groupi_n_1557 ,csa_tree_add_190_195_groupi_n_1989);
  nor csa_tree_add_190_195_groupi_g45693(csa_tree_add_190_195_groupi_n_3468 ,csa_tree_add_190_195_groupi_n_2661 ,csa_tree_add_190_195_groupi_n_2063);
  or csa_tree_add_190_195_groupi_g45694(csa_tree_add_190_195_groupi_n_3467 ,csa_tree_add_190_195_groupi_n_2487 ,csa_tree_add_190_195_groupi_n_1964);
  or csa_tree_add_190_195_groupi_g45695(csa_tree_add_190_195_groupi_n_3466 ,csa_tree_add_190_195_groupi_n_2455 ,csa_tree_add_190_195_groupi_n_1993);
  or csa_tree_add_190_195_groupi_g45696(csa_tree_add_190_195_groupi_n_3465 ,csa_tree_add_190_195_groupi_n_2505 ,csa_tree_add_190_195_groupi_n_762);
  or csa_tree_add_190_195_groupi_g45697(csa_tree_add_190_195_groupi_n_3464 ,csa_tree_add_190_195_groupi_n_673 ,csa_tree_add_190_195_groupi_n_1963);
  or csa_tree_add_190_195_groupi_g45698(csa_tree_add_190_195_groupi_n_3463 ,csa_tree_add_190_195_groupi_n_1475 ,csa_tree_add_190_195_groupi_n_1715);
  or csa_tree_add_190_195_groupi_g45699(csa_tree_add_190_195_groupi_n_3462 ,csa_tree_add_190_195_groupi_n_2642 ,csa_tree_add_190_195_groupi_n_1998);
  nor csa_tree_add_190_195_groupi_g45700(csa_tree_add_190_195_groupi_n_3461 ,csa_tree_add_190_195_groupi_n_2370 ,csa_tree_add_190_195_groupi_n_1996);
  or csa_tree_add_190_195_groupi_g45701(csa_tree_add_190_195_groupi_n_3460 ,csa_tree_add_190_195_groupi_n_733 ,csa_tree_add_190_195_groupi_n_1929);
  nor csa_tree_add_190_195_groupi_g45702(csa_tree_add_190_195_groupi_n_3459 ,csa_tree_add_190_195_groupi_n_2660 ,csa_tree_add_190_195_groupi_n_2158);
  or csa_tree_add_190_195_groupi_g45703(csa_tree_add_190_195_groupi_n_3458 ,csa_tree_add_190_195_groupi_n_702 ,csa_tree_add_190_195_groupi_n_1932);
  and csa_tree_add_190_195_groupi_g45704(csa_tree_add_190_195_groupi_n_3457 ,csa_tree_add_190_195_groupi_n_2091 ,csa_tree_add_190_195_groupi_n_681);
  nor csa_tree_add_190_195_groupi_g45705(csa_tree_add_190_195_groupi_n_3456 ,csa_tree_add_190_195_groupi_n_2371 ,csa_tree_add_190_195_groupi_n_859);
  or csa_tree_add_190_195_groupi_g45706(csa_tree_add_190_195_groupi_n_3455 ,csa_tree_add_190_195_groupi_n_691 ,csa_tree_add_190_195_groupi_n_1809);
  or csa_tree_add_190_195_groupi_g45707(csa_tree_add_190_195_groupi_n_3454 ,csa_tree_add_190_195_groupi_n_2631 ,csa_tree_add_190_195_groupi_n_1997);
  or csa_tree_add_190_195_groupi_g45708(csa_tree_add_190_195_groupi_n_3453 ,csa_tree_add_190_195_groupi_n_1493 ,csa_tree_add_190_195_groupi_n_407);
  nor csa_tree_add_190_195_groupi_g45709(csa_tree_add_190_195_groupi_n_3452 ,csa_tree_add_190_195_groupi_n_2444 ,csa_tree_add_190_195_groupi_n_1006);
  or csa_tree_add_190_195_groupi_g45710(csa_tree_add_190_195_groupi_n_3451 ,csa_tree_add_190_195_groupi_n_2474 ,csa_tree_add_190_195_groupi_n_2117);
  or csa_tree_add_190_195_groupi_g45711(csa_tree_add_190_195_groupi_n_3450 ,csa_tree_add_190_195_groupi_n_2489 ,csa_tree_add_190_195_groupi_n_1839);
  and csa_tree_add_190_195_groupi_g45712(csa_tree_add_190_195_groupi_n_3449 ,csa_tree_add_190_195_groupi_n_201 ,csa_tree_add_190_195_groupi_n_2634);
  nor csa_tree_add_190_195_groupi_g45713(csa_tree_add_190_195_groupi_n_3448 ,csa_tree_add_190_195_groupi_n_1442 ,csa_tree_add_190_195_groupi_n_2039);
  nor csa_tree_add_190_195_groupi_g45714(csa_tree_add_190_195_groupi_n_3447 ,csa_tree_add_190_195_groupi_n_586 ,csa_tree_add_190_195_groupi_n_1397);
  or csa_tree_add_190_195_groupi_g45715(csa_tree_add_190_195_groupi_n_3446 ,csa_tree_add_190_195_groupi_n_661 ,csa_tree_add_190_195_groupi_n_939);
  or csa_tree_add_190_195_groupi_g45716(csa_tree_add_190_195_groupi_n_3445 ,csa_tree_add_190_195_groupi_n_2646 ,csa_tree_add_190_195_groupi_n_1161);
  or csa_tree_add_190_195_groupi_g45717(csa_tree_add_190_195_groupi_n_3444 ,csa_tree_add_190_195_groupi_n_2491 ,csa_tree_add_190_195_groupi_n_883);
  or csa_tree_add_190_195_groupi_g45718(csa_tree_add_190_195_groupi_n_3443 ,csa_tree_add_190_195_groupi_n_1480 ,csa_tree_add_190_195_groupi_n_1000);
  nor csa_tree_add_190_195_groupi_g45719(csa_tree_add_190_195_groupi_n_3442 ,csa_tree_add_190_195_groupi_n_2487 ,csa_tree_add_190_195_groupi_n_2055);
  or csa_tree_add_190_195_groupi_g45720(csa_tree_add_190_195_groupi_n_3441 ,csa_tree_add_190_195_groupi_n_2448 ,csa_tree_add_190_195_groupi_n_2053);
  or csa_tree_add_190_195_groupi_g45721(csa_tree_add_190_195_groupi_n_3440 ,csa_tree_add_190_195_groupi_n_2495 ,csa_tree_add_190_195_groupi_n_1065);
  and csa_tree_add_190_195_groupi_g45722(csa_tree_add_190_195_groupi_n_3439 ,csa_tree_add_190_195_groupi_n_407 ,csa_tree_add_190_195_groupi_n_2650);
  nor csa_tree_add_190_195_groupi_g45723(csa_tree_add_190_195_groupi_n_3438 ,csa_tree_add_190_195_groupi_n_2641 ,csa_tree_add_190_195_groupi_n_1730);
  nor csa_tree_add_190_195_groupi_g45724(csa_tree_add_190_195_groupi_n_3437 ,csa_tree_add_190_195_groupi_n_566 ,csa_tree_add_190_195_groupi_n_1458);
  or csa_tree_add_190_195_groupi_g45725(csa_tree_add_190_195_groupi_n_3436 ,csa_tree_add_190_195_groupi_n_1493 ,csa_tree_add_190_195_groupi_n_1216);
  nor csa_tree_add_190_195_groupi_g45726(csa_tree_add_190_195_groupi_n_3435 ,csa_tree_add_190_195_groupi_n_1364 ,csa_tree_add_190_195_groupi_n_904);
  or csa_tree_add_190_195_groupi_g45727(csa_tree_add_190_195_groupi_n_3434 ,csa_tree_add_190_195_groupi_n_670 ,csa_tree_add_190_195_groupi_n_773);
  or csa_tree_add_190_195_groupi_g45728(csa_tree_add_190_195_groupi_n_3433 ,csa_tree_add_190_195_groupi_n_2654 ,csa_tree_add_190_195_groupi_n_972);
  or csa_tree_add_190_195_groupi_g45729(csa_tree_add_190_195_groupi_n_3432 ,csa_tree_add_190_195_groupi_n_2618 ,csa_tree_add_190_195_groupi_n_1056);
  nor csa_tree_add_190_195_groupi_g45730(csa_tree_add_190_195_groupi_n_3431 ,csa_tree_add_190_195_groupi_n_1397 ,csa_tree_add_190_195_groupi_n_1922);
  nor csa_tree_add_190_195_groupi_g45731(csa_tree_add_190_195_groupi_n_3430 ,csa_tree_add_190_195_groupi_n_1531 ,csa_tree_add_190_195_groupi_n_1745);
  or csa_tree_add_190_195_groupi_g45732(csa_tree_add_190_195_groupi_n_3429 ,csa_tree_add_190_195_groupi_n_664 ,csa_tree_add_190_195_groupi_n_1024);
  or csa_tree_add_190_195_groupi_g45733(csa_tree_add_190_195_groupi_n_3428 ,csa_tree_add_190_195_groupi_n_1353 ,csa_tree_add_190_195_groupi_n_437);
  nor csa_tree_add_190_195_groupi_g45734(csa_tree_add_190_195_groupi_n_3427 ,csa_tree_add_190_195_groupi_n_2496 ,csa_tree_add_190_195_groupi_n_1138);
  or csa_tree_add_190_195_groupi_g45735(csa_tree_add_190_195_groupi_n_3426 ,csa_tree_add_190_195_groupi_n_1350 ,csa_tree_add_190_195_groupi_n_758);
  or csa_tree_add_190_195_groupi_g45736(csa_tree_add_190_195_groupi_n_3425 ,csa_tree_add_190_195_groupi_n_1422 ,csa_tree_add_190_195_groupi_n_943);
  or csa_tree_add_190_195_groupi_g45737(csa_tree_add_190_195_groupi_n_3424 ,csa_tree_add_190_195_groupi_n_2482 ,csa_tree_add_190_195_groupi_n_1003);
  nor csa_tree_add_190_195_groupi_g45738(csa_tree_add_190_195_groupi_n_3423 ,csa_tree_add_190_195_groupi_n_2636 ,csa_tree_add_190_195_groupi_n_790);
  nor csa_tree_add_190_195_groupi_g45739(csa_tree_add_190_195_groupi_n_3422 ,csa_tree_add_190_195_groupi_n_767 ,csa_tree_add_190_195_groupi_n_1864);
  nor csa_tree_add_190_195_groupi_g45740(csa_tree_add_190_195_groupi_n_3421 ,csa_tree_add_190_195_groupi_n_1399 ,csa_tree_add_190_195_groupi_n_1924);
  nor csa_tree_add_190_195_groupi_g45741(csa_tree_add_190_195_groupi_n_3420 ,csa_tree_add_190_195_groupi_n_2658 ,csa_tree_add_190_195_groupi_n_937);
  and csa_tree_add_190_195_groupi_g45742(csa_tree_add_190_195_groupi_n_3419 ,csa_tree_add_190_195_groupi_n_913 ,csa_tree_add_190_195_groupi_n_1535);
  nor csa_tree_add_190_195_groupi_g45743(csa_tree_add_190_195_groupi_n_3418 ,csa_tree_add_190_195_groupi_n_2490 ,csa_tree_add_190_195_groupi_n_864);
  or csa_tree_add_190_195_groupi_g45744(csa_tree_add_190_195_groupi_n_3417 ,csa_tree_add_190_195_groupi_n_2638 ,csa_tree_add_190_195_groupi_n_2152);
  or csa_tree_add_190_195_groupi_g45745(csa_tree_add_190_195_groupi_n_3416 ,csa_tree_add_190_195_groupi_n_2654 ,csa_tree_add_190_195_groupi_n_958);
  and csa_tree_add_190_195_groupi_g45746(csa_tree_add_190_195_groupi_n_3415 ,csa_tree_add_190_195_groupi_n_940 ,csa_tree_add_190_195_groupi_n_660);
  or csa_tree_add_190_195_groupi_g45747(csa_tree_add_190_195_groupi_n_3414 ,csa_tree_add_190_195_groupi_n_2500 ,csa_tree_add_190_195_groupi_n_1977);
  nor csa_tree_add_190_195_groupi_g45748(csa_tree_add_190_195_groupi_n_3413 ,csa_tree_add_190_195_groupi_n_480 ,csa_tree_add_190_195_groupi_n_2497);
  and csa_tree_add_190_195_groupi_g45749(csa_tree_add_190_195_groupi_n_3412 ,csa_tree_add_190_195_groupi_n_1114 ,csa_tree_add_190_195_groupi_n_666);
  nor csa_tree_add_190_195_groupi_g45750(csa_tree_add_190_195_groupi_n_3411 ,csa_tree_add_190_195_groupi_n_1545 ,csa_tree_add_190_195_groupi_n_777);
  nor csa_tree_add_190_195_groupi_g45751(csa_tree_add_190_195_groupi_n_3410 ,csa_tree_add_190_195_groupi_n_2608 ,csa_tree_add_190_195_groupi_n_2050);
  or csa_tree_add_190_195_groupi_g45752(csa_tree_add_190_195_groupi_n_3409 ,csa_tree_add_190_195_groupi_n_1436 ,csa_tree_add_190_195_groupi_n_1831);
  or csa_tree_add_190_195_groupi_g45753(csa_tree_add_190_195_groupi_n_3408 ,csa_tree_add_190_195_groupi_n_2503 ,csa_tree_add_190_195_groupi_n_1053);
  and csa_tree_add_190_195_groupi_g45754(csa_tree_add_190_195_groupi_n_3407 ,csa_tree_add_190_195_groupi_n_1054 ,csa_tree_add_190_195_groupi_n_1460);
  and csa_tree_add_190_195_groupi_g45755(csa_tree_add_190_195_groupi_n_3406 ,csa_tree_add_190_195_groupi_n_1068 ,csa_tree_add_190_195_groupi_n_1466);
  nor csa_tree_add_190_195_groupi_g45756(csa_tree_add_190_195_groupi_n_3405 ,csa_tree_add_190_195_groupi_n_2499 ,csa_tree_add_190_195_groupi_n_794);
  or csa_tree_add_190_195_groupi_g45757(csa_tree_add_190_195_groupi_n_3404 ,csa_tree_add_190_195_groupi_n_1564 ,csa_tree_add_190_195_groupi_n_1994);
  nor csa_tree_add_190_195_groupi_g45758(csa_tree_add_190_195_groupi_n_3403 ,csa_tree_add_190_195_groupi_n_2498 ,csa_tree_add_190_195_groupi_n_790);
  nor csa_tree_add_190_195_groupi_g45759(csa_tree_add_190_195_groupi_n_3402 ,csa_tree_add_190_195_groupi_n_2465 ,csa_tree_add_190_195_groupi_n_1969);
  or csa_tree_add_190_195_groupi_g45760(csa_tree_add_190_195_groupi_n_3401 ,csa_tree_add_190_195_groupi_n_2458 ,csa_tree_add_190_195_groupi_n_1831);
  and csa_tree_add_190_195_groupi_g45761(csa_tree_add_190_195_groupi_n_3400 ,csa_tree_add_190_195_groupi_n_2211 ,csa_tree_add_190_195_groupi_n_664);
  or csa_tree_add_190_195_groupi_g45762(csa_tree_add_190_195_groupi_n_3399 ,csa_tree_add_190_195_groupi_n_2482 ,csa_tree_add_190_195_groupi_n_779);
  or csa_tree_add_190_195_groupi_g45763(csa_tree_add_190_195_groupi_n_3398 ,csa_tree_add_190_195_groupi_n_663 ,csa_tree_add_190_195_groupi_n_2211);
  nor csa_tree_add_190_195_groupi_g45764(csa_tree_add_190_195_groupi_n_3397 ,csa_tree_add_190_195_groupi_n_591 ,csa_tree_add_190_195_groupi_n_2436);
  or csa_tree_add_190_195_groupi_g45765(csa_tree_add_190_195_groupi_n_3396 ,csa_tree_add_190_195_groupi_n_1484 ,csa_tree_add_190_195_groupi_n_1996);
  or csa_tree_add_190_195_groupi_g45766(csa_tree_add_190_195_groupi_n_3395 ,csa_tree_add_190_195_groupi_n_2458 ,csa_tree_add_190_195_groupi_n_2041);
  or csa_tree_add_190_195_groupi_g45767(csa_tree_add_190_195_groupi_n_3394 ,csa_tree_add_190_195_groupi_n_1356 ,csa_tree_add_190_195_groupi_n_861);
  or csa_tree_add_190_195_groupi_g45768(csa_tree_add_190_195_groupi_n_3393 ,csa_tree_add_190_195_groupi_n_2615 ,csa_tree_add_190_195_groupi_n_480);
  and csa_tree_add_190_195_groupi_g45769(csa_tree_add_190_195_groupi_n_3392 ,csa_tree_add_190_195_groupi_n_928 ,csa_tree_add_190_195_groupi_n_669);
  nor csa_tree_add_190_195_groupi_g45770(csa_tree_add_190_195_groupi_n_3391 ,csa_tree_add_190_195_groupi_n_2458 ,csa_tree_add_190_195_groupi_n_1923);
  nor csa_tree_add_190_195_groupi_g45771(csa_tree_add_190_195_groupi_n_3390 ,csa_tree_add_190_195_groupi_n_2446 ,csa_tree_add_190_195_groupi_n_1114);
  nor csa_tree_add_190_195_groupi_g45772(csa_tree_add_190_195_groupi_n_3389 ,csa_tree_add_190_195_groupi_n_1440 ,csa_tree_add_190_195_groupi_n_1962);
  or csa_tree_add_190_195_groupi_g45773(csa_tree_add_190_195_groupi_n_3388 ,csa_tree_add_190_195_groupi_n_697 ,csa_tree_add_190_195_groupi_n_1180);
  or csa_tree_add_190_195_groupi_g45774(csa_tree_add_190_195_groupi_n_3387 ,csa_tree_add_190_195_groupi_n_1374 ,csa_tree_add_190_195_groupi_n_414);
  or csa_tree_add_190_195_groupi_g45775(csa_tree_add_190_195_groupi_n_3386 ,csa_tree_add_190_195_groupi_n_2602 ,in55[1]);
  nor csa_tree_add_190_195_groupi_g45776(csa_tree_add_190_195_groupi_n_3385 ,csa_tree_add_190_195_groupi_n_1503 ,csa_tree_add_190_195_groupi_n_416);
  nor csa_tree_add_190_195_groupi_g45777(csa_tree_add_190_195_groupi_n_3384 ,csa_tree_add_190_195_groupi_n_524 ,csa_tree_add_190_195_groupi_n_2456);
  nor csa_tree_add_190_195_groupi_g45778(csa_tree_add_190_195_groupi_n_3383 ,csa_tree_add_190_195_groupi_n_483 ,csa_tree_add_190_195_groupi_n_2628);
  nor csa_tree_add_190_195_groupi_g45779(csa_tree_add_190_195_groupi_n_3382 ,csa_tree_add_190_195_groupi_n_502 ,csa_tree_add_190_195_groupi_n_2455);
  nor csa_tree_add_190_195_groupi_g45780(csa_tree_add_190_195_groupi_n_3381 ,csa_tree_add_190_195_groupi_n_2632 ,csa_tree_add_190_195_groupi_n_2062);
  or csa_tree_add_190_195_groupi_g45781(csa_tree_add_190_195_groupi_n_3380 ,csa_tree_add_190_195_groupi_n_1406 ,csa_tree_add_190_195_groupi_n_1977);
  nor csa_tree_add_190_195_groupi_g45782(csa_tree_add_190_195_groupi_n_3379 ,csa_tree_add_190_195_groupi_n_2582 ,csa_tree_add_190_195_groupi_n_1053);
  or csa_tree_add_190_195_groupi_g45783(csa_tree_add_190_195_groupi_n_3378 ,csa_tree_add_190_195_groupi_n_688 ,csa_tree_add_190_195_groupi_n_380);
  nor csa_tree_add_190_195_groupi_g45784(csa_tree_add_190_195_groupi_n_3377 ,csa_tree_add_190_195_groupi_n_2419 ,csa_tree_add_190_195_groupi_n_1975);
  or csa_tree_add_190_195_groupi_g45785(csa_tree_add_190_195_groupi_n_3376 ,csa_tree_add_190_195_groupi_n_2476 ,csa_tree_add_190_195_groupi_n_960);
  nor csa_tree_add_190_195_groupi_g45786(csa_tree_add_190_195_groupi_n_3375 ,csa_tree_add_190_195_groupi_n_1432 ,csa_tree_add_190_195_groupi_n_1960);
  or csa_tree_add_190_195_groupi_g45787(csa_tree_add_190_195_groupi_n_3374 ,csa_tree_add_190_195_groupi_n_670 ,csa_tree_add_190_195_groupi_n_868);
  or csa_tree_add_190_195_groupi_g45788(csa_tree_add_190_195_groupi_n_3373 ,csa_tree_add_190_195_groupi_n_1395 ,csa_tree_add_190_195_groupi_n_2049);
  or csa_tree_add_190_195_groupi_g45789(csa_tree_add_190_195_groupi_n_3372 ,csa_tree_add_190_195_groupi_n_1528 ,csa_tree_add_190_195_groupi_n_879);
  and csa_tree_add_190_195_groupi_g45790(csa_tree_add_190_195_groupi_n_3371 ,csa_tree_add_190_195_groupi_n_901 ,csa_tree_add_190_195_groupi_n_979);
  or csa_tree_add_190_195_groupi_g45791(csa_tree_add_190_195_groupi_n_3370 ,csa_tree_add_190_195_groupi_n_831 ,csa_tree_add_190_195_groupi_n_1202);
  and csa_tree_add_190_195_groupi_g45792(csa_tree_add_190_195_groupi_n_3369 ,csa_tree_add_190_195_groupi_n_879 ,csa_tree_add_190_195_groupi_n_2473);
  or csa_tree_add_190_195_groupi_g45793(csa_tree_add_190_195_groupi_n_3368 ,csa_tree_add_190_195_groupi_n_2463 ,csa_tree_add_190_195_groupi_n_261);
  or csa_tree_add_190_195_groupi_g45794(csa_tree_add_190_195_groupi_n_3367 ,csa_tree_add_190_195_groupi_n_2448 ,csa_tree_add_190_195_groupi_n_558);
  nor csa_tree_add_190_195_groupi_g45795(csa_tree_add_190_195_groupi_n_3366 ,csa_tree_add_190_195_groupi_n_1418 ,csa_tree_add_190_195_groupi_n_1922);
  nor csa_tree_add_190_195_groupi_g45796(csa_tree_add_190_195_groupi_n_3365 ,csa_tree_add_190_195_groupi_n_2459 ,csa_tree_add_190_195_groupi_n_2158);
  nor csa_tree_add_190_195_groupi_g45797(csa_tree_add_190_195_groupi_n_3364 ,csa_tree_add_190_195_groupi_n_2625 ,csa_tree_add_190_195_groupi_n_1072);
  or csa_tree_add_190_195_groupi_g45798(csa_tree_add_190_195_groupi_n_3363 ,csa_tree_add_190_195_groupi_n_2605 ,csa_tree_add_190_195_groupi_n_411);
  or csa_tree_add_190_195_groupi_g45799(csa_tree_add_190_195_groupi_n_3362 ,csa_tree_add_190_195_groupi_n_2469 ,csa_tree_add_190_195_groupi_n_867);
  nor csa_tree_add_190_195_groupi_g45800(csa_tree_add_190_195_groupi_n_3361 ,csa_tree_add_190_195_groupi_n_1384 ,csa_tree_add_190_195_groupi_n_1921);
  or csa_tree_add_190_195_groupi_g45801(csa_tree_add_190_195_groupi_n_3360 ,csa_tree_add_190_195_groupi_n_1496 ,csa_tree_add_190_195_groupi_n_2049);
  nor csa_tree_add_190_195_groupi_g45802(csa_tree_add_190_195_groupi_n_3359 ,csa_tree_add_190_195_groupi_n_1533 ,csa_tree_add_190_195_groupi_n_788);
  nor csa_tree_add_190_195_groupi_g45803(csa_tree_add_190_195_groupi_n_3358 ,csa_tree_add_190_195_groupi_n_1401 ,csa_tree_add_190_195_groupi_n_1960);
  nor csa_tree_add_190_195_groupi_g45804(csa_tree_add_190_195_groupi_n_3357 ,csa_tree_add_190_195_groupi_n_348 ,csa_tree_add_190_195_groupi_n_2622);
  and csa_tree_add_190_195_groupi_g45805(csa_tree_add_190_195_groupi_n_3356 ,csa_tree_add_190_195_groupi_n_964 ,csa_tree_add_190_195_groupi_n_768);
  or csa_tree_add_190_195_groupi_g45806(csa_tree_add_190_195_groupi_n_3355 ,csa_tree_add_190_195_groupi_n_2619 ,csa_tree_add_190_195_groupi_n_840);
  or csa_tree_add_190_195_groupi_g45807(csa_tree_add_190_195_groupi_n_3354 ,csa_tree_add_190_195_groupi_n_1474 ,csa_tree_add_190_195_groupi_n_927);
  or csa_tree_add_190_195_groupi_g45808(csa_tree_add_190_195_groupi_n_3353 ,csa_tree_add_190_195_groupi_n_2577 ,csa_tree_add_190_195_groupi_n_2210);
  and csa_tree_add_190_195_groupi_g45809(csa_tree_add_190_195_groupi_n_3352 ,csa_tree_add_190_195_groupi_n_1269 ,csa_tree_add_190_195_groupi_n_697);
  or csa_tree_add_190_195_groupi_g45810(csa_tree_add_190_195_groupi_n_3351 ,csa_tree_add_190_195_groupi_n_1485 ,csa_tree_add_190_195_groupi_n_2063);
  or csa_tree_add_190_195_groupi_g45811(csa_tree_add_190_195_groupi_n_3350 ,csa_tree_add_190_195_groupi_n_739 ,csa_tree_add_190_195_groupi_n_2060);
  or csa_tree_add_190_195_groupi_g45812(csa_tree_add_190_195_groupi_n_3349 ,csa_tree_add_190_195_groupi_n_1366 ,csa_tree_add_190_195_groupi_n_904);
  nor csa_tree_add_190_195_groupi_g45813(csa_tree_add_190_195_groupi_n_3348 ,csa_tree_add_190_195_groupi_n_1424 ,csa_tree_add_190_195_groupi_n_393);
  nor csa_tree_add_190_195_groupi_g45814(csa_tree_add_190_195_groupi_n_3347 ,csa_tree_add_190_195_groupi_n_1564 ,csa_tree_add_190_195_groupi_n_2061);
  nor csa_tree_add_190_195_groupi_g45815(csa_tree_add_190_195_groupi_n_3346 ,csa_tree_add_190_195_groupi_n_526 ,csa_tree_add_190_195_groupi_n_1430);
  nor csa_tree_add_190_195_groupi_g45816(csa_tree_add_190_195_groupi_n_3345 ,csa_tree_add_190_195_groupi_n_343 ,csa_tree_add_190_195_groupi_n_2443);
  nor csa_tree_add_190_195_groupi_g45817(csa_tree_add_190_195_groupi_n_3344 ,csa_tree_add_190_195_groupi_n_504 ,csa_tree_add_190_195_groupi_n_2631);
  or csa_tree_add_190_195_groupi_g45818(csa_tree_add_190_195_groupi_n_3343 ,csa_tree_add_190_195_groupi_n_2476 ,csa_tree_add_190_195_groupi_n_295);
  or csa_tree_add_190_195_groupi_g45819(csa_tree_add_190_195_groupi_n_3342 ,csa_tree_add_190_195_groupi_n_2467 ,csa_tree_add_190_195_groupi_n_358);
  nor csa_tree_add_190_195_groupi_g45820(csa_tree_add_190_195_groupi_n_3341 ,csa_tree_add_190_195_groupi_n_516 ,csa_tree_add_190_195_groupi_n_2618);
  or csa_tree_add_190_195_groupi_g45821(csa_tree_add_190_195_groupi_n_3340 ,csa_tree_add_190_195_groupi_n_1360 ,csa_tree_add_190_195_groupi_n_910);
  nor csa_tree_add_190_195_groupi_g45822(csa_tree_add_190_195_groupi_n_3339 ,csa_tree_add_190_195_groupi_n_1560 ,csa_tree_add_190_195_groupi_n_1973);
  or csa_tree_add_190_195_groupi_g45823(csa_tree_add_190_195_groupi_n_3338 ,csa_tree_add_190_195_groupi_n_782 ,csa_tree_add_190_195_groupi_n_1988);
  or csa_tree_add_190_195_groupi_g45824(csa_tree_add_190_195_groupi_n_3337 ,csa_tree_add_190_195_groupi_n_2624 ,csa_tree_add_190_195_groupi_n_1922);
  or csa_tree_add_190_195_groupi_g45825(csa_tree_add_190_195_groupi_n_3336 ,csa_tree_add_190_195_groupi_n_2610 ,csa_tree_add_190_195_groupi_n_268);
  nor csa_tree_add_190_195_groupi_g45826(csa_tree_add_190_195_groupi_n_3335 ,csa_tree_add_190_195_groupi_n_2617 ,csa_tree_add_190_195_groupi_n_422);
  or csa_tree_add_190_195_groupi_g45827(csa_tree_add_190_195_groupi_n_3334 ,csa_tree_add_190_195_groupi_n_2457 ,csa_tree_add_190_195_groupi_n_2211);
  nor csa_tree_add_190_195_groupi_g45828(csa_tree_add_190_195_groupi_n_3333 ,csa_tree_add_190_195_groupi_n_2633 ,csa_tree_add_190_195_groupi_n_2214);
  or csa_tree_add_190_195_groupi_g45829(csa_tree_add_190_195_groupi_n_3332 ,csa_tree_add_190_195_groupi_n_1487 ,csa_tree_add_190_195_groupi_n_1026);
  nor csa_tree_add_190_195_groupi_g45830(csa_tree_add_190_195_groupi_n_3331 ,csa_tree_add_190_195_groupi_n_2479 ,csa_tree_add_190_195_groupi_n_892);
  nor csa_tree_add_190_195_groupi_g45831(csa_tree_add_190_195_groupi_n_3330 ,csa_tree_add_190_195_groupi_n_2611 ,csa_tree_add_190_195_groupi_n_485);
  nor csa_tree_add_190_195_groupi_g45832(csa_tree_add_190_195_groupi_n_3329 ,csa_tree_add_190_195_groupi_n_1520 ,csa_tree_add_190_195_groupi_n_1973);
  or csa_tree_add_190_195_groupi_g45833(csa_tree_add_190_195_groupi_n_3328 ,csa_tree_add_190_195_groupi_n_2612 ,csa_tree_add_190_195_groupi_n_2040);
  or csa_tree_add_190_195_groupi_g45834(csa_tree_add_190_195_groupi_n_3327 ,csa_tree_add_190_195_groupi_n_1531 ,csa_tree_add_190_195_groupi_n_1047);
  or csa_tree_add_190_195_groupi_g45835(csa_tree_add_190_195_groupi_n_3326 ,csa_tree_add_190_195_groupi_n_2624 ,csa_tree_add_190_195_groupi_n_991);
  or csa_tree_add_190_195_groupi_g45836(csa_tree_add_190_195_groupi_n_3325 ,csa_tree_add_190_195_groupi_n_675 ,csa_tree_add_190_195_groupi_n_880);
  nor csa_tree_add_190_195_groupi_g45837(csa_tree_add_190_195_groupi_n_3324 ,csa_tree_add_190_195_groupi_n_1368 ,csa_tree_add_190_195_groupi_n_877);
  or csa_tree_add_190_195_groupi_g45838(csa_tree_add_190_195_groupi_n_3323 ,csa_tree_add_190_195_groupi_n_704 ,csa_tree_add_190_195_groupi_n_710);
  or csa_tree_add_190_195_groupi_g45839(csa_tree_add_190_195_groupi_n_3322 ,csa_tree_add_190_195_groupi_n_1471 ,csa_tree_add_190_195_groupi_n_936);
  nor csa_tree_add_190_195_groupi_g45840(csa_tree_add_190_195_groupi_n_3321 ,csa_tree_add_190_195_groupi_n_2596 ,csa_tree_add_190_195_groupi_n_786);
  nor csa_tree_add_190_195_groupi_g45841(csa_tree_add_190_195_groupi_n_3320 ,csa_tree_add_190_195_groupi_n_2449 ,csa_tree_add_190_195_groupi_n_1923);
  or csa_tree_add_190_195_groupi_g45842(csa_tree_add_190_195_groupi_n_3319 ,csa_tree_add_190_195_groupi_n_2463 ,csa_tree_add_190_195_groupi_n_924);
  or csa_tree_add_190_195_groupi_g45843(csa_tree_add_190_195_groupi_n_3318 ,csa_tree_add_190_195_groupi_n_1488 ,csa_tree_add_190_195_groupi_n_1105);
  nor csa_tree_add_190_195_groupi_g45844(csa_tree_add_190_195_groupi_n_3317 ,csa_tree_add_190_195_groupi_n_508 ,csa_tree_add_190_195_groupi_n_2479);
  nor csa_tree_add_190_195_groupi_g45845(csa_tree_add_190_195_groupi_n_3316 ,csa_tree_add_190_195_groupi_n_2464 ,csa_tree_add_190_195_groupi_n_1255);
  or csa_tree_add_190_195_groupi_g45846(csa_tree_add_190_195_groupi_n_3315 ,csa_tree_add_190_195_groupi_n_2620 ,csa_tree_add_190_195_groupi_n_1214);
  or csa_tree_add_190_195_groupi_g45847(csa_tree_add_190_195_groupi_n_3314 ,csa_tree_add_190_195_groupi_n_2626 ,csa_tree_add_190_195_groupi_n_1051);
  nor csa_tree_add_190_195_groupi_g45848(csa_tree_add_190_195_groupi_n_3313 ,csa_tree_add_190_195_groupi_n_1358 ,csa_tree_add_190_195_groupi_n_1083);
  or csa_tree_add_190_195_groupi_g45849(csa_tree_add_190_195_groupi_n_3312 ,csa_tree_add_190_195_groupi_n_1415 ,csa_tree_add_190_195_groupi_n_1149);
  nor csa_tree_add_190_195_groupi_g45850(csa_tree_add_190_195_groupi_n_3311 ,csa_tree_add_190_195_groupi_n_2587 ,csa_tree_add_190_195_groupi_n_1918);
  nor csa_tree_add_190_195_groupi_g45851(csa_tree_add_190_195_groupi_n_3310 ,csa_tree_add_190_195_groupi_n_1408 ,csa_tree_add_190_195_groupi_n_1976);
  nor csa_tree_add_190_195_groupi_g45852(csa_tree_add_190_195_groupi_n_3309 ,csa_tree_add_190_195_groupi_n_1570 ,csa_tree_add_190_195_groupi_n_2055);
  or csa_tree_add_190_195_groupi_g45853(csa_tree_add_190_195_groupi_n_3308 ,csa_tree_add_190_195_groupi_n_694 ,csa_tree_add_190_195_groupi_n_2060);
  or csa_tree_add_190_195_groupi_g45854(csa_tree_add_190_195_groupi_n_3307 ,csa_tree_add_190_195_groupi_n_2600 ,in55[12]);
  nor csa_tree_add_190_195_groupi_g45855(csa_tree_add_190_195_groupi_n_3306 ,csa_tree_add_190_195_groupi_n_2600 ,in55[14]);
  nor csa_tree_add_190_195_groupi_g45856(csa_tree_add_190_195_groupi_n_3305 ,csa_tree_add_190_195_groupi_n_2595 ,in55[10]);
  or csa_tree_add_190_195_groupi_g45857(csa_tree_add_190_195_groupi_n_3304 ,csa_tree_add_190_195_groupi_n_1346 ,in55[10]);
  nor csa_tree_add_190_195_groupi_g45858(csa_tree_add_190_195_groupi_n_3303 ,csa_tree_add_190_195_groupi_n_2434 ,in55[8]);
  nor csa_tree_add_190_195_groupi_g45859(csa_tree_add_190_195_groupi_n_3302 ,csa_tree_add_190_195_groupi_n_2599 ,in55[11]);
  or csa_tree_add_190_195_groupi_g45860(csa_tree_add_190_195_groupi_n_3301 ,csa_tree_add_190_195_groupi_n_2593 ,in55[3]);
  nor csa_tree_add_190_195_groupi_g45861(csa_tree_add_190_195_groupi_n_3300 ,csa_tree_add_190_195_groupi_n_412 ,csa_tree_add_190_195_groupi_n_2212);
  or csa_tree_add_190_195_groupi_g45862(csa_tree_add_190_195_groupi_n_3299 ,csa_tree_add_190_195_groupi_n_2423 ,in55[13]);
  nor csa_tree_add_190_195_groupi_g45863(csa_tree_add_190_195_groupi_n_3298 ,csa_tree_add_190_195_groupi_n_519 ,in55[0]);
  nor csa_tree_add_190_195_groupi_g45864(csa_tree_add_190_195_groupi_n_3297 ,in55[12] ,in55[11]);
  or csa_tree_add_190_195_groupi_g45865(csa_tree_add_190_195_groupi_n_3296 ,csa_tree_add_190_195_groupi_n_2428 ,in55[1]);
  nor csa_tree_add_190_195_groupi_g45866(csa_tree_add_190_195_groupi_n_3295 ,csa_tree_add_190_195_groupi_n_2425 ,in55[5]);
  nor csa_tree_add_190_195_groupi_g45867(csa_tree_add_190_195_groupi_n_3294 ,csa_tree_add_190_195_groupi_n_1346 ,in55[12]);
  or csa_tree_add_190_195_groupi_g45868(csa_tree_add_190_195_groupi_n_3293 ,csa_tree_add_190_195_groupi_n_1336 ,in55[9]);
  or csa_tree_add_190_195_groupi_g45869(csa_tree_add_190_195_groupi_n_3292 ,csa_tree_add_190_195_groupi_n_2592 ,in55[7]);
  or csa_tree_add_190_195_groupi_g45870(csa_tree_add_190_195_groupi_n_3291 ,csa_tree_add_190_195_groupi_n_1523 ,csa_tree_add_190_195_groupi_n_319);
  and csa_tree_add_190_195_groupi_g45871(csa_tree_add_190_195_groupi_n_3290 ,csa_tree_add_190_195_groupi_n_360 ,csa_tree_add_190_195_groupi_n_1522);
  or csa_tree_add_190_195_groupi_g45872(csa_tree_add_190_195_groupi_n_3289 ,csa_tree_add_190_195_groupi_n_1340 ,in55[14]);
  or csa_tree_add_190_195_groupi_g45873(csa_tree_add_190_195_groupi_n_3288 ,csa_tree_add_190_195_groupi_n_1513 ,csa_tree_add_190_195_groupi_n_885);
  nor csa_tree_add_190_195_groupi_g45874(csa_tree_add_190_195_groupi_n_3287 ,csa_tree_add_190_195_groupi_n_2423 ,in55[9]);
  nor csa_tree_add_190_195_groupi_g45875(csa_tree_add_190_195_groupi_n_3286 ,csa_tree_add_190_195_groupi_n_2430 ,in55[7]);
  or csa_tree_add_190_195_groupi_g45876(csa_tree_add_190_195_groupi_n_3285 ,csa_tree_add_190_195_groupi_n_2431 ,in55[2]);
  or csa_tree_add_190_195_groupi_g45877(csa_tree_add_190_195_groupi_n_3284 ,csa_tree_add_190_195_groupi_n_2430 ,in55[11]);
  or csa_tree_add_190_195_groupi_g45878(csa_tree_add_190_195_groupi_n_3283 ,csa_tree_add_190_195_groupi_n_1667 ,csa_tree_add_190_195_groupi_n_2209);
  or csa_tree_add_190_195_groupi_g45879(csa_tree_add_190_195_groupi_n_3282 ,csa_tree_add_190_195_groupi_n_1487 ,csa_tree_add_190_195_groupi_n_837);
  nor csa_tree_add_190_195_groupi_g45880(csa_tree_add_190_195_groupi_n_3281 ,csa_tree_add_190_195_groupi_n_531 ,csa_tree_add_190_195_groupi_n_1468);
  nor csa_tree_add_190_195_groupi_g45881(csa_tree_add_190_195_groupi_n_3280 ,csa_tree_add_190_195_groupi_n_2590 ,in55[4]);
  nor csa_tree_add_190_195_groupi_g45882(csa_tree_add_190_195_groupi_n_3279 ,csa_tree_add_190_195_groupi_n_1469 ,csa_tree_add_190_195_groupi_n_1071);
  nor csa_tree_add_190_195_groupi_g45883(csa_tree_add_190_195_groupi_n_3278 ,csa_tree_add_190_195_groupi_n_2596 ,in55[6]);
  nor csa_tree_add_190_195_groupi_g45884(csa_tree_add_190_195_groupi_n_3277 ,csa_tree_add_190_195_groupi_n_1511 ,csa_tree_add_190_195_groupi_n_1283);
  nor csa_tree_add_190_195_groupi_g45885(csa_tree_add_190_195_groupi_n_3276 ,csa_tree_add_190_195_groupi_n_1344 ,in55[0]);
  or csa_tree_add_190_195_groupi_g45886(csa_tree_add_190_195_groupi_n_3275 ,csa_tree_add_190_195_groupi_n_1447 ,csa_tree_add_190_195_groupi_n_315);
  nor csa_tree_add_190_195_groupi_g45887(csa_tree_add_190_195_groupi_n_3274 ,csa_tree_add_190_195_groupi_n_1380 ,csa_tree_add_190_195_groupi_n_234);
  or csa_tree_add_190_195_groupi_g45888(csa_tree_add_190_195_groupi_n_3273 ,csa_tree_add_190_195_groupi_n_2589 ,in55[2]);
  or csa_tree_add_190_195_groupi_g45889(csa_tree_add_190_195_groupi_n_3272 ,csa_tree_add_190_195_groupi_n_1440 ,csa_tree_add_190_195_groupi_n_547);
  or csa_tree_add_190_195_groupi_g45890(csa_tree_add_190_195_groupi_n_3271 ,csa_tree_add_190_195_groupi_n_1453 ,in55[15]);
  or csa_tree_add_190_195_groupi_g45891(csa_tree_add_190_195_groupi_n_3270 ,csa_tree_add_190_195_groupi_n_1338 ,in55[15]);
  nor csa_tree_add_190_195_groupi_g45892(csa_tree_add_190_195_groupi_n_3269 ,csa_tree_add_190_195_groupi_n_708 ,in55[11]);
  nor csa_tree_add_190_195_groupi_g45893(csa_tree_add_190_195_groupi_n_3268 ,csa_tree_add_190_195_groupi_n_2424 ,csa_tree_add_190_195_groupi_n_1244);
  or csa_tree_add_190_195_groupi_g45894(csa_tree_add_190_195_groupi_n_3267 ,csa_tree_add_190_195_groupi_n_1525 ,csa_tree_add_190_195_groupi_n_235);
  nor csa_tree_add_190_195_groupi_g45895(csa_tree_add_190_195_groupi_n_3266 ,csa_tree_add_190_195_groupi_n_514 ,csa_tree_add_190_195_groupi_n_1453);
  nor csa_tree_add_190_195_groupi_g45896(csa_tree_add_190_195_groupi_n_3265 ,csa_tree_add_190_195_groupi_n_1514 ,csa_tree_add_190_195_groupi_n_1228);
  nor csa_tree_add_190_195_groupi_g45897(csa_tree_add_190_195_groupi_n_3264 ,csa_tree_add_190_195_groupi_n_564 ,csa_tree_add_190_195_groupi_n_1410);
  or csa_tree_add_190_195_groupi_g45898(csa_tree_add_190_195_groupi_n_3263 ,csa_tree_add_190_195_groupi_n_1415 ,csa_tree_add_190_195_groupi_n_1234);
  nor csa_tree_add_190_195_groupi_g45899(csa_tree_add_190_195_groupi_n_3262 ,csa_tree_add_190_195_groupi_n_458 ,csa_tree_add_190_195_groupi_n_689);
  or csa_tree_add_190_195_groupi_g45900(csa_tree_add_190_195_groupi_n_3261 ,csa_tree_add_190_195_groupi_n_215 ,csa_tree_add_190_195_groupi_n_627);
  or csa_tree_add_190_195_groupi_g45901(csa_tree_add_190_195_groupi_n_3260 ,csa_tree_add_190_195_groupi_n_2428 ,csa_tree_add_190_195_groupi_n_2557);
  and csa_tree_add_190_195_groupi_g45902(csa_tree_add_190_195_groupi_n_3259 ,csa_tree_add_190_195_groupi_n_615 ,csa_tree_add_190_195_groupi_n_1776);
  nor csa_tree_add_190_195_groupi_g45903(csa_tree_add_190_195_groupi_n_3258 ,csa_tree_add_190_195_groupi_n_1245 ,csa_tree_add_190_195_groupi_n_906);
  nor csa_tree_add_190_195_groupi_g45904(csa_tree_add_190_195_groupi_n_3257 ,csa_tree_add_190_195_groupi_n_798 ,csa_tree_add_190_195_groupi_n_1808);
  or csa_tree_add_190_195_groupi_g45905(csa_tree_add_190_195_groupi_n_3256 ,in61[15] ,in59[15]);
  and csa_tree_add_190_195_groupi_g45906(csa_tree_add_190_195_groupi_n_3255 ,csa_tree_add_190_195_groupi_n_1999 ,csa_tree_add_190_195_groupi_n_2064);
  nor csa_tree_add_190_195_groupi_g45907(csa_tree_add_190_195_groupi_n_3254 ,csa_tree_add_190_195_groupi_n_1108 ,csa_tree_add_190_195_groupi_n_477);
  and csa_tree_add_190_195_groupi_g45908(csa_tree_add_190_195_groupi_n_3253 ,csa_tree_add_190_195_groupi_n_529 ,csa_tree_add_190_195_groupi_n_997);
  or csa_tree_add_190_195_groupi_g45909(csa_tree_add_190_195_groupi_n_3252 ,csa_tree_add_190_195_groupi_n_328 ,csa_tree_add_190_195_groupi_n_1962);
  and csa_tree_add_190_195_groupi_g45910(csa_tree_add_190_195_groupi_n_3251 ,csa_tree_add_190_195_groupi_n_1242 ,csa_tree_add_190_195_groupi_n_1177);
  or csa_tree_add_190_195_groupi_g45911(csa_tree_add_190_195_groupi_n_3250 ,csa_tree_add_190_195_groupi_n_2438 ,csa_tree_add_190_195_groupi_n_2500);
  and csa_tree_add_190_195_groupi_g45912(csa_tree_add_190_195_groupi_n_3249 ,csa_tree_add_190_195_groupi_n_1153 ,csa_tree_add_190_195_groupi_n_1074);
  and csa_tree_add_190_195_groupi_g45913(csa_tree_add_190_195_groupi_n_3248 ,csa_tree_add_190_195_groupi_n_612 ,csa_tree_add_190_195_groupi_n_2213);
  or csa_tree_add_190_195_groupi_g45914(csa_tree_add_190_195_groupi_n_3247 ,csa_tree_add_190_195_groupi_n_1045 ,csa_tree_add_190_195_groupi_n_1818);
  or csa_tree_add_190_195_groupi_g45915(csa_tree_add_190_195_groupi_n_3246 ,csa_tree_add_190_195_groupi_n_473 ,csa_tree_add_190_195_groupi_n_1862);
  and csa_tree_add_190_195_groupi_g45916(csa_tree_add_190_195_groupi_n_3245 ,csa_tree_add_190_195_groupi_n_621 ,csa_tree_add_190_195_groupi_n_531);
  nor csa_tree_add_190_195_groupi_g45917(csa_tree_add_190_195_groupi_n_3244 ,csa_tree_add_190_195_groupi_n_1999 ,csa_tree_add_190_195_groupi_n_1837);
  nor csa_tree_add_190_195_groupi_g45918(csa_tree_add_190_195_groupi_n_3243 ,csa_tree_add_190_195_groupi_n_978 ,csa_tree_add_190_195_groupi_n_1554);
  or csa_tree_add_190_195_groupi_g45919(csa_tree_add_190_195_groupi_n_3242 ,csa_tree_add_190_195_groupi_n_1057 ,csa_tree_add_190_195_groupi_n_1777);
  or csa_tree_add_190_195_groupi_g45920(csa_tree_add_190_195_groupi_n_3241 ,csa_tree_add_190_195_groupi_n_691 ,csa_tree_add_190_195_groupi_n_2554);
  and csa_tree_add_190_195_groupi_g45921(csa_tree_add_190_195_groupi_n_3240 ,csa_tree_add_190_195_groupi_n_871 ,csa_tree_add_190_195_groupi_n_945);
  nor csa_tree_add_190_195_groupi_g45922(csa_tree_add_190_195_groupi_n_3239 ,csa_tree_add_190_195_groupi_n_1247 ,csa_tree_add_190_195_groupi_n_1048);
  nor csa_tree_add_190_195_groupi_g45923(csa_tree_add_190_195_groupi_n_3238 ,csa_tree_add_190_195_groupi_n_356 ,csa_tree_add_190_195_groupi_n_1876);
  or csa_tree_add_190_195_groupi_g45924(csa_tree_add_190_195_groupi_n_3237 ,csa_tree_add_190_195_groupi_n_2430 ,csa_tree_add_190_195_groupi_n_2561);
  nor csa_tree_add_190_195_groupi_g45925(csa_tree_add_190_195_groupi_n_3236 ,csa_tree_add_190_195_groupi_n_1961 ,csa_tree_add_190_195_groupi_n_1945);
  nor csa_tree_add_190_195_groupi_g45926(csa_tree_add_190_195_groupi_n_3235 ,csa_tree_add_190_195_groupi_n_423 ,csa_tree_add_190_195_groupi_n_806);
  nor csa_tree_add_190_195_groupi_g45927(csa_tree_add_190_195_groupi_n_3234 ,csa_tree_add_190_195_groupi_n_2082 ,csa_tree_add_190_195_groupi_n_1742);
  and csa_tree_add_190_195_groupi_g45928(csa_tree_add_190_195_groupi_n_3233 ,csa_tree_add_190_195_groupi_n_1888 ,csa_tree_add_190_195_groupi_n_1833);
  nor csa_tree_add_190_195_groupi_g45929(csa_tree_add_190_195_groupi_n_3232 ,csa_tree_add_190_195_groupi_n_853 ,csa_tree_add_190_195_groupi_n_304);
  or csa_tree_add_190_195_groupi_g45930(csa_tree_add_190_195_groupi_n_3231 ,csa_tree_add_190_195_groupi_n_2676 ,csa_tree_add_190_195_groupi_n_2449);
  and csa_tree_add_190_195_groupi_g45931(csa_tree_add_190_195_groupi_n_3230 ,csa_tree_add_190_195_groupi_n_457 ,csa_tree_add_190_195_groupi_n_1182);
  or csa_tree_add_190_195_groupi_g45932(csa_tree_add_190_195_groupi_n_3229 ,csa_tree_add_190_195_groupi_n_1071 ,csa_tree_add_190_195_groupi_n_2152);
  or csa_tree_add_190_195_groupi_g45933(csa_tree_add_190_195_groupi_n_3729 ,csa_tree_add_190_195_groupi_n_2526 ,csa_tree_add_190_195_groupi_n_1907);
  or csa_tree_add_190_195_groupi_g45934(csa_tree_add_190_195_groupi_n_3727 ,csa_tree_add_190_195_groupi_n_2706 ,csa_tree_add_190_195_groupi_n_2677);
  nor csa_tree_add_190_195_groupi_g45935(csa_tree_add_190_195_groupi_n_3228 ,csa_tree_add_190_195_groupi_n_2551 ,csa_tree_add_190_195_groupi_n_1916);
  or csa_tree_add_190_195_groupi_g45936(csa_tree_add_190_195_groupi_n_3227 ,csa_tree_add_190_195_groupi_n_2377 ,csa_tree_add_190_195_groupi_n_1842);
  and csa_tree_add_190_195_groupi_g45937(csa_tree_add_190_195_groupi_n_3726 ,csa_tree_add_190_195_groupi_n_1584 ,csa_tree_add_190_195_groupi_n_1450);
  and csa_tree_add_190_195_groupi_g45938(csa_tree_add_190_195_groupi_n_3724 ,csa_tree_add_190_195_groupi_n_1210 ,csa_tree_add_190_195_groupi_n_2716);
  and csa_tree_add_190_195_groupi_g45939(csa_tree_add_190_195_groupi_n_3723 ,csa_tree_add_190_195_groupi_n_1911 ,csa_tree_add_190_195_groupi_n_2512);
  or csa_tree_add_190_195_groupi_g45940(csa_tree_add_190_195_groupi_n_3722 ,csa_tree_add_190_195_groupi_n_2512 ,csa_tree_add_190_195_groupi_n_1911);
  and csa_tree_add_190_195_groupi_g45941(csa_tree_add_190_195_groupi_n_3720 ,csa_tree_add_190_195_groupi_n_1971 ,csa_tree_add_190_195_groupi_n_2521);
  and csa_tree_add_190_195_groupi_g45942(csa_tree_add_190_195_groupi_n_3718 ,csa_tree_add_190_195_groupi_n_1259 ,csa_tree_add_190_195_groupi_n_2522);
  or csa_tree_add_190_195_groupi_g45943(csa_tree_add_190_195_groupi_n_3716 ,csa_tree_add_190_195_groupi_n_2522 ,csa_tree_add_190_195_groupi_n_386);
  and csa_tree_add_190_195_groupi_g45944(csa_tree_add_190_195_groupi_n_3714 ,csa_tree_add_190_195_groupi_n_846 ,csa_tree_add_190_195_groupi_n_1378);
  and csa_tree_add_190_195_groupi_g45945(csa_tree_add_190_195_groupi_n_3713 ,csa_tree_add_190_195_groupi_n_1865 ,csa_tree_add_190_195_groupi_n_2692);
  or csa_tree_add_190_195_groupi_g45946(csa_tree_add_190_195_groupi_n_3711 ,csa_tree_add_190_195_groupi_n_1378 ,csa_tree_add_190_195_groupi_n_847);
  and csa_tree_add_190_195_groupi_g45947(csa_tree_add_190_195_groupi_n_3710 ,csa_tree_add_190_195_groupi_n_291 ,csa_tree_add_190_195_groupi_n_561);
  and csa_tree_add_190_195_groupi_g45948(csa_tree_add_190_195_groupi_n_3709 ,csa_tree_add_190_195_groupi_n_1907 ,csa_tree_add_190_195_groupi_n_2526);
  or csa_tree_add_190_195_groupi_g45949(csa_tree_add_190_195_groupi_n_3708 ,csa_tree_add_190_195_groupi_n_1449 ,csa_tree_add_190_195_groupi_n_1583);
  or csa_tree_add_190_195_groupi_g45950(csa_tree_add_190_195_groupi_n_3706 ,csa_tree_add_190_195_groupi_n_2716 ,csa_tree_add_190_195_groupi_n_340);
  or csa_tree_add_190_195_groupi_g45951(csa_tree_add_190_195_groupi_n_3705 ,csa_tree_add_190_195_groupi_n_2428 ,in55[4]);
  or csa_tree_add_190_195_groupi_g45952(csa_tree_add_190_195_groupi_n_3704 ,csa_tree_add_190_195_groupi_n_2434 ,in55[1]);
  and csa_tree_add_190_195_groupi_g45953(csa_tree_add_190_195_groupi_n_3702 ,in55[5] ,csa_tree_add_190_195_groupi_n_2434);
  and csa_tree_add_190_195_groupi_g45954(csa_tree_add_190_195_groupi_n_3701 ,csa_tree_add_190_195_groupi_n_1702 ,csa_tree_add_190_195_groupi_n_1376);
  and csa_tree_add_190_195_groupi_g45955(csa_tree_add_190_195_groupi_n_3699 ,in60[15] ,csa_tree_add_190_195_groupi_n_2731);
  and csa_tree_add_190_195_groupi_g45956(csa_tree_add_190_195_groupi_n_3697 ,in55[15] ,csa_tree_add_190_195_groupi_n_2599);
  or csa_tree_add_190_195_groupi_g45957(csa_tree_add_190_195_groupi_n_3696 ,csa_tree_add_190_195_groupi_n_2568 ,in55[9]);
  or csa_tree_add_190_195_groupi_g45958(csa_tree_add_190_195_groupi_n_3695 ,csa_tree_add_190_195_groupi_n_2572 ,in55[10]);
  and csa_tree_add_190_195_groupi_g45959(csa_tree_add_190_195_groupi_n_3694 ,in56[3] ,csa_tree_add_190_195_groupi_n_2571);
  and csa_tree_add_190_195_groupi_g45960(csa_tree_add_190_195_groupi_n_3693 ,csa_tree_add_190_195_groupi_n_1698 ,csa_tree_add_190_195_groupi_n_2718);
  and csa_tree_add_190_195_groupi_g45961(csa_tree_add_190_195_groupi_n_3690 ,csa_tree_add_190_195_groupi_n_1193 ,csa_tree_add_190_195_groupi_n_2733);
  not csa_tree_add_190_195_groupi_g45962(csa_tree_add_190_195_groupi_n_3224 ,csa_tree_add_190_195_groupi_n_3223);
  not csa_tree_add_190_195_groupi_g45963(csa_tree_add_190_195_groupi_n_3222 ,csa_tree_add_190_195_groupi_n_3221);
  not csa_tree_add_190_195_groupi_g45964(csa_tree_add_190_195_groupi_n_3220 ,csa_tree_add_190_195_groupi_n_3219);
  not csa_tree_add_190_195_groupi_g45965(csa_tree_add_190_195_groupi_n_3216 ,csa_tree_add_190_195_groupi_n_3215);
  not csa_tree_add_190_195_groupi_g45966(csa_tree_add_190_195_groupi_n_3214 ,csa_tree_add_190_195_groupi_n_3213);
  not csa_tree_add_190_195_groupi_g45967(csa_tree_add_190_195_groupi_n_3212 ,csa_tree_add_190_195_groupi_n_3211);
  not csa_tree_add_190_195_groupi_g45968(csa_tree_add_190_195_groupi_n_3204 ,csa_tree_add_190_195_groupi_n_3203);
  or csa_tree_add_190_195_groupi_g45971(csa_tree_add_190_195_groupi_n_3199 ,csa_tree_add_190_195_groupi_n_1490 ,csa_tree_add_190_195_groupi_n_1195);
  nor csa_tree_add_190_195_groupi_g45972(csa_tree_add_190_195_groupi_n_3198 ,csa_tree_add_190_195_groupi_n_1444 ,csa_tree_add_190_195_groupi_n_2441);
  or csa_tree_add_190_195_groupi_g45973(csa_tree_add_190_195_groupi_n_3197 ,csa_tree_add_190_195_groupi_n_2425 ,csa_tree_add_190_195_groupi_n_2724);
  nor csa_tree_add_190_195_groupi_g45974(csa_tree_add_190_195_groupi_n_3196 ,csa_tree_add_190_195_groupi_n_1828 ,csa_tree_add_190_195_groupi_n_991);
  or csa_tree_add_190_195_groupi_g45975(csa_tree_add_190_195_groupi_n_3195 ,csa_tree_add_190_195_groupi_n_188 ,csa_tree_add_190_195_groupi_n_999);
  or csa_tree_add_190_195_groupi_g45976(csa_tree_add_190_195_groupi_n_3194 ,csa_tree_add_190_195_groupi_n_1511 ,csa_tree_add_190_195_groupi_n_2459);
  nor csa_tree_add_190_195_groupi_g45977(csa_tree_add_190_195_groupi_n_3193 ,csa_tree_add_190_195_groupi_n_2578 ,csa_tree_add_190_195_groupi_n_679);
  nor csa_tree_add_190_195_groupi_g45978(csa_tree_add_190_195_groupi_n_3192 ,csa_tree_add_190_195_groupi_n_2406 ,csa_tree_add_190_195_groupi_n_2535);
  or csa_tree_add_190_195_groupi_g45979(csa_tree_add_190_195_groupi_n_3191 ,csa_tree_add_190_195_groupi_n_702 ,csa_tree_add_190_195_groupi_n_2697);
  nor csa_tree_add_190_195_groupi_g45980(csa_tree_add_190_195_groupi_n_3190 ,csa_tree_add_190_195_groupi_n_770 ,csa_tree_add_190_195_groupi_n_1541);
  and csa_tree_add_190_195_groupi_g45981(csa_tree_add_190_195_groupi_n_3189 ,csa_tree_add_190_195_groupi_n_429 ,csa_tree_add_190_195_groupi_n_1870);
  nor csa_tree_add_190_195_groupi_g45982(csa_tree_add_190_195_groupi_n_3188 ,csa_tree_add_190_195_groupi_n_1517 ,csa_tree_add_190_195_groupi_n_1408);
  and csa_tree_add_190_195_groupi_g45983(csa_tree_add_190_195_groupi_n_3187 ,csa_tree_add_190_195_groupi_n_1970 ,csa_tree_add_190_195_groupi_n_1966);
  nor csa_tree_add_190_195_groupi_g45984(csa_tree_add_190_195_groupi_n_3186 ,csa_tree_add_190_195_groupi_n_1948 ,csa_tree_add_190_195_groupi_n_2042);
  nor csa_tree_add_190_195_groupi_g45985(csa_tree_add_190_195_groupi_n_3185 ,csa_tree_add_190_195_groupi_n_2641 ,csa_tree_add_190_195_groupi_n_2710);
  nor csa_tree_add_190_195_groupi_g45986(csa_tree_add_190_195_groupi_n_3184 ,csa_tree_add_190_195_groupi_n_1530 ,csa_tree_add_190_195_groupi_n_2625);
  and csa_tree_add_190_195_groupi_g45987(csa_tree_add_190_195_groupi_n_3183 ,csa_tree_add_190_195_groupi_n_606 ,csa_tree_add_190_195_groupi_n_1101);
  nor csa_tree_add_190_195_groupi_g45988(csa_tree_add_190_195_groupi_n_3182 ,in55[4] ,in59[7]);
  or csa_tree_add_190_195_groupi_g45989(csa_tree_add_190_195_groupi_n_3181 ,csa_tree_add_190_195_groupi_n_1011 ,csa_tree_add_190_195_groupi_n_1829);
  and csa_tree_add_190_195_groupi_g45990(csa_tree_add_190_195_groupi_n_3180 ,csa_tree_add_190_195_groupi_n_414 ,csa_tree_add_190_195_groupi_n_2212);
  nor csa_tree_add_190_195_groupi_g45991(csa_tree_add_190_195_groupi_n_3179 ,csa_tree_add_190_195_groupi_n_560 ,csa_tree_add_190_195_groupi_n_1968);
  and csa_tree_add_190_195_groupi_g45992(csa_tree_add_190_195_groupi_n_3178 ,csa_tree_add_190_195_groupi_n_345 ,csa_tree_add_190_195_groupi_n_1126);
  and csa_tree_add_190_195_groupi_g45993(csa_tree_add_190_195_groupi_n_3177 ,in55[4] ,in60[8]);
  and csa_tree_add_190_195_groupi_g45994(csa_tree_add_190_195_groupi_n_3176 ,csa_tree_add_190_195_groupi_n_223 ,csa_tree_add_190_195_groupi_n_1906);
  nor csa_tree_add_190_195_groupi_g45995(csa_tree_add_190_195_groupi_n_3175 ,csa_tree_add_190_195_groupi_n_465 ,csa_tree_add_190_195_groupi_n_745);
  or csa_tree_add_190_195_groupi_g45996(csa_tree_add_190_195_groupi_n_3174 ,csa_tree_add_190_195_groupi_n_2675 ,csa_tree_add_190_195_groupi_n_2382);
  nor csa_tree_add_190_195_groupi_g45997(csa_tree_add_190_195_groupi_n_3173 ,csa_tree_add_190_195_groupi_n_768 ,csa_tree_add_190_195_groupi_n_2438);
  nor csa_tree_add_190_195_groupi_g45998(csa_tree_add_190_195_groupi_n_3172 ,csa_tree_add_190_195_groupi_n_1517 ,csa_tree_add_190_195_groupi_n_2439);
  or csa_tree_add_190_195_groupi_g45999(csa_tree_add_190_195_groupi_n_3171 ,csa_tree_add_190_195_groupi_n_1230 ,csa_tree_add_190_195_groupi_n_1859);
  nor csa_tree_add_190_195_groupi_g46000(csa_tree_add_190_195_groupi_n_3170 ,csa_tree_add_190_195_groupi_n_1222 ,csa_tree_add_190_195_groupi_n_1226);
  or csa_tree_add_190_195_groupi_g46001(csa_tree_add_190_195_groupi_n_3169 ,csa_tree_add_190_195_groupi_n_1937 ,csa_tree_add_190_195_groupi_n_1992);
  nand csa_tree_add_190_195_groupi_g46002(csa_tree_add_190_195_groupi_n_3168 ,in60[13] ,in58[13]);
  or csa_tree_add_190_195_groupi_g46003(csa_tree_add_190_195_groupi_n_3167 ,csa_tree_add_190_195_groupi_n_2620 ,csa_tree_add_190_195_groupi_n_1424);
  and csa_tree_add_190_195_groupi_g46004(csa_tree_add_190_195_groupi_n_3166 ,csa_tree_add_190_195_groupi_n_1273 ,csa_tree_add_190_195_groupi_n_570);
  or csa_tree_add_190_195_groupi_g46005(csa_tree_add_190_195_groupi_n_3165 ,csa_tree_add_190_195_groupi_n_1960 ,csa_tree_add_190_195_groupi_n_1780);
  and csa_tree_add_190_195_groupi_g46006(csa_tree_add_190_195_groupi_n_3164 ,csa_tree_add_190_195_groupi_n_240 ,csa_tree_add_190_195_groupi_n_289);
  nor csa_tree_add_190_195_groupi_g46007(csa_tree_add_190_195_groupi_n_3163 ,csa_tree_add_190_195_groupi_n_434 ,csa_tree_add_190_195_groupi_n_2213);
  or csa_tree_add_190_195_groupi_g46008(csa_tree_add_190_195_groupi_n_3162 ,csa_tree_add_190_195_groupi_n_835 ,csa_tree_add_190_195_groupi_n_1829);
  or csa_tree_add_190_195_groupi_g46009(csa_tree_add_190_195_groupi_n_3161 ,csa_tree_add_190_195_groupi_n_2667 ,csa_tree_add_190_195_groupi_n_2486);
  or csa_tree_add_190_195_groupi_g46010(csa_tree_add_190_195_groupi_n_3160 ,csa_tree_add_190_195_groupi_n_771 ,csa_tree_add_190_195_groupi_n_2533);
  nor csa_tree_add_190_195_groupi_g46011(csa_tree_add_190_195_groupi_n_3159 ,csa_tree_add_190_195_groupi_n_627 ,csa_tree_add_190_195_groupi_n_2156);
  or csa_tree_add_190_195_groupi_g46012(csa_tree_add_190_195_groupi_n_3158 ,csa_tree_add_190_195_groupi_n_1687 ,csa_tree_add_190_195_groupi_n_1941);
  and csa_tree_add_190_195_groupi_g46013(csa_tree_add_190_195_groupi_n_3157 ,csa_tree_add_190_195_groupi_n_1168 ,csa_tree_add_190_195_groupi_n_1834);
  and csa_tree_add_190_195_groupi_g46014(csa_tree_add_190_195_groupi_n_3156 ,csa_tree_add_190_195_groupi_n_1063 ,csa_tree_add_190_195_groupi_n_1038);
  nor csa_tree_add_190_195_groupi_g46015(csa_tree_add_190_195_groupi_n_3155 ,csa_tree_add_190_195_groupi_n_2501 ,csa_tree_add_190_195_groupi_n_1436);
  nor csa_tree_add_190_195_groupi_g46016(csa_tree_add_190_195_groupi_n_3154 ,csa_tree_add_190_195_groupi_n_533 ,csa_tree_add_190_195_groupi_n_1844);
  nor csa_tree_add_190_195_groupi_g46017(csa_tree_add_190_195_groupi_n_3153 ,csa_tree_add_190_195_groupi_n_1411 ,csa_tree_add_190_195_groupi_n_2462);
  or csa_tree_add_190_195_groupi_g46018(csa_tree_add_190_195_groupi_n_3152 ,csa_tree_add_190_195_groupi_n_254 ,csa_tree_add_190_195_groupi_n_1032);
  and csa_tree_add_190_195_groupi_g46019(csa_tree_add_190_195_groupi_n_3151 ,csa_tree_add_190_195_groupi_n_934 ,in58[1]);
  and csa_tree_add_190_195_groupi_g46020(csa_tree_add_190_195_groupi_n_3150 ,csa_tree_add_190_195_groupi_n_2051 ,csa_tree_add_190_195_groupi_n_420);
  nor csa_tree_add_190_195_groupi_g46021(csa_tree_add_190_195_groupi_n_3149 ,csa_tree_add_190_195_groupi_n_445 ,csa_tree_add_190_195_groupi_n_1962);
  nor csa_tree_add_190_195_groupi_g46022(csa_tree_add_190_195_groupi_n_3148 ,csa_tree_add_190_195_groupi_n_1734 ,csa_tree_add_190_195_groupi_n_1607);
  and csa_tree_add_190_195_groupi_g46023(csa_tree_add_190_195_groupi_n_3147 ,csa_tree_add_190_195_groupi_n_948 ,csa_tree_add_190_195_groupi_n_323);
  nor csa_tree_add_190_195_groupi_g46024(csa_tree_add_190_195_groupi_n_3146 ,csa_tree_add_190_195_groupi_n_464 ,csa_tree_add_190_195_groupi_n_1836);
  or csa_tree_add_190_195_groupi_g46025(csa_tree_add_190_195_groupi_n_3145 ,csa_tree_add_190_195_groupi_n_1808 ,csa_tree_add_190_195_groupi_n_1199);
  nor csa_tree_add_190_195_groupi_g46026(csa_tree_add_190_195_groupi_n_3144 ,csa_tree_add_190_195_groupi_n_535 ,csa_tree_add_190_195_groupi_n_479);
  nor csa_tree_add_190_195_groupi_g46027(csa_tree_add_190_195_groupi_n_3143 ,csa_tree_add_190_195_groupi_n_579 ,csa_tree_add_190_195_groupi_n_1162);
  nor csa_tree_add_190_195_groupi_g46028(csa_tree_add_190_195_groupi_n_3142 ,csa_tree_add_190_195_groupi_n_1554 ,csa_tree_add_190_195_groupi_n_2603);
  and csa_tree_add_190_195_groupi_g46029(csa_tree_add_190_195_groupi_n_3141 ,csa_tree_add_190_195_groupi_n_1702 ,csa_tree_add_190_195_groupi_n_802);
  or csa_tree_add_190_195_groupi_g46030(csa_tree_add_190_195_groupi_n_3140 ,csa_tree_add_190_195_groupi_n_925 ,csa_tree_add_190_195_groupi_n_2055);
  or csa_tree_add_190_195_groupi_g46031(csa_tree_add_190_195_groupi_n_3139 ,csa_tree_add_190_195_groupi_n_1344 ,csa_tree_add_190_195_groupi_n_2719);
  and csa_tree_add_190_195_groupi_g46033(csa_tree_add_190_195_groupi_n_3138 ,csa_tree_add_190_195_groupi_n_990 ,csa_tree_add_190_195_groupi_n_1829);
  or csa_tree_add_190_195_groupi_g46034(csa_tree_add_190_195_groupi_n_3137 ,csa_tree_add_190_195_groupi_n_403 ,csa_tree_add_190_195_groupi_n_2119);
  nor csa_tree_add_190_195_groupi_g46035(csa_tree_add_190_195_groupi_n_3136 ,in55[14] ,in55[13]);
  nor csa_tree_add_190_195_groupi_g46036(csa_tree_add_190_195_groupi_n_3135 ,csa_tree_add_190_195_groupi_n_549 ,csa_tree_add_190_195_groupi_n_2040);
  or csa_tree_add_190_195_groupi_g46037(csa_tree_add_190_195_groupi_n_3134 ,csa_tree_add_190_195_groupi_n_440 ,csa_tree_add_190_195_groupi_n_946);
  nor csa_tree_add_190_195_groupi_g46038(csa_tree_add_190_195_groupi_n_3133 ,csa_tree_add_190_195_groupi_n_588 ,csa_tree_add_190_195_groupi_n_1249);
  and csa_tree_add_190_195_groupi_g46039(csa_tree_add_190_195_groupi_n_3132 ,csa_tree_add_190_195_groupi_n_1014 ,csa_tree_add_190_195_groupi_n_1951);
  or csa_tree_add_190_195_groupi_g46040(csa_tree_add_190_195_groupi_n_3131 ,csa_tree_add_190_195_groupi_n_2049 ,csa_tree_add_190_195_groupi_n_1763);
  or csa_tree_add_190_195_groupi_g46041(csa_tree_add_190_195_groupi_n_3130 ,csa_tree_add_190_195_groupi_n_2057 ,csa_tree_add_190_195_groupi_n_1965);
  nor csa_tree_add_190_195_groupi_g46042(csa_tree_add_190_195_groupi_n_3129 ,csa_tree_add_190_195_groupi_n_1845 ,csa_tree_add_190_195_groupi_n_1096);
  nor csa_tree_add_190_195_groupi_g46043(csa_tree_add_190_195_groupi_n_3128 ,csa_tree_add_190_195_groupi_n_727 ,csa_tree_add_190_195_groupi_n_1539);
  or csa_tree_add_190_195_groupi_g46044(csa_tree_add_190_195_groupi_n_3127 ,csa_tree_add_190_195_groupi_n_736 ,csa_tree_add_190_195_groupi_n_2439);
  and csa_tree_add_190_195_groupi_g46045(csa_tree_add_190_195_groupi_n_3126 ,csa_tree_add_190_195_groupi_n_307 ,csa_tree_add_190_195_groupi_n_1915);
  or csa_tree_add_190_195_groupi_g46046(csa_tree_add_190_195_groupi_n_3125 ,csa_tree_add_190_195_groupi_n_1449 ,csa_tree_add_190_195_groupi_n_2342);
  or csa_tree_add_190_195_groupi_g46047(csa_tree_add_190_195_groupi_n_3124 ,csa_tree_add_190_195_groupi_n_1224 ,csa_tree_add_190_195_groupi_n_756);
  nor csa_tree_add_190_195_groupi_g46048(csa_tree_add_190_195_groupi_n_3123 ,in55[6] ,in60[10]);
  and csa_tree_add_190_195_groupi_g46049(csa_tree_add_190_195_groupi_n_3122 ,csa_tree_add_190_195_groupi_n_206 ,csa_tree_add_190_195_groupi_n_898);
  nor csa_tree_add_190_195_groupi_g46050(csa_tree_add_190_195_groupi_n_3121 ,csa_tree_add_190_195_groupi_n_543 ,csa_tree_add_190_195_groupi_n_1279);
  nor csa_tree_add_190_195_groupi_g46051(csa_tree_add_190_195_groupi_n_3120 ,csa_tree_add_190_195_groupi_n_1848 ,csa_tree_add_190_195_groupi_n_1847);
  nor csa_tree_add_190_195_groupi_g46052(csa_tree_add_190_195_groupi_n_3119 ,csa_tree_add_190_195_groupi_n_1552 ,csa_tree_add_190_195_groupi_n_2420);
  and csa_tree_add_190_195_groupi_g46053(csa_tree_add_190_195_groupi_n_3118 ,csa_tree_add_190_195_groupi_n_190 ,csa_tree_add_190_195_groupi_n_963);
  and csa_tree_add_190_195_groupi_g46054(csa_tree_add_190_195_groupi_n_3117 ,csa_tree_add_190_195_groupi_n_541 ,csa_tree_add_190_195_groupi_n_1218);
  nor csa_tree_add_190_195_groupi_g46055(csa_tree_add_190_195_groupi_n_3116 ,csa_tree_add_190_195_groupi_n_1516 ,csa_tree_add_190_195_groupi_n_686);
  nor csa_tree_add_190_195_groupi_g46056(csa_tree_add_190_195_groupi_n_3115 ,csa_tree_add_190_195_groupi_n_1368 ,csa_tree_add_190_195_groupi_n_1360);
  or csa_tree_add_190_195_groupi_g46057(csa_tree_add_190_195_groupi_n_3114 ,csa_tree_add_190_195_groupi_n_522 ,csa_tree_add_190_195_groupi_n_2155);
  or csa_tree_add_190_195_groupi_g46058(csa_tree_add_190_195_groupi_n_3113 ,csa_tree_add_190_195_groupi_n_1336 ,csa_tree_add_190_195_groupi_n_2553);
  nor csa_tree_add_190_195_groupi_g46059(csa_tree_add_190_195_groupi_n_3112 ,csa_tree_add_190_195_groupi_n_1236 ,csa_tree_add_190_195_groupi_n_1906);
  nor csa_tree_add_190_195_groupi_g46060(csa_tree_add_190_195_groupi_n_3111 ,csa_tree_add_190_195_groupi_n_2062 ,csa_tree_add_190_195_groupi_n_2060);
  nor csa_tree_add_190_195_groupi_g46061(csa_tree_add_190_195_groupi_n_3110 ,csa_tree_add_190_195_groupi_n_1514 ,csa_tree_add_190_195_groupi_n_1478);
  nor csa_tree_add_190_195_groupi_g46062(csa_tree_add_190_195_groupi_n_3109 ,csa_tree_add_190_195_groupi_n_1413 ,csa_tree_add_190_195_groupi_n_2497);
  nor csa_tree_add_190_195_groupi_g46063(csa_tree_add_190_195_groupi_n_3108 ,csa_tree_add_190_195_groupi_n_540 ,csa_tree_add_190_195_groupi_n_1748);
  nor csa_tree_add_190_195_groupi_g46064(csa_tree_add_190_195_groupi_n_3107 ,csa_tree_add_190_195_groupi_n_371 ,csa_tree_add_190_195_groupi_n_1974);
  nor csa_tree_add_190_195_groupi_g46065(csa_tree_add_190_195_groupi_n_3106 ,csa_tree_add_190_195_groupi_n_518 ,csa_tree_add_190_195_groupi_n_786);
  nor csa_tree_add_190_195_groupi_g46066(csa_tree_add_190_195_groupi_n_3105 ,csa_tree_add_190_195_groupi_n_2447 ,csa_tree_add_190_195_groupi_n_2471);
  nor csa_tree_add_190_195_groupi_g46067(csa_tree_add_190_195_groupi_n_3104 ,in58[12] ,in59[12]);
  nor csa_tree_add_190_195_groupi_g46068(csa_tree_add_190_195_groupi_n_3103 ,csa_tree_add_190_195_groupi_n_2440 ,csa_tree_add_190_195_groupi_n_2626);
  or csa_tree_add_190_195_groupi_g46069(csa_tree_add_190_195_groupi_n_3102 ,in55[5] ,in58[8]);
  or csa_tree_add_190_195_groupi_g46070(csa_tree_add_190_195_groupi_n_3101 ,csa_tree_add_190_195_groupi_n_426 ,csa_tree_add_190_195_groupi_n_2001);
  and csa_tree_add_190_195_groupi_g46071(csa_tree_add_190_195_groupi_n_3100 ,csa_tree_add_190_195_groupi_n_1078 ,csa_tree_add_190_195_groupi_n_1968);
  nor csa_tree_add_190_195_groupi_g46072(csa_tree_add_190_195_groupi_n_3099 ,csa_tree_add_190_195_groupi_n_2638 ,csa_tree_add_190_195_groupi_n_2489);
  nor csa_tree_add_190_195_groupi_g46073(csa_tree_add_190_195_groupi_n_3098 ,csa_tree_add_190_195_groupi_n_468 ,csa_tree_add_190_195_groupi_n_1186);
  or csa_tree_add_190_195_groupi_g46074(csa_tree_add_190_195_groupi_n_3097 ,csa_tree_add_190_195_groupi_n_948 ,csa_tree_add_190_195_groupi_n_886);
  and csa_tree_add_190_195_groupi_g46075(csa_tree_add_190_195_groupi_n_3096 ,csa_tree_add_190_195_groupi_n_286 ,csa_tree_add_190_195_groupi_n_2212);
  nor csa_tree_add_190_195_groupi_g46076(csa_tree_add_190_195_groupi_n_3095 ,csa_tree_add_190_195_groupi_n_1422 ,csa_tree_add_190_195_groupi_n_1495);
  nor csa_tree_add_190_195_groupi_g46077(csa_tree_add_190_195_groupi_n_3094 ,csa_tree_add_190_195_groupi_n_814 ,csa_tree_add_190_195_groupi_n_873);
  or csa_tree_add_190_195_groupi_g46078(csa_tree_add_190_195_groupi_n_3093 ,csa_tree_add_190_195_groupi_n_1426 ,csa_tree_add_190_195_groupi_n_2481);
  and csa_tree_add_190_195_groupi_g46079(csa_tree_add_190_195_groupi_n_3092 ,csa_tree_add_190_195_groupi_n_279 ,csa_tree_add_190_195_groupi_n_1889);
  and csa_tree_add_190_195_groupi_g46080(csa_tree_add_190_195_groupi_n_3091 ,csa_tree_add_190_195_groupi_n_213 ,csa_tree_add_190_195_groupi_n_2015);
  nor csa_tree_add_190_195_groupi_g46081(csa_tree_add_190_195_groupi_n_3090 ,csa_tree_add_190_195_groupi_n_2462 ,csa_tree_add_190_195_groupi_n_2532);
  nor csa_tree_add_190_195_groupi_g46082(csa_tree_add_190_195_groupi_n_3089 ,csa_tree_add_190_195_groupi_n_277 ,csa_tree_add_190_195_groupi_n_1707);
  and csa_tree_add_190_195_groupi_g46083(csa_tree_add_190_195_groupi_n_3088 ,csa_tree_add_190_195_groupi_n_375 ,csa_tree_add_190_195_groupi_n_252);
  or csa_tree_add_190_195_groupi_g46084(csa_tree_add_190_195_groupi_n_3087 ,csa_tree_add_190_195_groupi_n_281 ,csa_tree_add_190_195_groupi_n_1843);
  nor csa_tree_add_190_195_groupi_g46085(csa_tree_add_190_195_groupi_n_3086 ,csa_tree_add_190_195_groupi_n_1978 ,in58[5]);
  or csa_tree_add_190_195_groupi_g46086(csa_tree_add_190_195_groupi_n_3085 ,csa_tree_add_190_195_groupi_n_1350 ,csa_tree_add_190_195_groupi_n_2536);
  or csa_tree_add_190_195_groupi_g46087(csa_tree_add_190_195_groupi_n_3084 ,csa_tree_add_190_195_groupi_n_816 ,csa_tree_add_190_195_groupi_n_1703);
  nor csa_tree_add_190_195_groupi_g46088(csa_tree_add_190_195_groupi_n_3083 ,csa_tree_add_190_195_groupi_n_1508 ,csa_tree_add_190_195_groupi_n_2687);
  or csa_tree_add_190_195_groupi_g46089(csa_tree_add_190_195_groupi_n_3082 ,csa_tree_add_190_195_groupi_n_1840 ,csa_tree_add_190_195_groupi_n_1916);
  or csa_tree_add_190_195_groupi_g46090(csa_tree_add_190_195_groupi_n_3081 ,csa_tree_add_190_195_groupi_n_1257 ,csa_tree_add_190_195_groupi_n_1968);
  nor csa_tree_add_190_195_groupi_g46091(csa_tree_add_190_195_groupi_n_3080 ,csa_tree_add_190_195_groupi_n_1499 ,csa_tree_add_190_195_groupi_n_2660);
  or csa_tree_add_190_195_groupi_g46092(csa_tree_add_190_195_groupi_n_3079 ,csa_tree_add_190_195_groupi_n_952 ,csa_tree_add_190_195_groupi_n_1125);
  nor csa_tree_add_190_195_groupi_g46093(csa_tree_add_190_195_groupi_n_3078 ,csa_tree_add_190_195_groupi_n_814 ,csa_tree_add_190_195_groupi_n_1921);
  nor csa_tree_add_190_195_groupi_g46094(csa_tree_add_190_195_groupi_n_3077 ,csa_tree_add_190_195_groupi_n_1549 ,csa_tree_add_190_195_groupi_n_2573);
  nor csa_tree_add_190_195_groupi_g46095(csa_tree_add_190_195_groupi_n_3076 ,csa_tree_add_190_195_groupi_n_1238 ,csa_tree_add_190_195_groupi_n_2051);
  nor csa_tree_add_190_195_groupi_g46096(csa_tree_add_190_195_groupi_n_3075 ,csa_tree_add_190_195_groupi_n_2091 ,csa_tree_add_190_195_groupi_n_2154);
  or csa_tree_add_190_195_groupi_g46097(csa_tree_add_190_195_groupi_n_3074 ,csa_tree_add_190_195_groupi_n_1863 ,csa_tree_add_190_195_groupi_n_915);
  nor csa_tree_add_190_195_groupi_g46098(csa_tree_add_190_195_groupi_n_3073 ,csa_tree_add_190_195_groupi_n_616 ,csa_tree_add_190_195_groupi_n_2118);
  nor csa_tree_add_190_195_groupi_g46099(csa_tree_add_190_195_groupi_n_3072 ,csa_tree_add_190_195_groupi_n_1301 ,csa_tree_add_190_195_groupi_n_1749);
  and csa_tree_add_190_195_groupi_g46100(csa_tree_add_190_195_groupi_n_3071 ,in55[6] ,in60[10]);
  or csa_tree_add_190_195_groupi_g46101(csa_tree_add_190_195_groupi_n_3070 ,csa_tree_add_190_195_groupi_n_370 ,csa_tree_add_190_195_groupi_n_1170);
  or csa_tree_add_190_195_groupi_g46102(csa_tree_add_190_195_groupi_n_3069 ,in55[8] ,in60[12]);
  nor csa_tree_add_190_195_groupi_g46103(csa_tree_add_190_195_groupi_n_3068 ,csa_tree_add_190_195_groupi_n_432 ,csa_tree_add_190_195_groupi_n_453);
  and csa_tree_add_190_195_groupi_g46104(csa_tree_add_190_195_groupi_n_3067 ,csa_tree_add_190_195_groupi_n_825 ,csa_tree_add_190_195_groupi_n_459);
  or csa_tree_add_190_195_groupi_g46105(csa_tree_add_190_195_groupi_n_3066 ,csa_tree_add_190_195_groupi_n_1850 ,csa_tree_add_190_195_groupi_n_1847);
  nor csa_tree_add_190_195_groupi_g46106(csa_tree_add_190_195_groupi_n_3065 ,csa_tree_add_190_195_groupi_n_2461 ,csa_tree_add_190_195_groupi_n_1364);
  nor csa_tree_add_190_195_groupi_g46107(csa_tree_add_190_195_groupi_n_3064 ,csa_tree_add_190_195_groupi_n_734 ,csa_tree_add_190_195_groupi_n_1388);
  nor csa_tree_add_190_195_groupi_g46108(csa_tree_add_190_195_groupi_n_3063 ,csa_tree_add_190_195_groupi_n_613 ,csa_tree_add_190_195_groupi_n_2088);
  nor csa_tree_add_190_195_groupi_g46109(csa_tree_add_190_195_groupi_n_3062 ,csa_tree_add_190_195_groupi_n_554 ,csa_tree_add_190_195_groupi_n_472);
  and csa_tree_add_190_195_groupi_g46110(csa_tree_add_190_195_groupi_n_3061 ,csa_tree_add_190_195_groupi_n_1143 ,csa_tree_add_190_195_groupi_n_1032);
  nor csa_tree_add_190_195_groupi_g46111(csa_tree_add_190_195_groupi_n_3060 ,csa_tree_add_190_195_groupi_n_436 ,csa_tree_add_190_195_groupi_n_241);
  or csa_tree_add_190_195_groupi_g46112(csa_tree_add_190_195_groupi_n_3059 ,csa_tree_add_190_195_groupi_n_1484 ,csa_tree_add_190_195_groupi_n_2631);
  nor csa_tree_add_190_195_groupi_g46113(csa_tree_add_190_195_groupi_n_3058 ,csa_tree_add_190_195_groupi_n_2578 ,csa_tree_add_190_195_groupi_n_1485);
  nor csa_tree_add_190_195_groupi_g46114(csa_tree_add_190_195_groupi_n_3057 ,csa_tree_add_190_195_groupi_n_1281 ,csa_tree_add_190_195_groupi_n_1934);
  or csa_tree_add_190_195_groupi_g46115(csa_tree_add_190_195_groupi_n_3056 ,csa_tree_add_190_195_groupi_n_2424 ,csa_tree_add_190_195_groupi_n_2418);
  or csa_tree_add_190_195_groupi_g46116(csa_tree_add_190_195_groupi_n_3055 ,csa_tree_add_190_195_groupi_n_368 ,csa_tree_add_190_195_groupi_n_1961);
  nor csa_tree_add_190_195_groupi_g46117(csa_tree_add_190_195_groupi_n_3054 ,csa_tree_add_190_195_groupi_n_1809 ,csa_tree_add_190_195_groupi_n_1705);
  nor csa_tree_add_190_195_groupi_g46118(csa_tree_add_190_195_groupi_n_3053 ,csa_tree_add_190_195_groupi_n_313 ,csa_tree_add_190_195_groupi_n_1257);
  nor csa_tree_add_190_195_groupi_g46119(csa_tree_add_190_195_groupi_n_3052 ,csa_tree_add_190_195_groupi_n_1482 ,csa_tree_add_190_195_groupi_n_1557);
  and csa_tree_add_190_195_groupi_g46120(csa_tree_add_190_195_groupi_n_3051 ,in55[0] ,in61[4]);
  nor csa_tree_add_190_195_groupi_g46121(csa_tree_add_190_195_groupi_n_3050 ,csa_tree_add_190_195_groupi_n_2630 ,csa_tree_add_190_195_groupi_n_2663);
  nor csa_tree_add_190_195_groupi_g46122(csa_tree_add_190_195_groupi_n_3049 ,csa_tree_add_190_195_groupi_n_2214 ,csa_tree_add_190_195_groupi_n_1744);
  and csa_tree_add_190_195_groupi_g46123(csa_tree_add_190_195_groupi_n_3048 ,csa_tree_add_190_195_groupi_n_1891 ,csa_tree_add_190_195_groupi_n_1887);
  or csa_tree_add_190_195_groupi_g46124(csa_tree_add_190_195_groupi_n_3047 ,csa_tree_add_190_195_groupi_n_694 ,csa_tree_add_190_195_groupi_n_2642);
  nor csa_tree_add_190_195_groupi_g46125(csa_tree_add_190_195_groupi_n_3046 ,csa_tree_add_190_195_groupi_n_442 ,csa_tree_add_190_195_groupi_n_1839);
  nor csa_tree_add_190_195_groupi_g46126(csa_tree_add_190_195_groupi_n_3045 ,csa_tree_add_190_195_groupi_n_558 ,csa_tree_add_190_195_groupi_n_1761);
  nor csa_tree_add_190_195_groupi_g46127(csa_tree_add_190_195_groupi_n_3044 ,csa_tree_add_190_195_groupi_n_1471 ,csa_tree_add_190_195_groupi_n_2605);
  or csa_tree_add_190_195_groupi_g46128(csa_tree_add_190_195_groupi_n_3043 ,csa_tree_add_190_195_groupi_n_2086 ,csa_tree_add_190_195_groupi_n_849);
  or csa_tree_add_190_195_groupi_g46129(csa_tree_add_190_195_groupi_n_3042 ,csa_tree_add_190_195_groupi_n_729 ,csa_tree_add_190_195_groupi_n_1376);
  nor csa_tree_add_190_195_groupi_g46130(csa_tree_add_190_195_groupi_n_3041 ,csa_tree_add_190_195_groupi_n_1253 ,csa_tree_add_190_195_groupi_n_1935);
  nor csa_tree_add_190_195_groupi_g46131(csa_tree_add_190_195_groupi_n_3040 ,csa_tree_add_190_195_groupi_n_495 ,csa_tree_add_190_195_groupi_n_1210);
  or csa_tree_add_190_195_groupi_g46132(csa_tree_add_190_195_groupi_n_3039 ,csa_tree_add_190_195_groupi_n_1750 ,csa_tree_add_190_195_groupi_n_1929);
  and csa_tree_add_190_195_groupi_g46133(csa_tree_add_190_195_groupi_n_3038 ,csa_tree_add_190_195_groupi_n_988 ,csa_tree_add_190_195_groupi_n_840);
  nor csa_tree_add_190_195_groupi_g46134(csa_tree_add_190_195_groupi_n_3037 ,csa_tree_add_190_195_groupi_n_2537 ,csa_tree_add_190_195_groupi_n_2464);
  nor csa_tree_add_190_195_groupi_g46135(csa_tree_add_190_195_groupi_n_3036 ,csa_tree_add_190_195_groupi_n_1520 ,csa_tree_add_190_195_groupi_n_2528);
  or csa_tree_add_190_195_groupi_g46136(csa_tree_add_190_195_groupi_n_3035 ,csa_tree_add_190_195_groupi_n_2442 ,csa_tree_add_190_195_groupi_n_2463);
  nor csa_tree_add_190_195_groupi_g46137(csa_tree_add_190_195_groupi_n_3034 ,csa_tree_add_190_195_groupi_n_1568 ,csa_tree_add_190_195_groupi_n_1556);
  or csa_tree_add_190_195_groupi_g46138(csa_tree_add_190_195_groupi_n_3033 ,csa_tree_add_190_195_groupi_n_628 ,csa_tree_add_190_195_groupi_n_1903);
  nor csa_tree_add_190_195_groupi_g46139(csa_tree_add_190_195_groupi_n_3032 ,csa_tree_add_190_195_groupi_n_1167 ,csa_tree_add_190_195_groupi_n_2153);
  and csa_tree_add_190_195_groupi_g46140(csa_tree_add_190_195_groupi_n_3031 ,csa_tree_add_190_195_groupi_n_556 ,csa_tree_add_190_195_groupi_n_2001);
  nor csa_tree_add_190_195_groupi_g46141(csa_tree_add_190_195_groupi_n_3030 ,csa_tree_add_190_195_groupi_n_2615 ,csa_tree_add_190_195_groupi_n_2436);
  nor csa_tree_add_190_195_groupi_g46142(csa_tree_add_190_195_groupi_n_3029 ,csa_tree_add_190_195_groupi_n_576 ,csa_tree_add_190_195_groupi_n_988);
  nor csa_tree_add_190_195_groupi_g46143(csa_tree_add_190_195_groupi_n_3028 ,csa_tree_add_190_195_groupi_n_563 ,csa_tree_add_190_195_groupi_n_1144);
  or csa_tree_add_190_195_groupi_g46144(csa_tree_add_190_195_groupi_n_3027 ,csa_tree_add_190_195_groupi_n_2521 ,csa_tree_add_190_195_groupi_n_1420);
  nor csa_tree_add_190_195_groupi_g46145(csa_tree_add_190_195_groupi_n_3026 ,csa_tree_add_190_195_groupi_n_829 ,csa_tree_add_190_195_groupi_n_705);
  or csa_tree_add_190_195_groupi_g46146(csa_tree_add_190_195_groupi_n_3025 ,csa_tree_add_190_195_groupi_n_353 ,csa_tree_add_190_195_groupi_n_1750);
  nor csa_tree_add_190_195_groupi_g46147(csa_tree_add_190_195_groupi_n_3024 ,csa_tree_add_190_195_groupi_n_2040 ,csa_tree_add_190_195_groupi_n_2158);
  or csa_tree_add_190_195_groupi_g46148(csa_tree_add_190_195_groupi_n_3023 ,csa_tree_add_190_195_groupi_n_2116 ,csa_tree_add_190_195_groupi_n_1141);
  or csa_tree_add_190_195_groupi_g46149(csa_tree_add_190_195_groupi_n_3022 ,csa_tree_add_190_195_groupi_n_1888 ,csa_tree_add_190_195_groupi_n_1833);
  and csa_tree_add_190_195_groupi_g46150(csa_tree_add_190_195_groupi_n_3021 ,csa_tree_add_190_195_groupi_n_458 ,csa_tree_add_190_195_groupi_n_1287);
  and csa_tree_add_190_195_groupi_g46151(csa_tree_add_190_195_groupi_n_3020 ,csa_tree_add_190_195_groupi_n_1155 ,csa_tree_add_190_195_groupi_n_1814);
  or csa_tree_add_190_195_groupi_g46152(csa_tree_add_190_195_groupi_n_3019 ,csa_tree_add_190_195_groupi_n_1446 ,csa_tree_add_190_195_groupi_n_1370);
  nor csa_tree_add_190_195_groupi_g46153(csa_tree_add_190_195_groupi_n_3018 ,csa_tree_add_190_195_groupi_n_287 ,csa_tree_add_190_195_groupi_n_2212);
  or csa_tree_add_190_195_groupi_g46154(csa_tree_add_190_195_groupi_n_3017 ,csa_tree_add_190_195_groupi_n_843 ,csa_tree_add_190_195_groupi_n_193);
  and csa_tree_add_190_195_groupi_g46155(csa_tree_add_190_195_groupi_n_3016 ,csa_tree_add_190_195_groupi_n_396 ,csa_tree_add_190_195_groupi_n_1135);
  nor csa_tree_add_190_195_groupi_g46156(csa_tree_add_190_195_groupi_n_3015 ,csa_tree_add_190_195_groupi_n_1299 ,csa_tree_add_190_195_groupi_n_1832);
  nor csa_tree_add_190_195_groupi_g46157(csa_tree_add_190_195_groupi_n_3014 ,csa_tree_add_190_195_groupi_n_2525 ,csa_tree_add_190_195_groupi_n_2450);
  and csa_tree_add_190_195_groupi_g46158(csa_tree_add_190_195_groupi_n_3013 ,csa_tree_add_190_195_groupi_n_443 ,csa_tree_add_190_195_groupi_n_1839);
  or csa_tree_add_190_195_groupi_g46159(csa_tree_add_190_195_groupi_n_3012 ,csa_tree_add_190_195_groupi_n_1403 ,csa_tree_add_190_195_groupi_n_1370);
  nor csa_tree_add_190_195_groupi_g46160(csa_tree_add_190_195_groupi_n_3011 ,csa_tree_add_190_195_groupi_n_2715 ,csa_tree_add_190_195_groupi_n_2508);
  and csa_tree_add_190_195_groupi_g46161(csa_tree_add_190_195_groupi_n_3010 ,csa_tree_add_190_195_groupi_n_338 ,csa_tree_add_190_195_groupi_n_1971);
  or csa_tree_add_190_195_groupi_g46162(csa_tree_add_190_195_groupi_n_3009 ,csa_tree_add_190_195_groupi_n_364 ,csa_tree_add_190_195_groupi_n_1674);
  nor csa_tree_add_190_195_groupi_g46163(csa_tree_add_190_195_groupi_n_3008 ,csa_tree_add_190_195_groupi_n_1430 ,csa_tree_add_190_195_groupi_n_2526);
  and csa_tree_add_190_195_groupi_g46164(csa_tree_add_190_195_groupi_n_3007 ,csa_tree_add_190_195_groupi_n_488 ,csa_tree_add_190_195_groupi_n_1749);
  and csa_tree_add_190_195_groupi_g46165(csa_tree_add_190_195_groupi_n_3006 ,csa_tree_add_190_195_groupi_n_373 ,csa_tree_add_190_195_groupi_n_297);
  nor csa_tree_add_190_195_groupi_g46166(csa_tree_add_190_195_groupi_n_3005 ,csa_tree_add_190_195_groupi_n_2637 ,csa_tree_add_190_195_groupi_n_2435);
  or csa_tree_add_190_195_groupi_g46167(csa_tree_add_190_195_groupi_n_3004 ,csa_tree_add_190_195_groupi_n_1510 ,csa_tree_add_190_195_groupi_n_2457);
  nor csa_tree_add_190_195_groupi_g46168(csa_tree_add_190_195_groupi_n_3003 ,csa_tree_add_190_195_groupi_n_1159 ,csa_tree_add_190_195_groupi_n_808);
  and csa_tree_add_190_195_groupi_g46169(csa_tree_add_190_195_groupi_n_3002 ,csa_tree_add_190_195_groupi_n_401 ,csa_tree_add_190_195_groupi_n_1275);
  or csa_tree_add_190_195_groupi_g46171(csa_tree_add_190_195_groupi_n_3001 ,csa_tree_add_190_195_groupi_n_2466 ,csa_tree_add_190_195_groupi_n_2339);
  and csa_tree_add_190_195_groupi_g46172(csa_tree_add_190_195_groupi_n_3000 ,csa_tree_add_190_195_groupi_n_345 ,csa_tree_add_190_195_groupi_n_1821);
  or csa_tree_add_190_195_groupi_g46173(csa_tree_add_190_195_groupi_n_2999 ,csa_tree_add_190_195_groupi_n_673 ,csa_tree_add_190_195_groupi_n_2539);
  nor csa_tree_add_190_195_groupi_g46174(csa_tree_add_190_195_groupi_n_2998 ,csa_tree_add_190_195_groupi_n_2550 ,csa_tree_add_190_195_groupi_n_2703);
  and csa_tree_add_190_195_groupi_g46175(csa_tree_add_190_195_groupi_n_2997 ,csa_tree_add_190_195_groupi_n_364 ,csa_tree_add_190_195_groupi_n_1081);
  or csa_tree_add_190_195_groupi_g46176(csa_tree_add_190_195_groupi_n_2996 ,csa_tree_add_190_195_groupi_n_389 ,csa_tree_add_190_195_groupi_n_1867);
  nor csa_tree_add_190_195_groupi_g46177(csa_tree_add_190_195_groupi_n_2995 ,csa_tree_add_190_195_groupi_n_521 ,csa_tree_add_190_195_groupi_n_901);
  or csa_tree_add_190_195_groupi_g46178(csa_tree_add_190_195_groupi_n_2994 ,csa_tree_add_190_195_groupi_n_1456 ,csa_tree_add_190_195_groupi_n_1428);
  or csa_tree_add_190_195_groupi_g46179(csa_tree_add_190_195_groupi_n_2993 ,csa_tree_add_190_195_groupi_n_2016 ,csa_tree_add_190_195_groupi_n_1965);
  nor csa_tree_add_190_195_groupi_g46180(csa_tree_add_190_195_groupi_n_2992 ,csa_tree_add_190_195_groupi_n_1240 ,csa_tree_add_190_195_groupi_n_439);
  or csa_tree_add_190_195_groupi_g46181(csa_tree_add_190_195_groupi_n_2991 ,csa_tree_add_190_195_groupi_n_2209 ,csa_tree_add_190_195_groupi_n_2215);
  nor csa_tree_add_190_195_groupi_g46182(csa_tree_add_190_195_groupi_n_2990 ,csa_tree_add_190_195_groupi_n_448 ,csa_tree_add_190_195_groupi_n_475);
  or csa_tree_add_190_195_groupi_g46183(csa_tree_add_190_195_groupi_n_2989 ,csa_tree_add_190_195_groupi_n_1516 ,csa_tree_add_190_195_groupi_n_1495);
  nor csa_tree_add_190_195_groupi_g46184(csa_tree_add_190_195_groupi_n_2988 ,csa_tree_add_190_195_groupi_n_751 ,csa_tree_add_190_195_groupi_n_1604);
  nor csa_tree_add_190_195_groupi_g46185(csa_tree_add_190_195_groupi_n_2987 ,csa_tree_add_190_195_groupi_n_2506 ,csa_tree_add_190_195_groupi_n_2471);
  nor csa_tree_add_190_195_groupi_g46186(csa_tree_add_190_195_groupi_n_2986 ,csa_tree_add_190_195_groupi_n_782 ,csa_tree_add_190_195_groupi_n_1444);
  and csa_tree_add_190_195_groupi_g46187(csa_tree_add_190_195_groupi_n_2985 ,csa_tree_add_190_195_groupi_n_1840 ,csa_tree_add_190_195_groupi_n_1916);
  nor csa_tree_add_190_195_groupi_g46188(csa_tree_add_190_195_groupi_n_2984 ,csa_tree_add_190_195_groupi_n_601 ,csa_tree_add_190_195_groupi_n_257);
  or csa_tree_add_190_195_groupi_g46189(csa_tree_add_190_195_groupi_n_2983 ,csa_tree_add_190_195_groupi_n_600 ,csa_tree_add_190_195_groupi_n_1942);
  or csa_tree_add_190_195_groupi_g46190(csa_tree_add_190_195_groupi_n_2982 ,csa_tree_add_190_195_groupi_n_1474 ,csa_tree_add_190_195_groupi_n_704);
  or csa_tree_add_190_195_groupi_g46191(csa_tree_add_190_195_groupi_n_2981 ,csa_tree_add_190_195_groupi_n_2589 ,csa_tree_add_190_195_groupi_n_1404);
  nor csa_tree_add_190_195_groupi_g46192(csa_tree_add_190_195_groupi_n_2980 ,csa_tree_add_190_195_groupi_n_1904 ,csa_tree_add_190_195_groupi_n_1906);
  nor csa_tree_add_190_195_groupi_g46193(csa_tree_add_190_195_groupi_n_2979 ,csa_tree_add_190_195_groupi_n_1526 ,csa_tree_add_190_195_groupi_n_2655);
  and csa_tree_add_190_195_groupi_g46194(csa_tree_add_190_195_groupi_n_2978 ,csa_tree_add_190_195_groupi_n_299 ,in60[2]);
  or csa_tree_add_190_195_groupi_g46195(csa_tree_add_190_195_groupi_n_2977 ,csa_tree_add_190_195_groupi_n_1212 ,csa_tree_add_190_195_groupi_n_2015);
  and csa_tree_add_190_195_groupi_g46196(csa_tree_add_190_195_groupi_n_2976 ,csa_tree_add_190_195_groupi_n_2116 ,csa_tree_add_190_195_groupi_n_1140);
  nor csa_tree_add_190_195_groupi_g46197(csa_tree_add_190_195_groupi_n_2975 ,csa_tree_add_190_195_groupi_n_501 ,csa_tree_add_190_195_groupi_n_1996);
  or csa_tree_add_190_195_groupi_g46199(csa_tree_add_190_195_groupi_n_2973 ,csa_tree_add_190_195_groupi_n_1455 ,csa_tree_add_190_195_groupi_n_2679);
  and csa_tree_add_190_195_groupi_g46200(csa_tree_add_190_195_groupi_n_2972 ,csa_tree_add_190_195_groupi_n_624 ,csa_tree_add_190_195_groupi_n_2088);
  nor csa_tree_add_190_195_groupi_g46201(csa_tree_add_190_195_groupi_n_2971 ,in55[2] ,in59[5]);
  nor csa_tree_add_190_195_groupi_g46202(csa_tree_add_190_195_groupi_n_2970 ,csa_tree_add_190_195_groupi_n_1845 ,csa_tree_add_190_195_groupi_n_1931);
  or csa_tree_add_190_195_groupi_g46203(csa_tree_add_190_195_groupi_n_2969 ,csa_tree_add_190_195_groupi_n_2061 ,csa_tree_add_190_195_groupi_n_976);
  nor csa_tree_add_190_195_groupi_g46204(csa_tree_add_190_195_groupi_n_2968 ,csa_tree_add_190_195_groupi_n_1432 ,csa_tree_add_190_195_groupi_n_2605);
  nor csa_tree_add_190_195_groupi_g46205(csa_tree_add_190_195_groupi_n_2967 ,csa_tree_add_190_195_groupi_n_498 ,csa_tree_add_190_195_groupi_n_2054);
  or csa_tree_add_190_195_groupi_g46206(csa_tree_add_190_195_groupi_n_2966 ,csa_tree_add_190_195_groupi_n_1976 ,csa_tree_add_190_195_groupi_n_1758);
  nor csa_tree_add_190_195_groupi_g46207(csa_tree_add_190_195_groupi_n_2965 ,csa_tree_add_190_195_groupi_n_610 ,csa_tree_add_190_195_groupi_n_1087);
  nor csa_tree_add_190_195_groupi_g46208(csa_tree_add_190_195_groupi_n_2964 ,csa_tree_add_190_195_groupi_n_2474 ,csa_tree_add_190_195_groupi_n_2507);
  or csa_tree_add_190_195_groupi_g46209(csa_tree_add_190_195_groupi_n_2963 ,csa_tree_add_190_195_groupi_n_1530 ,csa_tree_add_190_195_groupi_n_2529);
  nor csa_tree_add_190_195_groupi_g46210(csa_tree_add_190_195_groupi_n_2962 ,csa_tree_add_190_195_groupi_n_2476 ,csa_tree_add_190_195_groupi_n_2524);
  or csa_tree_add_190_195_groupi_g46211(csa_tree_add_190_195_groupi_n_2961 ,csa_tree_add_190_195_groupi_n_619 ,csa_tree_add_190_195_groupi_n_2090);
  nor csa_tree_add_190_195_groupi_g46212(csa_tree_add_190_195_groupi_n_2960 ,csa_tree_add_190_195_groupi_n_823 ,csa_tree_add_190_195_groupi_n_2478);
  nor csa_tree_add_190_195_groupi_g46213(csa_tree_add_190_195_groupi_n_2959 ,csa_tree_add_190_195_groupi_n_949 ,csa_tree_add_190_195_groupi_n_897);
  nor csa_tree_add_190_195_groupi_g46214(csa_tree_add_190_195_groupi_n_2958 ,csa_tree_add_190_195_groupi_n_592 ,csa_tree_add_190_195_groupi_n_2063);
  and csa_tree_add_190_195_groupi_g46215(csa_tree_add_190_195_groupi_n_2957 ,csa_tree_add_190_195_groupi_n_1191 ,csa_tree_add_190_195_groupi_n_800);
  or csa_tree_add_190_195_groupi_g46216(csa_tree_add_190_195_groupi_n_2956 ,csa_tree_add_190_195_groupi_n_1167 ,csa_tree_add_190_195_groupi_n_1834);
  or csa_tree_add_190_195_groupi_g46217(csa_tree_add_190_195_groupi_n_2955 ,csa_tree_add_190_195_groupi_n_1934 ,csa_tree_add_190_195_groupi_n_1994);
  nor csa_tree_add_190_195_groupi_g46218(csa_tree_add_190_195_groupi_n_2954 ,in55[1] ,csa_tree_add_190_195_groupi_n_1193);
  nor csa_tree_add_190_195_groupi_g46219(csa_tree_add_190_195_groupi_n_2953 ,in55[2] ,in60[6]);
  nor csa_tree_add_190_195_groupi_g46220(csa_tree_add_190_195_groupi_n_2952 ,in60[13] ,in58[13]);
  or csa_tree_add_190_195_groupi_g46221(csa_tree_add_190_195_groupi_n_2951 ,csa_tree_add_190_195_groupi_n_817 ,csa_tree_add_190_195_groupi_n_918);
  nor csa_tree_add_190_195_groupi_g46222(csa_tree_add_190_195_groupi_n_2950 ,csa_tree_add_190_195_groupi_n_2589 ,csa_tree_add_190_195_groupi_n_692);
  and csa_tree_add_190_195_groupi_g46223(csa_tree_add_190_195_groupi_n_2949 ,csa_tree_add_190_195_groupi_n_358 ,csa_tree_add_190_195_groupi_n_1942);
  or csa_tree_add_190_195_groupi_g46225(csa_tree_add_190_195_groupi_n_2948 ,csa_tree_add_190_195_groupi_n_191 ,csa_tree_add_190_195_groupi_n_1971);
  or csa_tree_add_190_195_groupi_g46226(csa_tree_add_190_195_groupi_n_2947 ,csa_tree_add_190_195_groupi_n_302 ,csa_tree_add_190_195_groupi_n_250);
  nor csa_tree_add_190_195_groupi_g46227(csa_tree_add_190_195_groupi_n_2946 ,csa_tree_add_190_195_groupi_n_1416 ,csa_tree_add_190_195_groupi_n_2635);
  and csa_tree_add_190_195_groupi_g46228(csa_tree_add_190_195_groupi_n_2945 ,csa_tree_add_190_195_groupi_n_389 ,csa_tree_add_190_195_groupi_n_2059);
  nor csa_tree_add_190_195_groupi_g46229(csa_tree_add_190_195_groupi_n_2944 ,csa_tree_add_190_195_groupi_n_1244 ,csa_tree_add_190_195_groupi_n_1165);
  nor csa_tree_add_190_195_groupi_g46230(csa_tree_add_190_195_groupi_n_2943 ,csa_tree_add_190_195_groupi_n_716 ,csa_tree_add_190_195_groupi_n_2509);
  or csa_tree_add_190_195_groupi_g46231(csa_tree_add_190_195_groupi_n_2942 ,csa_tree_add_190_195_groupi_n_1089 ,csa_tree_add_190_195_groupi_n_2059);
  nor csa_tree_add_190_195_groupi_g46233(csa_tree_add_190_195_groupi_n_2941 ,csa_tree_add_190_195_groupi_n_1273 ,csa_tree_add_190_195_groupi_n_238);
  and csa_tree_add_190_195_groupi_g46234(csa_tree_add_190_195_groupi_n_2940 ,in55[3] ,in58[6]);
  and csa_tree_add_190_195_groupi_g46235(csa_tree_add_190_195_groupi_n_2939 ,csa_tree_add_190_195_groupi_n_2155 ,csa_tree_add_190_195_groupi_n_1754);
  and csa_tree_add_190_195_groupi_g46236(csa_tree_add_190_195_groupi_n_2938 ,in55[5] ,in58[8]);
  nor csa_tree_add_190_195_groupi_g46237(csa_tree_add_190_195_groupi_n_2937 ,csa_tree_add_190_195_groupi_n_765 ,csa_tree_add_190_195_groupi_n_1393);
  or csa_tree_add_190_195_groupi_g46238(csa_tree_add_190_195_groupi_n_2936 ,csa_tree_add_190_195_groupi_n_1384 ,csa_tree_add_190_195_groupi_n_720);
  or csa_tree_add_190_195_groupi_g46239(csa_tree_add_190_195_groupi_n_2935 ,csa_tree_add_190_195_groupi_n_2595 ,csa_tree_add_190_195_groupi_n_1338);
  and csa_tree_add_190_195_groupi_g46240(csa_tree_add_190_195_groupi_n_2934 ,csa_tree_add_190_195_groupi_n_469 ,csa_tree_add_190_195_groupi_n_1134);
  or csa_tree_add_190_195_groupi_g46241(csa_tree_add_190_195_groupi_n_2933 ,csa_tree_add_190_195_groupi_n_1891 ,csa_tree_add_190_195_groupi_n_1887);
  nor csa_tree_add_190_195_groupi_g46242(csa_tree_add_190_195_groupi_n_2932 ,csa_tree_add_190_195_groupi_n_622 ,csa_tree_add_190_195_groupi_n_244);
  nor csa_tree_add_190_195_groupi_g46243(csa_tree_add_190_195_groupi_n_2931 ,csa_tree_add_190_195_groupi_n_1488 ,csa_tree_add_190_195_groupi_n_1442);
  nor csa_tree_add_190_195_groupi_g46244(csa_tree_add_190_195_groupi_n_2930 ,csa_tree_add_190_195_groupi_n_1496 ,csa_tree_add_190_195_groupi_n_1559);
  or csa_tree_add_190_195_groupi_g46245(csa_tree_add_190_195_groupi_n_2929 ,csa_tree_add_190_195_groupi_n_2345 ,csa_tree_add_190_195_groupi_n_2621);
  and csa_tree_add_190_195_groupi_g46246(csa_tree_add_190_195_groupi_n_2928 ,in55[8] ,in60[12]);
  or csa_tree_add_190_195_groupi_g46247(csa_tree_add_190_195_groupi_n_2927 ,csa_tree_add_190_195_groupi_n_736 ,csa_tree_add_190_195_groupi_n_2629);
  nor csa_tree_add_190_195_groupi_g46248(csa_tree_add_190_195_groupi_n_2926 ,csa_tree_add_190_195_groupi_n_1568 ,csa_tree_add_190_195_groupi_n_695);
  and csa_tree_add_190_195_groupi_g46249(csa_tree_add_190_195_groupi_n_2925 ,csa_tree_add_190_195_groupi_n_1808 ,csa_tree_add_190_195_groupi_n_820);
  nor csa_tree_add_190_195_groupi_g46250(csa_tree_add_190_195_groupi_n_2924 ,in55[7] ,in60[11]);
  and csa_tree_add_190_195_groupi_g46251(csa_tree_add_190_195_groupi_n_2923 ,csa_tree_add_190_195_groupi_n_1849 ,csa_tree_add_190_195_groupi_n_888);
  or csa_tree_add_190_195_groupi_g46252(csa_tree_add_190_195_groupi_n_2922 ,csa_tree_add_190_195_groupi_n_1505 ,csa_tree_add_190_195_groupi_n_2368);
  nor csa_tree_add_190_195_groupi_g46253(csa_tree_add_190_195_groupi_n_2921 ,csa_tree_add_190_195_groupi_n_1865 ,csa_tree_add_190_195_groupi_n_2057);
  nor csa_tree_add_190_195_groupi_g46254(csa_tree_add_190_195_groupi_n_2920 ,csa_tree_add_190_195_groupi_n_1491 ,csa_tree_add_190_195_groupi_n_1382);
  and csa_tree_add_190_195_groupi_g46255(csa_tree_add_190_195_groupi_n_2919 ,csa_tree_add_190_195_groupi_n_1204 ,in61[3]);
  nor csa_tree_add_190_195_groupi_g46256(csa_tree_add_190_195_groupi_n_2918 ,csa_tree_add_190_195_groupi_n_1393 ,csa_tree_add_190_195_groupi_n_2698);
  or csa_tree_add_190_195_groupi_g46257(csa_tree_add_190_195_groupi_n_2917 ,csa_tree_add_190_195_groupi_n_1137 ,csa_tree_add_190_195_groupi_n_1905);
  or csa_tree_add_190_195_groupi_g46258(csa_tree_add_190_195_groupi_n_2916 ,csa_tree_add_190_195_groupi_n_987 ,csa_tree_add_190_195_groupi_n_841);
  and csa_tree_add_190_195_groupi_g46259(csa_tree_add_190_195_groupi_n_2915 ,csa_tree_add_190_195_groupi_n_362 ,csa_tree_add_190_195_groupi_n_210);
  or csa_tree_add_190_195_groupi_g46260(csa_tree_add_190_195_groupi_n_2914 ,csa_tree_add_190_195_groupi_n_1849 ,csa_tree_add_190_195_groupi_n_844);
  or csa_tree_add_190_195_groupi_g46261(csa_tree_add_190_195_groupi_n_2913 ,csa_tree_add_190_195_groupi_n_1475 ,csa_tree_add_190_195_groupi_n_2341);
  nor csa_tree_add_190_195_groupi_g46262(csa_tree_add_190_195_groupi_n_2912 ,csa_tree_add_190_195_groupi_n_598 ,csa_tree_add_190_195_groupi_n_1915);
  nor csa_tree_add_190_195_groupi_g46263(csa_tree_add_190_195_groupi_n_2911 ,csa_tree_add_190_195_groupi_n_440 ,csa_tree_add_190_195_groupi_n_1129);
  nor csa_tree_add_190_195_groupi_g46264(csa_tree_add_190_195_groupi_n_2910 ,csa_tree_add_190_195_groupi_n_456 ,csa_tree_add_190_195_groupi_n_1183);
  or csa_tree_add_190_195_groupi_g46265(csa_tree_add_190_195_groupi_n_2909 ,csa_tree_add_190_195_groupi_n_1131 ,csa_tree_add_190_195_groupi_n_1033);
  and csa_tree_add_190_195_groupi_g46266(csa_tree_add_190_195_groupi_n_2908 ,in61[14] ,in58[14]);
  or csa_tree_add_190_195_groupi_g46267(csa_tree_add_190_195_groupi_n_2907 ,csa_tree_add_190_195_groupi_n_1893 ,csa_tree_add_190_195_groupi_n_1835);
  nor csa_tree_add_190_195_groupi_g46268(csa_tree_add_190_195_groupi_n_2906 ,csa_tree_add_190_195_groupi_n_1510 ,csa_tree_add_190_195_groupi_n_2700);
  or csa_tree_add_190_195_groupi_g46269(csa_tree_add_190_195_groupi_n_2905 ,csa_tree_add_190_195_groupi_n_2431 ,csa_tree_add_190_195_groupi_n_2728);
  nor csa_tree_add_190_195_groupi_g46270(csa_tree_add_190_195_groupi_n_2904 ,csa_tree_add_190_195_groupi_n_1513 ,csa_tree_add_190_195_groupi_n_2680);
  nor csa_tree_add_190_195_groupi_g46271(csa_tree_add_190_195_groupi_n_2903 ,csa_tree_add_190_195_groupi_n_271 ,csa_tree_add_190_195_groupi_n_1826);
  nor csa_tree_add_190_195_groupi_g46272(csa_tree_add_190_195_groupi_n_2902 ,csa_tree_add_190_195_groupi_n_568 ,csa_tree_add_190_195_groupi_n_227);
  nor csa_tree_add_190_195_groupi_g46273(csa_tree_add_190_195_groupi_n_2901 ,csa_tree_add_190_195_groupi_n_1295 ,csa_tree_add_190_195_groupi_n_2054);
  or csa_tree_add_190_195_groupi_g46274(csa_tree_add_190_195_groupi_n_2900 ,csa_tree_add_190_195_groupi_n_330 ,csa_tree_add_190_195_groupi_n_1977);
  and csa_tree_add_190_195_groupi_g46275(csa_tree_add_190_195_groupi_n_2899 ,csa_tree_add_190_195_groupi_n_889 ,csa_tree_add_190_195_groupi_n_849);
  or csa_tree_add_190_195_groupi_g46276(csa_tree_add_190_195_groupi_n_2898 ,in55[0] ,in61[4]);
  and csa_tree_add_190_195_groupi_g46277(csa_tree_add_190_195_groupi_n_2897 ,csa_tree_add_190_195_groupi_n_1967 ,csa_tree_add_190_195_groupi_n_1035);
  nor csa_tree_add_190_195_groupi_g46278(csa_tree_add_190_195_groupi_n_2896 ,csa_tree_add_190_195_groupi_n_2050 ,csa_tree_add_190_195_groupi_n_1059);
  or csa_tree_add_190_195_groupi_g46279(csa_tree_add_190_195_groupi_n_2895 ,csa_tree_add_190_195_groupi_n_1452 ,csa_tree_add_190_195_groupi_n_1374);
  and csa_tree_add_190_195_groupi_g46280(csa_tree_add_190_195_groupi_n_2894 ,csa_tree_add_190_195_groupi_n_2214 ,csa_tree_add_190_195_groupi_n_1744);
  or csa_tree_add_190_195_groupi_g46281(csa_tree_add_190_195_groupi_n_2893 ,csa_tree_add_190_195_groupi_n_2596 ,csa_tree_add_190_195_groupi_n_1446);
  or csa_tree_add_190_195_groupi_g46282(csa_tree_add_190_195_groupi_n_2892 ,csa_tree_add_190_195_groupi_n_321 ,csa_tree_add_190_195_groupi_n_1164);
  and csa_tree_add_190_195_groupi_g46283(csa_tree_add_190_195_groupi_n_2891 ,csa_tree_add_190_195_groupi_n_350 ,csa_tree_add_190_195_groupi_n_1859);
  or csa_tree_add_190_195_groupi_g46284(csa_tree_add_190_195_groupi_n_2890 ,csa_tree_add_190_195_groupi_n_831 ,csa_tree_add_190_195_groupi_n_1362);
  nor csa_tree_add_190_195_groupi_g46285(csa_tree_add_190_195_groupi_n_2889 ,csa_tree_add_190_195_groupi_n_284 ,csa_tree_add_190_195_groupi_n_788);
  or csa_tree_add_190_195_groupi_g46286(csa_tree_add_190_195_groupi_n_2888 ,csa_tree_add_190_195_groupi_n_1450 ,csa_tree_add_190_195_groupi_n_2469);
  nor csa_tree_add_190_195_groupi_g46287(csa_tree_add_190_195_groupi_n_2887 ,csa_tree_add_190_195_groupi_n_1570 ,csa_tree_add_190_195_groupi_n_2619);
  and csa_tree_add_190_195_groupi_g46288(csa_tree_add_190_195_groupi_n_2886 ,csa_tree_add_190_195_groupi_n_949 ,csa_tree_add_190_195_groupi_n_838);
  or csa_tree_add_190_195_groupi_g46289(csa_tree_add_190_195_groupi_n_2885 ,csa_tree_add_190_195_groupi_n_289 ,in60[2]);
  or csa_tree_add_190_195_groupi_g46290(csa_tree_add_190_195_groupi_n_2884 ,in55[8] ,in58[11]);
  nor csa_tree_add_190_195_groupi_g46291(csa_tree_add_190_195_groupi_n_2883 ,csa_tree_add_190_195_groupi_n_1305 ,csa_tree_add_190_195_groupi_n_1991);
  or csa_tree_add_190_195_groupi_g46292(csa_tree_add_190_195_groupi_n_2882 ,csa_tree_add_190_195_groupi_n_1877 ,csa_tree_add_190_195_groupi_n_1810);
  or csa_tree_add_190_195_groupi_g46293(csa_tree_add_190_195_groupi_n_2881 ,csa_tree_add_190_195_groupi_n_618 ,csa_tree_add_190_195_groupi_n_1271);
  and csa_tree_add_190_195_groupi_g46294(csa_tree_add_190_195_groupi_n_2880 ,csa_tree_add_190_195_groupi_n_226 ,csa_tree_add_190_195_groupi_n_568);
  nor csa_tree_add_190_195_groupi_g46295(csa_tree_add_190_195_groupi_n_2879 ,csa_tree_add_190_195_groupi_n_537 ,csa_tree_add_190_195_groupi_n_2062);
  or csa_tree_add_190_195_groupi_g46296(csa_tree_add_190_195_groupi_n_2878 ,csa_tree_add_190_195_groupi_n_2633 ,csa_tree_add_190_195_groupi_n_2686);
  or csa_tree_add_190_195_groupi_g46297(csa_tree_add_190_195_groupi_n_2877 ,csa_tree_add_190_195_groupi_n_1179 ,csa_tree_add_190_195_groupi_n_1027);
  and csa_tree_add_190_195_groupi_g46298(csa_tree_add_190_195_groupi_n_2876 ,csa_tree_add_190_195_groupi_n_219 ,csa_tree_add_190_195_groupi_n_916);
  or csa_tree_add_190_195_groupi_g46299(csa_tree_add_190_195_groupi_n_2875 ,in55[3] ,in58[6]);
  or csa_tree_add_190_195_groupi_g46300(csa_tree_add_190_195_groupi_n_2874 ,csa_tree_add_190_195_groupi_n_391 ,csa_tree_add_190_195_groupi_n_1062);
  nor csa_tree_add_190_195_groupi_g46301(csa_tree_add_190_195_groupi_n_2873 ,csa_tree_add_190_195_groupi_n_1123 ,in60[4]);
  nor csa_tree_add_190_195_groupi_g46302(csa_tree_add_190_195_groupi_n_2872 ,csa_tree_add_190_195_groupi_n_572 ,csa_tree_add_190_195_groupi_n_1281);
  or csa_tree_add_190_195_groupi_g46303(csa_tree_add_190_195_groupi_n_2871 ,csa_tree_add_190_195_groupi_n_2590 ,csa_tree_add_190_195_groupi_n_2552);
  or csa_tree_add_190_195_groupi_g46304(csa_tree_add_190_195_groupi_n_2870 ,csa_tree_add_190_195_groupi_n_2157 ,csa_tree_add_190_195_groupi_n_1206);
  and csa_tree_add_190_195_groupi_g46305(csa_tree_add_190_195_groupi_n_2869 ,csa_tree_add_190_195_groupi_n_295 ,csa_tree_add_190_195_groupi_n_1111);
  and csa_tree_add_190_195_groupi_g46306(csa_tree_add_190_195_groupi_n_2868 ,csa_tree_add_190_195_groupi_n_188 ,csa_tree_add_190_195_groupi_n_202);
  nor csa_tree_add_190_195_groupi_g46307(csa_tree_add_190_195_groupi_n_2867 ,in55[7] ,in58[10]);
  nor csa_tree_add_190_195_groupi_g46308(csa_tree_add_190_195_groupi_n_2866 ,csa_tree_add_190_195_groupi_n_737 ,csa_tree_add_190_195_groupi_n_2543);
  or csa_tree_add_190_195_groupi_g46309(csa_tree_add_190_195_groupi_n_2865 ,csa_tree_add_190_195_groupi_n_2468 ,csa_tree_add_190_195_groupi_n_2723);
  and csa_tree_add_190_195_groupi_g46310(csa_tree_add_190_195_groupi_n_2864 ,csa_tree_add_190_195_groupi_n_1850 ,csa_tree_add_190_195_groupi_n_1847);
  nor csa_tree_add_190_195_groupi_g46311(csa_tree_add_190_195_groupi_n_2863 ,csa_tree_add_190_195_groupi_n_781 ,csa_tree_add_190_195_groupi_n_1413);
  nor csa_tree_add_190_195_groupi_g46312(csa_tree_add_190_195_groupi_n_2862 ,csa_tree_add_190_195_groupi_n_808 ,csa_tree_add_190_195_groupi_n_1681);
  nor csa_tree_add_190_195_groupi_g46313(csa_tree_add_190_195_groupi_n_2861 ,csa_tree_add_190_195_groupi_n_351 ,csa_tree_add_190_195_groupi_n_891);
  or csa_tree_add_190_195_groupi_g46314(csa_tree_add_190_195_groupi_n_2860 ,csa_tree_add_190_195_groupi_n_1969 ,csa_tree_add_190_195_groupi_n_373);
  nor csa_tree_add_190_195_groupi_g46315(csa_tree_add_190_195_groupi_n_2859 ,csa_tree_add_190_195_groupi_n_1261 ,csa_tree_add_190_195_groupi_n_1144);
  and csa_tree_add_190_195_groupi_g46316(csa_tree_add_190_195_groupi_n_2858 ,csa_tree_add_190_195_groupi_n_622 ,csa_tree_add_190_195_groupi_n_243);
  or csa_tree_add_190_195_groupi_g46317(csa_tree_add_190_195_groupi_n_2857 ,csa_tree_add_190_195_groupi_n_301 ,csa_tree_add_190_195_groupi_n_826);
  or csa_tree_add_190_195_groupi_g46318(csa_tree_add_190_195_groupi_n_2856 ,csa_tree_add_190_195_groupi_n_597 ,csa_tree_add_190_195_groupi_n_984);
  or csa_tree_add_190_195_groupi_g46319(csa_tree_add_190_195_groupi_n_2855 ,csa_tree_add_190_195_groupi_n_256 ,csa_tree_add_190_195_groupi_n_1176);
  nor csa_tree_add_190_195_groupi_g46320(csa_tree_add_190_195_groupi_n_2854 ,csa_tree_add_190_195_groupi_n_1386 ,csa_tree_add_190_195_groupi_n_2478);
  or csa_tree_add_190_195_groupi_g46321(csa_tree_add_190_195_groupi_n_2853 ,csa_tree_add_190_195_groupi_n_2459 ,csa_tree_add_190_195_groupi_n_2612);
  or csa_tree_add_190_195_groupi_g46322(csa_tree_add_190_195_groupi_n_2852 ,csa_tree_add_190_195_groupi_n_1059 ,csa_tree_add_190_195_groupi_n_1039);
  nor csa_tree_add_190_195_groupi_g46323(csa_tree_add_190_195_groupi_n_2851 ,csa_tree_add_190_195_groupi_n_490 ,csa_tree_add_190_195_groupi_n_1195);
  and csa_tree_add_190_195_groupi_g46324(csa_tree_add_190_195_groupi_n_2850 ,csa_tree_add_190_195_groupi_n_933 ,csa_tree_add_190_195_groupi_n_819);
  and csa_tree_add_190_195_groupi_g46325(csa_tree_add_190_195_groupi_n_2849 ,csa_tree_add_190_195_groupi_n_2086 ,csa_tree_add_190_195_groupi_n_850);
  or csa_tree_add_190_195_groupi_g46326(csa_tree_add_190_195_groupi_n_2848 ,csa_tree_add_190_195_groupi_n_2039 ,csa_tree_add_190_195_groupi_n_1924);
  or csa_tree_add_190_195_groupi_g46327(csa_tree_add_190_195_groupi_n_2847 ,csa_tree_add_190_195_groupi_n_342 ,csa_tree_add_190_195_groupi_n_1102);
  or csa_tree_add_190_195_groupi_g46328(csa_tree_add_190_195_groupi_n_2846 ,csa_tree_add_190_195_groupi_n_398 ,csa_tree_add_190_195_groupi_n_1146);
  nor csa_tree_add_190_195_groupi_g46329(csa_tree_add_190_195_groupi_n_2845 ,csa_tree_add_190_195_groupi_n_744 ,csa_tree_add_190_195_groupi_n_1382);
  nor csa_tree_add_190_195_groupi_g46330(csa_tree_add_190_195_groupi_n_2844 ,csa_tree_add_190_195_groupi_n_2211 ,csa_tree_add_190_195_groupi_n_1832);
  nor csa_tree_add_190_195_groupi_g46331(csa_tree_add_190_195_groupi_n_2843 ,csa_tree_add_190_195_groupi_n_2575 ,csa_tree_add_190_195_groupi_n_1522);
  or csa_tree_add_190_195_groupi_g46332(csa_tree_add_190_195_groupi_n_2842 ,csa_tree_add_190_195_groupi_n_2051 ,csa_tree_add_190_195_groupi_n_297);
  nor csa_tree_add_190_195_groupi_g46333(csa_tree_add_190_195_groupi_n_2841 ,csa_tree_add_190_195_groupi_n_1480 ,csa_tree_add_190_195_groupi_n_1428);
  or csa_tree_add_190_195_groupi_g46334(csa_tree_add_190_195_groupi_n_2840 ,csa_tree_add_190_195_groupi_n_1208 ,csa_tree_add_190_195_groupi_n_1220);
  nor csa_tree_add_190_195_groupi_g46335(csa_tree_add_190_195_groupi_n_2839 ,csa_tree_add_190_195_groupi_n_1975 ,csa_tree_add_190_195_groupi_n_1150);
  nor csa_tree_add_190_195_groupi_g46336(csa_tree_add_190_195_groupi_n_2838 ,csa_tree_add_190_195_groupi_n_1153 ,csa_tree_add_190_195_groupi_n_1814);
  or csa_tree_add_190_195_groupi_g46337(csa_tree_add_190_195_groupi_n_2837 ,csa_tree_add_190_195_groupi_n_1967 ,csa_tree_add_190_195_groupi_n_1036);
  nor csa_tree_add_190_195_groupi_g46338(csa_tree_add_190_195_groupi_n_2836 ,csa_tree_add_190_195_groupi_n_552 ,csa_tree_add_190_195_groupi_n_1135);
  and csa_tree_add_190_195_groupi_g46339(csa_tree_add_190_195_groupi_n_2835 ,csa_tree_add_190_195_groupi_n_1263 ,csa_tree_add_190_195_groupi_n_1867);
  nor csa_tree_add_190_195_groupi_g46340(csa_tree_add_190_195_groupi_n_2834 ,csa_tree_add_190_195_groupi_n_589 ,csa_tree_add_190_195_groupi_n_1930);
  nor csa_tree_add_190_195_groupi_g46341(csa_tree_add_190_195_groupi_n_2833 ,csa_tree_add_190_195_groupi_n_1128 ,csa_tree_add_190_195_groupi_n_1706);
  nor csa_tree_add_190_195_groupi_g46342(csa_tree_add_190_195_groupi_n_2832 ,csa_tree_add_190_195_groupi_n_437 ,csa_tree_add_190_195_groupi_n_876);
  nor csa_tree_add_190_195_groupi_g46343(csa_tree_add_190_195_groupi_n_2831 ,csa_tree_add_190_195_groupi_n_274 ,csa_tree_add_190_195_groupi_n_1838);
  or csa_tree_add_190_195_groupi_g46344(csa_tree_add_190_195_groupi_n_2830 ,csa_tree_add_190_195_groupi_n_1462 ,csa_tree_add_190_195_groupi_n_2354);
  and csa_tree_add_190_195_groupi_g46345(csa_tree_add_190_195_groupi_n_2829 ,csa_tree_add_190_195_groupi_n_435 ,csa_tree_add_190_195_groupi_n_2088);
  nor csa_tree_add_190_195_groupi_g46346(csa_tree_add_190_195_groupi_n_2828 ,csa_tree_add_190_195_groupi_n_1420 ,csa_tree_add_190_195_groupi_n_2437);
  nor csa_tree_add_190_195_groupi_g46347(csa_tree_add_190_195_groupi_n_2827 ,csa_tree_add_190_195_groupi_n_428 ,csa_tree_add_190_195_groupi_n_1870);
  or csa_tree_add_190_195_groupi_g46348(csa_tree_add_190_195_groupi_n_2826 ,csa_tree_add_190_195_groupi_n_336 ,csa_tree_add_190_195_groupi_n_1877);
  or csa_tree_add_190_195_groupi_g46349(csa_tree_add_190_195_groupi_n_2825 ,csa_tree_add_190_195_groupi_n_2610 ,csa_tree_add_190_195_groupi_n_2456);
  nor csa_tree_add_190_195_groupi_g46350(csa_tree_add_190_195_groupi_n_2824 ,csa_tree_add_190_195_groupi_n_764 ,csa_tree_add_190_195_groupi_n_1366);
  or csa_tree_add_190_195_groupi_g46351(csa_tree_add_190_195_groupi_n_2823 ,csa_tree_add_190_195_groupi_n_286 ,csa_tree_add_190_195_groupi_n_1048);
  nor csa_tree_add_190_195_groupi_g46352(csa_tree_add_190_195_groupi_n_2822 ,csa_tree_add_190_195_groupi_n_546 ,csa_tree_add_190_195_groupi_n_1218);
  or csa_tree_add_190_195_groupi_g46353(csa_tree_add_190_195_groupi_n_2821 ,csa_tree_add_190_195_groupi_n_861 ,csa_tree_add_190_195_groupi_n_1083);
  nor csa_tree_add_190_195_groupi_g46354(csa_tree_add_190_195_groupi_n_2820 ,csa_tree_add_190_195_groupi_n_1438 ,csa_tree_add_190_195_groupi_n_2609);
  and csa_tree_add_190_195_groupi_g46355(csa_tree_add_190_195_groupi_n_2819 ,csa_tree_add_190_195_groupi_n_1012 ,csa_tree_add_190_195_groupi_n_1829);
  nor csa_tree_add_190_195_groupi_g46356(csa_tree_add_190_195_groupi_n_2818 ,csa_tree_add_190_195_groupi_n_1434 ,csa_tree_add_190_195_groupi_n_1501);
  nor csa_tree_add_190_195_groupi_g46357(csa_tree_add_190_195_groupi_n_2817 ,csa_tree_add_190_195_groupi_n_2041 ,csa_tree_add_190_195_groupi_n_1827);
  nor csa_tree_add_190_195_groupi_g46358(csa_tree_add_190_195_groupi_n_2816 ,csa_tree_add_190_195_groupi_n_1548 ,csa_tree_add_190_195_groupi_n_2512);
  and csa_tree_add_190_195_groupi_g46359(csa_tree_add_190_195_groupi_n_2815 ,csa_tree_add_190_195_groupi_n_307 ,csa_tree_add_190_195_groupi_n_1843);
  nor csa_tree_add_190_195_groupi_g46360(csa_tree_add_190_195_groupi_n_2814 ,csa_tree_add_190_195_groupi_n_1289 ,csa_tree_add_190_195_groupi_n_1995);
  and csa_tree_add_190_195_groupi_g46361(csa_tree_add_190_195_groupi_n_2813 ,csa_tree_add_190_195_groupi_n_281 ,csa_tree_add_190_195_groupi_n_981);
  and csa_tree_add_190_195_groupi_g46362(csa_tree_add_190_195_groupi_n_2812 ,csa_tree_add_190_195_groupi_n_1120 ,csa_tree_add_190_195_groupi_n_1777);
  or csa_tree_add_190_195_groupi_g46363(csa_tree_add_190_195_groupi_n_2811 ,csa_tree_add_190_195_groupi_n_1970 ,csa_tree_add_190_195_groupi_n_1966);
  nor csa_tree_add_190_195_groupi_g46364(csa_tree_add_190_195_groupi_n_2810 ,csa_tree_add_190_195_groupi_n_310 ,in61[2]);
  nor csa_tree_add_190_195_groupi_g46365(csa_tree_add_190_195_groupi_n_2809 ,csa_tree_add_190_195_groupi_n_724 ,csa_tree_add_190_195_groupi_n_1388);
  nor csa_tree_add_190_195_groupi_g46366(csa_tree_add_190_195_groupi_n_2808 ,csa_tree_add_190_195_groupi_n_399 ,csa_tree_add_190_195_groupi_n_2007);
  nor csa_tree_add_190_195_groupi_g46367(csa_tree_add_190_195_groupi_n_2807 ,csa_tree_add_190_195_groupi_n_1267 ,csa_tree_add_190_195_groupi_n_1973);
  or csa_tree_add_190_195_groupi_g46368(csa_tree_add_190_195_groupi_n_2806 ,csa_tree_add_190_195_groupi_n_1380 ,csa_tree_add_190_195_groupi_n_2696);
  and csa_tree_add_190_195_groupi_g46369(csa_tree_add_190_195_groupi_n_2805 ,csa_tree_add_190_195_groupi_n_609 ,csa_tree_add_190_195_groupi_n_1261);
  nor csa_tree_add_190_195_groupi_g46370(csa_tree_add_190_195_groupi_n_2804 ,csa_tree_add_190_195_groupi_n_1240 ,csa_tree_add_190_195_groupi_n_1614);
  or csa_tree_add_190_195_groupi_g46371(csa_tree_add_190_195_groupi_n_2803 ,csa_tree_add_190_195_groupi_n_453 ,csa_tree_add_190_195_groupi_n_1776);
  and csa_tree_add_190_195_groupi_g46372(csa_tree_add_190_195_groupi_n_2802 ,csa_tree_add_190_195_groupi_n_2209 ,csa_tree_add_190_195_groupi_n_2215);
  or csa_tree_add_190_195_groupi_g46373(csa_tree_add_190_195_groupi_n_2801 ,csa_tree_add_190_195_groupi_n_1197 ,csa_tree_add_190_195_groupi_n_1675);
  nor csa_tree_add_190_195_groupi_g46374(csa_tree_add_190_195_groupi_n_2800 ,csa_tree_add_190_195_groupi_n_832 ,csa_tree_add_190_195_groupi_n_2606);
  nor csa_tree_add_190_195_groupi_g46375(csa_tree_add_190_195_groupi_n_2799 ,in55[6] ,in58[9]);
  and csa_tree_add_190_195_groupi_g46376(csa_tree_add_190_195_groupi_n_2798 ,csa_tree_add_190_195_groupi_n_1185 ,csa_tree_add_190_195_groupi_n_212);
  nor csa_tree_add_190_195_groupi_g46377(csa_tree_add_190_195_groupi_n_2797 ,csa_tree_add_190_195_groupi_n_1498 ,csa_tree_add_190_195_groupi_n_2613);
  or csa_tree_add_190_195_groupi_g46378(csa_tree_add_190_195_groupi_n_2796 ,csa_tree_add_190_195_groupi_n_966 ,csa_tree_add_190_195_groupi_n_1597);
  nor csa_tree_add_190_195_groupi_g46379(csa_tree_add_190_195_groupi_n_2795 ,csa_tree_add_190_195_groupi_n_1552 ,csa_tree_add_190_195_groupi_n_2630);
  or csa_tree_add_190_195_groupi_g46380(csa_tree_add_190_195_groupi_n_2794 ,csa_tree_add_190_195_groupi_n_726 ,csa_tree_add_190_195_groupi_n_2470);
  or csa_tree_add_190_195_groupi_g46381(csa_tree_add_190_195_groupi_n_2793 ,csa_tree_add_190_195_groupi_n_360 ,csa_tree_add_190_195_groupi_n_1267);
  and csa_tree_add_190_195_groupi_g46382(csa_tree_add_190_195_groupi_n_2792 ,csa_tree_add_190_195_groupi_n_323 ,csa_tree_add_190_195_groupi_n_196);
  or csa_tree_add_190_195_groupi_g46383(csa_tree_add_190_195_groupi_n_2791 ,csa_tree_add_190_195_groupi_n_1104 ,csa_tree_add_190_195_groupi_n_1018);
  or csa_tree_add_190_195_groupi_g46384(csa_tree_add_190_195_groupi_n_2790 ,csa_tree_add_190_195_groupi_n_1506 ,csa_tree_add_190_195_groupi_n_2620);
  nor csa_tree_add_190_195_groupi_g46385(csa_tree_add_190_195_groupi_n_2789 ,csa_tree_add_190_195_groupi_n_1251 ,csa_tree_add_190_195_groupi_n_1751);
  nor csa_tree_add_190_195_groupi_g46386(csa_tree_add_190_195_groupi_n_2788 ,csa_tree_add_190_195_groupi_n_420 ,csa_tree_add_190_195_groupi_n_1242);
  nor csa_tree_add_190_195_groupi_g46387(csa_tree_add_190_195_groupi_n_2787 ,csa_tree_add_190_195_groupi_n_2042 ,csa_tree_add_190_195_groupi_n_1860);
  or csa_tree_add_190_195_groupi_g46388(csa_tree_add_190_195_groupi_n_2786 ,csa_tree_add_190_195_groupi_n_2508 ,csa_tree_add_190_195_groupi_n_2712);
  and csa_tree_add_190_195_groupi_g46389(csa_tree_add_190_195_groupi_n_2785 ,in61[15] ,in59[15]);
  and csa_tree_add_190_195_groupi_g46390(csa_tree_add_190_195_groupi_n_2784 ,in55[8] ,in58[11]);
  or csa_tree_add_190_195_groupi_g46391(csa_tree_add_190_195_groupi_n_2783 ,csa_tree_add_190_195_groupi_n_279 ,csa_tree_add_190_195_groupi_n_1889);
  or csa_tree_add_190_195_groupi_g46392(csa_tree_add_190_195_groupi_n_2782 ,csa_tree_add_190_195_groupi_n_731 ,csa_tree_add_190_195_groupi_n_1356);
  or csa_tree_add_190_195_groupi_g46393(csa_tree_add_190_195_groupi_n_2781 ,csa_tree_add_190_195_groupi_n_1232 ,csa_tree_add_190_195_groupi_n_321);
  and csa_tree_add_190_195_groupi_g46394(csa_tree_add_190_195_groupi_n_2780 ,csa_tree_add_190_195_groupi_n_191 ,csa_tree_add_190_195_groupi_n_1970);
  or csa_tree_add_190_195_groupi_g46395(csa_tree_add_190_195_groupi_n_2779 ,csa_tree_add_190_195_groupi_n_2607 ,csa_tree_add_190_195_groupi_n_2540);
  and csa_tree_add_190_195_groupi_g46396(csa_tree_add_190_195_groupi_n_2778 ,csa_tree_add_190_195_groupi_n_246 ,csa_tree_add_190_195_groupi_n_1746);
  or csa_tree_add_190_195_groupi_g46397(csa_tree_add_190_195_groupi_n_2777 ,csa_tree_add_190_195_groupi_n_315 ,in61[3]);
  and csa_tree_add_190_195_groupi_g46398(csa_tree_add_190_195_groupi_n_2776 ,csa_tree_add_190_195_groupi_n_1122 ,in60[4]);
  or csa_tree_add_190_195_groupi_g46399(csa_tree_add_190_195_groupi_n_2775 ,csa_tree_add_190_195_groupi_n_582 ,csa_tree_add_190_195_groupi_n_2088);
  and csa_tree_add_190_195_groupi_g46400(csa_tree_add_190_195_groupi_n_2774 ,csa_tree_add_190_195_groupi_n_604 ,csa_tree_add_190_195_groupi_n_222);
  nor csa_tree_add_190_195_groupi_g46401(csa_tree_add_190_195_groupi_n_2773 ,csa_tree_add_190_195_groupi_n_1519 ,csa_tree_add_190_195_groupi_n_2448);
  or csa_tree_add_190_195_groupi_g46402(csa_tree_add_190_195_groupi_n_2772 ,in55[0] ,csa_tree_add_190_195_groupi_n_325);
  nor csa_tree_add_190_195_groupi_g46403(csa_tree_add_190_195_groupi_n_2771 ,csa_tree_add_190_195_groupi_n_740 ,csa_tree_add_190_195_groupi_n_2455);
  or csa_tree_add_190_195_groupi_g46404(csa_tree_add_190_195_groupi_n_2770 ,csa_tree_add_190_195_groupi_n_1015 ,csa_tree_add_190_195_groupi_n_1951);
  or csa_tree_add_190_195_groupi_g46405(csa_tree_add_190_195_groupi_n_2769 ,csa_tree_add_190_195_groupi_n_2216 ,csa_tree_add_190_195_groupi_n_1920);
  or csa_tree_add_190_195_groupi_g46406(csa_tree_add_190_195_groupi_n_2768 ,csa_tree_add_190_195_groupi_n_1477 ,csa_tree_add_190_195_groupi_n_2666);
  nor csa_tree_add_190_195_groupi_g46407(csa_tree_add_190_195_groupi_n_2767 ,in55[4] ,in60[8]);
  or csa_tree_add_190_195_groupi_g46408(csa_tree_add_190_195_groupi_n_2766 ,csa_tree_add_190_195_groupi_n_2585 ,csa_tree_add_190_195_groupi_n_2702);
  or csa_tree_add_190_195_groupi_g46409(csa_tree_add_190_195_groupi_n_2765 ,csa_tree_add_190_195_groupi_n_822 ,csa_tree_add_190_195_groupi_n_2629);
  and csa_tree_add_190_195_groupi_g46410(csa_tree_add_190_195_groupi_n_2764 ,csa_tree_add_190_195_groupi_n_233 ,csa_tree_add_190_195_groupi_n_299);
  nor csa_tree_add_190_195_groupi_g46411(csa_tree_add_190_195_groupi_n_2763 ,csa_tree_add_190_195_groupi_n_1108 ,csa_tree_add_190_195_groupi_n_909);
  or csa_tree_add_190_195_groupi_g46412(csa_tree_add_190_195_groupi_n_2762 ,csa_tree_add_190_195_groupi_n_1372 ,csa_tree_add_190_195_groupi_n_2516);
  or csa_tree_add_190_195_groupi_g46413(csa_tree_add_190_195_groupi_n_2761 ,csa_tree_add_190_195_groupi_n_676 ,csa_tree_add_190_195_groupi_n_2523);
  nor csa_tree_add_190_195_groupi_g46414(csa_tree_add_190_195_groupi_n_2760 ,csa_tree_add_190_195_groupi_n_583 ,csa_tree_add_190_195_groupi_n_2214);
  nor csa_tree_add_190_195_groupi_g46415(csa_tree_add_190_195_groupi_n_2759 ,csa_tree_add_190_195_groupi_n_528 ,csa_tree_add_190_195_groupi_n_894);
  or csa_tree_add_190_195_groupi_g46416(csa_tree_add_190_195_groupi_n_2758 ,csa_tree_add_190_195_groupi_n_2369 ,csa_tree_add_190_195_groupi_n_2445);
  and csa_tree_add_190_195_groupi_g46417(csa_tree_add_190_195_groupi_n_2757 ,csa_tree_add_190_195_groupi_n_1848 ,csa_tree_add_190_195_groupi_n_1847);
  or csa_tree_add_190_195_groupi_g46418(csa_tree_add_190_195_groupi_n_2756 ,csa_tree_add_190_195_groupi_n_2155 ,csa_tree_add_190_195_groupi_n_1754);
  nor csa_tree_add_190_195_groupi_g46419(csa_tree_add_190_195_groupi_n_2755 ,csa_tree_add_190_195_groupi_n_2577 ,csa_tree_add_190_195_groupi_n_2443);
  and csa_tree_add_190_195_groupi_g46420(csa_tree_add_190_195_groupi_n_2754 ,csa_tree_add_190_195_groupi_n_2157 ,csa_tree_add_190_195_groupi_n_194);
  or csa_tree_add_190_195_groupi_g46421(csa_tree_add_190_195_groupi_n_2753 ,csa_tree_add_190_195_groupi_n_512 ,csa_tree_add_190_195_groupi_n_1746);
  nor csa_tree_add_190_195_groupi_g46422(csa_tree_add_190_195_groupi_n_2752 ,csa_tree_add_190_195_groupi_n_1411 ,csa_tree_add_190_195_groupi_n_698);
  nor csa_tree_add_190_195_groupi_g46423(csa_tree_add_190_195_groupi_n_2751 ,csa_tree_add_190_195_groupi_n_771 ,csa_tree_add_190_195_groupi_n_2453);
  nor csa_tree_add_190_195_groupi_g46424(csa_tree_add_190_195_groupi_n_2750 ,csa_tree_add_190_195_groupi_n_1406 ,csa_tree_add_190_195_groupi_n_2542);
  and csa_tree_add_190_195_groupi_g46425(csa_tree_add_190_195_groupi_n_2749 ,csa_tree_add_190_195_groupi_n_825 ,csa_tree_add_190_195_groupi_n_1675);
  or csa_tree_add_190_195_groupi_g46426(csa_tree_add_190_195_groupi_n_2748 ,csa_tree_add_190_195_groupi_n_1395 ,csa_tree_add_190_195_groupi_n_2645);
  or csa_tree_add_190_195_groupi_g46427(csa_tree_add_190_195_groupi_n_2747 ,csa_tree_add_190_195_groupi_n_338 ,csa_tree_add_190_195_groupi_n_1970);
  nor csa_tree_add_190_195_groupi_g46428(csa_tree_add_190_195_groupi_n_2746 ,csa_tree_add_190_195_groupi_n_1171 ,csa_tree_add_190_195_groupi_n_1966);
  or csa_tree_add_190_195_groupi_g46429(csa_tree_add_190_195_groupi_n_2745 ,csa_tree_add_190_195_groupi_n_1702 ,csa_tree_add_190_195_groupi_n_921);
  and csa_tree_add_190_195_groupi_g46430(csa_tree_add_190_195_groupi_n_2744 ,csa_tree_add_190_195_groupi_n_496 ,csa_tree_add_190_195_groupi_n_1832);
  nor csa_tree_add_190_195_groupi_g46431(csa_tree_add_190_195_groupi_n_2743 ,csa_tree_add_190_195_groupi_n_581 ,csa_tree_add_190_195_groupi_n_2153);
  or csa_tree_add_190_195_groupi_g46432(csa_tree_add_190_195_groupi_n_2742 ,csa_tree_add_190_195_groupi_n_454 ,csa_tree_add_190_195_groupi_n_891);
  nor csa_tree_add_190_195_groupi_g46433(csa_tree_add_190_195_groupi_n_2741 ,in55[5] ,in60[9]);
  or csa_tree_add_190_195_groupi_g46434(csa_tree_add_190_195_groupi_n_2740 ,csa_tree_add_190_195_groupi_n_1358 ,csa_tree_add_190_195_groupi_n_2534);
  or csa_tree_add_190_195_groupi_g46435(csa_tree_add_190_195_groupi_n_2739 ,csa_tree_add_190_195_groupi_n_209 ,csa_tree_add_190_195_groupi_n_246);
  or csa_tree_add_190_195_groupi_g46436(csa_tree_add_190_195_groupi_n_2738 ,csa_tree_add_190_195_groupi_n_1708 ,csa_tree_add_190_195_groupi_n_1999);
  and csa_tree_add_190_195_groupi_g46437(csa_tree_add_190_195_groupi_n_2737 ,csa_tree_add_190_195_groupi_n_204 ,csa_tree_add_190_195_groupi_n_1703);
  nor csa_tree_add_190_195_groupi_g46438(csa_tree_add_190_195_groupi_n_2736 ,csa_tree_add_190_195_groupi_n_1907 ,csa_tree_add_190_195_groupi_n_1090);
  or csa_tree_add_190_195_groupi_g46439(csa_tree_add_190_195_groupi_n_2735 ,csa_tree_add_190_195_groupi_n_2486 ,csa_tree_add_190_195_groupi_n_2531);
  or csa_tree_add_190_195_groupi_g46440(csa_tree_add_190_195_groupi_n_2734 ,csa_tree_add_190_195_groupi_n_603 ,csa_tree_add_190_195_groupi_n_2210);
  and csa_tree_add_190_195_groupi_g46441(csa_tree_add_190_195_groupi_n_3226 ,csa_tree_add_190_195_groupi_n_1077 ,csa_tree_add_190_195_groupi_n_2052);
  and csa_tree_add_190_195_groupi_g46442(csa_tree_add_190_195_groupi_n_3225 ,csa_tree_add_190_195_groupi_n_2706 ,csa_tree_add_190_195_groupi_n_2677);
  or csa_tree_add_190_195_groupi_g46443(csa_tree_add_190_195_groupi_n_3223 ,csa_tree_add_190_195_groupi_n_347 ,csa_tree_add_190_195_groupi_n_382);
  or csa_tree_add_190_195_groupi_g46444(csa_tree_add_190_195_groupi_n_3221 ,csa_tree_add_190_195_groupi_n_1865 ,csa_tree_add_190_195_groupi_n_1971);
  and csa_tree_add_190_195_groupi_g46445(csa_tree_add_190_195_groupi_n_3219 ,csa_tree_add_190_195_groupi_n_1455 ,csa_tree_add_190_195_groupi_n_2725);
  and csa_tree_add_190_195_groupi_g46446(csa_tree_add_190_195_groupi_n_3218 ,csa_tree_add_190_195_groupi_n_822 ,csa_tree_add_190_195_groupi_n_2562);
  and csa_tree_add_190_195_groupi_g46447(csa_tree_add_190_195_groupi_n_3217 ,csa_tree_add_190_195_groupi_n_1452 ,csa_tree_add_190_195_groupi_n_2676);
  or csa_tree_add_190_195_groupi_g46448(csa_tree_add_190_195_groupi_n_3215 ,csa_tree_add_190_195_groupi_n_823 ,csa_tree_add_190_195_groupi_n_2562);
  or csa_tree_add_190_195_groupi_g46449(csa_tree_add_190_195_groupi_n_3213 ,csa_tree_add_190_195_groupi_n_1456 ,csa_tree_add_190_195_groupi_n_2725);
  and csa_tree_add_190_195_groupi_g46450(csa_tree_add_190_195_groupi_n_3211 ,csa_tree_add_190_195_groupi_n_685 ,csa_tree_add_190_195_groupi_n_2373);
  or csa_tree_add_190_195_groupi_g46451(csa_tree_add_190_195_groupi_n_3210 ,csa_tree_add_190_195_groupi_n_2521 ,csa_tree_add_190_195_groupi_n_2692);
  and csa_tree_add_190_195_groupi_g46452(csa_tree_add_190_195_groupi_n_3209 ,csa_tree_add_190_195_groupi_n_248 ,csa_tree_add_190_195_groupi_n_1828);
  and csa_tree_add_190_195_groupi_g46453(csa_tree_add_190_195_groupi_n_3208 ,csa_tree_add_190_195_groupi_n_1342 ,csa_tree_add_190_195_groupi_n_1340);
  or csa_tree_add_190_195_groupi_g46454(csa_tree_add_190_195_groupi_n_3207 ,csa_tree_add_190_195_groupi_n_1334 ,csa_tree_add_190_195_groupi_n_2567);
  or csa_tree_add_190_195_groupi_g46455(csa_tree_add_190_195_groupi_n_3206 ,csa_tree_add_190_195_groupi_n_707 ,csa_tree_add_190_195_groupi_n_2591);
  or csa_tree_add_190_195_groupi_g46456(csa_tree_add_190_195_groupi_n_3205 ,csa_tree_add_190_195_groupi_n_2593 ,csa_tree_add_190_195_groupi_n_2564);
  and csa_tree_add_190_195_groupi_g46457(csa_tree_add_190_195_groupi_n_3203 ,csa_tree_add_190_195_groupi_n_707 ,csa_tree_add_190_195_groupi_n_2418);
  and csa_tree_add_190_195_groupi_g46458(csa_tree_add_190_195_groupi_n_3202 ,csa_tree_add_190_195_groupi_n_1447 ,csa_tree_add_190_195_groupi_n_1404);
  and csa_tree_add_190_195_groupi_g46459(csa_tree_add_190_195_groupi_n_3201 ,csa_tree_add_190_195_groupi_n_2504 ,csa_tree_add_190_195_groupi_n_2732);
  or csa_tree_add_190_195_groupi_g46460(csa_tree_add_190_195_groupi_n_3200 ,csa_tree_add_190_195_groupi_n_1615 ,csa_tree_add_190_195_groupi_n_1809);
  not csa_tree_add_190_195_groupi_g46461(csa_tree_add_190_195_groupi_n_2733 ,in60[0]);
  not csa_tree_add_190_195_groupi_g46462(csa_tree_add_190_195_groupi_n_2732 ,in58[1]);
  not csa_tree_add_190_195_groupi_g46463(csa_tree_add_190_195_groupi_n_2731 ,in57[15]);
  not csa_tree_add_190_195_groupi_g46464(csa_tree_add_190_195_groupi_n_2730 ,in59[9]);
  not csa_tree_add_190_195_groupi_g46465(csa_tree_add_190_195_groupi_n_2729 ,in56[7]);
  not csa_tree_add_190_195_groupi_g46466(csa_tree_add_190_195_groupi_n_2728 ,in59[7]);
  not csa_tree_add_190_195_groupi_g46467(csa_tree_add_190_195_groupi_n_2727 ,in60[9]);
  not csa_tree_add_190_195_groupi_g46468(csa_tree_add_190_195_groupi_n_2726 ,in60[14]);
  not csa_tree_add_190_195_groupi_g46469(csa_tree_add_190_195_groupi_n_2725 ,csa_tree_add_190_195_groupi_n_1572);
  not csa_tree_add_190_195_groupi_g46470(csa_tree_add_190_195_groupi_n_2724 ,in58[10]);
  not csa_tree_add_190_195_groupi_g46471(csa_tree_add_190_195_groupi_n_2723 ,in58[5]);
  not csa_tree_add_190_195_groupi_g46472(csa_tree_add_190_195_groupi_n_2722 ,csa_tree_add_190_195_groupi_n_1543);
  not csa_tree_add_190_195_groupi_g46473(csa_tree_add_190_195_groupi_n_2721 ,in56[11]);
  not csa_tree_add_190_195_groupi_g46474(csa_tree_add_190_195_groupi_n_2720 ,in59[2]);
  not csa_tree_add_190_195_groupi_g46475(csa_tree_add_190_195_groupi_n_2719 ,in59[5]);
  not csa_tree_add_190_195_groupi_g46476(csa_tree_add_190_195_groupi_n_2718 ,csa_tree_add_190_195_groupi_n_1585);
  not csa_tree_add_190_195_groupi_g46479(csa_tree_add_190_195_groupi_n_2717 ,csa_tree_add_190_195_groupi_n_1581);
  not csa_tree_add_190_195_groupi_g46481(csa_tree_add_190_195_groupi_n_2716 ,csa_tree_add_190_195_groupi_n_1609);
  not csa_tree_add_190_195_groupi_g46484(csa_tree_add_190_195_groupi_n_2715 ,csa_tree_add_190_195_groupi_n_1614);
  not csa_tree_add_190_195_groupi_g46488(csa_tree_add_190_195_groupi_n_2714 ,csa_tree_add_190_195_groupi_n_1700);
  not csa_tree_add_190_195_groupi_g46494(csa_tree_add_190_195_groupi_n_2713 ,csa_tree_add_190_195_groupi_n_1664);
  not csa_tree_add_190_195_groupi_g46496(csa_tree_add_190_195_groupi_n_2712 ,csa_tree_add_190_195_groupi_n_1705);
  not csa_tree_add_190_195_groupi_g46497(csa_tree_add_190_195_groupi_n_2711 ,csa_tree_add_190_195_groupi_n_1711);
  not csa_tree_add_190_195_groupi_g46498(csa_tree_add_190_195_groupi_n_2710 ,csa_tree_add_190_195_groupi_n_1598);
  not csa_tree_add_190_195_groupi_g46503(csa_tree_add_190_195_groupi_n_2709 ,csa_tree_add_190_195_groupi_n_1868);
  not csa_tree_add_190_195_groupi_g46504(csa_tree_add_190_195_groupi_n_2708 ,csa_tree_add_190_195_groupi_n_1571);
  not csa_tree_add_190_195_groupi_g46505(csa_tree_add_190_195_groupi_n_2707 ,csa_tree_add_190_195_groupi_n_1951);
  not csa_tree_add_190_195_groupi_g46506(csa_tree_add_190_195_groupi_n_2706 ,csa_tree_add_190_195_groupi_n_1695);
  not csa_tree_add_190_195_groupi_g46507(csa_tree_add_190_195_groupi_n_2705 ,csa_tree_add_190_195_groupi_n_1936);
  not csa_tree_add_190_195_groupi_g46508(csa_tree_add_190_195_groupi_n_2704 ,csa_tree_add_190_195_groupi_n_1830);
  not csa_tree_add_190_195_groupi_g46509(csa_tree_add_190_195_groupi_n_2703 ,csa_tree_add_190_195_groupi_n_1941);
  not csa_tree_add_190_195_groupi_g46510(csa_tree_add_190_195_groupi_n_2702 ,csa_tree_add_190_195_groupi_n_1968);
  not csa_tree_add_190_195_groupi_g46511(csa_tree_add_190_195_groupi_n_2701 ,csa_tree_add_190_195_groupi_n_2087);
  not csa_tree_add_190_195_groupi_g46512(csa_tree_add_190_195_groupi_n_2700 ,csa_tree_add_190_195_groupi_n_1748);
  not csa_tree_add_190_195_groupi_g46513(csa_tree_add_190_195_groupi_n_2699 ,csa_tree_add_190_195_groupi_n_1950);
  not csa_tree_add_190_195_groupi_g46514(csa_tree_add_190_195_groupi_n_2698 ,csa_tree_add_190_195_groupi_n_1674);
  not csa_tree_add_190_195_groupi_g46515(csa_tree_add_190_195_groupi_n_2697 ,csa_tree_add_190_195_groupi_n_1935);
  not csa_tree_add_190_195_groupi_g46516(csa_tree_add_190_195_groupi_n_2696 ,csa_tree_add_190_195_groupi_n_1707);
  not csa_tree_add_190_195_groupi_g46517(csa_tree_add_190_195_groupi_n_2695 ,csa_tree_add_190_195_groupi_n_1702);
  not csa_tree_add_190_195_groupi_g46518(csa_tree_add_190_195_groupi_n_2694 ,csa_tree_add_190_195_groupi_n_1869);
  not csa_tree_add_190_195_groupi_g46519(csa_tree_add_190_195_groupi_n_2693 ,csa_tree_add_190_195_groupi_n_1890);
  not csa_tree_add_190_195_groupi_g46520(csa_tree_add_190_195_groupi_n_2692 ,csa_tree_add_190_195_groupi_n_1971);
  not csa_tree_add_190_195_groupi_g46521(csa_tree_add_190_195_groupi_n_2691 ,csa_tree_add_190_195_groupi_n_1967);
  not csa_tree_add_190_195_groupi_g46522(csa_tree_add_190_195_groupi_n_2690 ,csa_tree_add_190_195_groupi_n_1944);
  not csa_tree_add_190_195_groupi_g46523(csa_tree_add_190_195_groupi_n_2689 ,csa_tree_add_190_195_groupi_n_1841);
  not csa_tree_add_190_195_groupi_g46524(csa_tree_add_190_195_groupi_n_2688 ,csa_tree_add_190_195_groupi_n_1848);
  not csa_tree_add_190_195_groupi_g46525(csa_tree_add_190_195_groupi_n_2687 ,csa_tree_add_190_195_groupi_n_1835);
  not csa_tree_add_190_195_groupi_g46526(csa_tree_add_190_195_groupi_n_2686 ,csa_tree_add_190_195_groupi_n_1832);
  not csa_tree_add_190_195_groupi_g46528(csa_tree_add_190_195_groupi_n_2685 ,csa_tree_add_190_195_groupi_n_1677);
  not csa_tree_add_190_195_groupi_g46529(csa_tree_add_190_195_groupi_n_2684 ,csa_tree_add_190_195_groupi_n_1992);
  not csa_tree_add_190_195_groupi_g46530(csa_tree_add_190_195_groupi_n_2683 ,csa_tree_add_190_195_groupi_n_1866);
  not csa_tree_add_190_195_groupi_g46531(csa_tree_add_190_195_groupi_n_2682 ,csa_tree_add_190_195_groupi_n_1849);
  not csa_tree_add_190_195_groupi_g46532(csa_tree_add_190_195_groupi_n_2681 ,csa_tree_add_190_195_groupi_n_1850);
  not csa_tree_add_190_195_groupi_g46533(csa_tree_add_190_195_groupi_n_2680 ,csa_tree_add_190_195_groupi_n_1862);
  not csa_tree_add_190_195_groupi_g46534(csa_tree_add_190_195_groupi_n_2679 ,csa_tree_add_190_195_groupi_n_1706);
  not csa_tree_add_190_195_groupi_g46535(csa_tree_add_190_195_groupi_n_2678 ,csa_tree_add_190_195_groupi_n_1774);
  not csa_tree_add_190_195_groupi_g46536(csa_tree_add_190_195_groupi_n_2677 ,csa_tree_add_190_195_groupi_n_1825);
  not csa_tree_add_190_195_groupi_g46539(csa_tree_add_190_195_groupi_n_2676 ,csa_tree_add_190_195_groupi_n_1828);
  not csa_tree_add_190_195_groupi_g46540(csa_tree_add_190_195_groupi_n_2675 ,csa_tree_add_190_195_groupi_n_2082);
  not csa_tree_add_190_195_groupi_g46541(csa_tree_add_190_195_groupi_n_2674 ,csa_tree_add_190_195_groupi_n_1817);
  not csa_tree_add_190_195_groupi_g46542(csa_tree_add_190_195_groupi_n_2673 ,csa_tree_add_190_195_groupi_n_1915);
  not csa_tree_add_190_195_groupi_g46543(csa_tree_add_190_195_groupi_n_2672 ,csa_tree_add_190_195_groupi_n_1920);
  not csa_tree_add_190_195_groupi_g46544(csa_tree_add_190_195_groupi_n_2671 ,csa_tree_add_190_195_groupi_n_1909);
  not csa_tree_add_190_195_groupi_g46545(csa_tree_add_190_195_groupi_n_2670 ,csa_tree_add_190_195_groupi_n_2056);
  not csa_tree_add_190_195_groupi_g46546(csa_tree_add_190_195_groupi_n_2669 ,csa_tree_add_190_195_groupi_n_1964);
  not csa_tree_add_190_195_groupi_g46547(csa_tree_add_190_195_groupi_n_2668 ,csa_tree_add_190_195_groupi_n_1827);
  not csa_tree_add_190_195_groupi_g46548(csa_tree_add_190_195_groupi_n_2667 ,csa_tree_add_190_195_groupi_n_1948);
  not csa_tree_add_190_195_groupi_g46549(csa_tree_add_190_195_groupi_n_2666 ,csa_tree_add_190_195_groupi_n_1844);
  not csa_tree_add_190_195_groupi_g46551(csa_tree_add_190_195_groupi_n_2665 ,csa_tree_add_190_195_groupi_n_1932);
  not csa_tree_add_190_195_groupi_g46552(csa_tree_add_190_195_groupi_n_2664 ,csa_tree_add_190_195_groupi_n_1989);
  not csa_tree_add_190_195_groupi_g46553(csa_tree_add_190_195_groupi_n_2663 ,csa_tree_add_190_195_groupi_n_1810);
  not csa_tree_add_190_195_groupi_g46554(csa_tree_add_190_195_groupi_n_2662 ,csa_tree_add_190_195_groupi_n_2006);
  not csa_tree_add_190_195_groupi_g46555(csa_tree_add_190_195_groupi_n_2661 ,csa_tree_add_190_195_groupi_n_1993);
  not csa_tree_add_190_195_groupi_g46557(csa_tree_add_190_195_groupi_n_2660 ,csa_tree_add_190_195_groupi_n_2155);
  not csa_tree_add_190_195_groupi_g46558(csa_tree_add_190_195_groupi_n_2659 ,csa_tree_add_190_195_groupi_n_1836);
  not csa_tree_add_190_195_groupi_g46559(csa_tree_add_190_195_groupi_n_2658 ,csa_tree_add_190_195_groupi_n_1057);
  not csa_tree_add_190_195_groupi_g46560(csa_tree_add_190_195_groupi_n_2657 ,csa_tree_add_190_195_groupi_n_1724);
  not csa_tree_add_190_195_groupi_g46561(csa_tree_add_190_195_groupi_n_2656 ,csa_tree_add_190_195_groupi_n_1839);
  not csa_tree_add_190_195_groupi_g46562(csa_tree_add_190_195_groupi_n_2655 ,csa_tree_add_190_195_groupi_n_2119);
  not csa_tree_add_190_195_groupi_g46563(csa_tree_add_190_195_groupi_n_2654 ,csa_tree_add_190_195_groupi_n_1006);
  not csa_tree_add_190_195_groupi_g46564(csa_tree_add_190_195_groupi_n_2653 ,csa_tree_add_190_195_groupi_n_1969);
  not csa_tree_add_190_195_groupi_g46565(csa_tree_add_190_195_groupi_n_2652 ,csa_tree_add_190_195_groupi_n_1824);
  not csa_tree_add_190_195_groupi_g46566(csa_tree_add_190_195_groupi_n_2651 ,csa_tree_add_190_195_groupi_n_1066);
  not csa_tree_add_190_195_groupi_g46567(csa_tree_add_190_195_groupi_n_2650 ,csa_tree_add_190_195_groupi_n_1864);
  not csa_tree_add_190_195_groupi_g46568(csa_tree_add_190_195_groupi_n_2649 ,csa_tree_add_190_195_groupi_n_1934);
  not csa_tree_add_190_195_groupi_g46569(csa_tree_add_190_195_groupi_n_2648 ,csa_tree_add_190_195_groupi_n_1846);
  not csa_tree_add_190_195_groupi_g46570(csa_tree_add_190_195_groupi_n_2647 ,csa_tree_add_190_195_groupi_n_1745);
  not csa_tree_add_190_195_groupi_g46571(csa_tree_add_190_195_groupi_n_2646 ,csa_tree_add_190_195_groupi_n_1691);
  not csa_tree_add_190_195_groupi_g46572(csa_tree_add_190_195_groupi_n_2645 ,csa_tree_add_190_195_groupi_n_2051);
  not csa_tree_add_190_195_groupi_g46573(csa_tree_add_190_195_groupi_n_2644 ,csa_tree_add_190_195_groupi_n_1638);
  not csa_tree_add_190_195_groupi_g46574(csa_tree_add_190_195_groupi_n_2643 ,csa_tree_add_190_195_groupi_n_1831);
  not csa_tree_add_190_195_groupi_g46575(csa_tree_add_190_195_groupi_n_2642 ,csa_tree_add_190_195_groupi_n_1995);
  not csa_tree_add_190_195_groupi_g46576(csa_tree_add_190_195_groupi_n_2641 ,csa_tree_add_190_195_groupi_n_1782);
  not csa_tree_add_190_195_groupi_g46577(csa_tree_add_190_195_groupi_n_2640 ,csa_tree_add_190_195_groupi_n_2086);
  not csa_tree_add_190_195_groupi_g46578(csa_tree_add_190_195_groupi_n_2639 ,csa_tree_add_190_195_groupi_n_1688);
  not csa_tree_add_190_195_groupi_g46579(csa_tree_add_190_195_groupi_n_2638 ,csa_tree_add_190_195_groupi_n_2039);
  not csa_tree_add_190_195_groupi_g46580(csa_tree_add_190_195_groupi_n_2637 ,csa_tree_add_190_195_groupi_n_1708);
  not csa_tree_add_190_195_groupi_g46581(csa_tree_add_190_195_groupi_n_2636 ,csa_tree_add_190_195_groupi_n_779);
  not csa_tree_add_190_195_groupi_g46582(csa_tree_add_190_195_groupi_n_2635 ,csa_tree_add_190_195_groupi_n_1974);
  not csa_tree_add_190_195_groupi_g46583(csa_tree_add_190_195_groupi_n_2634 ,csa_tree_add_190_195_groupi_n_1838);
  not csa_tree_add_190_195_groupi_g46584(csa_tree_add_190_195_groupi_n_2633 ,csa_tree_add_190_195_groupi_n_2211);
  not csa_tree_add_190_195_groupi_g46585(csa_tree_add_190_195_groupi_n_2632 ,csa_tree_add_190_195_groupi_n_1000);
  not csa_tree_add_190_195_groupi_g46586(csa_tree_add_190_195_groupi_n_2631 ,csa_tree_add_190_195_groupi_n_1996);
  not csa_tree_add_190_195_groupi_g46587(csa_tree_add_190_195_groupi_n_2630 ,csa_tree_add_190_195_groupi_n_1877);
  not csa_tree_add_190_195_groupi_g46588(csa_tree_add_190_195_groupi_n_2629 ,csa_tree_add_190_195_groupi_n_1096);
  not csa_tree_add_190_195_groupi_g46589(csa_tree_add_190_195_groupi_n_2628 ,csa_tree_add_190_195_groupi_n_812);
  not csa_tree_add_190_195_groupi_g46590(csa_tree_add_190_195_groupi_n_2627 ,csa_tree_add_190_195_groupi_n_2041);
  not csa_tree_add_190_195_groupi_g46591(csa_tree_add_190_195_groupi_n_2626 ,csa_tree_add_190_195_groupi_n_1921);
  not csa_tree_add_190_195_groupi_g46592(csa_tree_add_190_195_groupi_n_2625 ,csa_tree_add_190_195_groupi_n_1105);
  not csa_tree_add_190_195_groupi_g46593(csa_tree_add_190_195_groupi_n_2624 ,csa_tree_add_190_195_groupi_n_1923);
  not csa_tree_add_190_195_groupi_g46594(csa_tree_add_190_195_groupi_n_2623 ,csa_tree_add_190_195_groupi_n_2057);
  not csa_tree_add_190_195_groupi_g46595(csa_tree_add_190_195_groupi_n_2622 ,csa_tree_add_190_195_groupi_n_2049);
  not csa_tree_add_190_195_groupi_g46596(csa_tree_add_190_195_groupi_n_2621 ,csa_tree_add_190_195_groupi_n_1090);
  not csa_tree_add_190_195_groupi_g46597(csa_tree_add_190_195_groupi_n_2620 ,csa_tree_add_190_195_groupi_n_2062);
  not csa_tree_add_190_195_groupi_g46598(csa_tree_add_190_195_groupi_n_2619 ,csa_tree_add_190_195_groupi_n_1162);
  not csa_tree_add_190_195_groupi_g46599(csa_tree_add_190_195_groupi_n_2618 ,csa_tree_add_190_195_groupi_n_936);
  not csa_tree_add_190_195_groupi_g46600(csa_tree_add_190_195_groupi_n_2617 ,csa_tree_add_190_195_groupi_n_1726);
  not csa_tree_add_190_195_groupi_g46601(csa_tree_add_190_195_groupi_n_2616 ,csa_tree_add_190_195_groupi_n_1930);
  not csa_tree_add_190_195_groupi_g46602(csa_tree_add_190_195_groupi_n_2615 ,csa_tree_add_190_195_groupi_n_2061);
  not csa_tree_add_190_195_groupi_g46603(csa_tree_add_190_195_groupi_n_2614 ,csa_tree_add_190_195_groupi_n_820);
  not csa_tree_add_190_195_groupi_g46604(csa_tree_add_190_195_groupi_n_2613 ,csa_tree_add_190_195_groupi_n_804);
  not csa_tree_add_190_195_groupi_g46606(csa_tree_add_190_195_groupi_n_2612 ,csa_tree_add_190_195_groupi_n_2158);
  not csa_tree_add_190_195_groupi_g46607(csa_tree_add_190_195_groupi_n_2611 ,csa_tree_add_190_195_groupi_n_2060);
  not csa_tree_add_190_195_groupi_g46608(csa_tree_add_190_195_groupi_n_2610 ,csa_tree_add_190_195_groupi_n_1975);
  not csa_tree_add_190_195_groupi_g46609(csa_tree_add_190_195_groupi_n_2609 ,csa_tree_add_190_195_groupi_n_931);
  not csa_tree_add_190_195_groupi_g46610(csa_tree_add_190_195_groupi_n_2608 ,csa_tree_add_190_195_groupi_n_1977);
  not csa_tree_add_190_195_groupi_g46611(csa_tree_add_190_195_groupi_n_2607 ,csa_tree_add_190_195_groupi_n_1171);
  not csa_tree_add_190_195_groupi_g46612(csa_tree_add_190_195_groupi_n_2606 ,csa_tree_add_190_195_groupi_n_748);
  not csa_tree_add_190_195_groupi_g46613(csa_tree_add_190_195_groupi_n_2605 ,csa_tree_add_190_195_groupi_n_1962);
  not csa_tree_add_190_195_groupi_g46614(csa_tree_add_190_195_groupi_n_2604 ,csa_tree_add_190_195_groupi_n_2152);
  not csa_tree_add_190_195_groupi_g46615(csa_tree_add_190_195_groupi_n_2603 ,csa_tree_add_190_195_groupi_n_1084);
  not csa_tree_add_190_195_groupi_g46616(csa_tree_add_190_195_groupi_n_2602 ,csa_tree_add_190_195_groupi_n_1029);
  not csa_tree_add_190_195_groupi_g46617(csa_tree_add_190_195_groupi_n_2601 ,csa_tree_add_190_195_groupi_n_871);
  not csa_tree_add_190_195_groupi_g46618(csa_tree_add_190_195_groupi_n_2600 ,in55[10]);
  not csa_tree_add_190_195_groupi_g46619(csa_tree_add_190_195_groupi_n_2599 ,in55[13]);
  not csa_tree_add_190_195_groupi_g46620(csa_tree_add_190_195_groupi_n_2598 ,csa_tree_add_190_195_groupi_n_796);
  not csa_tree_add_190_195_groupi_g46621(csa_tree_add_190_195_groupi_n_2597 ,csa_tree_add_190_195_groupi_n_1132);
  not csa_tree_add_190_195_groupi_g46622(csa_tree_add_190_195_groupi_n_2596 ,in55[1]);
  not csa_tree_add_190_195_groupi_g46623(csa_tree_add_190_195_groupi_n_2595 ,in55[12]);
  not csa_tree_add_190_195_groupi_g46624(csa_tree_add_190_195_groupi_n_2594 ,csa_tree_add_190_195_groupi_n_2090);
  not csa_tree_add_190_195_groupi_g46625(csa_tree_add_190_195_groupi_n_2593 ,in55[8]);
  not csa_tree_add_190_195_groupi_g46626(csa_tree_add_190_195_groupi_n_2592 ,in55[5]);
  not csa_tree_add_190_195_groupi_g46627(csa_tree_add_190_195_groupi_n_2591 ,in55[14]);
  not csa_tree_add_190_195_groupi_g46628(csa_tree_add_190_195_groupi_n_2590 ,in55[2]);
  not csa_tree_add_190_195_groupi_g46629(csa_tree_add_190_195_groupi_n_2589 ,in55[0]);
  not csa_tree_add_190_195_groupi_g46630(csa_tree_add_190_195_groupi_n_2588 ,csa_tree_add_190_195_groupi_n_874);
  not csa_tree_add_190_195_groupi_g46631(csa_tree_add_190_195_groupi_n_2587 ,csa_tree_add_190_195_groupi_n_1285);
  not csa_tree_add_190_195_groupi_g46633(csa_tree_add_190_195_groupi_n_2586 ,csa_tree_add_190_195_groupi_n_1078);
  not csa_tree_add_190_195_groupi_g46634(csa_tree_add_190_195_groupi_n_2585 ,csa_tree_add_190_195_groupi_n_457);
  not csa_tree_add_190_195_groupi_g46640(csa_tree_add_190_195_groupi_n_2584 ,csa_tree_add_190_195_groupi_n_1295);
  not csa_tree_add_190_195_groupi_g46641(csa_tree_add_190_195_groupi_n_2583 ,csa_tree_add_190_195_groupi_n_305);
  not csa_tree_add_190_195_groupi_g46643(csa_tree_add_190_195_groupi_n_2582 ,csa_tree_add_190_195_groupi_n_446);
  not csa_tree_add_190_195_groupi_g46644(csa_tree_add_190_195_groupi_n_2581 ,csa_tree_add_190_195_groupi_n_394);
  not csa_tree_add_190_195_groupi_g46646(csa_tree_add_190_195_groupi_n_2580 ,csa_tree_add_190_195_groupi_n_482);
  not csa_tree_add_190_195_groupi_g46647(csa_tree_add_190_195_groupi_n_2579 ,csa_tree_add_190_195_groupi_n_1208);
  not csa_tree_add_190_195_groupi_g46649(csa_tree_add_190_195_groupi_n_2578 ,csa_tree_add_190_195_groupi_n_426);
  not csa_tree_add_190_195_groupi_g46650(csa_tree_add_190_195_groupi_n_2577 ,csa_tree_add_190_195_groupi_n_435);
  not csa_tree_add_190_195_groupi_g46652(csa_tree_add_190_195_groupi_n_2576 ,csa_tree_add_190_195_groupi_n_1216);
  not csa_tree_add_190_195_groupi_g46653(csa_tree_add_190_195_groupi_n_2575 ,csa_tree_add_190_195_groupi_n_469);
  not csa_tree_add_190_195_groupi_g46654(csa_tree_add_190_195_groupi_n_2574 ,csa_tree_add_190_195_groupi_n_429);
  not csa_tree_add_190_195_groupi_g46655(csa_tree_add_190_195_groupi_n_2573 ,csa_tree_add_190_195_groupi_n_595);
  not csa_tree_add_190_195_groupi_g46656(csa_tree_add_190_195_groupi_n_2572 ,in57[14]);
  not csa_tree_add_190_195_groupi_g46657(csa_tree_add_190_195_groupi_n_2571 ,in60[3]);
  not csa_tree_add_190_195_groupi_g46658(csa_tree_add_190_195_groupi_n_2570 ,in59[1]);
  not csa_tree_add_190_195_groupi_g46659(csa_tree_add_190_195_groupi_n_2569 ,in60[1]);
  not csa_tree_add_190_195_groupi_g46660(csa_tree_add_190_195_groupi_n_2568 ,in57[12]);
  not csa_tree_add_190_195_groupi_g46661(csa_tree_add_190_195_groupi_n_2567 ,in61[7]);
  not csa_tree_add_190_195_groupi_g46662(csa_tree_add_190_195_groupi_n_2566 ,in56[15]);
  not csa_tree_add_190_195_groupi_g46663(csa_tree_add_190_195_groupi_n_2565 ,in59[10]);
  not csa_tree_add_190_195_groupi_g46664(csa_tree_add_190_195_groupi_n_2564 ,in61[5]);
  not csa_tree_add_190_195_groupi_g46665(csa_tree_add_190_195_groupi_n_2563 ,in56[10]);
  not csa_tree_add_190_195_groupi_g46666(csa_tree_add_190_195_groupi_n_2562 ,csa_tree_add_190_195_groupi_n_1550);
  not csa_tree_add_190_195_groupi_g46667(csa_tree_add_190_195_groupi_n_2561 ,in61[13]);
  not csa_tree_add_190_195_groupi_g46668(csa_tree_add_190_195_groupi_n_2560 ,in58[7]);
  not csa_tree_add_190_195_groupi_g46669(csa_tree_add_190_195_groupi_n_2559 ,in61[1]);
  not csa_tree_add_190_195_groupi_g46670(csa_tree_add_190_195_groupi_n_2558 ,in58[0]);
  not csa_tree_add_190_195_groupi_g46671(csa_tree_add_190_195_groupi_n_2557 ,in58[9]);
  not csa_tree_add_190_195_groupi_g46672(csa_tree_add_190_195_groupi_n_2556 ,in56[9]);
  not csa_tree_add_190_195_groupi_g46673(csa_tree_add_190_195_groupi_n_2555 ,in56[0]);
  not csa_tree_add_190_195_groupi_g46674(csa_tree_add_190_195_groupi_n_2554 ,in61[2]);
  not csa_tree_add_190_195_groupi_g46675(csa_tree_add_190_195_groupi_n_2553 ,in60[11]);
  not csa_tree_add_190_195_groupi_g46676(csa_tree_add_190_195_groupi_n_2552 ,in60[6]);
  not csa_tree_add_190_195_groupi_g46677(csa_tree_add_190_195_groupi_n_2551 ,csa_tree_add_190_195_groupi_n_1842);
  not csa_tree_add_190_195_groupi_g46678(csa_tree_add_190_195_groupi_n_2550 ,csa_tree_add_190_195_groupi_n_1687);
  not csa_tree_add_190_195_groupi_g46679(csa_tree_add_190_195_groupi_n_2549 ,csa_tree_add_190_195_groupi_n_1586);
  not csa_tree_add_190_195_groupi_g46682(csa_tree_add_190_195_groupi_n_2548 ,csa_tree_add_190_195_groupi_n_1620);
  not csa_tree_add_190_195_groupi_g46683(csa_tree_add_190_195_groupi_n_2547 ,csa_tree_add_190_195_groupi_n_1595);
  not csa_tree_add_190_195_groupi_g46684(csa_tree_add_190_195_groupi_n_2546 ,csa_tree_add_190_195_groupi_n_1694);
  not csa_tree_add_190_195_groupi_g46685(csa_tree_add_190_195_groupi_n_2545 ,csa_tree_add_190_195_groupi_n_1679);
  not csa_tree_add_190_195_groupi_g46687(csa_tree_add_190_195_groupi_n_2544 ,csa_tree_add_190_195_groupi_n_1760);
  not csa_tree_add_190_195_groupi_g46688(csa_tree_add_190_195_groupi_n_2543 ,csa_tree_add_190_195_groupi_n_1761);
  not csa_tree_add_190_195_groupi_g46689(csa_tree_add_190_195_groupi_n_2542 ,csa_tree_add_190_195_groupi_n_1758);
  not csa_tree_add_190_195_groupi_g46694(csa_tree_add_190_195_groupi_n_2541 ,csa_tree_add_190_195_groupi_n_1678);
  not csa_tree_add_190_195_groupi_g46700(csa_tree_add_190_195_groupi_n_2540 ,csa_tree_add_190_195_groupi_n_1966);
  not csa_tree_add_190_195_groupi_g46702(csa_tree_add_190_195_groupi_n_2539 ,csa_tree_add_190_195_groupi_n_1906);
  not csa_tree_add_190_195_groupi_g46703(csa_tree_add_190_195_groupi_n_2538 ,csa_tree_add_190_195_groupi_n_1819);
  not csa_tree_add_190_195_groupi_g46704(csa_tree_add_190_195_groupi_n_2537 ,csa_tree_add_190_195_groupi_n_1863);
  not csa_tree_add_190_195_groupi_g46705(csa_tree_add_190_195_groupi_n_2536 ,csa_tree_add_190_195_groupi_n_1604);
  not csa_tree_add_190_195_groupi_g46706(csa_tree_add_190_195_groupi_n_2535 ,csa_tree_add_190_195_groupi_n_1903);
  not csa_tree_add_190_195_groupi_g46707(csa_tree_add_190_195_groupi_n_2534 ,csa_tree_add_190_195_groupi_n_1607);
  not csa_tree_add_190_195_groupi_g46708(csa_tree_add_190_195_groupi_n_2533 ,csa_tree_add_190_195_groupi_n_1751);
  not csa_tree_add_190_195_groupi_g46709(csa_tree_add_190_195_groupi_n_2532 ,csa_tree_add_190_195_groupi_n_1945);
  not csa_tree_add_190_195_groupi_g46710(csa_tree_add_190_195_groupi_n_2531 ,csa_tree_add_190_195_groupi_n_1860);
  not csa_tree_add_190_195_groupi_g46711(csa_tree_add_190_195_groupi_n_2530 ,csa_tree_add_190_195_groupi_n_1823);
  not csa_tree_add_190_195_groupi_g46712(csa_tree_add_190_195_groupi_n_2529 ,csa_tree_add_190_195_groupi_n_2007);
  not csa_tree_add_190_195_groupi_g46713(csa_tree_add_190_195_groupi_n_2528 ,csa_tree_add_190_195_groupi_n_1818);
  not csa_tree_add_190_195_groupi_g46714(csa_tree_add_190_195_groupi_n_2527 ,csa_tree_add_190_195_groupi_n_1812);
  not csa_tree_add_190_195_groupi_g46715(csa_tree_add_190_195_groupi_n_2526 ,csa_tree_add_190_195_groupi_n_1763);
  not csa_tree_add_190_195_groupi_g46717(csa_tree_add_190_195_groupi_n_2525 ,csa_tree_add_190_195_groupi_n_1668);
  not csa_tree_add_190_195_groupi_g46718(csa_tree_add_190_195_groupi_n_2524 ,csa_tree_add_190_195_groupi_n_1780);
  not csa_tree_add_190_195_groupi_g46719(csa_tree_add_190_195_groupi_n_2523 ,csa_tree_add_190_195_groupi_n_1991);
  not csa_tree_add_190_195_groupi_g46720(csa_tree_add_190_195_groupi_n_2522 ,csa_tree_add_190_195_groupi_n_1855);
  not csa_tree_add_190_195_groupi_g46721(csa_tree_add_190_195_groupi_n_2521 ,csa_tree_add_190_195_groupi_n_1865);
  not csa_tree_add_190_195_groupi_g46722(csa_tree_add_190_195_groupi_n_2520 ,csa_tree_add_190_195_groupi_n_2084);
  not csa_tree_add_190_195_groupi_g46723(csa_tree_add_190_195_groupi_n_2519 ,csa_tree_add_190_195_groupi_n_1910);
  not csa_tree_add_190_195_groupi_g46724(csa_tree_add_190_195_groupi_n_2518 ,csa_tree_add_190_195_groupi_n_1851);
  not csa_tree_add_190_195_groupi_g46725(csa_tree_add_190_195_groupi_n_2517 ,csa_tree_add_190_195_groupi_n_2089);
  not csa_tree_add_190_195_groupi_g46726(csa_tree_add_190_195_groupi_n_2516 ,csa_tree_add_190_195_groupi_n_1808);
  not csa_tree_add_190_195_groupi_g46727(csa_tree_add_190_195_groupi_n_2515 ,csa_tree_add_190_195_groupi_n_1990);
  not csa_tree_add_190_195_groupi_g46728(csa_tree_add_190_195_groupi_n_2514 ,csa_tree_add_190_195_groupi_n_1972);
  not csa_tree_add_190_195_groupi_g46729(csa_tree_add_190_195_groupi_n_2513 ,csa_tree_add_190_195_groupi_n_1987);
  not csa_tree_add_190_195_groupi_g46730(csa_tree_add_190_195_groupi_n_2512 ,csa_tree_add_190_195_groupi_n_1826);
  not csa_tree_add_190_195_groupi_g46733(csa_tree_add_190_195_groupi_n_2511 ,csa_tree_add_190_195_groupi_n_810);
  not csa_tree_add_190_195_groupi_g46734(csa_tree_add_190_195_groupi_n_2510 ,csa_tree_add_190_195_groupi_n_2058);
  not csa_tree_add_190_195_groupi_g46735(csa_tree_add_190_195_groupi_n_2509 ,csa_tree_add_190_195_groupi_n_1929);
  not csa_tree_add_190_195_groupi_g46736(csa_tree_add_190_195_groupi_n_2508 ,csa_tree_add_190_195_groupi_n_1809);
  not csa_tree_add_190_195_groupi_g46737(csa_tree_add_190_195_groupi_n_2507 ,csa_tree_add_190_195_groupi_n_1905);
  not csa_tree_add_190_195_groupi_g46738(csa_tree_add_190_195_groupi_n_2506 ,csa_tree_add_190_195_groupi_n_2091);
  not csa_tree_add_190_195_groupi_g46739(csa_tree_add_190_195_groupi_n_2505 ,csa_tree_add_190_195_groupi_n_1715);
  not csa_tree_add_190_195_groupi_g46740(csa_tree_add_190_195_groupi_n_2504 ,csa_tree_add_190_195_groupi_n_934);
  not csa_tree_add_190_195_groupi_g46742(csa_tree_add_190_195_groupi_n_2503 ,csa_tree_add_190_195_groupi_n_1775);
  not csa_tree_add_190_195_groupi_g46743(csa_tree_add_190_195_groupi_n_2502 ,csa_tree_add_190_195_groupi_n_2216);
  not csa_tree_add_190_195_groupi_g46744(csa_tree_add_190_195_groupi_n_2501 ,csa_tree_add_190_195_groupi_n_2156);
  not csa_tree_add_190_195_groupi_g46745(csa_tree_add_190_195_groupi_n_2500 ,csa_tree_add_190_195_groupi_n_2050);
  not csa_tree_add_190_195_groupi_g46746(csa_tree_add_190_195_groupi_n_2499 ,csa_tree_add_190_195_groupi_n_1806);
  not csa_tree_add_190_195_groupi_g46747(csa_tree_add_190_195_groupi_n_2498 ,csa_tree_add_190_195_groupi_n_792);
  not csa_tree_add_190_195_groupi_g46748(csa_tree_add_190_195_groupi_n_2497 ,csa_tree_add_190_195_groupi_n_1994);
  not csa_tree_add_190_195_groupi_g46749(csa_tree_add_190_195_groupi_n_2496 ,csa_tree_add_190_195_groupi_n_2117);
  not csa_tree_add_190_195_groupi_g46750(csa_tree_add_190_195_groupi_n_2495 ,csa_tree_add_190_195_groupi_n_1820);
  not csa_tree_add_190_195_groupi_g46751(csa_tree_add_190_195_groupi_n_2494 ,csa_tree_add_190_195_groupi_n_1141);
  not csa_tree_add_190_195_groupi_g46752(csa_tree_add_190_195_groupi_n_2493 ,csa_tree_add_190_195_groupi_n_773);
  not csa_tree_add_190_195_groupi_g46753(csa_tree_add_190_195_groupi_n_2492 ,csa_tree_add_190_195_groupi_n_2016);
  not csa_tree_add_190_195_groupi_g46754(csa_tree_add_190_195_groupi_n_2491 ,csa_tree_add_190_195_groupi_n_1042);
  not csa_tree_add_190_195_groupi_g46755(csa_tree_add_190_195_groupi_n_2490 ,csa_tree_add_190_195_groupi_n_1798);
  not csa_tree_add_190_195_groupi_g46756(csa_tree_add_190_195_groupi_n_2489 ,csa_tree_add_190_195_groupi_n_1924);
  not csa_tree_add_190_195_groupi_g46757(csa_tree_add_190_195_groupi_n_2488 ,csa_tree_add_190_195_groupi_n_1893);
  not csa_tree_add_190_195_groupi_g46758(csa_tree_add_190_195_groupi_n_2487 ,csa_tree_add_190_195_groupi_n_2053);
  not csa_tree_add_190_195_groupi_g46759(csa_tree_add_190_195_groupi_n_2486 ,csa_tree_add_190_195_groupi_n_2042);
  not csa_tree_add_190_195_groupi_g46760(csa_tree_add_190_195_groupi_n_2485 ,csa_tree_add_190_195_groupi_n_1843);
  not csa_tree_add_190_195_groupi_g46761(csa_tree_add_190_195_groupi_n_2484 ,csa_tree_add_190_195_groupi_n_984);
  not csa_tree_add_190_195_groupi_g46762(csa_tree_add_190_195_groupi_n_2483 ,csa_tree_add_190_195_groupi_n_847);
  not csa_tree_add_190_195_groupi_g46763(csa_tree_add_190_195_groupi_n_2482 ,csa_tree_add_190_195_groupi_n_969);
  not csa_tree_add_190_195_groupi_g46764(csa_tree_add_190_195_groupi_n_2481 ,csa_tree_add_190_195_groupi_n_2118);
  not csa_tree_add_190_195_groupi_g46765(csa_tree_add_190_195_groupi_n_2480 ,csa_tree_add_190_195_groupi_n_858);
  not csa_tree_add_190_195_groupi_g46766(csa_tree_add_190_195_groupi_n_2479 ,csa_tree_add_190_195_groupi_n_868);
  not csa_tree_add_190_195_groupi_g46768(csa_tree_add_190_195_groupi_n_2478 ,csa_tree_add_190_195_groupi_n_1931);
  not csa_tree_add_190_195_groupi_g46769(csa_tree_add_190_195_groupi_n_2477 ,csa_tree_add_190_195_groupi_n_817);
  not csa_tree_add_190_195_groupi_g46770(csa_tree_add_190_195_groupi_n_2476 ,csa_tree_add_190_195_groupi_n_1960);
  not csa_tree_add_190_195_groupi_g46771(csa_tree_add_190_195_groupi_n_2475 ,csa_tree_add_190_195_groupi_n_742);
  not csa_tree_add_190_195_groupi_g46772(csa_tree_add_190_195_groupi_n_2474 ,csa_tree_add_190_195_groupi_n_1189);
  not csa_tree_add_190_195_groupi_g46773(csa_tree_add_190_195_groupi_n_2473 ,csa_tree_add_190_195_groupi_n_2083);
  not csa_tree_add_190_195_groupi_g46774(csa_tree_add_190_195_groupi_n_2472 ,csa_tree_add_190_195_groupi_n_1020);
  not csa_tree_add_190_195_groupi_g46775(csa_tree_add_190_195_groupi_n_2471 ,csa_tree_add_190_195_groupi_n_2154);
  not csa_tree_add_190_195_groupi_g46776(csa_tree_add_190_195_groupi_n_2470 ,csa_tree_add_190_195_groupi_n_1012);
  not csa_tree_add_190_195_groupi_g46777(csa_tree_add_190_195_groupi_n_2469 ,csa_tree_add_190_195_groupi_n_892);
  not csa_tree_add_190_195_groupi_g46778(csa_tree_add_190_195_groupi_n_2468 ,csa_tree_add_190_195_groupi_n_1978);
  not csa_tree_add_190_195_groupi_g46779(csa_tree_add_190_195_groupi_n_2467 ,csa_tree_add_190_195_groupi_n_1117);
  not csa_tree_add_190_195_groupi_g46780(csa_tree_add_190_195_groupi_n_2466 ,csa_tree_add_190_195_groupi_n_1110);
  not csa_tree_add_190_195_groupi_g46781(csa_tree_add_190_195_groupi_n_2465 ,csa_tree_add_190_195_groupi_n_1075);
  not csa_tree_add_190_195_groupi_g46782(csa_tree_add_190_195_groupi_n_2464 ,csa_tree_add_190_195_groupi_n_916);
  not csa_tree_add_190_195_groupi_g46783(csa_tree_add_190_195_groupi_n_2463 ,csa_tree_add_190_195_groupi_n_1973);
  not csa_tree_add_190_195_groupi_g46784(csa_tree_add_190_195_groupi_n_2462 ,csa_tree_add_190_195_groupi_n_1961);
  not csa_tree_add_190_195_groupi_g46785(csa_tree_add_190_195_groupi_n_2461 ,csa_tree_add_190_195_groupi_n_955);
  not csa_tree_add_190_195_groupi_g46786(csa_tree_add_190_195_groupi_n_2460 ,csa_tree_add_190_195_groupi_n_1988);
  not csa_tree_add_190_195_groupi_g46787(csa_tree_add_190_195_groupi_n_2459 ,csa_tree_add_190_195_groupi_n_2040);
  not csa_tree_add_190_195_groupi_g46788(csa_tree_add_190_195_groupi_n_2458 ,csa_tree_add_190_195_groupi_n_1922);
  not csa_tree_add_190_195_groupi_g46789(csa_tree_add_190_195_groupi_n_2457 ,csa_tree_add_190_195_groupi_n_2214);
  not csa_tree_add_190_195_groupi_g46790(csa_tree_add_190_195_groupi_n_2456 ,csa_tree_add_190_195_groupi_n_1150);
  not csa_tree_add_190_195_groupi_g46791(csa_tree_add_190_195_groupi_n_2455 ,csa_tree_add_190_195_groupi_n_2063);
  not csa_tree_add_190_195_groupi_g46792(csa_tree_add_190_195_groupi_n_2454 ,csa_tree_add_190_195_groupi_n_1928);
  not csa_tree_add_190_195_groupi_g46793(csa_tree_add_190_195_groupi_n_2453 ,csa_tree_add_190_195_groupi_n_1750);
  not csa_tree_add_190_195_groupi_g46794(csa_tree_add_190_195_groupi_n_2452 ,csa_tree_add_190_195_groupi_n_913);
  not csa_tree_add_190_195_groupi_g46795(csa_tree_add_190_195_groupi_n_2451 ,csa_tree_add_190_195_groupi_n_1976);
  not csa_tree_add_190_195_groupi_g46796(csa_tree_add_190_195_groupi_n_2450 ,csa_tree_add_190_195_groupi_n_2209);
  not csa_tree_add_190_195_groupi_g46797(csa_tree_add_190_195_groupi_n_2449 ,csa_tree_add_190_195_groupi_n_835);
  not csa_tree_add_190_195_groupi_g46798(csa_tree_add_190_195_groupi_n_2448 ,csa_tree_add_190_195_groupi_n_2055);
  not csa_tree_add_190_195_groupi_g46799(csa_tree_add_190_195_groupi_n_2447 ,csa_tree_add_190_195_groupi_n_2213);
  not csa_tree_add_190_195_groupi_g46800(csa_tree_add_190_195_groupi_n_2446 ,csa_tree_add_190_195_groupi_n_841);
  not csa_tree_add_190_195_groupi_g46801(csa_tree_add_190_195_groupi_n_2445 ,csa_tree_add_190_195_groupi_n_1087);
  not csa_tree_add_190_195_groupi_g46802(csa_tree_add_190_195_groupi_n_2444 ,csa_tree_add_190_195_groupi_n_958);
  not csa_tree_add_190_195_groupi_g46803(csa_tree_add_190_195_groupi_n_2443 ,csa_tree_add_190_195_groupi_n_2210);
  not csa_tree_add_190_195_groupi_g46804(csa_tree_add_190_195_groupi_n_2442 ,csa_tree_add_190_195_groupi_n_964);
  not csa_tree_add_190_195_groupi_g46805(csa_tree_add_190_195_groupi_n_2441 ,csa_tree_add_190_195_groupi_n_2153);
  not csa_tree_add_190_195_groupi_g46806(csa_tree_add_190_195_groupi_n_2440 ,csa_tree_add_190_195_groupi_n_1051);
  not csa_tree_add_190_195_groupi_g46807(csa_tree_add_190_195_groupi_n_2439 ,csa_tree_add_190_195_groupi_n_2054);
  not csa_tree_add_190_195_groupi_g46808(csa_tree_add_190_195_groupi_n_2438 ,csa_tree_add_190_195_groupi_n_1062);
  not csa_tree_add_190_195_groupi_g46809(csa_tree_add_190_195_groupi_n_2437 ,csa_tree_add_190_195_groupi_n_1965);
  not csa_tree_add_190_195_groupi_g46810(csa_tree_add_190_195_groupi_n_2436 ,csa_tree_add_190_195_groupi_n_880);
  not csa_tree_add_190_195_groupi_g46811(csa_tree_add_190_195_groupi_n_2435 ,csa_tree_add_190_195_groupi_n_1999);
  not csa_tree_add_190_195_groupi_g46812(csa_tree_add_190_195_groupi_n_2434 ,in55[3]);
  not csa_tree_add_190_195_groupi_g46813(csa_tree_add_190_195_groupi_n_2433 ,csa_tree_add_190_195_groupi_n_925);
  not csa_tree_add_190_195_groupi_g46814(csa_tree_add_190_195_groupi_n_2432 ,csa_tree_add_190_195_groupi_n_1904);
  not csa_tree_add_190_195_groupi_g46815(csa_tree_add_190_195_groupi_n_2431 ,in55[4]);
  not csa_tree_add_190_195_groupi_g46816(csa_tree_add_190_195_groupi_n_2430 ,in55[9]);
  not csa_tree_add_190_195_groupi_g46817(csa_tree_add_190_195_groupi_n_2429 ,csa_tree_add_190_195_groupi_n_961);
  not csa_tree_add_190_195_groupi_g46818(csa_tree_add_190_195_groupi_n_2428 ,in55[6]);
  not csa_tree_add_190_195_groupi_g46819(csa_tree_add_190_195_groupi_n_2427 ,csa_tree_add_190_195_groupi_n_838);
  not csa_tree_add_190_195_groupi_g46820(csa_tree_add_190_195_groupi_n_2426 ,csa_tree_add_190_195_groupi_n_1845);
  not csa_tree_add_190_195_groupi_g46821(csa_tree_add_190_195_groupi_n_2425 ,in55[7]);
  not csa_tree_add_190_195_groupi_g46822(csa_tree_add_190_195_groupi_n_2424 ,in55[15]);
  not csa_tree_add_190_195_groupi_g46823(csa_tree_add_190_195_groupi_n_2423 ,in55[11]);
  not csa_tree_add_190_195_groupi_g46824(csa_tree_add_190_195_groupi_n_2422 ,csa_tree_add_190_195_groupi_n_1072);
  not csa_tree_add_190_195_groupi_g46826(csa_tree_add_190_195_groupi_n_2421 ,csa_tree_add_190_195_groupi_n_253);
  not csa_tree_add_190_195_groupi_g46829(csa_tree_add_190_195_groupi_n_2420 ,csa_tree_add_190_195_groupi_n_1204);
  not csa_tree_add_190_195_groupi_g46831(csa_tree_add_190_195_groupi_n_2419 ,csa_tree_add_190_195_groupi_n_1238);
  not csa_tree_add_190_195_groupi_g46833(csa_tree_add_190_195_groupi_n_2418 ,csa_tree_add_190_195_groupi_n_443);
  not csa_tree_add_190_195_groupi_g46835(csa_tree_add_190_195_groupi_n_2417 ,csa_tree_add_190_195_groupi_n_1307);
  not csa_tree_add_190_195_groupi_g46836(csa_tree_add_190_195_groupi_n_2416 ,csa_tree_add_190_195_groupi_n_1291);
  not csa_tree_add_190_195_groupi_g46838(csa_tree_add_190_195_groupi_n_2415 ,csa_tree_add_190_195_groupi_n_1247);
  not csa_tree_add_190_195_groupi_g46839(csa_tree_add_190_195_groupi_n_2414 ,csa_tree_add_190_195_groupi_n_431);
  not csa_tree_add_190_195_groupi_g46840(csa_tree_add_190_195_groupi_n_2413 ,csa_tree_add_190_195_groupi_n_463);
  not csa_tree_add_190_195_groupi_g46842(csa_tree_add_190_195_groupi_n_2412 ,csa_tree_add_190_195_groupi_n_451);
  not csa_tree_add_190_195_groupi_g46844(csa_tree_add_190_195_groupi_n_2411 ,csa_tree_add_190_195_groupi_n_852);
  not csa_tree_add_190_195_groupi_g46845(csa_tree_add_190_195_groupi_n_2410 ,csa_tree_add_190_195_groupi_n_1158);
  not csa_tree_add_190_195_groupi_g46847(csa_tree_add_190_195_groupi_n_2409 ,csa_tree_add_190_195_groupi_n_449);
  not csa_tree_add_190_195_groupi_g46851(csa_tree_add_190_195_groupi_n_2408 ,csa_tree_add_190_195_groupi_n_1251);
  not csa_tree_add_190_195_groupi_g46852(csa_tree_add_190_195_groupi_n_2407 ,csa_tree_add_190_195_groupi_n_1309);
  not csa_tree_add_190_195_groupi_g46853(csa_tree_add_190_195_groupi_n_2406 ,csa_tree_add_190_195_groupi_n_585);
  not csa_tree_add_190_195_groupi_drc_bufs(csa_tree_add_190_195_groupi_n_2327 ,csa_tree_add_190_195_groupi_n_2325);
  not csa_tree_add_190_195_groupi_drc_bufs46854(csa_tree_add_190_195_groupi_n_2326 ,csa_tree_add_190_195_groupi_n_2325);
  not csa_tree_add_190_195_groupi_drc_bufs46855(csa_tree_add_190_195_groupi_n_2325 ,n_454);
  not csa_tree_add_190_195_groupi_drc_bufs46859(csa_tree_add_190_195_groupi_n_2324 ,csa_tree_add_190_195_groupi_n_2322);
  not csa_tree_add_190_195_groupi_drc_bufs46860(csa_tree_add_190_195_groupi_n_2323 ,csa_tree_add_190_195_groupi_n_2322);
  not csa_tree_add_190_195_groupi_drc_bufs46861(csa_tree_add_190_195_groupi_n_2322 ,n_447);
  not csa_tree_add_190_195_groupi_drc_bufs46865(csa_tree_add_190_195_groupi_n_2321 ,csa_tree_add_190_195_groupi_n_2319);
  not csa_tree_add_190_195_groupi_drc_bufs46866(csa_tree_add_190_195_groupi_n_2320 ,csa_tree_add_190_195_groupi_n_2319);
  not csa_tree_add_190_195_groupi_drc_bufs46867(csa_tree_add_190_195_groupi_n_2319 ,n_362);
  not csa_tree_add_190_195_groupi_drc_bufs46871(csa_tree_add_190_195_groupi_n_2318 ,csa_tree_add_190_195_groupi_n_2316);
  not csa_tree_add_190_195_groupi_drc_bufs46872(csa_tree_add_190_195_groupi_n_2317 ,csa_tree_add_190_195_groupi_n_2316);
  not csa_tree_add_190_195_groupi_drc_bufs46873(csa_tree_add_190_195_groupi_n_2316 ,n_369);
  not csa_tree_add_190_195_groupi_drc_bufs46877(csa_tree_add_190_195_groupi_n_2315 ,csa_tree_add_190_195_groupi_n_2313);
  not csa_tree_add_190_195_groupi_drc_bufs46878(csa_tree_add_190_195_groupi_n_2314 ,csa_tree_add_190_195_groupi_n_2313);
  not csa_tree_add_190_195_groupi_drc_bufs46879(csa_tree_add_190_195_groupi_n_2313 ,n_430);
  not csa_tree_add_190_195_groupi_drc_bufs46883(csa_tree_add_190_195_groupi_n_2312 ,csa_tree_add_190_195_groupi_n_2310);
  not csa_tree_add_190_195_groupi_drc_bufs46884(csa_tree_add_190_195_groupi_n_2311 ,csa_tree_add_190_195_groupi_n_2310);
  not csa_tree_add_190_195_groupi_drc_bufs46885(csa_tree_add_190_195_groupi_n_2310 ,n_437);
  not csa_tree_add_190_195_groupi_drc_bufs46889(csa_tree_add_190_195_groupi_n_2309 ,csa_tree_add_190_195_groupi_n_2307);
  not csa_tree_add_190_195_groupi_drc_bufs46890(csa_tree_add_190_195_groupi_n_2308 ,csa_tree_add_190_195_groupi_n_2307);
  not csa_tree_add_190_195_groupi_drc_bufs46891(csa_tree_add_190_195_groupi_n_2307 ,n_452);
  not csa_tree_add_190_195_groupi_drc_bufs46895(csa_tree_add_190_195_groupi_n_2306 ,csa_tree_add_190_195_groupi_n_2304);
  not csa_tree_add_190_195_groupi_drc_bufs46896(csa_tree_add_190_195_groupi_n_2305 ,csa_tree_add_190_195_groupi_n_2304);
  not csa_tree_add_190_195_groupi_drc_bufs46897(csa_tree_add_190_195_groupi_n_2304 ,n_367);
  not csa_tree_add_190_195_groupi_drc_bufs46901(csa_tree_add_190_195_groupi_n_2303 ,csa_tree_add_190_195_groupi_n_2301);
  not csa_tree_add_190_195_groupi_drc_bufs46902(csa_tree_add_190_195_groupi_n_2302 ,csa_tree_add_190_195_groupi_n_2301);
  not csa_tree_add_190_195_groupi_drc_bufs46903(csa_tree_add_190_195_groupi_n_2301 ,n_442);
  not csa_tree_add_190_195_groupi_drc_bufs46907(csa_tree_add_190_195_groupi_n_2300 ,csa_tree_add_190_195_groupi_n_2298);
  not csa_tree_add_190_195_groupi_drc_bufs46908(csa_tree_add_190_195_groupi_n_2299 ,csa_tree_add_190_195_groupi_n_2298);
  not csa_tree_add_190_195_groupi_drc_bufs46909(csa_tree_add_190_195_groupi_n_2298 ,n_359);
  not csa_tree_add_190_195_groupi_drc_bufs46913(csa_tree_add_190_195_groupi_n_2297 ,csa_tree_add_190_195_groupi_n_2295);
  not csa_tree_add_190_195_groupi_drc_bufs46914(csa_tree_add_190_195_groupi_n_2296 ,csa_tree_add_190_195_groupi_n_2295);
  not csa_tree_add_190_195_groupi_drc_bufs46915(csa_tree_add_190_195_groupi_n_2295 ,n_435);
  not csa_tree_add_190_195_groupi_drc_bufs46919(csa_tree_add_190_195_groupi_n_2294 ,csa_tree_add_190_195_groupi_n_2292);
  not csa_tree_add_190_195_groupi_drc_bufs46920(csa_tree_add_190_195_groupi_n_2293 ,csa_tree_add_190_195_groupi_n_2292);
  not csa_tree_add_190_195_groupi_drc_bufs46921(csa_tree_add_190_195_groupi_n_2292 ,n_335);
  not csa_tree_add_190_195_groupi_drc_bufs46924(csa_tree_add_190_195_groupi_n_2291 ,csa_tree_add_190_195_groupi_n_2289);
  not csa_tree_add_190_195_groupi_drc_bufs46925(csa_tree_add_190_195_groupi_n_2290 ,csa_tree_add_190_195_groupi_n_2289);
  not csa_tree_add_190_195_groupi_drc_bufs46926(csa_tree_add_190_195_groupi_n_2289 ,n_441);
  not csa_tree_add_190_195_groupi_drc_bufs46930(csa_tree_add_190_195_groupi_n_2288 ,csa_tree_add_190_195_groupi_n_2286);
  not csa_tree_add_190_195_groupi_drc_bufs46931(csa_tree_add_190_195_groupi_n_2287 ,csa_tree_add_190_195_groupi_n_2286);
  not csa_tree_add_190_195_groupi_drc_bufs46932(csa_tree_add_190_195_groupi_n_2286 ,n_326);
  not csa_tree_add_190_195_groupi_drc_bufs46936(csa_tree_add_190_195_groupi_n_2285 ,csa_tree_add_190_195_groupi_n_2283);
  not csa_tree_add_190_195_groupi_drc_bufs46937(csa_tree_add_190_195_groupi_n_2284 ,csa_tree_add_190_195_groupi_n_2283);
  not csa_tree_add_190_195_groupi_drc_bufs46938(csa_tree_add_190_195_groupi_n_2283 ,n_440);
  not csa_tree_add_190_195_groupi_drc_bufs46942(csa_tree_add_190_195_groupi_n_2282 ,csa_tree_add_190_195_groupi_n_2280);
  not csa_tree_add_190_195_groupi_drc_bufs46943(csa_tree_add_190_195_groupi_n_2281 ,csa_tree_add_190_195_groupi_n_2280);
  not csa_tree_add_190_195_groupi_drc_bufs46944(csa_tree_add_190_195_groupi_n_2280 ,n_445);
  not csa_tree_add_190_195_groupi_drc_bufs46948(csa_tree_add_190_195_groupi_n_2279 ,csa_tree_add_190_195_groupi_n_2277);
  not csa_tree_add_190_195_groupi_drc_bufs46949(csa_tree_add_190_195_groupi_n_2278 ,csa_tree_add_190_195_groupi_n_2277);
  not csa_tree_add_190_195_groupi_drc_bufs46950(csa_tree_add_190_195_groupi_n_2277 ,n_332);
  not csa_tree_add_190_195_groupi_drc_bufs46954(csa_tree_add_190_195_groupi_n_2276 ,csa_tree_add_190_195_groupi_n_2274);
  not csa_tree_add_190_195_groupi_drc_bufs46955(csa_tree_add_190_195_groupi_n_2275 ,csa_tree_add_190_195_groupi_n_2274);
  not csa_tree_add_190_195_groupi_drc_bufs46956(csa_tree_add_190_195_groupi_n_2274 ,n_451);
  not csa_tree_add_190_195_groupi_drc_bufs46960(csa_tree_add_190_195_groupi_n_2273 ,csa_tree_add_190_195_groupi_n_2271);
  not csa_tree_add_190_195_groupi_drc_bufs46961(csa_tree_add_190_195_groupi_n_2272 ,csa_tree_add_190_195_groupi_n_2271);
  not csa_tree_add_190_195_groupi_drc_bufs46962(csa_tree_add_190_195_groupi_n_2271 ,n_450);
  not csa_tree_add_190_195_groupi_drc_bufs46966(csa_tree_add_190_195_groupi_n_2270 ,csa_tree_add_190_195_groupi_n_2268);
  not csa_tree_add_190_195_groupi_drc_bufs46967(csa_tree_add_190_195_groupi_n_2269 ,csa_tree_add_190_195_groupi_n_2268);
  not csa_tree_add_190_195_groupi_drc_bufs46968(csa_tree_add_190_195_groupi_n_2268 ,n_365);
  not csa_tree_add_190_195_groupi_drc_bufs46972(csa_tree_add_190_195_groupi_n_2267 ,csa_tree_add_190_195_groupi_n_2265);
  not csa_tree_add_190_195_groupi_drc_bufs46973(csa_tree_add_190_195_groupi_n_2266 ,csa_tree_add_190_195_groupi_n_2265);
  not csa_tree_add_190_195_groupi_drc_bufs46974(csa_tree_add_190_195_groupi_n_2265 ,n_429);
  not csa_tree_add_190_195_groupi_drc_bufs46978(csa_tree_add_190_195_groupi_n_2264 ,csa_tree_add_190_195_groupi_n_2262);
  not csa_tree_add_190_195_groupi_drc_bufs46979(csa_tree_add_190_195_groupi_n_2263 ,csa_tree_add_190_195_groupi_n_2262);
  not csa_tree_add_190_195_groupi_drc_bufs46980(csa_tree_add_190_195_groupi_n_2262 ,n_373);
  not csa_tree_add_190_195_groupi_drc_bufs46984(csa_tree_add_190_195_groupi_n_2261 ,csa_tree_add_190_195_groupi_n_2259);
  not csa_tree_add_190_195_groupi_drc_bufs46985(csa_tree_add_190_195_groupi_n_2260 ,csa_tree_add_190_195_groupi_n_2259);
  not csa_tree_add_190_195_groupi_drc_bufs46986(csa_tree_add_190_195_groupi_n_2259 ,n_370);
  not csa_tree_add_190_195_groupi_drc_bufs46990(csa_tree_add_190_195_groupi_n_2258 ,csa_tree_add_190_195_groupi_n_2256);
  not csa_tree_add_190_195_groupi_drc_bufs46991(csa_tree_add_190_195_groupi_n_2257 ,csa_tree_add_190_195_groupi_n_2256);
  not csa_tree_add_190_195_groupi_drc_bufs46992(csa_tree_add_190_195_groupi_n_2256 ,n_438);
  not csa_tree_add_190_195_groupi_drc_bufs46996(csa_tree_add_190_195_groupi_n_2255 ,csa_tree_add_190_195_groupi_n_2253);
  not csa_tree_add_190_195_groupi_drc_bufs46997(csa_tree_add_190_195_groupi_n_2254 ,csa_tree_add_190_195_groupi_n_2253);
  not csa_tree_add_190_195_groupi_drc_bufs46998(csa_tree_add_190_195_groupi_n_2253 ,n_455);
  not csa_tree_add_190_195_groupi_drc_bufs47002(csa_tree_add_190_195_groupi_n_2252 ,csa_tree_add_190_195_groupi_n_2250);
  not csa_tree_add_190_195_groupi_drc_bufs47003(csa_tree_add_190_195_groupi_n_2251 ,csa_tree_add_190_195_groupi_n_2250);
  not csa_tree_add_190_195_groupi_drc_bufs47004(csa_tree_add_190_195_groupi_n_2250 ,n_426);
  not csa_tree_add_190_195_groupi_drc_bufs47008(csa_tree_add_190_195_groupi_n_2249 ,csa_tree_add_190_195_groupi_n_2247);
  not csa_tree_add_190_195_groupi_drc_bufs47009(csa_tree_add_190_195_groupi_n_2248 ,csa_tree_add_190_195_groupi_n_2247);
  not csa_tree_add_190_195_groupi_drc_bufs47010(csa_tree_add_190_195_groupi_n_2247 ,n_330);
  not csa_tree_add_190_195_groupi_drc_bufs47014(csa_tree_add_190_195_groupi_n_2246 ,csa_tree_add_190_195_groupi_n_2244);
  not csa_tree_add_190_195_groupi_drc_bufs47015(csa_tree_add_190_195_groupi_n_2245 ,csa_tree_add_190_195_groupi_n_2244);
  not csa_tree_add_190_195_groupi_drc_bufs47016(csa_tree_add_190_195_groupi_n_2244 ,n_420);
  not csa_tree_add_190_195_groupi_drc_bufs47019(csa_tree_add_190_195_groupi_n_2243 ,csa_tree_add_190_195_groupi_n_2241);
  not csa_tree_add_190_195_groupi_drc_bufs47020(csa_tree_add_190_195_groupi_n_2242 ,csa_tree_add_190_195_groupi_n_2241);
  not csa_tree_add_190_195_groupi_drc_bufs47021(csa_tree_add_190_195_groupi_n_2241 ,n_250);
  not csa_tree_add_190_195_groupi_drc_bufs47024(csa_tree_add_190_195_groupi_n_2240 ,csa_tree_add_190_195_groupi_n_2238);
  not csa_tree_add_190_195_groupi_drc_bufs47025(csa_tree_add_190_195_groupi_n_2239 ,csa_tree_add_190_195_groupi_n_2238);
  not csa_tree_add_190_195_groupi_drc_bufs47026(csa_tree_add_190_195_groupi_n_2238 ,n_243);
  not csa_tree_add_190_195_groupi_drc_bufs47029(csa_tree_add_190_195_groupi_n_2237 ,csa_tree_add_190_195_groupi_n_2235);
  not csa_tree_add_190_195_groupi_drc_bufs47030(csa_tree_add_190_195_groupi_n_2236 ,csa_tree_add_190_195_groupi_n_2235);
  not csa_tree_add_190_195_groupi_drc_bufs47031(csa_tree_add_190_195_groupi_n_2235 ,n_360);
  not csa_tree_add_190_195_groupi_drc_bufs47034(csa_tree_add_190_195_groupi_n_2234 ,csa_tree_add_190_195_groupi_n_2232);
  not csa_tree_add_190_195_groupi_drc_bufs47035(csa_tree_add_190_195_groupi_n_2233 ,csa_tree_add_190_195_groupi_n_2232);
  not csa_tree_add_190_195_groupi_drc_bufs47036(csa_tree_add_190_195_groupi_n_2232 ,n_366);
  not csa_tree_add_190_195_groupi_drc_bufs47039(csa_tree_add_190_195_groupi_n_2231 ,csa_tree_add_190_195_groupi_n_2229);
  not csa_tree_add_190_195_groupi_drc_bufs47040(csa_tree_add_190_195_groupi_n_2230 ,csa_tree_add_190_195_groupi_n_2229);
  not csa_tree_add_190_195_groupi_drc_bufs47041(csa_tree_add_190_195_groupi_n_2229 ,n_433);
  not csa_tree_add_190_195_groupi_drc_bufs47044(csa_tree_add_190_195_groupi_n_2228 ,csa_tree_add_190_195_groupi_n_2226);
  not csa_tree_add_190_195_groupi_drc_bufs47045(csa_tree_add_190_195_groupi_n_2227 ,csa_tree_add_190_195_groupi_n_2226);
  not csa_tree_add_190_195_groupi_drc_bufs47046(csa_tree_add_190_195_groupi_n_2226 ,n_428);
  not csa_tree_add_190_195_groupi_drc_bufs47049(csa_tree_add_190_195_groupi_n_2225 ,csa_tree_add_190_195_groupi_n_2223);
  not csa_tree_add_190_195_groupi_drc_bufs47050(csa_tree_add_190_195_groupi_n_2224 ,csa_tree_add_190_195_groupi_n_2223);
  not csa_tree_add_190_195_groupi_drc_bufs47051(csa_tree_add_190_195_groupi_n_2223 ,n_299);
  not csa_tree_add_190_195_groupi_drc_bufs47054(csa_tree_add_190_195_groupi_n_2222 ,csa_tree_add_190_195_groupi_n_2220);
  not csa_tree_add_190_195_groupi_drc_bufs47055(csa_tree_add_190_195_groupi_n_2221 ,csa_tree_add_190_195_groupi_n_2220);
  not csa_tree_add_190_195_groupi_drc_bufs47056(csa_tree_add_190_195_groupi_n_2220 ,n_418);
  not csa_tree_add_190_195_groupi_drc_bufs47059(csa_tree_add_190_195_groupi_n_2219 ,csa_tree_add_190_195_groupi_n_2217);
  not csa_tree_add_190_195_groupi_drc_bufs47060(csa_tree_add_190_195_groupi_n_2218 ,csa_tree_add_190_195_groupi_n_2217);
  not csa_tree_add_190_195_groupi_drc_bufs47061(csa_tree_add_190_195_groupi_n_2217 ,n_401);
  not csa_tree_add_190_195_groupi_drc_bufs47104(csa_tree_add_190_195_groupi_n_2208 ,csa_tree_add_190_195_groupi_n_2206);
  not csa_tree_add_190_195_groupi_drc_bufs47105(csa_tree_add_190_195_groupi_n_2207 ,csa_tree_add_190_195_groupi_n_2206);
  not csa_tree_add_190_195_groupi_drc_bufs47106(csa_tree_add_190_195_groupi_n_2206 ,n_361);
  not csa_tree_add_190_195_groupi_drc_bufs47109(csa_tree_add_190_195_groupi_n_2205 ,csa_tree_add_190_195_groupi_n_2203);
  not csa_tree_add_190_195_groupi_drc_bufs47110(csa_tree_add_190_195_groupi_n_2204 ,csa_tree_add_190_195_groupi_n_2203);
  not csa_tree_add_190_195_groupi_drc_bufs47111(csa_tree_add_190_195_groupi_n_2203 ,n_446);
  not csa_tree_add_190_195_groupi_drc_bufs47114(csa_tree_add_190_195_groupi_n_2202 ,csa_tree_add_190_195_groupi_n_2200);
  not csa_tree_add_190_195_groupi_drc_bufs47115(csa_tree_add_190_195_groupi_n_2201 ,csa_tree_add_190_195_groupi_n_2200);
  not csa_tree_add_190_195_groupi_drc_bufs47116(csa_tree_add_190_195_groupi_n_2200 ,n_371);
  not csa_tree_add_190_195_groupi_drc_bufs47119(csa_tree_add_190_195_groupi_n_2199 ,csa_tree_add_190_195_groupi_n_2197);
  not csa_tree_add_190_195_groupi_drc_bufs47120(csa_tree_add_190_195_groupi_n_2198 ,csa_tree_add_190_195_groupi_n_2197);
  not csa_tree_add_190_195_groupi_drc_bufs47121(csa_tree_add_190_195_groupi_n_2197 ,n_444);
  not csa_tree_add_190_195_groupi_drc_bufs47124(csa_tree_add_190_195_groupi_n_2196 ,csa_tree_add_190_195_groupi_n_2194);
  not csa_tree_add_190_195_groupi_drc_bufs47125(csa_tree_add_190_195_groupi_n_2195 ,csa_tree_add_190_195_groupi_n_2194);
  not csa_tree_add_190_195_groupi_drc_bufs47126(csa_tree_add_190_195_groupi_n_2194 ,n_449);
  not csa_tree_add_190_195_groupi_drc_bufs47129(csa_tree_add_190_195_groupi_n_2193 ,csa_tree_add_190_195_groupi_n_2191);
  not csa_tree_add_190_195_groupi_drc_bufs47130(csa_tree_add_190_195_groupi_n_2192 ,csa_tree_add_190_195_groupi_n_2191);
  not csa_tree_add_190_195_groupi_drc_bufs47131(csa_tree_add_190_195_groupi_n_2191 ,n_364);
  not csa_tree_add_190_195_groupi_drc_bufs47134(csa_tree_add_190_195_groupi_n_2190 ,csa_tree_add_190_195_groupi_n_2188);
  not csa_tree_add_190_195_groupi_drc_bufs47135(csa_tree_add_190_195_groupi_n_2189 ,csa_tree_add_190_195_groupi_n_2188);
  not csa_tree_add_190_195_groupi_drc_bufs47136(csa_tree_add_190_195_groupi_n_2188 ,n_436);
  not csa_tree_add_190_195_groupi_drc_bufs47139(csa_tree_add_190_195_groupi_n_2187 ,csa_tree_add_190_195_groupi_n_2185);
  not csa_tree_add_190_195_groupi_drc_bufs47140(csa_tree_add_190_195_groupi_n_2186 ,csa_tree_add_190_195_groupi_n_2185);
  not csa_tree_add_190_195_groupi_drc_bufs47141(csa_tree_add_190_195_groupi_n_2185 ,n_453);
  not csa_tree_add_190_195_groupi_drc_bufs47144(csa_tree_add_190_195_groupi_n_2184 ,csa_tree_add_190_195_groupi_n_2182);
  not csa_tree_add_190_195_groupi_drc_bufs47145(csa_tree_add_190_195_groupi_n_2183 ,csa_tree_add_190_195_groupi_n_2182);
  not csa_tree_add_190_195_groupi_drc_bufs47146(csa_tree_add_190_195_groupi_n_2182 ,n_358);
  not csa_tree_add_190_195_groupi_drc_bufs47149(csa_tree_add_190_195_groupi_n_2181 ,csa_tree_add_190_195_groupi_n_2179);
  not csa_tree_add_190_195_groupi_drc_bufs47150(csa_tree_add_190_195_groupi_n_2180 ,csa_tree_add_190_195_groupi_n_2179);
  not csa_tree_add_190_195_groupi_drc_bufs47151(csa_tree_add_190_195_groupi_n_2179 ,n_434);
  not csa_tree_add_190_195_groupi_drc_bufs47154(csa_tree_add_190_195_groupi_n_2178 ,csa_tree_add_190_195_groupi_n_2176);
  not csa_tree_add_190_195_groupi_drc_bufs47155(csa_tree_add_190_195_groupi_n_2177 ,csa_tree_add_190_195_groupi_n_2176);
  not csa_tree_add_190_195_groupi_drc_bufs47156(csa_tree_add_190_195_groupi_n_2176 ,n_399);
  not csa_tree_add_190_195_groupi_drc_bufs47159(csa_tree_add_190_195_groupi_n_2175 ,csa_tree_add_190_195_groupi_n_2174);
  not csa_tree_add_190_195_groupi_drc_bufs47161(csa_tree_add_190_195_groupi_n_2174 ,n_197);
  not csa_tree_add_190_195_groupi_drc_bufs47164(csa_tree_add_190_195_groupi_n_2173 ,csa_tree_add_190_195_groupi_n_2172);
  not csa_tree_add_190_195_groupi_drc_bufs47166(csa_tree_add_190_195_groupi_n_2172 ,n_265);
  not csa_tree_add_190_195_groupi_drc_bufs47169(csa_tree_add_190_195_groupi_n_2171 ,csa_tree_add_190_195_groupi_n_2170);
  not csa_tree_add_190_195_groupi_drc_bufs47171(csa_tree_add_190_195_groupi_n_2170 ,n_248);
  not csa_tree_add_190_195_groupi_drc_bufs47174(csa_tree_add_190_195_groupi_n_2169 ,csa_tree_add_190_195_groupi_n_2168);
  not csa_tree_add_190_195_groupi_drc_bufs47176(csa_tree_add_190_195_groupi_n_2168 ,n_333);
  not csa_tree_add_190_195_groupi_drc_bufs47179(csa_tree_add_190_195_groupi_n_2167 ,csa_tree_add_190_195_groupi_n_2165);
  not csa_tree_add_190_195_groupi_drc_bufs47180(csa_tree_add_190_195_groupi_n_2166 ,csa_tree_add_190_195_groupi_n_2165);
  not csa_tree_add_190_195_groupi_drc_bufs47181(csa_tree_add_190_195_groupi_n_2165 ,n_387);
  not csa_tree_add_190_195_groupi_drc_bufs47184(csa_tree_add_190_195_groupi_n_2164 ,csa_tree_add_190_195_groupi_n_2162);
  not csa_tree_add_190_195_groupi_drc_bufs47185(csa_tree_add_190_195_groupi_n_2163 ,csa_tree_add_190_195_groupi_n_2162);
  not csa_tree_add_190_195_groupi_drc_bufs47186(csa_tree_add_190_195_groupi_n_2162 ,n_421);
  not csa_tree_add_190_195_groupi_drc_bufs47189(csa_tree_add_190_195_groupi_n_2161 ,csa_tree_add_190_195_groupi_n_2159);
  not csa_tree_add_190_195_groupi_drc_bufs47190(csa_tree_add_190_195_groupi_n_2160 ,csa_tree_add_190_195_groupi_n_2159);
  not csa_tree_add_190_195_groupi_drc_bufs47191(csa_tree_add_190_195_groupi_n_2159 ,n_336);
  not csa_tree_add_190_195_groupi_drc_bufs47222(csa_tree_add_190_195_groupi_n_2151 ,csa_tree_add_190_195_groupi_n_2149);
  not csa_tree_add_190_195_groupi_drc_bufs47223(csa_tree_add_190_195_groupi_n_2150 ,csa_tree_add_190_195_groupi_n_2149);
  not csa_tree_add_190_195_groupi_drc_bufs47224(csa_tree_add_190_195_groupi_n_2149 ,n_432);
  not csa_tree_add_190_195_groupi_drc_bufs47227(csa_tree_add_190_195_groupi_n_2148 ,csa_tree_add_190_195_groupi_n_2147);
  not csa_tree_add_190_195_groupi_drc_bufs47229(csa_tree_add_190_195_groupi_n_2147 ,n_394);
  not csa_tree_add_190_195_groupi_drc_bufs47232(csa_tree_add_190_195_groupi_n_2146 ,csa_tree_add_190_195_groupi_n_2144);
  not csa_tree_add_190_195_groupi_drc_bufs47233(csa_tree_add_190_195_groupi_n_2145 ,csa_tree_add_190_195_groupi_n_2144);
  not csa_tree_add_190_195_groupi_drc_bufs47234(csa_tree_add_190_195_groupi_n_2144 ,n_157);
  not csa_tree_add_190_195_groupi_drc_bufs47237(csa_tree_add_190_195_groupi_n_2143 ,csa_tree_add_190_195_groupi_n_2142);
  not csa_tree_add_190_195_groupi_drc_bufs47239(csa_tree_add_190_195_groupi_n_2142 ,n_331);
  not csa_tree_add_190_195_groupi_drc_bufs47242(csa_tree_add_190_195_groupi_n_2141 ,csa_tree_add_190_195_groupi_n_2140);
  not csa_tree_add_190_195_groupi_drc_bufs47244(csa_tree_add_190_195_groupi_n_2140 ,n_162);
  not csa_tree_add_190_195_groupi_drc_bufs47247(csa_tree_add_190_195_groupi_n_2139 ,csa_tree_add_190_195_groupi_n_2138);
  not csa_tree_add_190_195_groupi_drc_bufs47249(csa_tree_add_190_195_groupi_n_2138 ,n_382);
  not csa_tree_add_190_195_groupi_drc_bufs47252(csa_tree_add_190_195_groupi_n_2137 ,csa_tree_add_190_195_groupi_n_2136);
  not csa_tree_add_190_195_groupi_drc_bufs47254(csa_tree_add_190_195_groupi_n_2136 ,n_264);
  not csa_tree_add_190_195_groupi_drc_bufs47257(csa_tree_add_190_195_groupi_n_2135 ,csa_tree_add_190_195_groupi_n_2134);
  not csa_tree_add_190_195_groupi_drc_bufs47259(csa_tree_add_190_195_groupi_n_2134 ,n_230);
  not csa_tree_add_190_195_groupi_drc_bufs47262(csa_tree_add_190_195_groupi_n_2133 ,csa_tree_add_190_195_groupi_n_2132);
  not csa_tree_add_190_195_groupi_drc_bufs47264(csa_tree_add_190_195_groupi_n_2132 ,n_166);
  not csa_tree_add_190_195_groupi_drc_bufs47267(csa_tree_add_190_195_groupi_n_2131 ,csa_tree_add_190_195_groupi_n_2130);
  not csa_tree_add_190_195_groupi_drc_bufs47269(csa_tree_add_190_195_groupi_n_2130 ,n_149);
  not csa_tree_add_190_195_groupi_drc_bufs47272(csa_tree_add_190_195_groupi_n_2129 ,csa_tree_add_190_195_groupi_n_2128);
  not csa_tree_add_190_195_groupi_drc_bufs47274(csa_tree_add_190_195_groupi_n_2128 ,n_302);
  not csa_tree_add_190_195_groupi_drc_bufs47277(csa_tree_add_190_195_groupi_n_2127 ,csa_tree_add_190_195_groupi_n_2126);
  not csa_tree_add_190_195_groupi_drc_bufs47279(csa_tree_add_190_195_groupi_n_2126 ,n_268);
  not csa_tree_add_190_195_groupi_drc_bufs47282(csa_tree_add_190_195_groupi_n_2125 ,csa_tree_add_190_195_groupi_n_2123);
  not csa_tree_add_190_195_groupi_drc_bufs47283(csa_tree_add_190_195_groupi_n_2124 ,csa_tree_add_190_195_groupi_n_2123);
  not csa_tree_add_190_195_groupi_drc_bufs47284(csa_tree_add_190_195_groupi_n_2123 ,n_427);
  not csa_tree_add_190_195_groupi_drc_bufs47287(csa_tree_add_190_195_groupi_n_2122 ,csa_tree_add_190_195_groupi_n_2120);
  not csa_tree_add_190_195_groupi_drc_bufs47288(csa_tree_add_190_195_groupi_n_2121 ,csa_tree_add_190_195_groupi_n_2120);
  not csa_tree_add_190_195_groupi_drc_bufs47289(csa_tree_add_190_195_groupi_n_2120 ,n_372);
  not csa_tree_add_190_195_groupi_drc_bufs47308(csa_tree_add_190_195_groupi_n_2115 ,csa_tree_add_190_195_groupi_n_2113);
  not csa_tree_add_190_195_groupi_drc_bufs47309(csa_tree_add_190_195_groupi_n_2114 ,csa_tree_add_190_195_groupi_n_2113);
  not csa_tree_add_190_195_groupi_drc_bufs47310(csa_tree_add_190_195_groupi_n_2113 ,n_228);
  not csa_tree_add_190_195_groupi_drc_bufs47313(csa_tree_add_190_195_groupi_n_2112 ,csa_tree_add_190_195_groupi_n_2110);
  not csa_tree_add_190_195_groupi_drc_bufs47314(csa_tree_add_190_195_groupi_n_2111 ,csa_tree_add_190_195_groupi_n_2110);
  not csa_tree_add_190_195_groupi_drc_bufs47315(csa_tree_add_190_195_groupi_n_2110 ,n_398);
  not csa_tree_add_190_195_groupi_drc_bufs47318(csa_tree_add_190_195_groupi_n_2109 ,csa_tree_add_190_195_groupi_n_2107);
  not csa_tree_add_190_195_groupi_drc_bufs47319(csa_tree_add_190_195_groupi_n_2108 ,csa_tree_add_190_195_groupi_n_2107);
  not csa_tree_add_190_195_groupi_drc_bufs47320(csa_tree_add_190_195_groupi_n_2107 ,n_385);
  not csa_tree_add_190_195_groupi_drc_bufs47323(csa_tree_add_190_195_groupi_n_2106 ,csa_tree_add_190_195_groupi_n_2104);
  not csa_tree_add_190_195_groupi_drc_bufs47324(csa_tree_add_190_195_groupi_n_2105 ,csa_tree_add_190_195_groupi_n_2104);
  not csa_tree_add_190_195_groupi_drc_bufs47325(csa_tree_add_190_195_groupi_n_2104 ,n_368);
  not csa_tree_add_190_195_groupi_drc_bufs47328(csa_tree_add_190_195_groupi_n_2103 ,csa_tree_add_190_195_groupi_n_2101);
  not csa_tree_add_190_195_groupi_drc_bufs47329(csa_tree_add_190_195_groupi_n_2102 ,csa_tree_add_190_195_groupi_n_2101);
  not csa_tree_add_190_195_groupi_drc_bufs47330(csa_tree_add_190_195_groupi_n_2101 ,n_363);
  not csa_tree_add_190_195_groupi_drc_bufs47333(csa_tree_add_190_195_groupi_n_2100 ,csa_tree_add_190_195_groupi_n_2098);
  not csa_tree_add_190_195_groupi_drc_bufs47334(csa_tree_add_190_195_groupi_n_2099 ,csa_tree_add_190_195_groupi_n_2098);
  not csa_tree_add_190_195_groupi_drc_bufs47335(csa_tree_add_190_195_groupi_n_2098 ,n_448);
  not csa_tree_add_190_195_groupi_drc_bufs47338(csa_tree_add_190_195_groupi_n_2097 ,csa_tree_add_190_195_groupi_n_2095);
  not csa_tree_add_190_195_groupi_drc_bufs47339(csa_tree_add_190_195_groupi_n_2096 ,csa_tree_add_190_195_groupi_n_2095);
  not csa_tree_add_190_195_groupi_drc_bufs47340(csa_tree_add_190_195_groupi_n_2095 ,n_458);
  not csa_tree_add_190_195_groupi_drc_bufs47343(csa_tree_add_190_195_groupi_n_2094 ,csa_tree_add_190_195_groupi_n_2092);
  not csa_tree_add_190_195_groupi_drc_bufs47344(csa_tree_add_190_195_groupi_n_2093 ,csa_tree_add_190_195_groupi_n_2092);
  not csa_tree_add_190_195_groupi_drc_bufs47345(csa_tree_add_190_195_groupi_n_2092 ,n_439);
  not csa_tree_add_190_195_groupi_drc_bufs47388(csa_tree_add_190_195_groupi_n_2081 ,csa_tree_add_190_195_groupi_n_2079);
  not csa_tree_add_190_195_groupi_drc_bufs47389(csa_tree_add_190_195_groupi_n_2080 ,csa_tree_add_190_195_groupi_n_2079);
  not csa_tree_add_190_195_groupi_drc_bufs47390(csa_tree_add_190_195_groupi_n_2079 ,n_459);
  not csa_tree_add_190_195_groupi_drc_bufs47393(csa_tree_add_190_195_groupi_n_2078 ,csa_tree_add_190_195_groupi_n_2076);
  not csa_tree_add_190_195_groupi_drc_bufs47394(csa_tree_add_190_195_groupi_n_2077 ,csa_tree_add_190_195_groupi_n_2076);
  not csa_tree_add_190_195_groupi_drc_bufs47395(csa_tree_add_190_195_groupi_n_2076 ,n_374);
  not csa_tree_add_190_195_groupi_drc_bufs47398(csa_tree_add_190_195_groupi_n_2075 ,csa_tree_add_190_195_groupi_n_2073);
  not csa_tree_add_190_195_groupi_drc_bufs47399(csa_tree_add_190_195_groupi_n_2074 ,csa_tree_add_190_195_groupi_n_2073);
  not csa_tree_add_190_195_groupi_drc_bufs47400(csa_tree_add_190_195_groupi_n_2073 ,n_337);
  not csa_tree_add_190_195_groupi_drc_bufs47403(csa_tree_add_190_195_groupi_n_2072 ,csa_tree_add_190_195_groupi_n_2070);
  not csa_tree_add_190_195_groupi_drc_bufs47404(csa_tree_add_190_195_groupi_n_2071 ,csa_tree_add_190_195_groupi_n_2070);
  not csa_tree_add_190_195_groupi_drc_bufs47405(csa_tree_add_190_195_groupi_n_2070 ,n_443);
  not csa_tree_add_190_195_groupi_drc_bufs47408(csa_tree_add_190_195_groupi_n_2069 ,csa_tree_add_190_195_groupi_n_2067);
  not csa_tree_add_190_195_groupi_drc_bufs47409(csa_tree_add_190_195_groupi_n_2068 ,csa_tree_add_190_195_groupi_n_2067);
  not csa_tree_add_190_195_groupi_drc_bufs47410(csa_tree_add_190_195_groupi_n_2067 ,n_324);
  not csa_tree_add_190_195_groupi_drc_bufs47413(csa_tree_add_190_195_groupi_n_2066 ,csa_tree_add_190_195_groupi_n_2065);
  not csa_tree_add_190_195_groupi_drc_bufs47415(csa_tree_add_190_195_groupi_n_2065 ,n_242);
  not csa_tree_add_190_195_groupi_drc_bufs47482(csa_tree_add_190_195_groupi_n_2048 ,csa_tree_add_190_195_groupi_n_2047);
  not csa_tree_add_190_195_groupi_drc_bufs47484(csa_tree_add_190_195_groupi_n_2047 ,n_325);
  not csa_tree_add_190_195_groupi_drc_bufs47487(csa_tree_add_190_195_groupi_n_2046 ,csa_tree_add_190_195_groupi_n_2045);
  not csa_tree_add_190_195_groupi_drc_bufs47489(csa_tree_add_190_195_groupi_n_2045 ,n_257);
  not csa_tree_add_190_195_groupi_drc_bufs47492(csa_tree_add_190_195_groupi_n_2044 ,csa_tree_add_190_195_groupi_n_2043);
  not csa_tree_add_190_195_groupi_drc_bufs47494(csa_tree_add_190_195_groupi_n_2043 ,n_240);
  not csa_tree_add_190_195_groupi_drc_bufs47513(csa_tree_add_190_195_groupi_n_2038 ,csa_tree_add_190_195_groupi_n_2037);
  not csa_tree_add_190_195_groupi_drc_bufs47515(csa_tree_add_190_195_groupi_n_2037 ,n_160);
  not csa_tree_add_190_195_groupi_drc_bufs47518(csa_tree_add_190_195_groupi_n_2036 ,csa_tree_add_190_195_groupi_n_2035);
  not csa_tree_add_190_195_groupi_drc_bufs47520(csa_tree_add_190_195_groupi_n_2035 ,n_381);
  not csa_tree_add_190_195_groupi_drc_bufs47523(csa_tree_add_190_195_groupi_n_2034 ,csa_tree_add_190_195_groupi_n_2033);
  not csa_tree_add_190_195_groupi_drc_bufs47525(csa_tree_add_190_195_groupi_n_2033 ,n_198);
  not csa_tree_add_190_195_groupi_drc_bufs47528(csa_tree_add_190_195_groupi_n_2032 ,csa_tree_add_190_195_groupi_n_2031);
  not csa_tree_add_190_195_groupi_drc_bufs47530(csa_tree_add_190_195_groupi_n_2031 ,n_164);
  not csa_tree_add_190_195_groupi_drc_bufs47533(csa_tree_add_190_195_groupi_n_2030 ,csa_tree_add_190_195_groupi_n_2029);
  not csa_tree_add_190_195_groupi_drc_bufs47535(csa_tree_add_190_195_groupi_n_2029 ,n_266);
  not csa_tree_add_190_195_groupi_drc_bufs47538(csa_tree_add_190_195_groupi_n_2028 ,csa_tree_add_190_195_groupi_n_2026);
  not csa_tree_add_190_195_groupi_drc_bufs47539(csa_tree_add_190_195_groupi_n_2027 ,csa_tree_add_190_195_groupi_n_2026);
  not csa_tree_add_190_195_groupi_drc_bufs47540(csa_tree_add_190_195_groupi_n_2026 ,n_142);
  not csa_tree_add_190_195_groupi_drc_bufs47543(csa_tree_add_190_195_groupi_n_2025 ,csa_tree_add_190_195_groupi_n_2023);
  not csa_tree_add_190_195_groupi_drc_bufs47544(csa_tree_add_190_195_groupi_n_2024 ,csa_tree_add_190_195_groupi_n_2023);
  not csa_tree_add_190_195_groupi_drc_bufs47545(csa_tree_add_190_195_groupi_n_2023 ,n_407);
  not csa_tree_add_190_195_groupi_drc_bufs47548(csa_tree_add_190_195_groupi_n_2022 ,csa_tree_add_190_195_groupi_n_2020);
  not csa_tree_add_190_195_groupi_drc_bufs47549(csa_tree_add_190_195_groupi_n_2021 ,csa_tree_add_190_195_groupi_n_2020);
  not csa_tree_add_190_195_groupi_drc_bufs47550(csa_tree_add_190_195_groupi_n_2020 ,n_237);
  not csa_tree_add_190_195_groupi_drc_bufs47553(csa_tree_add_190_195_groupi_n_2019 ,csa_tree_add_190_195_groupi_n_2017);
  not csa_tree_add_190_195_groupi_drc_bufs47554(csa_tree_add_190_195_groupi_n_2018 ,csa_tree_add_190_195_groupi_n_2017);
  not csa_tree_add_190_195_groupi_drc_bufs47555(csa_tree_add_190_195_groupi_n_2017 ,n_425);
  not csa_tree_add_190_195_groupi_drc_bufs47566(csa_tree_add_190_195_groupi_n_2014 ,csa_tree_add_190_195_groupi_n_2012);
  not csa_tree_add_190_195_groupi_drc_bufs47567(csa_tree_add_190_195_groupi_n_2013 ,csa_tree_add_190_195_groupi_n_2012);
  not csa_tree_add_190_195_groupi_drc_bufs47568(csa_tree_add_190_195_groupi_n_2012 ,n_256);
  not csa_tree_add_190_195_groupi_drc_bufs47571(csa_tree_add_190_195_groupi_n_2011 ,csa_tree_add_190_195_groupi_n_2009);
  not csa_tree_add_190_195_groupi_drc_bufs47572(csa_tree_add_190_195_groupi_n_2010 ,csa_tree_add_190_195_groupi_n_2009);
  not csa_tree_add_190_195_groupi_drc_bufs47573(csa_tree_add_190_195_groupi_n_2009 ,n_205);
  not csa_tree_add_190_195_groupi_drc_bufs47594(csa_tree_add_190_195_groupi_n_2375 ,csa_tree_add_190_195_groupi_n_2004);
  not csa_tree_add_190_195_groupi_drc_bufs47602(csa_tree_add_190_195_groupi_n_2350 ,csa_tree_add_190_195_groupi_n_2002);
  not csa_tree_add_190_195_groupi_drc_bufs47610(csa_tree_add_190_195_groupi_n_2376 ,csa_tree_add_190_195_groupi_n_2000);
  not csa_tree_add_190_195_groupi_drc_bufs47664(csa_tree_add_190_195_groupi_n_1986 ,csa_tree_add_190_195_groupi_n_1985);
  not csa_tree_add_190_195_groupi_drc_bufs47666(csa_tree_add_190_195_groupi_n_1985 ,n_329);
  not csa_tree_add_190_195_groupi_drc_bufs47669(csa_tree_add_190_195_groupi_n_1984 ,csa_tree_add_190_195_groupi_n_1983);
  not csa_tree_add_190_195_groupi_drc_bufs47671(csa_tree_add_190_195_groupi_n_1983 ,n_159);
  not csa_tree_add_190_195_groupi_drc_bufs47674(csa_tree_add_190_195_groupi_n_1982 ,csa_tree_add_190_195_groupi_n_1981);
  not csa_tree_add_190_195_groupi_drc_bufs47676(csa_tree_add_190_195_groupi_n_1981 ,n_295);
  not csa_tree_add_190_195_groupi_drc_bufs47679(csa_tree_add_190_195_groupi_n_1980 ,csa_tree_add_190_195_groupi_n_1979);
  not csa_tree_add_190_195_groupi_drc_bufs47681(csa_tree_add_190_195_groupi_n_1979 ,n_346);
  not csa_tree_add_190_195_groupi_drc_bufs47760(csa_tree_add_190_195_groupi_n_1959 ,csa_tree_add_190_195_groupi_n_1958);
  not csa_tree_add_190_195_groupi_drc_bufs47762(csa_tree_add_190_195_groupi_n_1958 ,n_271);
  not csa_tree_add_190_195_groupi_drc_bufs47765(csa_tree_add_190_195_groupi_n_1957 ,csa_tree_add_190_195_groupi_n_1956);
  not csa_tree_add_190_195_groupi_drc_bufs47767(csa_tree_add_190_195_groupi_n_1956 ,n_339);
  not csa_tree_add_190_195_groupi_drc_bufs47770(csa_tree_add_190_195_groupi_n_1955 ,csa_tree_add_190_195_groupi_n_1954);
  not csa_tree_add_190_195_groupi_drc_bufs47772(csa_tree_add_190_195_groupi_n_1954 ,n_170);
  not csa_tree_add_190_195_groupi_drc_bufs47775(csa_tree_add_190_195_groupi_n_1953 ,csa_tree_add_190_195_groupi_n_1952);
  not csa_tree_add_190_195_groupi_drc_bufs47777(csa_tree_add_190_195_groupi_n_1952 ,n_340);
  not csa_tree_add_190_195_groupi_drc_bufs47796(csa_tree_add_190_195_groupi_n_1947 ,csa_tree_add_190_195_groupi_n_1946);
  not csa_tree_add_190_195_groupi_drc_bufs47798(csa_tree_add_190_195_groupi_n_1946 ,n_392);
  not csa_tree_add_190_195_groupi_drc_bufs47821(csa_tree_add_190_195_groupi_n_1940 ,csa_tree_add_190_195_groupi_n_1938);
  not csa_tree_add_190_195_groupi_drc_bufs47822(csa_tree_add_190_195_groupi_n_1939 ,csa_tree_add_190_195_groupi_n_1938);
  not csa_tree_add_190_195_groupi_drc_bufs47823(csa_tree_add_190_195_groupi_n_1938 ,n_456);
  not csa_tree_add_190_195_groupi_drc_bufs47866(csa_tree_add_190_195_groupi_n_1927 ,csa_tree_add_190_195_groupi_n_1925);
  not csa_tree_add_190_195_groupi_drc_bufs47867(csa_tree_add_190_195_groupi_n_1926 ,csa_tree_add_190_195_groupi_n_1925);
  not csa_tree_add_190_195_groupi_drc_bufs47868(csa_tree_add_190_195_groupi_n_1925 ,n_424);
  not csa_tree_add_190_195_groupi_drc_bufs47890(csa_tree_add_190_195_groupi_n_1919 ,csa_tree_add_190_195_groupi_n_1917);
  not csa_tree_add_190_195_groupi_drc_bufs47891(csa_tree_add_190_195_groupi_n_1918 ,csa_tree_add_190_195_groupi_n_1917);
  not csa_tree_add_190_195_groupi_drc_bufs47892(csa_tree_add_190_195_groupi_n_1917 ,n_272);
  not csa_tree_add_190_195_groupi_drc_bufs47902(csa_tree_add_190_195_groupi_n_1914 ,csa_tree_add_190_195_groupi_n_1912);
  not csa_tree_add_190_195_groupi_drc_bufs47903(csa_tree_add_190_195_groupi_n_1913 ,csa_tree_add_190_195_groupi_n_1912);
  not csa_tree_add_190_195_groupi_drc_bufs47904(csa_tree_add_190_195_groupi_n_1912 ,n_238);
  not csa_tree_add_190_195_groupi_drc_bufs47953(csa_tree_add_190_195_groupi_n_2390 ,csa_tree_add_190_195_groupi_n_1901);
  not csa_tree_add_190_195_groupi_drc_bufs47969(csa_tree_add_190_195_groupi_n_2356 ,csa_tree_add_190_195_groupi_n_1897);
  not csa_tree_add_190_195_groupi_drc_bufs47989(csa_tree_add_190_195_groupi_n_2383 ,csa_tree_add_190_195_groupi_n_1892);
  not csa_tree_add_190_195_groupi_drc_bufs48001(csa_tree_add_190_195_groupi_n_2381 ,csa_tree_add_190_195_groupi_n_1889);
  not csa_tree_add_190_195_groupi_drc_bufs48011(csa_tree_add_190_195_groupi_n_1886 ,csa_tree_add_190_195_groupi_n_1884);
  not csa_tree_add_190_195_groupi_drc_bufs48012(csa_tree_add_190_195_groupi_n_1885 ,csa_tree_add_190_195_groupi_n_1884);
  not csa_tree_add_190_195_groupi_drc_bufs48013(csa_tree_add_190_195_groupi_n_1884 ,n_188);
  not csa_tree_add_190_195_groupi_drc_bufs48015(csa_tree_add_190_195_groupi_n_1883 ,csa_tree_add_190_195_groupi_n_1881);
  not csa_tree_add_190_195_groupi_drc_bufs48016(csa_tree_add_190_195_groupi_n_1882 ,csa_tree_add_190_195_groupi_n_1881);
  not csa_tree_add_190_195_groupi_drc_bufs48017(csa_tree_add_190_195_groupi_n_1881 ,n_154);
  not csa_tree_add_190_195_groupi_drc_bufs48019(csa_tree_add_190_195_groupi_n_1880 ,csa_tree_add_190_195_groupi_n_1878);
  not csa_tree_add_190_195_groupi_drc_bufs48020(csa_tree_add_190_195_groupi_n_1879 ,csa_tree_add_190_195_groupi_n_1878);
  not csa_tree_add_190_195_groupi_drc_bufs48021(csa_tree_add_190_195_groupi_n_1878 ,n_290);
  not csa_tree_add_190_195_groupi_drc_bufs48027(csa_tree_add_190_195_groupi_n_1876 ,csa_tree_add_190_195_groupi_n_1874);
  not csa_tree_add_190_195_groupi_drc_bufs48028(csa_tree_add_190_195_groupi_n_1875 ,csa_tree_add_190_195_groupi_n_1874);
  not csa_tree_add_190_195_groupi_drc_bufs48029(csa_tree_add_190_195_groupi_n_1874 ,n_341);
  not csa_tree_add_190_195_groupi_drc_bufs48041(csa_tree_add_190_195_groupi_n_2380 ,csa_tree_add_190_195_groupi_n_1871);
  not csa_tree_add_190_195_groupi_drc_bufs48081(csa_tree_add_190_195_groupi_n_2385 ,csa_tree_add_190_195_groupi_n_1861);
  not csa_tree_add_190_195_groupi_drc_bufs48091(csa_tree_add_190_195_groupi_n_1858 ,csa_tree_add_190_195_groupi_n_1857);
  not csa_tree_add_190_195_groupi_drc_bufs48093(csa_tree_add_190_195_groupi_n_1857 ,n_388);
  not csa_tree_add_190_195_groupi_drc_bufs48106(csa_tree_add_190_195_groupi_n_2392 ,csa_tree_add_190_195_groupi_n_1854);
  not csa_tree_add_190_195_groupi_drc_bufs48292(csa_tree_add_190_195_groupi_n_1807 ,csa_tree_add_190_195_groupi_n_1805);
  not csa_tree_add_190_195_groupi_drc_bufs48293(csa_tree_add_190_195_groupi_n_1806 ,csa_tree_add_190_195_groupi_n_1805);
  not csa_tree_add_190_195_groupi_drc_bufs48294(csa_tree_add_190_195_groupi_n_1805 ,n_201);
  not csa_tree_add_190_195_groupi_drc_bufs48296(csa_tree_add_190_195_groupi_n_1804 ,csa_tree_add_190_195_groupi_n_1802);
  not csa_tree_add_190_195_groupi_drc_bufs48297(csa_tree_add_190_195_groupi_n_1803 ,csa_tree_add_190_195_groupi_n_1802);
  not csa_tree_add_190_195_groupi_drc_bufs48298(csa_tree_add_190_195_groupi_n_1802 ,n_167);
  not csa_tree_add_190_195_groupi_drc_bufs48300(csa_tree_add_190_195_groupi_n_1801 ,csa_tree_add_190_195_groupi_n_1799);
  not csa_tree_add_190_195_groupi_drc_bufs48301(csa_tree_add_190_195_groupi_n_1800 ,csa_tree_add_190_195_groupi_n_1799);
  not csa_tree_add_190_195_groupi_drc_bufs48302(csa_tree_add_190_195_groupi_n_1799 ,n_422);
  not csa_tree_add_190_195_groupi_drc_bufs48304(csa_tree_add_190_195_groupi_n_1798 ,csa_tree_add_190_195_groupi_n_1796);
  not csa_tree_add_190_195_groupi_drc_bufs48305(csa_tree_add_190_195_groupi_n_1797 ,csa_tree_add_190_195_groupi_n_1796);
  not csa_tree_add_190_195_groupi_drc_bufs48306(csa_tree_add_190_195_groupi_n_1796 ,n_150);
  not csa_tree_add_190_195_groupi_drc_bufs48308(csa_tree_add_190_195_groupi_n_1795 ,csa_tree_add_190_195_groupi_n_1793);
  not csa_tree_add_190_195_groupi_drc_bufs48309(csa_tree_add_190_195_groupi_n_1794 ,csa_tree_add_190_195_groupi_n_1793);
  not csa_tree_add_190_195_groupi_drc_bufs48310(csa_tree_add_190_195_groupi_n_1793 ,n_252);
  not csa_tree_add_190_195_groupi_drc_bufs48312(csa_tree_add_190_195_groupi_n_1792 ,csa_tree_add_190_195_groupi_n_1790);
  not csa_tree_add_190_195_groupi_drc_bufs48313(csa_tree_add_190_195_groupi_n_1791 ,csa_tree_add_190_195_groupi_n_1790);
  not csa_tree_add_190_195_groupi_drc_bufs48314(csa_tree_add_190_195_groupi_n_1790 ,n_354);
  not csa_tree_add_190_195_groupi_drc_bufs48316(csa_tree_add_190_195_groupi_n_1789 ,csa_tree_add_190_195_groupi_n_1787);
  not csa_tree_add_190_195_groupi_drc_bufs48317(csa_tree_add_190_195_groupi_n_1788 ,csa_tree_add_190_195_groupi_n_1787);
  not csa_tree_add_190_195_groupi_drc_bufs48318(csa_tree_add_190_195_groupi_n_1787 ,n_405);
  not csa_tree_add_190_195_groupi_drc_bufs48320(csa_tree_add_190_195_groupi_n_1786 ,csa_tree_add_190_195_groupi_n_1784);
  not csa_tree_add_190_195_groupi_drc_bufs48321(csa_tree_add_190_195_groupi_n_1785 ,csa_tree_add_190_195_groupi_n_1784);
  not csa_tree_add_190_195_groupi_drc_bufs48322(csa_tree_add_190_195_groupi_n_1784 ,n_235);
  not csa_tree_add_190_195_groupi_drc_bufs48324(csa_tree_add_190_195_groupi_n_1783 ,csa_tree_add_190_195_groupi_n_1781);
  not csa_tree_add_190_195_groupi_drc_bufs48325(csa_tree_add_190_195_groupi_n_1782 ,csa_tree_add_190_195_groupi_n_1781);
  not csa_tree_add_190_195_groupi_drc_bufs48326(csa_tree_add_190_195_groupi_n_1781 ,n_218);
  not csa_tree_add_190_195_groupi_drc_bufs48334(csa_tree_add_190_195_groupi_n_2353 ,csa_tree_add_190_195_groupi_n_1779);
  not csa_tree_add_190_195_groupi_drc_bufs48338(csa_tree_add_190_195_groupi_n_2389 ,csa_tree_add_190_195_groupi_n_1778);
  not csa_tree_add_190_195_groupi_drc_bufs48356(csa_tree_add_190_195_groupi_n_1773 ,csa_tree_add_190_195_groupi_n_1772);
  not csa_tree_add_190_195_groupi_drc_bufs48358(csa_tree_add_190_195_groupi_n_1772 ,n_270);
  not csa_tree_add_190_195_groupi_drc_bufs48361(csa_tree_add_190_195_groupi_n_1771 ,csa_tree_add_190_195_groupi_n_1770);
  not csa_tree_add_190_195_groupi_drc_bufs48363(csa_tree_add_190_195_groupi_n_1770 ,n_457);
  not csa_tree_add_190_195_groupi_drc_bufs48366(csa_tree_add_190_195_groupi_n_1769 ,csa_tree_add_190_195_groupi_n_1768);
  not csa_tree_add_190_195_groupi_drc_bufs48368(csa_tree_add_190_195_groupi_n_1768 ,n_219);
  not csa_tree_add_190_195_groupi_drc_bufs48377(csa_tree_add_190_195_groupi_n_2391 ,csa_tree_add_190_195_groupi_n_1766);
  not csa_tree_add_190_195_groupi_drc_bufs48413(csa_tree_add_190_195_groupi_n_2357 ,csa_tree_add_190_195_groupi_n_1757);
  not csa_tree_add_190_195_groupi_drc_bufs48483(csa_tree_add_190_195_groupi_n_1741 ,csa_tree_add_190_195_groupi_n_1739);
  not csa_tree_add_190_195_groupi_drc_bufs48484(csa_tree_add_190_195_groupi_n_1740 ,csa_tree_add_190_195_groupi_n_1739);
  not csa_tree_add_190_195_groupi_drc_bufs48485(csa_tree_add_190_195_groupi_n_1739 ,n_202);
  not csa_tree_add_190_195_groupi_drc_bufs48487(csa_tree_add_190_195_groupi_n_1738 ,csa_tree_add_190_195_groupi_n_1736);
  not csa_tree_add_190_195_groupi_drc_bufs48488(csa_tree_add_190_195_groupi_n_1737 ,csa_tree_add_190_195_groupi_n_1736);
  not csa_tree_add_190_195_groupi_drc_bufs48489(csa_tree_add_190_195_groupi_n_1736 ,n_168);
  not csa_tree_add_190_195_groupi_drc_bufs48491(csa_tree_add_190_195_groupi_n_1735 ,csa_tree_add_190_195_groupi_n_1733);
  not csa_tree_add_190_195_groupi_drc_bufs48492(csa_tree_add_190_195_groupi_n_1734 ,csa_tree_add_190_195_groupi_n_1733);
  not csa_tree_add_190_195_groupi_drc_bufs48493(csa_tree_add_190_195_groupi_n_1733 ,n_423);
  not csa_tree_add_190_195_groupi_drc_bufs48495(csa_tree_add_190_195_groupi_n_1732 ,csa_tree_add_190_195_groupi_n_1731);
  not csa_tree_add_190_195_groupi_drc_bufs48497(csa_tree_add_190_195_groupi_n_1731 ,n_151);
  not csa_tree_add_190_195_groupi_drc_bufs48499(csa_tree_add_190_195_groupi_n_1730 ,csa_tree_add_190_195_groupi_n_1728);
  not csa_tree_add_190_195_groupi_drc_bufs48500(csa_tree_add_190_195_groupi_n_1729 ,csa_tree_add_190_195_groupi_n_1728);
  not csa_tree_add_190_195_groupi_drc_bufs48501(csa_tree_add_190_195_groupi_n_1728 ,n_304);
  not csa_tree_add_190_195_groupi_drc_bufs48503(csa_tree_add_190_195_groupi_n_1727 ,csa_tree_add_190_195_groupi_n_1725);
  not csa_tree_add_190_195_groupi_drc_bufs48504(csa_tree_add_190_195_groupi_n_1726 ,csa_tree_add_190_195_groupi_n_1725);
  not csa_tree_add_190_195_groupi_drc_bufs48505(csa_tree_add_190_195_groupi_n_1725 ,n_253);
  not csa_tree_add_190_195_groupi_drc_bufs48507(csa_tree_add_190_195_groupi_n_1724 ,csa_tree_add_190_195_groupi_n_1722);
  not csa_tree_add_190_195_groupi_drc_bufs48508(csa_tree_add_190_195_groupi_n_1723 ,csa_tree_add_190_195_groupi_n_1722);
  not csa_tree_add_190_195_groupi_drc_bufs48509(csa_tree_add_190_195_groupi_n_1722 ,n_355);
  not csa_tree_add_190_195_groupi_drc_bufs48511(csa_tree_add_190_195_groupi_n_1721 ,csa_tree_add_190_195_groupi_n_1719);
  not csa_tree_add_190_195_groupi_drc_bufs48512(csa_tree_add_190_195_groupi_n_1720 ,csa_tree_add_190_195_groupi_n_1719);
  not csa_tree_add_190_195_groupi_drc_bufs48513(csa_tree_add_190_195_groupi_n_1719 ,n_236);
  not csa_tree_add_190_195_groupi_drc_bufs48515(csa_tree_add_190_195_groupi_n_1718 ,csa_tree_add_190_195_groupi_n_1716);
  not csa_tree_add_190_195_groupi_drc_bufs48516(csa_tree_add_190_195_groupi_n_1717 ,csa_tree_add_190_195_groupi_n_1716);
  not csa_tree_add_190_195_groupi_drc_bufs48517(csa_tree_add_190_195_groupi_n_1716 ,n_338);
  not csa_tree_add_190_195_groupi_drc_bufs48523(csa_tree_add_190_195_groupi_n_1714 ,csa_tree_add_190_195_groupi_n_1712);
  not csa_tree_add_190_195_groupi_drc_bufs48524(csa_tree_add_190_195_groupi_n_1713 ,csa_tree_add_190_195_groupi_n_1712);
  not csa_tree_add_190_195_groupi_drc_bufs48525(csa_tree_add_190_195_groupi_n_1712 ,n_269);
  not csa_tree_add_190_195_groupi_drc_bufs48557(csa_tree_add_190_195_groupi_n_2384 ,csa_tree_add_190_195_groupi_n_1704);
  not csa_tree_add_190_195_groupi_drc_bufs48613(csa_tree_add_190_195_groupi_n_2358 ,csa_tree_add_190_195_groupi_n_1690);
  not csa_tree_add_190_195_groupi_drc_bufs48631(csa_tree_add_190_195_groupi_n_1685 ,csa_tree_add_190_195_groupi_n_1683);
  not csa_tree_add_190_195_groupi_drc_bufs48632(csa_tree_add_190_195_groupi_n_1684 ,csa_tree_add_190_195_groupi_n_1683);
  not csa_tree_add_190_195_groupi_drc_bufs48633(csa_tree_add_190_195_groupi_n_1683 ,n_389);
  not csa_tree_add_190_195_groupi_drc_bufs48635(csa_tree_add_190_195_groupi_n_1682 ,csa_tree_add_190_195_groupi_n_1680);
  not csa_tree_add_190_195_groupi_drc_bufs48636(csa_tree_add_190_195_groupi_n_1681 ,csa_tree_add_190_195_groupi_n_1680);
  not csa_tree_add_190_195_groupi_drc_bufs48637(csa_tree_add_190_195_groupi_n_1680 ,n_406);
  not csa_tree_add_190_195_groupi_drc_bufs48653(csa_tree_add_190_195_groupi_n_2378 ,csa_tree_add_190_195_groupi_n_1676);
  not csa_tree_add_190_195_groupi_drc_bufs48671(csa_tree_add_190_195_groupi_n_1671 ,csa_tree_add_190_195_groupi_n_658);
  not csa_tree_add_190_195_groupi_drc_bufs48672(csa_tree_add_190_195_groupi_n_1670 ,csa_tree_add_190_195_groupi_n_658);
  not csa_tree_add_190_195_groupi_drc_bufs48673(csa_tree_add_190_195_groupi_n_1669 ,n_176);
  not csa_tree_add_190_195_groupi_drc_bufs48675(csa_tree_add_190_195_groupi_n_1668 ,csa_tree_add_190_195_groupi_n_644);
  not csa_tree_add_190_195_groupi_drc_bufs48676(csa_tree_add_190_195_groupi_n_1667 ,csa_tree_add_190_195_groupi_n_644);
  not csa_tree_add_190_195_groupi_drc_bufs48677(csa_tree_add_190_195_groupi_n_1666 ,n_261);
  not csa_tree_add_190_195_groupi_drc_bufs48679(csa_tree_add_190_195_groupi_n_1665 ,csa_tree_add_190_195_groupi_n_654);
  not csa_tree_add_190_195_groupi_drc_bufs48680(csa_tree_add_190_195_groupi_n_1664 ,csa_tree_add_190_195_groupi_n_654);
  not csa_tree_add_190_195_groupi_drc_bufs48681(csa_tree_add_190_195_groupi_n_1663 ,n_40);
  not csa_tree_add_190_195_groupi_drc_bufs48683(csa_tree_add_190_195_groupi_n_1662 ,csa_tree_add_190_195_groupi_n_656);
  not csa_tree_add_190_195_groupi_drc_bufs48684(csa_tree_add_190_195_groupi_n_1661 ,csa_tree_add_190_195_groupi_n_656);
  not csa_tree_add_190_195_groupi_drc_bufs48685(csa_tree_add_190_195_groupi_n_1660 ,n_6);
  not csa_tree_add_190_195_groupi_drc_bufs48687(csa_tree_add_190_195_groupi_n_1659 ,csa_tree_add_190_195_groupi_n_642);
  not csa_tree_add_190_195_groupi_drc_bufs48688(csa_tree_add_190_195_groupi_n_1658 ,csa_tree_add_190_195_groupi_n_642);
  not csa_tree_add_190_195_groupi_drc_bufs48689(csa_tree_add_190_195_groupi_n_1657 ,n_186);
  not csa_tree_add_190_195_groupi_drc_bufs48691(csa_tree_add_190_195_groupi_n_1656 ,csa_tree_add_190_195_groupi_n_652);
  not csa_tree_add_190_195_groupi_drc_bufs48692(csa_tree_add_190_195_groupi_n_1655 ,csa_tree_add_190_195_groupi_n_652);
  not csa_tree_add_190_195_groupi_drc_bufs48693(csa_tree_add_190_195_groupi_n_1654 ,n_135);
  not csa_tree_add_190_195_groupi_drc_bufs48695(csa_tree_add_190_195_groupi_n_1653 ,csa_tree_add_190_195_groupi_n_646);
  not csa_tree_add_190_195_groupi_drc_bufs48696(csa_tree_add_190_195_groupi_n_1652 ,csa_tree_add_190_195_groupi_n_646);
  not csa_tree_add_190_195_groupi_drc_bufs48697(csa_tree_add_190_195_groupi_n_1651 ,n_101);
  not csa_tree_add_190_195_groupi_drc_bufs48699(csa_tree_add_190_195_groupi_n_1650 ,csa_tree_add_190_195_groupi_n_650);
  not csa_tree_add_190_195_groupi_drc_bufs48700(csa_tree_add_190_195_groupi_n_1649 ,csa_tree_add_190_195_groupi_n_650);
  not csa_tree_add_190_195_groupi_drc_bufs48701(csa_tree_add_190_195_groupi_n_1648 ,n_50);
  not csa_tree_add_190_195_groupi_drc_bufs48703(csa_tree_add_190_195_groupi_n_1647 ,csa_tree_add_190_195_groupi_n_648);
  not csa_tree_add_190_195_groupi_drc_bufs48704(csa_tree_add_190_195_groupi_n_1646 ,csa_tree_add_190_195_groupi_n_648);
  not csa_tree_add_190_195_groupi_drc_bufs48705(csa_tree_add_190_195_groupi_n_1645 ,n_33);
  not csa_tree_add_190_195_groupi_drc_bufs48707(csa_tree_add_190_195_groupi_n_1644 ,csa_tree_add_190_195_groupi_n_640);
  not csa_tree_add_190_195_groupi_drc_bufs48708(csa_tree_add_190_195_groupi_n_1643 ,csa_tree_add_190_195_groupi_n_640);
  not csa_tree_add_190_195_groupi_drc_bufs48709(csa_tree_add_190_195_groupi_n_1642 ,n_16);
  not csa_tree_add_190_195_groupi_drc_bufs48711(csa_tree_add_190_195_groupi_n_1641 ,csa_tree_add_190_195_groupi_n_638);
  not csa_tree_add_190_195_groupi_drc_bufs48712(csa_tree_add_190_195_groupi_n_1640 ,csa_tree_add_190_195_groupi_n_638);
  not csa_tree_add_190_195_groupi_drc_bufs48713(csa_tree_add_190_195_groupi_n_1639 ,n_187);
  not csa_tree_add_190_195_groupi_drc_bufs48715(csa_tree_add_190_195_groupi_n_1638 ,csa_tree_add_190_195_groupi_n_1636);
  not csa_tree_add_190_195_groupi_drc_bufs48716(csa_tree_add_190_195_groupi_n_1637 ,csa_tree_add_190_195_groupi_n_1636);
  not csa_tree_add_190_195_groupi_drc_bufs48717(csa_tree_add_190_195_groupi_n_1636 ,n_391);
  not csa_tree_add_190_195_groupi_drc_bufs48719(csa_tree_add_190_195_groupi_n_1635 ,csa_tree_add_190_195_groupi_n_630);
  not csa_tree_add_190_195_groupi_drc_bufs48721(csa_tree_add_190_195_groupi_n_1634 ,n_119);
  not csa_tree_add_190_195_groupi_drc_bufs48723(csa_tree_add_190_195_groupi_n_1633 ,csa_tree_add_190_195_groupi_n_636);
  not csa_tree_add_190_195_groupi_drc_bufs48724(csa_tree_add_190_195_groupi_n_1632 ,csa_tree_add_190_195_groupi_n_636);
  not csa_tree_add_190_195_groupi_drc_bufs48725(csa_tree_add_190_195_groupi_n_1631 ,n_102);
  not csa_tree_add_190_195_groupi_drc_bufs48727(csa_tree_add_190_195_groupi_n_1630 ,csa_tree_add_190_195_groupi_n_632);
  not csa_tree_add_190_195_groupi_drc_bufs48728(csa_tree_add_190_195_groupi_n_1629 ,csa_tree_add_190_195_groupi_n_632);
  not csa_tree_add_190_195_groupi_drc_bufs48729(csa_tree_add_190_195_groupi_n_1628 ,n_34);
  not csa_tree_add_190_195_groupi_drc_bufs48731(csa_tree_add_190_195_groupi_n_1627 ,csa_tree_add_190_195_groupi_n_634);
  not csa_tree_add_190_195_groupi_drc_bufs48732(csa_tree_add_190_195_groupi_n_1626 ,csa_tree_add_190_195_groupi_n_634);
  not csa_tree_add_190_195_groupi_drc_bufs48733(csa_tree_add_190_195_groupi_n_1625 ,n_17);
  not csa_tree_add_190_195_groupi_drc_bufs48739(csa_tree_add_190_195_groupi_n_1624 ,csa_tree_add_190_195_groupi_n_1622);
  not csa_tree_add_190_195_groupi_drc_bufs48740(csa_tree_add_190_195_groupi_n_1623 ,csa_tree_add_190_195_groupi_n_1622);
  not csa_tree_add_190_195_groupi_drc_bufs48741(csa_tree_add_190_195_groupi_n_1622 ,n_120);
  not csa_tree_add_190_195_groupi_drc_bufs48743(csa_tree_add_190_195_groupi_n_1621 ,csa_tree_add_190_195_groupi_n_1619);
  not csa_tree_add_190_195_groupi_drc_bufs48744(csa_tree_add_190_195_groupi_n_1620 ,csa_tree_add_190_195_groupi_n_1619);
  not csa_tree_add_190_195_groupi_drc_bufs48745(csa_tree_add_190_195_groupi_n_1619 ,n_86);
  not csa_tree_add_190_195_groupi_drc_bufs48747(csa_tree_add_190_195_groupi_n_1618 ,csa_tree_add_190_195_groupi_n_1616);
  not csa_tree_add_190_195_groupi_drc_bufs48748(csa_tree_add_190_195_groupi_n_1617 ,csa_tree_add_190_195_groupi_n_1616);
  not csa_tree_add_190_195_groupi_drc_bufs48749(csa_tree_add_190_195_groupi_n_1616 ,n_52);
  not csa_tree_add_190_195_groupi_drc_bufs48751(csa_tree_add_190_195_groupi_n_1615 ,csa_tree_add_190_195_groupi_n_1613);
  not csa_tree_add_190_195_groupi_drc_bufs48752(csa_tree_add_190_195_groupi_n_1614 ,csa_tree_add_190_195_groupi_n_1613);
  not csa_tree_add_190_195_groupi_drc_bufs48753(csa_tree_add_190_195_groupi_n_1613 ,n_409);
  not csa_tree_add_190_195_groupi_drc_bufs48755(csa_tree_add_190_195_groupi_n_1612 ,csa_tree_add_190_195_groupi_n_1610);
  not csa_tree_add_190_195_groupi_drc_bufs48756(csa_tree_add_190_195_groupi_n_1611 ,csa_tree_add_190_195_groupi_n_1610);
  not csa_tree_add_190_195_groupi_drc_bufs48757(csa_tree_add_190_195_groupi_n_1610 ,n_1);
  not csa_tree_add_190_195_groupi_drc_bufs48785(csa_tree_add_190_195_groupi_n_2348 ,csa_tree_add_190_195_groupi_n_1605);
  not csa_tree_add_190_195_groupi_drc_bufs48797(csa_tree_add_190_195_groupi_n_2352 ,csa_tree_add_190_195_groupi_n_1602);
  not csa_tree_add_190_195_groupi_drc_bufs48811(csa_tree_add_190_195_groupi_n_1601 ,csa_tree_add_190_195_groupi_n_1599);
  not csa_tree_add_190_195_groupi_drc_bufs48812(csa_tree_add_190_195_groupi_n_1600 ,csa_tree_add_190_195_groupi_n_1599);
  not csa_tree_add_190_195_groupi_drc_bufs48813(csa_tree_add_190_195_groupi_n_1599 ,n_116);
  not csa_tree_add_190_195_groupi_drc_bufs48815(csa_tree_add_190_195_groupi_n_1598 ,csa_tree_add_190_195_groupi_n_1596);
  not csa_tree_add_190_195_groupi_drc_bufs48816(csa_tree_add_190_195_groupi_n_1597 ,csa_tree_add_190_195_groupi_n_1596);
  not csa_tree_add_190_195_groupi_drc_bufs48817(csa_tree_add_190_195_groupi_n_1596 ,n_99);
  not csa_tree_add_190_195_groupi_drc_bufs48819(csa_tree_add_190_195_groupi_n_1595 ,csa_tree_add_190_195_groupi_n_1593);
  not csa_tree_add_190_195_groupi_drc_bufs48820(csa_tree_add_190_195_groupi_n_1594 ,csa_tree_add_190_195_groupi_n_1593);
  not csa_tree_add_190_195_groupi_drc_bufs48821(csa_tree_add_190_195_groupi_n_1593 ,n_48);
  not csa_tree_add_190_195_groupi_drc_bufs48823(csa_tree_add_190_195_groupi_n_1592 ,csa_tree_add_190_195_groupi_n_1590);
  not csa_tree_add_190_195_groupi_drc_bufs48824(csa_tree_add_190_195_groupi_n_1591 ,csa_tree_add_190_195_groupi_n_1590);
  not csa_tree_add_190_195_groupi_drc_bufs48825(csa_tree_add_190_195_groupi_n_1590 ,n_31);
  not csa_tree_add_190_195_groupi_drc_bufs48827(csa_tree_add_190_195_groupi_n_1589 ,csa_tree_add_190_195_groupi_n_1587);
  not csa_tree_add_190_195_groupi_drc_bufs48828(csa_tree_add_190_195_groupi_n_1588 ,csa_tree_add_190_195_groupi_n_1587);
  not csa_tree_add_190_195_groupi_drc_bufs48829(csa_tree_add_190_195_groupi_n_1587 ,n_14);
  not csa_tree_add_190_195_groupi_drc_bufs48839(csa_tree_add_190_195_groupi_n_1584 ,csa_tree_add_190_195_groupi_n_1582);
  not csa_tree_add_190_195_groupi_drc_bufs48840(csa_tree_add_190_195_groupi_n_1583 ,csa_tree_add_190_195_groupi_n_1582);
  not csa_tree_add_190_195_groupi_drc_bufs48841(csa_tree_add_190_195_groupi_n_1582 ,n_185);
  not csa_tree_add_190_195_groupi_drc_bufs48843(csa_tree_add_190_195_groupi_n_1581 ,csa_tree_add_190_195_groupi_n_1579);
  not csa_tree_add_190_195_groupi_drc_bufs48844(csa_tree_add_190_195_groupi_n_1580 ,csa_tree_add_190_195_groupi_n_1579);
  not csa_tree_add_190_195_groupi_drc_bufs48845(csa_tree_add_190_195_groupi_n_1579 ,n_66);
  not csa_tree_add_190_195_groupi_drc_bufs48847(csa_tree_add_190_195_groupi_n_1578 ,csa_tree_add_190_195_groupi_n_1576);
  not csa_tree_add_190_195_groupi_drc_bufs48848(csa_tree_add_190_195_groupi_n_1577 ,csa_tree_add_190_195_groupi_n_1576);
  not csa_tree_add_190_195_groupi_drc_bufs48849(csa_tree_add_190_195_groupi_n_1576 ,n_32);
  not csa_tree_add_190_195_groupi_drc_bufs48851(csa_tree_add_190_195_groupi_n_1575 ,csa_tree_add_190_195_groupi_n_1573);
  not csa_tree_add_190_195_groupi_drc_bufs48852(csa_tree_add_190_195_groupi_n_1574 ,csa_tree_add_190_195_groupi_n_1573);
  not csa_tree_add_190_195_groupi_drc_bufs48853(csa_tree_add_190_195_groupi_n_1573 ,n_15);
  not csa_tree_add_190_195_groupi_drc_bufs48863(csa_tree_add_190_195_groupi_n_1570 ,csa_tree_add_190_195_groupi_n_1569);
  not csa_tree_add_190_195_groupi_drc_bufs48865(csa_tree_add_190_195_groupi_n_1569 ,csa_tree_add_190_195_groupi_n_2584);
  not csa_tree_add_190_195_groupi_drc_bufs48868(csa_tree_add_190_195_groupi_n_1568 ,csa_tree_add_190_195_groupi_n_1567);
  not csa_tree_add_190_195_groupi_drc_bufs48869(csa_tree_add_190_195_groupi_n_1567 ,csa_tree_add_190_195_groupi_n_2409);
  not csa_tree_add_190_195_groupi_drc_bufs48872(csa_tree_add_190_195_groupi_n_1566 ,csa_tree_add_190_195_groupi_n_1565);
  not csa_tree_add_190_195_groupi_drc_bufs48873(csa_tree_add_190_195_groupi_n_1565 ,csa_tree_add_190_195_groupi_n_2637);
  not csa_tree_add_190_195_groupi_drc_bufs48876(csa_tree_add_190_195_groupi_n_1564 ,csa_tree_add_190_195_groupi_n_1563);
  not csa_tree_add_190_195_groupi_drc_bufs48877(csa_tree_add_190_195_groupi_n_1563 ,csa_tree_add_190_195_groupi_n_2581);
  not csa_tree_add_190_195_groupi_drc_bufs48880(csa_tree_add_190_195_groupi_n_1562 ,csa_tree_add_190_195_groupi_n_1561);
  not csa_tree_add_190_195_groupi_drc_bufs48881(csa_tree_add_190_195_groupi_n_1561 ,csa_tree_add_190_195_groupi_n_2586);
  not csa_tree_add_190_195_groupi_drc_bufs48887(csa_tree_add_190_195_groupi_n_1560 ,csa_tree_add_190_195_groupi_n_1558);
  not csa_tree_add_190_195_groupi_drc_bufs48888(csa_tree_add_190_195_groupi_n_1559 ,csa_tree_add_190_195_groupi_n_1558);
  not csa_tree_add_190_195_groupi_drc_bufs48889(csa_tree_add_190_195_groupi_n_1558 ,csa_tree_add_190_195_groupi_n_2361);
  not csa_tree_add_190_195_groupi_drc_bufs48891(csa_tree_add_190_195_groupi_n_1557 ,csa_tree_add_190_195_groupi_n_1555);
  not csa_tree_add_190_195_groupi_drc_bufs48892(csa_tree_add_190_195_groupi_n_1556 ,csa_tree_add_190_195_groupi_n_1555);
  not csa_tree_add_190_195_groupi_drc_bufs48893(csa_tree_add_190_195_groupi_n_1555 ,csa_tree_add_190_195_groupi_n_2333);
  not csa_tree_add_190_195_groupi_drc_bufs48895(csa_tree_add_190_195_groupi_n_1554 ,csa_tree_add_190_195_groupi_n_1553);
  not csa_tree_add_190_195_groupi_drc_bufs48897(csa_tree_add_190_195_groupi_n_1553 ,csa_tree_add_190_195_groupi_n_2583);
  not csa_tree_add_190_195_groupi_drc_bufs48899(csa_tree_add_190_195_groupi_n_1552 ,csa_tree_add_190_195_groupi_n_1551);
  not csa_tree_add_190_195_groupi_drc_bufs48901(csa_tree_add_190_195_groupi_n_1551 ,csa_tree_add_190_195_groupi_n_2579);
  not csa_tree_add_190_195_groupi_drc_bufs48907(csa_tree_add_190_195_groupi_n_1549 ,csa_tree_add_190_195_groupi_n_1547);
  not csa_tree_add_190_195_groupi_drc_bufs48908(csa_tree_add_190_195_groupi_n_1548 ,csa_tree_add_190_195_groupi_n_1547);
  not csa_tree_add_190_195_groupi_drc_bufs48909(csa_tree_add_190_195_groupi_n_1547 ,csa_tree_add_190_195_groupi_n_2362);
  not csa_tree_add_190_195_groupi_drc_bufs48911(csa_tree_add_190_195_groupi_n_1546 ,csa_tree_add_190_195_groupi_n_1544);
  not csa_tree_add_190_195_groupi_drc_bufs48912(csa_tree_add_190_195_groupi_n_1545 ,csa_tree_add_190_195_groupi_n_1544);
  not csa_tree_add_190_195_groupi_drc_bufs48913(csa_tree_add_190_195_groupi_n_1544 ,csa_tree_add_190_195_groupi_n_2335);
  not csa_tree_add_190_195_groupi_drc_bufs48915(csa_tree_add_190_195_groupi_n_1543 ,csa_tree_add_190_195_groupi_n_1542);
  not csa_tree_add_190_195_groupi_drc_bufs48917(csa_tree_add_190_195_groupi_n_1542 ,n_83);
  not csa_tree_add_190_195_groupi_drc_bufs48927(csa_tree_add_190_195_groupi_n_1541 ,csa_tree_add_190_195_groupi_n_1540);
  not csa_tree_add_190_195_groupi_drc_bufs48929(csa_tree_add_190_195_groupi_n_1540 ,csa_tree_add_190_195_groupi_n_2417);
  not csa_tree_add_190_195_groupi_drc_bufs48931(csa_tree_add_190_195_groupi_n_1539 ,csa_tree_add_190_195_groupi_n_1538);
  not csa_tree_add_190_195_groupi_drc_bufs48933(csa_tree_add_190_195_groupi_n_1538 ,csa_tree_add_190_195_groupi_n_2416);
  not csa_tree_add_190_195_groupi_drc_bufs48936(csa_tree_add_190_195_groupi_n_1537 ,csa_tree_add_190_195_groupi_n_1536);
  not csa_tree_add_190_195_groupi_drc_bufs48937(csa_tree_add_190_195_groupi_n_1536 ,csa_tree_add_190_195_groupi_n_2588);
  not csa_tree_add_190_195_groupi_drc_bufs48943(csa_tree_add_190_195_groupi_n_1535 ,csa_tree_add_190_195_groupi_n_1534);
  not csa_tree_add_190_195_groupi_drc_bufs48945(csa_tree_add_190_195_groupi_n_1534 ,csa_tree_add_190_195_groupi_n_2644);
  not csa_tree_add_190_195_groupi_drc_bufs48947(csa_tree_add_190_195_groupi_n_1533 ,csa_tree_add_190_195_groupi_n_1532);
  not csa_tree_add_190_195_groupi_drc_bufs48949(csa_tree_add_190_195_groupi_n_1532 ,csa_tree_add_190_195_groupi_n_2598);
  not csa_tree_add_190_195_groupi_drc_bufs48951(csa_tree_add_190_195_groupi_n_1531 ,csa_tree_add_190_195_groupi_n_1529);
  not csa_tree_add_190_195_groupi_drc_bufs48952(csa_tree_add_190_195_groupi_n_1530 ,csa_tree_add_190_195_groupi_n_1529);
  not csa_tree_add_190_195_groupi_drc_bufs48953(csa_tree_add_190_195_groupi_n_1529 ,csa_tree_add_190_195_groupi_n_2580);
  not csa_tree_add_190_195_groupi_drc_bufs48956(csa_tree_add_190_195_groupi_n_1528 ,csa_tree_add_190_195_groupi_n_1527);
  not csa_tree_add_190_195_groupi_drc_bufs48957(csa_tree_add_190_195_groupi_n_1527 ,csa_tree_add_190_195_groupi_n_2473);
  not csa_tree_add_190_195_groupi_drc_bufs48959(csa_tree_add_190_195_groupi_n_1526 ,csa_tree_add_190_195_groupi_n_1524);
  not csa_tree_add_190_195_groupi_drc_bufs48960(csa_tree_add_190_195_groupi_n_1525 ,csa_tree_add_190_195_groupi_n_1524);
  not csa_tree_add_190_195_groupi_drc_bufs48961(csa_tree_add_190_195_groupi_n_1524 ,csa_tree_add_190_195_groupi_n_2414);
  not csa_tree_add_190_195_groupi_drc_bufs48963(csa_tree_add_190_195_groupi_n_1523 ,csa_tree_add_190_195_groupi_n_1521);
  not csa_tree_add_190_195_groupi_drc_bufs48964(csa_tree_add_190_195_groupi_n_1522 ,csa_tree_add_190_195_groupi_n_1521);
  not csa_tree_add_190_195_groupi_drc_bufs48965(csa_tree_add_190_195_groupi_n_1521 ,csa_tree_add_190_195_groupi_n_2597);
  not csa_tree_add_190_195_groupi_drc_bufs48967(csa_tree_add_190_195_groupi_n_1520 ,csa_tree_add_190_195_groupi_n_1518);
  not csa_tree_add_190_195_groupi_drc_bufs48968(csa_tree_add_190_195_groupi_n_1519 ,csa_tree_add_190_195_groupi_n_1518);
  not csa_tree_add_190_195_groupi_drc_bufs48969(csa_tree_add_190_195_groupi_n_1518 ,csa_tree_add_190_195_groupi_n_2433);
  not csa_tree_add_190_195_groupi_drc_bufs48971(csa_tree_add_190_195_groupi_n_1517 ,csa_tree_add_190_195_groupi_n_1515);
  not csa_tree_add_190_195_groupi_drc_bufs48972(csa_tree_add_190_195_groupi_n_1516 ,csa_tree_add_190_195_groupi_n_1515);
  not csa_tree_add_190_195_groupi_drc_bufs48973(csa_tree_add_190_195_groupi_n_1515 ,csa_tree_add_190_195_groupi_n_2574);
  not csa_tree_add_190_195_groupi_drc_bufs48975(csa_tree_add_190_195_groupi_n_1514 ,csa_tree_add_190_195_groupi_n_1512);
  not csa_tree_add_190_195_groupi_drc_bufs48976(csa_tree_add_190_195_groupi_n_1513 ,csa_tree_add_190_195_groupi_n_1512);
  not csa_tree_add_190_195_groupi_drc_bufs48977(csa_tree_add_190_195_groupi_n_1512 ,csa_tree_add_190_195_groupi_n_2329);
  not csa_tree_add_190_195_groupi_drc_bufs48979(csa_tree_add_190_195_groupi_n_1511 ,csa_tree_add_190_195_groupi_n_1509);
  not csa_tree_add_190_195_groupi_drc_bufs48980(csa_tree_add_190_195_groupi_n_1510 ,csa_tree_add_190_195_groupi_n_1509);
  not csa_tree_add_190_195_groupi_drc_bufs48981(csa_tree_add_190_195_groupi_n_1509 ,csa_tree_add_190_195_groupi_n_2363);
  not csa_tree_add_190_195_groupi_drc_bufs48984(csa_tree_add_190_195_groupi_n_1508 ,csa_tree_add_190_195_groupi_n_1507);
  not csa_tree_add_190_195_groupi_drc_bufs48985(csa_tree_add_190_195_groupi_n_1507 ,csa_tree_add_190_195_groupi_n_2488);
  not csa_tree_add_190_195_groupi_drc_bufs48987(csa_tree_add_190_195_groupi_n_1506 ,csa_tree_add_190_195_groupi_n_1504);
  not csa_tree_add_190_195_groupi_drc_bufs48988(csa_tree_add_190_195_groupi_n_1505 ,csa_tree_add_190_195_groupi_n_1504);
  not csa_tree_add_190_195_groupi_drc_bufs48989(csa_tree_add_190_195_groupi_n_1504 ,csa_tree_add_190_195_groupi_n_2331);
  not csa_tree_add_190_195_groupi_drc_bufs48992(csa_tree_add_190_195_groupi_n_1503 ,csa_tree_add_190_195_groupi_n_1502);
  not csa_tree_add_190_195_groupi_drc_bufs48993(csa_tree_add_190_195_groupi_n_1502 ,csa_tree_add_190_195_groupi_n_2460);
  not csa_tree_add_190_195_groupi_drc_bufs48995(csa_tree_add_190_195_groupi_n_1501 ,csa_tree_add_190_195_groupi_n_1500);
  not csa_tree_add_190_195_groupi_drc_bufs48997(csa_tree_add_190_195_groupi_n_1500 ,csa_tree_add_190_195_groupi_n_2437);
  not csa_tree_add_190_195_groupi_drc_bufs48999(csa_tree_add_190_195_groupi_n_1499 ,csa_tree_add_190_195_groupi_n_1497);
  not csa_tree_add_190_195_groupi_drc_bufs49000(csa_tree_add_190_195_groupi_n_1498 ,csa_tree_add_190_195_groupi_n_1497);
  not csa_tree_add_190_195_groupi_drc_bufs49001(csa_tree_add_190_195_groupi_n_1497 ,csa_tree_add_190_195_groupi_n_2360);
  not csa_tree_add_190_195_groupi_drc_bufs49003(csa_tree_add_190_195_groupi_n_1496 ,csa_tree_add_190_195_groupi_n_1494);
  not csa_tree_add_190_195_groupi_drc_bufs49004(csa_tree_add_190_195_groupi_n_1495 ,csa_tree_add_190_195_groupi_n_1494);
  not csa_tree_add_190_195_groupi_drc_bufs49005(csa_tree_add_190_195_groupi_n_1494 ,csa_tree_add_190_195_groupi_n_2328);
  not csa_tree_add_190_195_groupi_drc_bufs49008(csa_tree_add_190_195_groupi_n_1493 ,csa_tree_add_190_195_groupi_n_1492);
  not csa_tree_add_190_195_groupi_drc_bufs49009(csa_tree_add_190_195_groupi_n_1492 ,csa_tree_add_190_195_groupi_n_2650);
  not csa_tree_add_190_195_groupi_drc_bufs49011(csa_tree_add_190_195_groupi_n_1491 ,csa_tree_add_190_195_groupi_n_1489);
  not csa_tree_add_190_195_groupi_drc_bufs49012(csa_tree_add_190_195_groupi_n_1490 ,csa_tree_add_190_195_groupi_n_1489);
  not csa_tree_add_190_195_groupi_drc_bufs49013(csa_tree_add_190_195_groupi_n_1489 ,csa_tree_add_190_195_groupi_n_2334);
  not csa_tree_add_190_195_groupi_drc_bufs49015(csa_tree_add_190_195_groupi_n_1488 ,csa_tree_add_190_195_groupi_n_1486);
  not csa_tree_add_190_195_groupi_drc_bufs49016(csa_tree_add_190_195_groupi_n_1487 ,csa_tree_add_190_195_groupi_n_1486);
  not csa_tree_add_190_195_groupi_drc_bufs49017(csa_tree_add_190_195_groupi_n_1486 ,csa_tree_add_190_195_groupi_n_2422);
  not csa_tree_add_190_195_groupi_drc_bufs49019(csa_tree_add_190_195_groupi_n_1485 ,csa_tree_add_190_195_groupi_n_1483);
  not csa_tree_add_190_195_groupi_drc_bufs49020(csa_tree_add_190_195_groupi_n_1484 ,csa_tree_add_190_195_groupi_n_1483);
  not csa_tree_add_190_195_groupi_drc_bufs49021(csa_tree_add_190_195_groupi_n_1483 ,csa_tree_add_190_195_groupi_n_2332);
  not csa_tree_add_190_195_groupi_drc_bufs49024(csa_tree_add_190_195_groupi_n_1482 ,csa_tree_add_190_195_groupi_n_1481);
  not csa_tree_add_190_195_groupi_drc_bufs49025(csa_tree_add_190_195_groupi_n_1481 ,csa_tree_add_190_195_groupi_n_2659);
  not csa_tree_add_190_195_groupi_drc_bufs49028(csa_tree_add_190_195_groupi_n_1480 ,csa_tree_add_190_195_groupi_n_1479);
  not csa_tree_add_190_195_groupi_drc_bufs49029(csa_tree_add_190_195_groupi_n_1479 ,csa_tree_add_190_195_groupi_n_2634);
  not csa_tree_add_190_195_groupi_drc_bufs49031(csa_tree_add_190_195_groupi_n_1478 ,csa_tree_add_190_195_groupi_n_1476);
  not csa_tree_add_190_195_groupi_drc_bufs49032(csa_tree_add_190_195_groupi_n_1477 ,csa_tree_add_190_195_groupi_n_1476);
  not csa_tree_add_190_195_groupi_drc_bufs49033(csa_tree_add_190_195_groupi_n_1476 ,csa_tree_add_190_195_groupi_n_2359);
  not csa_tree_add_190_195_groupi_drc_bufs49035(csa_tree_add_190_195_groupi_n_1475 ,csa_tree_add_190_195_groupi_n_1473);
  not csa_tree_add_190_195_groupi_drc_bufs49036(csa_tree_add_190_195_groupi_n_1474 ,csa_tree_add_190_195_groupi_n_1473);
  not csa_tree_add_190_195_groupi_drc_bufs49037(csa_tree_add_190_195_groupi_n_1473 ,csa_tree_add_190_195_groupi_n_2330);
  not csa_tree_add_190_195_groupi_drc_bufs49039(csa_tree_add_190_195_groupi_n_1472 ,csa_tree_add_190_195_groupi_n_1470);
  not csa_tree_add_190_195_groupi_drc_bufs49040(csa_tree_add_190_195_groupi_n_1471 ,csa_tree_add_190_195_groupi_n_1470);
  not csa_tree_add_190_195_groupi_drc_bufs49041(csa_tree_add_190_195_groupi_n_1470 ,csa_tree_add_190_195_groupi_n_2365);
  not csa_tree_add_190_195_groupi_drc_bufs49043(csa_tree_add_190_195_groupi_n_1469 ,csa_tree_add_190_195_groupi_n_1467);
  not csa_tree_add_190_195_groupi_drc_bufs49044(csa_tree_add_190_195_groupi_n_1468 ,csa_tree_add_190_195_groupi_n_1467);
  not csa_tree_add_190_195_groupi_drc_bufs49045(csa_tree_add_190_195_groupi_n_1467 ,csa_tree_add_190_195_groupi_n_2427);
  not csa_tree_add_190_195_groupi_drc_bufs49048(csa_tree_add_190_195_groupi_n_1466 ,csa_tree_add_190_195_groupi_n_1465);
  not csa_tree_add_190_195_groupi_drc_bufs49049(csa_tree_add_190_195_groupi_n_1465 ,csa_tree_add_190_195_groupi_n_2495);
  not csa_tree_add_190_195_groupi_drc_bufs49052(csa_tree_add_190_195_groupi_n_1464 ,csa_tree_add_190_195_groupi_n_1463);
  not csa_tree_add_190_195_groupi_drc_bufs49053(csa_tree_add_190_195_groupi_n_1463 ,csa_tree_add_190_195_groupi_n_2652);
  not csa_tree_add_190_195_groupi_drc_bufs49056(csa_tree_add_190_195_groupi_n_1462 ,csa_tree_add_190_195_groupi_n_1461);
  not csa_tree_add_190_195_groupi_drc_bufs49057(csa_tree_add_190_195_groupi_n_1461 ,csa_tree_add_190_195_groupi_n_2435);
  not csa_tree_add_190_195_groupi_drc_bufs49060(csa_tree_add_190_195_groupi_n_1460 ,csa_tree_add_190_195_groupi_n_1459);
  not csa_tree_add_190_195_groupi_drc_bufs49061(csa_tree_add_190_195_groupi_n_1459 ,csa_tree_add_190_195_groupi_n_2503);
  not csa_tree_add_190_195_groupi_drc_bufs49064(csa_tree_add_190_195_groupi_n_1458 ,csa_tree_add_190_195_groupi_n_1457);
  not csa_tree_add_190_195_groupi_drc_bufs49065(csa_tree_add_190_195_groupi_n_1457 ,csa_tree_add_190_195_groupi_n_2647);
  not csa_tree_add_190_195_groupi_drc_bufs49067(csa_tree_add_190_195_groupi_n_1456 ,csa_tree_add_190_195_groupi_n_1454);
  not csa_tree_add_190_195_groupi_drc_bufs49068(csa_tree_add_190_195_groupi_n_1455 ,csa_tree_add_190_195_groupi_n_1454);
  not csa_tree_add_190_195_groupi_drc_bufs49069(csa_tree_add_190_195_groupi_n_1454 ,csa_tree_add_190_195_groupi_n_2421);
  not csa_tree_add_190_195_groupi_drc_bufs49071(csa_tree_add_190_195_groupi_n_1453 ,csa_tree_add_190_195_groupi_n_1451);
  not csa_tree_add_190_195_groupi_drc_bufs49072(csa_tree_add_190_195_groupi_n_1452 ,csa_tree_add_190_195_groupi_n_1451);
  not csa_tree_add_190_195_groupi_drc_bufs49073(csa_tree_add_190_195_groupi_n_1451 ,csa_tree_add_190_195_groupi_n_2336);
  not csa_tree_add_190_195_groupi_drc_bufs49075(csa_tree_add_190_195_groupi_n_1450 ,csa_tree_add_190_195_groupi_n_1448);
  not csa_tree_add_190_195_groupi_drc_bufs49076(csa_tree_add_190_195_groupi_n_1449 ,csa_tree_add_190_195_groupi_n_1448);
  not csa_tree_add_190_195_groupi_drc_bufs49077(csa_tree_add_190_195_groupi_n_1448 ,csa_tree_add_190_195_groupi_n_2337);
  not csa_tree_add_190_195_groupi_drc_bufs49079(csa_tree_add_190_195_groupi_n_1447 ,csa_tree_add_190_195_groupi_n_1445);
  not csa_tree_add_190_195_groupi_drc_bufs49080(csa_tree_add_190_195_groupi_n_1446 ,csa_tree_add_190_195_groupi_n_1445);
  not csa_tree_add_190_195_groupi_drc_bufs49081(csa_tree_add_190_195_groupi_n_1445 ,csa_tree_add_190_195_groupi_n_2338);
  not csa_tree_add_190_195_groupi_drc_bufs49087(csa_tree_add_190_195_groupi_n_1444 ,csa_tree_add_190_195_groupi_n_1443);
  not csa_tree_add_190_195_groupi_drc_bufs49089(csa_tree_add_190_195_groupi_n_1443 ,csa_tree_add_190_195_groupi_n_2412);
  not csa_tree_add_190_195_groupi_drc_bufs49091(csa_tree_add_190_195_groupi_n_1442 ,csa_tree_add_190_195_groupi_n_1441);
  not csa_tree_add_190_195_groupi_drc_bufs49093(csa_tree_add_190_195_groupi_n_1441 ,csa_tree_add_190_195_groupi_n_2604);
  not csa_tree_add_190_195_groupi_drc_bufs49095(csa_tree_add_190_195_groupi_n_1440 ,csa_tree_add_190_195_groupi_n_1439);
  not csa_tree_add_190_195_groupi_drc_bufs49097(csa_tree_add_190_195_groupi_n_1439 ,csa_tree_add_190_195_groupi_n_2587);
  not csa_tree_add_190_195_groupi_drc_bufs49103(csa_tree_add_190_195_groupi_n_1438 ,csa_tree_add_190_195_groupi_n_1437);
  not csa_tree_add_190_195_groupi_drc_bufs49105(csa_tree_add_190_195_groupi_n_1437 ,csa_tree_add_190_195_groupi_n_2441);
  not csa_tree_add_190_195_groupi_drc_bufs49107(csa_tree_add_190_195_groupi_n_1436 ,csa_tree_add_190_195_groupi_n_1435);
  not csa_tree_add_190_195_groupi_drc_bufs49109(csa_tree_add_190_195_groupi_n_1435 ,csa_tree_add_190_195_groupi_n_2406);
  not csa_tree_add_190_195_groupi_drc_bufs49123(csa_tree_add_190_195_groupi_n_1434 ,csa_tree_add_190_195_groupi_n_1433);
  not csa_tree_add_190_195_groupi_drc_bufs49125(csa_tree_add_190_195_groupi_n_1433 ,csa_tree_add_190_195_groupi_n_2492);
  not csa_tree_add_190_195_groupi_drc_bufs49127(csa_tree_add_190_195_groupi_n_1432 ,csa_tree_add_190_195_groupi_n_1431);
  not csa_tree_add_190_195_groupi_drc_bufs49129(csa_tree_add_190_195_groupi_n_1431 ,csa_tree_add_190_195_groupi_n_2582);
  not csa_tree_add_190_195_groupi_drc_bufs49139(csa_tree_add_190_195_groupi_n_1430 ,csa_tree_add_190_195_groupi_n_1429);
  not csa_tree_add_190_195_groupi_drc_bufs49141(csa_tree_add_190_195_groupi_n_1429 ,csa_tree_add_190_195_groupi_n_2622);
  not csa_tree_add_190_195_groupi_drc_bufs49147(csa_tree_add_190_195_groupi_n_1428 ,csa_tree_add_190_195_groupi_n_1427);
  not csa_tree_add_190_195_groupi_drc_bufs49149(csa_tree_add_190_195_groupi_n_1427 ,csa_tree_add_190_195_groupi_n_2573);
  not csa_tree_add_190_195_groupi_drc_bufs49152(csa_tree_add_190_195_groupi_n_1426 ,csa_tree_add_190_195_groupi_n_1425);
  not csa_tree_add_190_195_groupi_drc_bufs49153(csa_tree_add_190_195_groupi_n_1425 ,csa_tree_add_190_195_groupi_n_2575);
  not csa_tree_add_190_195_groupi_drc_bufs49155(csa_tree_add_190_195_groupi_n_1424 ,csa_tree_add_190_195_groupi_n_1423);
  not csa_tree_add_190_195_groupi_drc_bufs49157(csa_tree_add_190_195_groupi_n_1423 ,csa_tree_add_190_195_groupi_n_2611);
  not csa_tree_add_190_195_groupi_drc_bufs49159(csa_tree_add_190_195_groupi_n_1422 ,csa_tree_add_190_195_groupi_n_1421);
  not csa_tree_add_190_195_groupi_drc_bufs49161(csa_tree_add_190_195_groupi_n_1421 ,csa_tree_add_190_195_groupi_n_2653);
  not csa_tree_add_190_195_groupi_drc_bufs49163(csa_tree_add_190_195_groupi_n_1420 ,csa_tree_add_190_195_groupi_n_1419);
  not csa_tree_add_190_195_groupi_drc_bufs49165(csa_tree_add_190_195_groupi_n_1419 ,csa_tree_add_190_195_groupi_n_2623);
  not csa_tree_add_190_195_groupi_drc_bufs49167(csa_tree_add_190_195_groupi_n_1418 ,csa_tree_add_190_195_groupi_n_1417);
  not csa_tree_add_190_195_groupi_drc_bufs49169(csa_tree_add_190_195_groupi_n_1417 ,csa_tree_add_190_195_groupi_n_2627);
  not csa_tree_add_190_195_groupi_drc_bufs49183(csa_tree_add_190_195_groupi_n_1416 ,csa_tree_add_190_195_groupi_n_1414);
  not csa_tree_add_190_195_groupi_drc_bufs49184(csa_tree_add_190_195_groupi_n_1415 ,csa_tree_add_190_195_groupi_n_1414);
  not csa_tree_add_190_195_groupi_drc_bufs49185(csa_tree_add_190_195_groupi_n_1414 ,csa_tree_add_190_195_groupi_n_2364);
  not csa_tree_add_190_195_groupi_drc_bufs49191(csa_tree_add_190_195_groupi_n_1413 ,csa_tree_add_190_195_groupi_n_1412);
  not csa_tree_add_190_195_groupi_drc_bufs49193(csa_tree_add_190_195_groupi_n_1412 ,csa_tree_add_190_195_groupi_n_2649);
  not csa_tree_add_190_195_groupi_drc_bufs49195(csa_tree_add_190_195_groupi_n_1411 ,csa_tree_add_190_195_groupi_n_1409);
  not csa_tree_add_190_195_groupi_drc_bufs49196(csa_tree_add_190_195_groupi_n_1410 ,csa_tree_add_190_195_groupi_n_1409);
  not csa_tree_add_190_195_groupi_drc_bufs49197(csa_tree_add_190_195_groupi_n_1409 ,csa_tree_add_190_195_groupi_n_2367);
  not csa_tree_add_190_195_groupi_drc_bufs49207(csa_tree_add_190_195_groupi_n_1408 ,csa_tree_add_190_195_groupi_n_1407);
  not csa_tree_add_190_195_groupi_drc_bufs49209(csa_tree_add_190_195_groupi_n_1407 ,csa_tree_add_190_195_groupi_n_2608);
  not csa_tree_add_190_195_groupi_drc_bufs49219(csa_tree_add_190_195_groupi_n_1406 ,csa_tree_add_190_195_groupi_n_1405);
  not csa_tree_add_190_195_groupi_drc_bufs49221(csa_tree_add_190_195_groupi_n_1405 ,csa_tree_add_190_195_groupi_n_2451);
  not csa_tree_add_190_195_groupi_drc_bufs49223(csa_tree_add_190_195_groupi_n_1404 ,csa_tree_add_190_195_groupi_n_1402);
  not csa_tree_add_190_195_groupi_drc_bufs49224(csa_tree_add_190_195_groupi_n_1403 ,csa_tree_add_190_195_groupi_n_1402);
  not csa_tree_add_190_195_groupi_drc_bufs49225(csa_tree_add_190_195_groupi_n_1402 ,csa_tree_add_190_195_groupi_n_2366);
  not csa_tree_add_190_195_groupi_drc_bufs49235(csa_tree_add_190_195_groupi_n_1401 ,csa_tree_add_190_195_groupi_n_1400);
  not csa_tree_add_190_195_groupi_drc_bufs49237(csa_tree_add_190_195_groupi_n_1400 ,csa_tree_add_190_195_groupi_n_2429);
  not csa_tree_add_190_195_groupi_drc_bufs49247(csa_tree_add_190_195_groupi_n_1399 ,csa_tree_add_190_195_groupi_n_1398);
  not csa_tree_add_190_195_groupi_drc_bufs49249(csa_tree_add_190_195_groupi_n_1398 ,csa_tree_add_190_195_groupi_n_2656);
  not csa_tree_add_190_195_groupi_drc_bufs49251(csa_tree_add_190_195_groupi_n_1397 ,csa_tree_add_190_195_groupi_n_1396);
  not csa_tree_add_190_195_groupi_drc_bufs49253(csa_tree_add_190_195_groupi_n_1396 ,csa_tree_add_190_195_groupi_n_2643);
  not csa_tree_add_190_195_groupi_drc_bufs49256(csa_tree_add_190_195_groupi_n_1395 ,csa_tree_add_190_195_groupi_n_1394);
  not csa_tree_add_190_195_groupi_drc_bufs49257(csa_tree_add_190_195_groupi_n_1394 ,csa_tree_add_190_195_groupi_n_2419);
  not csa_tree_add_190_195_groupi_drc_bufs49275(csa_tree_add_190_195_groupi_n_1393 ,csa_tree_add_190_195_groupi_n_1391);
  not csa_tree_add_190_195_groupi_drc_bufs49276(csa_tree_add_190_195_groupi_n_1392 ,csa_tree_add_190_195_groupi_n_1391);
  not csa_tree_add_190_195_groupi_drc_bufs49277(csa_tree_add_190_195_groupi_n_1391 ,csa_tree_add_190_195_groupi_n_2340);
  not csa_tree_add_190_195_groupi_drc_bufs49283(csa_tree_add_190_195_groupi_n_1390 ,csa_tree_add_190_195_groupi_n_1389);
  not csa_tree_add_190_195_groupi_drc_bufs49285(csa_tree_add_190_195_groupi_n_1389 ,csa_tree_add_190_195_groupi_n_2648);
  not csa_tree_add_190_195_groupi_drc_bufs49287(csa_tree_add_190_195_groupi_n_1388 ,csa_tree_add_190_195_groupi_n_1387);
  not csa_tree_add_190_195_groupi_drc_bufs49289(csa_tree_add_190_195_groupi_n_1387 ,csa_tree_add_190_195_groupi_n_2616);
  not csa_tree_add_190_195_groupi_drc_bufs49291(csa_tree_add_190_195_groupi_n_1386 ,csa_tree_add_190_195_groupi_n_1385);
  not csa_tree_add_190_195_groupi_drc_bufs49293(csa_tree_add_190_195_groupi_n_1385 ,csa_tree_add_190_195_groupi_n_2454);
  not csa_tree_add_190_195_groupi_drc_bufs49295(csa_tree_add_190_195_groupi_n_1384 ,csa_tree_add_190_195_groupi_n_1383);
  not csa_tree_add_190_195_groupi_drc_bufs49297(csa_tree_add_190_195_groupi_n_1383 ,csa_tree_add_190_195_groupi_n_2440);
  not csa_tree_add_190_195_groupi_drc_bufs49299(csa_tree_add_190_195_groupi_n_1382 ,csa_tree_add_190_195_groupi_n_1381);
  not csa_tree_add_190_195_groupi_drc_bufs49301(csa_tree_add_190_195_groupi_n_1381 ,csa_tree_add_190_195_groupi_n_2628);
  not csa_tree_add_190_195_groupi_drc_bufs49319(csa_tree_add_190_195_groupi_n_1380 ,csa_tree_add_190_195_groupi_n_1379);
  not csa_tree_add_190_195_groupi_drc_bufs49321(csa_tree_add_190_195_groupi_n_1379 ,csa_tree_add_190_195_groupi_n_2420);
  not csa_tree_add_190_195_groupi_drc_bufs49328(csa_tree_add_190_195_groupi_n_1378 ,csa_tree_add_190_195_groupi_n_1377);
  not csa_tree_add_190_195_groupi_drc_bufs49329(csa_tree_add_190_195_groupi_n_1377 ,csa_tree_add_190_195_groupi_n_2525);
  not csa_tree_add_190_195_groupi_drc_bufs49344(csa_tree_add_190_195_groupi_n_1376 ,csa_tree_add_190_195_groupi_n_1375);
  not csa_tree_add_190_195_groupi_drc_bufs49345(csa_tree_add_190_195_groupi_n_1375 ,csa_tree_add_190_195_groupi_n_2715);
  not csa_tree_add_190_195_groupi_drc_bufs49352(csa_tree_add_190_195_groupi_n_1374 ,csa_tree_add_190_195_groupi_n_1373);
  not csa_tree_add_190_195_groupi_drc_bufs49353(csa_tree_add_190_195_groupi_n_1373 ,csa_tree_add_190_195_groupi_n_2613);
  not csa_tree_add_190_195_groupi_drc_bufs49359(csa_tree_add_190_195_groupi_n_1372 ,csa_tree_add_190_195_groupi_n_1371);
  not csa_tree_add_190_195_groupi_drc_bufs49361(csa_tree_add_190_195_groupi_n_1371 ,csa_tree_add_190_195_groupi_n_2472);
  not csa_tree_add_190_195_groupi_drc_bufs49363(csa_tree_add_190_195_groupi_n_1370 ,csa_tree_add_190_195_groupi_n_1369);
  not csa_tree_add_190_195_groupi_drc_bufs49365(csa_tree_add_190_195_groupi_n_1369 ,csa_tree_add_190_195_groupi_n_2602);
  not csa_tree_add_190_195_groupi_drc_bufs49367(csa_tree_add_190_195_groupi_n_1368 ,csa_tree_add_190_195_groupi_n_1367);
  not csa_tree_add_190_195_groupi_drc_bufs49369(csa_tree_add_190_195_groupi_n_1367 ,csa_tree_add_190_195_groupi_n_2617);
  not csa_tree_add_190_195_groupi_drc_bufs49371(csa_tree_add_190_195_groupi_n_1366 ,csa_tree_add_190_195_groupi_n_1365);
  not csa_tree_add_190_195_groupi_drc_bufs49373(csa_tree_add_190_195_groupi_n_1365 ,csa_tree_add_190_195_groupi_n_2444);
  not csa_tree_add_190_195_groupi_drc_bufs49375(csa_tree_add_190_195_groupi_n_1364 ,csa_tree_add_190_195_groupi_n_1363);
  not csa_tree_add_190_195_groupi_drc_bufs49377(csa_tree_add_190_195_groupi_n_1363 ,csa_tree_add_190_195_groupi_n_2493);
  not csa_tree_add_190_195_groupi_drc_bufs49384(csa_tree_add_190_195_groupi_n_1362 ,csa_tree_add_190_195_groupi_n_1361);
  not csa_tree_add_190_195_groupi_drc_bufs49385(csa_tree_add_190_195_groupi_n_1361 ,csa_tree_add_190_195_groupi_n_2461);
  not csa_tree_add_190_195_groupi_drc_bufs49387(csa_tree_add_190_195_groupi_n_1360 ,csa_tree_add_190_195_groupi_n_1359);
  not csa_tree_add_190_195_groupi_drc_bufs49389(csa_tree_add_190_195_groupi_n_1359 ,csa_tree_add_190_195_groupi_n_2603);
  not csa_tree_add_190_195_groupi_drc_bufs49391(csa_tree_add_190_195_groupi_n_1358 ,csa_tree_add_190_195_groupi_n_1357);
  not csa_tree_add_190_195_groupi_drc_bufs49393(csa_tree_add_190_195_groupi_n_1357 ,csa_tree_add_190_195_groupi_n_2606);
  not csa_tree_add_190_195_groupi_drc_bufs49395(csa_tree_add_190_195_groupi_n_1356 ,csa_tree_add_190_195_groupi_n_1355);
  not csa_tree_add_190_195_groupi_drc_bufs49397(csa_tree_add_190_195_groupi_n_1355 ,csa_tree_add_190_195_groupi_n_2475);
  not csa_tree_add_190_195_groupi_drc_bufs49400(csa_tree_add_190_195_groupi_n_1354 ,csa_tree_add_190_195_groupi_n_2393);
  not csa_tree_add_190_195_groupi_drc_bufs49401(csa_tree_add_190_195_groupi_n_2393 ,csa_tree_add_190_195_groupi_n_3202);
  not csa_tree_add_190_195_groupi_drc_bufs49404(csa_tree_add_190_195_groupi_n_1353 ,csa_tree_add_190_195_groupi_n_1352);
  not csa_tree_add_190_195_groupi_drc_bufs49405(csa_tree_add_190_195_groupi_n_1352 ,csa_tree_add_190_195_groupi_n_2636);
  not csa_tree_add_190_195_groupi_drc_bufs49408(csa_tree_add_190_195_groupi_n_1351 ,csa_tree_add_190_195_groupi_n_2394);
  not csa_tree_add_190_195_groupi_drc_bufs49409(csa_tree_add_190_195_groupi_n_2394 ,csa_tree_add_190_195_groupi_n_3695);
  not csa_tree_add_190_195_groupi_drc_bufs49411(csa_tree_add_190_195_groupi_n_1350 ,csa_tree_add_190_195_groupi_n_1349);
  not csa_tree_add_190_195_groupi_drc_bufs49413(csa_tree_add_190_195_groupi_n_1349 ,csa_tree_add_190_195_groupi_n_2480);
  not csa_tree_add_190_195_groupi_drc_bufs49416(csa_tree_add_190_195_groupi_n_1348 ,csa_tree_add_190_195_groupi_n_1347);
  not csa_tree_add_190_195_groupi_drc_bufs49417(csa_tree_add_190_195_groupi_n_1347 ,csa_tree_add_190_195_groupi_n_3201);
  not csa_tree_add_190_195_groupi_drc_bufs49420(csa_tree_add_190_195_groupi_n_1346 ,csa_tree_add_190_195_groupi_n_1345);
  not csa_tree_add_190_195_groupi_drc_bufs49421(csa_tree_add_190_195_groupi_n_1345 ,csa_tree_add_190_195_groupi_n_2591);
  not csa_tree_add_190_195_groupi_drc_bufs49424(csa_tree_add_190_195_groupi_n_1344 ,csa_tree_add_190_195_groupi_n_1343);
  not csa_tree_add_190_195_groupi_drc_bufs49425(csa_tree_add_190_195_groupi_n_1343 ,csa_tree_add_190_195_groupi_n_2590);
  not csa_tree_add_190_195_groupi_drc_bufs49428(csa_tree_add_190_195_groupi_n_1342 ,csa_tree_add_190_195_groupi_n_1341);
  not csa_tree_add_190_195_groupi_drc_bufs49429(csa_tree_add_190_195_groupi_n_1341 ,csa_tree_add_190_195_groupi_n_2599);
  not csa_tree_add_190_195_groupi_drc_bufs49432(csa_tree_add_190_195_groupi_n_1340 ,csa_tree_add_190_195_groupi_n_1339);
  not csa_tree_add_190_195_groupi_drc_bufs49433(csa_tree_add_190_195_groupi_n_1339 ,csa_tree_add_190_195_groupi_n_2595);
  not csa_tree_add_190_195_groupi_drc_bufs49436(csa_tree_add_190_195_groupi_n_1338 ,csa_tree_add_190_195_groupi_n_1337);
  not csa_tree_add_190_195_groupi_drc_bufs49437(csa_tree_add_190_195_groupi_n_1337 ,csa_tree_add_190_195_groupi_n_2423);
  not csa_tree_add_190_195_groupi_drc_bufs49440(csa_tree_add_190_195_groupi_n_1336 ,csa_tree_add_190_195_groupi_n_1335);
  not csa_tree_add_190_195_groupi_drc_bufs49441(csa_tree_add_190_195_groupi_n_1335 ,csa_tree_add_190_195_groupi_n_2425);
  not csa_tree_add_190_195_groupi_drc_bufs49444(csa_tree_add_190_195_groupi_n_1334 ,csa_tree_add_190_195_groupi_n_1333);
  not csa_tree_add_190_195_groupi_drc_bufs49445(csa_tree_add_190_195_groupi_n_1333 ,csa_tree_add_190_195_groupi_n_2600);
  not csa_tree_add_190_195_groupi_drc_bufs49552(csa_tree_add_190_195_groupi_n_1332 ,csa_tree_add_190_195_groupi_n_1331);
  not csa_tree_add_190_195_groupi_drc_bufs49553(csa_tree_add_190_195_groupi_n_1331 ,csa_tree_add_190_195_groupi_n_8313);
  not csa_tree_add_190_195_groupi_drc_bufs49582(csa_tree_add_190_195_groupi_n_1330 ,csa_tree_add_190_195_groupi_n_4114);
  not csa_tree_add_190_195_groupi_drc_bufs49596(csa_tree_add_190_195_groupi_n_1329 ,csa_tree_add_190_195_groupi_n_3200);
  buf csa_tree_add_190_195_groupi_drc_bufs49603(out1[12] ,csa_tree_add_190_195_groupi_n_184);
  buf csa_tree_add_190_195_groupi_drc_bufs49604(out1[19] ,csa_tree_add_190_195_groupi_n_185);
  buf csa_tree_add_190_195_groupi_drc_bufs49605(out1[23] ,csa_tree_add_190_195_groupi_n_12597);
  buf csa_tree_add_190_195_groupi_drc_bufs49606(out1[20] ,csa_tree_add_190_195_groupi_n_12589);
  buf csa_tree_add_190_195_groupi_drc_bufs49607(out1[25] ,csa_tree_add_190_195_groupi_n_12603);
  buf csa_tree_add_190_195_groupi_drc_bufs49608(out1[26] ,csa_tree_add_190_195_groupi_n_12606);
  buf csa_tree_add_190_195_groupi_drc_bufs49609(out1[27] ,csa_tree_add_190_195_groupi_n_12609);
  buf csa_tree_add_190_195_groupi_drc_bufs49610(out1[13] ,csa_tree_add_190_195_groupi_n_12566);
  buf csa_tree_add_190_195_groupi_drc_bufs49611(out1[24] ,csa_tree_add_190_195_groupi_n_12600);
  buf csa_tree_add_190_195_groupi_drc_bufs49612(out1[21] ,csa_tree_add_190_195_groupi_n_186);
  buf csa_tree_add_190_195_groupi_drc_bufs49613(out1[22] ,csa_tree_add_190_195_groupi_n_12594);
  buf csa_tree_add_190_195_groupi_drc_bufs49614(out1[17] ,csa_tree_add_190_195_groupi_n_12580);
  buf csa_tree_add_190_195_groupi_drc_bufs49615(out1[14] ,csa_tree_add_190_195_groupi_n_12570);
  buf csa_tree_add_190_195_groupi_drc_bufs49616(out1[15] ,csa_tree_add_190_195_groupi_n_12573);
  not csa_tree_add_190_195_groupi_drc_bufs49618(csa_tree_add_190_195_groupi_n_1314 ,csa_tree_add_190_195_groupi_n_3690);
  not csa_tree_add_190_195_groupi_drc_bufs49628(csa_tree_add_190_195_groupi_n_2396 ,csa_tree_add_190_195_groupi_n_5257);
  not csa_tree_add_190_195_groupi_drc_bufs49632(csa_tree_add_190_195_groupi_n_2401 ,csa_tree_add_190_195_groupi_n_5550);
  not csa_tree_add_190_195_groupi_drc_bufs49635(csa_tree_add_190_195_groupi_n_1313 ,csa_tree_add_190_195_groupi_n_2395);
  not csa_tree_add_190_195_groupi_drc_bufs49636(csa_tree_add_190_195_groupi_n_2395 ,csa_tree_add_190_195_groupi_n_5210);
  not csa_tree_add_190_195_groupi_drc_bufs49640(csa_tree_add_190_195_groupi_n_2403 ,csa_tree_add_190_195_groupi_n_37);
  not csa_tree_add_190_195_groupi_drc_bufs49644(csa_tree_add_190_195_groupi_n_2397 ,csa_tree_add_190_195_groupi_n_5286);
  not csa_tree_add_190_195_groupi_drc_bufs49653(csa_tree_add_190_195_groupi_n_2398 ,csa_tree_add_190_195_groupi_n_5329);
  not csa_tree_add_190_195_groupi_drc_bufs49661(csa_tree_add_190_195_groupi_n_2404 ,csa_tree_add_190_195_groupi_n_5916);
  not csa_tree_add_190_195_groupi_drc_bufs49664(csa_tree_add_190_195_groupi_n_1312 ,csa_tree_add_190_195_groupi_n_2400);
  not csa_tree_add_190_195_groupi_drc_bufs49665(csa_tree_add_190_195_groupi_n_2400 ,csa_tree_add_190_195_groupi_n_5520);
  not csa_tree_add_190_195_groupi_drc_bufs49669(csa_tree_add_190_195_groupi_n_2399 ,csa_tree_add_190_195_groupi_n_5422);
  not csa_tree_add_190_195_groupi_drc_bufs49672(csa_tree_add_190_195_groupi_n_1311 ,csa_tree_add_190_195_groupi_n_2402);
  not csa_tree_add_190_195_groupi_drc_bufs49673(csa_tree_add_190_195_groupi_n_2402 ,csa_tree_add_190_195_groupi_n_5900);
  not csa_tree_add_190_195_groupi_drc_bufs49676(csa_tree_add_190_195_groupi_n_1310 ,csa_tree_add_190_195_groupi_n_2405);
  not csa_tree_add_190_195_groupi_drc_bufs49677(csa_tree_add_190_195_groupi_n_2405 ,csa_tree_add_190_195_groupi_n_9897);
  buf csa_tree_add_190_195_groupi_drc_bufs49935(csa_tree_add_190_195_groupi_n_1903 ,n_114);
  buf csa_tree_add_190_195_groupi_drc_bufs49936(csa_tree_add_190_195_groupi_n_1900 ,n_80);
  buf csa_tree_add_190_195_groupi_drc_bufs49937(csa_tree_add_190_195_groupi_n_1899 ,n_73);
  buf csa_tree_add_190_195_groupi_drc_bufs49938(csa_tree_add_190_195_groupi_n_1898 ,n_63);
  buf csa_tree_add_190_195_groupi_drc_bufs49939(csa_tree_add_190_195_groupi_n_1896 ,n_22);
  buf csa_tree_add_190_195_groupi_drc_bufs49940(csa_tree_add_190_195_groupi_n_1895 ,n_12);
  buf csa_tree_add_190_195_groupi_drc_bufs49941(csa_tree_add_190_195_groupi_n_1894 ,n_5);
  buf csa_tree_add_190_195_groupi_drc_bufs49942(csa_tree_add_190_195_groupi_n_1901 ,n_97);
  buf csa_tree_add_190_195_groupi_drc_bufs49943(csa_tree_add_190_195_groupi_n_1897 ,n_56);
  buf csa_tree_add_190_195_groupi_drc_bufs49944(csa_tree_add_190_195_groupi_n_1902 ,n_284);
  buf csa_tree_add_190_195_groupi_drc_bufs49945(csa_tree_add_190_195_groupi_n_1694 ,n_44);
  not csa_tree_add_190_195_groupi_drc_bufs49947(csa_tree_add_190_195_groupi_n_1309 ,csa_tree_add_190_195_groupi_n_1308);
  not csa_tree_add_190_195_groupi_drc_bufs49948(csa_tree_add_190_195_groupi_n_1308 ,csa_tree_add_190_195_groupi_n_2228);
  not csa_tree_add_190_195_groupi_drc_bufs49951(csa_tree_add_190_195_groupi_n_1307 ,csa_tree_add_190_195_groupi_n_1306);
  not csa_tree_add_190_195_groupi_drc_bufs49952(csa_tree_add_190_195_groupi_n_1306 ,csa_tree_add_190_195_groupi_n_2103);
  not csa_tree_add_190_195_groupi_drc_bufs49955(csa_tree_add_190_195_groupi_n_1305 ,csa_tree_add_190_195_groupi_n_1304);
  not csa_tree_add_190_195_groupi_drc_bufs49956(csa_tree_add_190_195_groupi_n_1304 ,csa_tree_add_190_195_groupi_n_2227);
  not csa_tree_add_190_195_groupi_drc_bufs49959(csa_tree_add_190_195_groupi_n_1303 ,csa_tree_add_190_195_groupi_n_1302);
  not csa_tree_add_190_195_groupi_drc_bufs49960(csa_tree_add_190_195_groupi_n_1302 ,csa_tree_add_190_195_groupi_n_2121);
  not csa_tree_add_190_195_groupi_drc_bufs49963(csa_tree_add_190_195_groupi_n_1301 ,csa_tree_add_190_195_groupi_n_1300);
  not csa_tree_add_190_195_groupi_drc_bufs49964(csa_tree_add_190_195_groupi_n_1300 ,csa_tree_add_190_195_groupi_n_2102);
  not csa_tree_add_190_195_groupi_drc_bufs49967(csa_tree_add_190_195_groupi_n_1299 ,csa_tree_add_190_195_groupi_n_1298);
  not csa_tree_add_190_195_groupi_drc_bufs49968(csa_tree_add_190_195_groupi_n_1298 ,csa_tree_add_190_195_groupi_n_2077);
  not csa_tree_add_190_195_groupi_drc_bufs49971(csa_tree_add_190_195_groupi_n_1297 ,csa_tree_add_190_195_groupi_n_1296);
  not csa_tree_add_190_195_groupi_drc_bufs49972(csa_tree_add_190_195_groupi_n_1296 ,csa_tree_add_190_195_groupi_n_2234);
  not csa_tree_add_190_195_groupi_drc_bufs49975(csa_tree_add_190_195_groupi_n_1295 ,csa_tree_add_190_195_groupi_n_1294);
  not csa_tree_add_190_195_groupi_drc_bufs49976(csa_tree_add_190_195_groupi_n_1294 ,csa_tree_add_190_195_groupi_n_2230);
  not csa_tree_add_190_195_groupi_drc_bufs49979(csa_tree_add_190_195_groupi_n_1293 ,csa_tree_add_190_195_groupi_n_1292);
  not csa_tree_add_190_195_groupi_drc_bufs49980(csa_tree_add_190_195_groupi_n_1292 ,csa_tree_add_190_195_groupi_n_2122);
  not csa_tree_add_190_195_groupi_drc_bufs49983(csa_tree_add_190_195_groupi_n_1291 ,csa_tree_add_190_195_groupi_n_1290);
  not csa_tree_add_190_195_groupi_drc_bufs49984(csa_tree_add_190_195_groupi_n_1290 ,csa_tree_add_190_195_groupi_n_2078);
  not csa_tree_add_190_195_groupi_drc_bufs49987(csa_tree_add_190_195_groupi_n_1289 ,csa_tree_add_190_195_groupi_n_1288);
  not csa_tree_add_190_195_groupi_drc_bufs49988(csa_tree_add_190_195_groupi_n_1288 ,csa_tree_add_190_195_groupi_n_2237);
  not csa_tree_add_190_195_groupi_drc_bufs49991(csa_tree_add_190_195_groupi_n_1287 ,csa_tree_add_190_195_groupi_n_1286);
  not csa_tree_add_190_195_groupi_drc_bufs49992(csa_tree_add_190_195_groupi_n_1286 ,csa_tree_add_190_195_groupi_n_2177);
  not csa_tree_add_190_195_groupi_drc_bufs49995(csa_tree_add_190_195_groupi_n_1285 ,csa_tree_add_190_195_groupi_n_1284);
  not csa_tree_add_190_195_groupi_drc_bufs49996(csa_tree_add_190_195_groupi_n_1284 ,csa_tree_add_190_195_groupi_n_2294);
  not csa_tree_add_190_195_groupi_drc_bufs49999(csa_tree_add_190_195_groupi_n_1283 ,csa_tree_add_190_195_groupi_n_1282);
  not csa_tree_add_190_195_groupi_drc_bufs50000(csa_tree_add_190_195_groupi_n_1282 ,csa_tree_add_190_195_groupi_n_2293);
  not csa_tree_add_190_195_groupi_drc_bufs50003(csa_tree_add_190_195_groupi_n_1281 ,csa_tree_add_190_195_groupi_n_1280);
  not csa_tree_add_190_195_groupi_drc_bufs50004(csa_tree_add_190_195_groupi_n_1280 ,csa_tree_add_190_195_groupi_n_2204);
  not csa_tree_add_190_195_groupi_drc_bufs50007(csa_tree_add_190_195_groupi_n_1279 ,csa_tree_add_190_195_groupi_n_1278);
  not csa_tree_add_190_195_groupi_drc_bufs50008(csa_tree_add_190_195_groupi_n_1278 ,csa_tree_add_190_195_groupi_n_2201);
  not csa_tree_add_190_195_groupi_drc_bufs50010(csa_tree_add_190_195_groupi_n_1277 ,csa_tree_add_190_195_groupi_n_1276);
  not csa_tree_add_190_195_groupi_drc_bufs50012(csa_tree_add_190_195_groupi_n_1276 ,csa_tree_add_190_195_groupi_n_2193);
  not csa_tree_add_190_195_groupi_drc_bufs50015(csa_tree_add_190_195_groupi_n_1275 ,csa_tree_add_190_195_groupi_n_1274);
  not csa_tree_add_190_195_groupi_drc_bufs50016(csa_tree_add_190_195_groupi_n_1274 ,csa_tree_add_190_195_groupi_n_2218);
  not csa_tree_add_190_195_groupi_drc_bufs50018(csa_tree_add_190_195_groupi_n_1273 ,csa_tree_add_190_195_groupi_n_1272);
  not csa_tree_add_190_195_groupi_drc_bufs50020(csa_tree_add_190_195_groupi_n_1272 ,csa_tree_add_190_195_groupi_n_2246);
  not csa_tree_add_190_195_groupi_drc_bufs50022(csa_tree_add_190_195_groupi_n_1271 ,csa_tree_add_190_195_groupi_n_1270);
  not csa_tree_add_190_195_groupi_drc_bufs50024(csa_tree_add_190_195_groupi_n_1270 ,csa_tree_add_190_195_groupi_n_2240);
  not csa_tree_add_190_195_groupi_drc_bufs50026(csa_tree_add_190_195_groupi_n_1269 ,csa_tree_add_190_195_groupi_n_1268);
  not csa_tree_add_190_195_groupi_drc_bufs50028(csa_tree_add_190_195_groupi_n_1268 ,csa_tree_add_190_195_groupi_n_2242);
  buf csa_tree_add_190_195_groupi_drc_bufs50030(csa_tree_add_190_195_groupi_n_2007 ,n_318);
  not csa_tree_add_190_195_groupi_drc_bufs50032(csa_tree_add_190_195_groupi_n_1267 ,csa_tree_add_190_195_groupi_n_1266);
  not csa_tree_add_190_195_groupi_drc_bufs50033(csa_tree_add_190_195_groupi_n_1266 ,csa_tree_add_190_195_groupi_n_2115);
  not csa_tree_add_190_195_groupi_drc_bufs50035(csa_tree_add_190_195_groupi_n_1265 ,csa_tree_add_190_195_groupi_n_1264);
  not csa_tree_add_190_195_groupi_drc_bufs50037(csa_tree_add_190_195_groupi_n_1264 ,csa_tree_add_190_195_groupi_n_2124);
  not csa_tree_add_190_195_groupi_drc_bufs50040(csa_tree_add_190_195_groupi_n_1263 ,csa_tree_add_190_195_groupi_n_1262);
  not csa_tree_add_190_195_groupi_drc_bufs50041(csa_tree_add_190_195_groupi_n_1262 ,csa_tree_add_190_195_groupi_n_2111);
  not csa_tree_add_190_195_groupi_drc_bufs50044(csa_tree_add_190_195_groupi_n_1261 ,csa_tree_add_190_195_groupi_n_1260);
  not csa_tree_add_190_195_groupi_drc_bufs50045(csa_tree_add_190_195_groupi_n_1260 ,csa_tree_add_190_195_groupi_n_2108);
  not csa_tree_add_190_195_groupi_drc_bufs50048(csa_tree_add_190_195_groupi_n_1259 ,csa_tree_add_190_195_groupi_n_1258);
  not csa_tree_add_190_195_groupi_drc_bufs50049(csa_tree_add_190_195_groupi_n_1258 ,csa_tree_add_190_195_groupi_n_2106);
  buf csa_tree_add_190_195_groupi_drc_bufs50051(csa_tree_add_190_195_groupi_n_2005 ,n_124);
  not csa_tree_add_190_195_groupi_drc_bufs50053(csa_tree_add_190_195_groupi_n_1257 ,csa_tree_add_190_195_groupi_n_1256);
  not csa_tree_add_190_195_groupi_drc_bufs50054(csa_tree_add_190_195_groupi_n_1256 ,csa_tree_add_190_195_groupi_n_2181);
  not csa_tree_add_190_195_groupi_drc_bufs50057(csa_tree_add_190_195_groupi_n_1255 ,csa_tree_add_190_195_groupi_n_1254);
  not csa_tree_add_190_195_groupi_drc_bufs50058(csa_tree_add_190_195_groupi_n_1254 ,csa_tree_add_190_195_groupi_n_2161);
  not csa_tree_add_190_195_groupi_drc_bufs50060(csa_tree_add_190_195_groupi_n_1253 ,csa_tree_add_190_195_groupi_n_1252);
  not csa_tree_add_190_195_groupi_drc_bufs50062(csa_tree_add_190_195_groupi_n_1252 ,csa_tree_add_190_195_groupi_n_2207);
  buf csa_tree_add_190_195_groupi_drc_bufs50064(csa_tree_add_190_195_groupi_n_2003 ,n_90);
  buf csa_tree_add_190_195_groupi_drc_bufs50065(csa_tree_add_190_195_groupi_n_2001 ,n_39);
  not csa_tree_add_190_195_groupi_drc_bufs50066(csa_tree_add_190_195_groupi_n_1251 ,csa_tree_add_190_195_groupi_n_1250);
  not csa_tree_add_190_195_groupi_drc_bufs50068(csa_tree_add_190_195_groupi_n_1250 ,csa_tree_add_190_195_groupi_n_2100);
  not csa_tree_add_190_195_groupi_drc_bufs50070(csa_tree_add_190_195_groupi_n_1249 ,csa_tree_add_190_195_groupi_n_1248);
  not csa_tree_add_190_195_groupi_drc_bufs50072(csa_tree_add_190_195_groupi_n_1248 ,csa_tree_add_190_195_groupi_n_2099);
  not csa_tree_add_190_195_groupi_drc_bufs50074(csa_tree_add_190_195_groupi_n_1247 ,csa_tree_add_190_195_groupi_n_1246);
  not csa_tree_add_190_195_groupi_drc_bufs50076(csa_tree_add_190_195_groupi_n_1246 ,csa_tree_add_190_195_groupi_n_2097);
  not csa_tree_add_190_195_groupi_drc_bufs50078(csa_tree_add_190_195_groupi_n_1245 ,csa_tree_add_190_195_groupi_n_2337);
  not csa_tree_add_190_195_groupi_drc_bufs50080(csa_tree_add_190_195_groupi_n_2337 ,csa_tree_add_190_195_groupi_n_2094);
  not csa_tree_add_190_195_groupi_drc_bufs50082(csa_tree_add_190_195_groupi_n_1244 ,csa_tree_add_190_195_groupi_n_1243);
  not csa_tree_add_190_195_groupi_drc_bufs50084(csa_tree_add_190_195_groupi_n_1243 ,csa_tree_add_190_195_groupi_n_2080);
  not csa_tree_add_190_195_groupi_drc_bufs50087(csa_tree_add_190_195_groupi_n_1242 ,csa_tree_add_190_195_groupi_n_1241);
  not csa_tree_add_190_195_groupi_drc_bufs50088(csa_tree_add_190_195_groupi_n_1241 ,csa_tree_add_190_195_groupi_n_2222);
  not csa_tree_add_190_195_groupi_drc_bufs50090(csa_tree_add_190_195_groupi_n_1240 ,csa_tree_add_190_195_groupi_n_1239);
  not csa_tree_add_190_195_groupi_drc_bufs50092(csa_tree_add_190_195_groupi_n_1239 ,csa_tree_add_190_195_groupi_n_2199);
  not csa_tree_add_190_195_groupi_drc_bufs50094(csa_tree_add_190_195_groupi_n_1238 ,csa_tree_add_190_195_groupi_n_1237);
  not csa_tree_add_190_195_groupi_drc_bufs50096(csa_tree_add_190_195_groupi_n_1237 ,csa_tree_add_190_195_groupi_n_2196);
  not csa_tree_add_190_195_groupi_drc_bufs50098(csa_tree_add_190_195_groupi_n_1236 ,csa_tree_add_190_195_groupi_n_1235);
  not csa_tree_add_190_195_groupi_drc_bufs50100(csa_tree_add_190_195_groupi_n_1235 ,csa_tree_add_190_195_groupi_n_2189);
  not csa_tree_add_190_195_groupi_drc_bufs50103(csa_tree_add_190_195_groupi_n_1234 ,csa_tree_add_190_195_groupi_n_1233);
  not csa_tree_add_190_195_groupi_drc_bufs50104(csa_tree_add_190_195_groupi_n_1233 ,csa_tree_add_190_195_groupi_n_2150);
  buf csa_tree_add_190_195_groupi_drc_bufs50106(csa_tree_add_190_195_groupi_n_1572 ,n_104);
  buf csa_tree_add_190_195_groupi_drc_bufs50107(csa_tree_add_190_195_groupi_n_2002 ,n_46);
  buf csa_tree_add_190_195_groupi_drc_bufs50108(csa_tree_add_190_195_groupi_n_2000 ,n_29);
  buf csa_tree_add_190_195_groupi_drc_bufs50109(csa_tree_add_190_195_groupi_n_1679 ,n_25);
  buf csa_tree_add_190_195_groupi_drc_bufs50110(csa_tree_add_190_195_groupi_n_2004 ,n_107);
  buf csa_tree_add_190_195_groupi_drc_bufs50111(csa_tree_add_190_195_groupi_n_1571 ,n_313);
  buf csa_tree_add_190_195_groupi_drc_bufs50112(csa_tree_add_190_195_groupi_n_1854 ,n_61);
  buf csa_tree_add_190_195_groupi_drc_bufs50113(csa_tree_add_190_195_groupi_n_1853 ,n_27);
  buf csa_tree_add_190_195_groupi_drc_bufs50114(csa_tree_add_190_195_groupi_n_1852 ,n_10);
  buf csa_tree_add_190_195_groupi_drc_bufs50115(csa_tree_add_190_195_groupi_n_1856 ,n_180);
  buf csa_tree_add_190_195_groupi_drc_bufs50116(csa_tree_add_190_195_groupi_n_2008 ,n_182);
  not csa_tree_add_190_195_groupi_drc_bufs50117(csa_tree_add_190_195_groupi_n_1232 ,csa_tree_add_190_195_groupi_n_1231);
  not csa_tree_add_190_195_groupi_drc_bufs50119(csa_tree_add_190_195_groupi_n_1231 ,csa_tree_add_190_195_groupi_n_2164);
  buf csa_tree_add_190_195_groupi_drc_bufs50121(csa_tree_add_190_195_groupi_n_1855 ,n_163);
  buf csa_tree_add_190_195_groupi_drc_bufs50122(csa_tree_add_190_195_groupi_n_2006 ,n_148);
  not csa_tree_add_190_195_groupi_drc_bufs50124(csa_tree_add_190_195_groupi_n_1230 ,csa_tree_add_190_195_groupi_n_1229);
  not csa_tree_add_190_195_groupi_drc_bufs50125(csa_tree_add_190_195_groupi_n_1229 ,csa_tree_add_190_195_groupi_n_2093);
  not csa_tree_add_190_195_groupi_drc_bufs50127(csa_tree_add_190_195_groupi_n_1228 ,csa_tree_add_190_195_groupi_n_1227);
  not csa_tree_add_190_195_groupi_drc_bufs50129(csa_tree_add_190_195_groupi_n_1227 ,csa_tree_add_190_195_groupi_n_2081);
  not csa_tree_add_190_195_groupi_drc_bufs50131(csa_tree_add_190_195_groupi_n_1226 ,csa_tree_add_190_195_groupi_n_1225);
  not csa_tree_add_190_195_groupi_drc_bufs50133(csa_tree_add_190_195_groupi_n_1225 ,csa_tree_add_190_195_groupi_n_2075);
  not csa_tree_add_190_195_groupi_drc_bufs50136(csa_tree_add_190_195_groupi_n_1224 ,csa_tree_add_190_195_groupi_n_1223);
  not csa_tree_add_190_195_groupi_drc_bufs50137(csa_tree_add_190_195_groupi_n_1223 ,csa_tree_add_190_195_groupi_n_2074);
  not csa_tree_add_190_195_groupi_drc_bufs50140(csa_tree_add_190_195_groupi_n_1222 ,csa_tree_add_190_195_groupi_n_1221);
  not csa_tree_add_190_195_groupi_drc_bufs50141(csa_tree_add_190_195_groupi_n_1221 ,csa_tree_add_190_195_groupi_n_1940);
  not csa_tree_add_190_195_groupi_drc_bufs50144(csa_tree_add_190_195_groupi_n_1220 ,csa_tree_add_190_195_groupi_n_1219);
  not csa_tree_add_190_195_groupi_drc_bufs50145(csa_tree_add_190_195_groupi_n_1219 ,csa_tree_add_190_195_groupi_n_2068);
  not csa_tree_add_190_195_groupi_drc_bufs50148(csa_tree_add_190_195_groupi_n_1218 ,csa_tree_add_190_195_groupi_n_1217);
  not csa_tree_add_190_195_groupi_drc_bufs50149(csa_tree_add_190_195_groupi_n_1217 ,csa_tree_add_190_195_groupi_n_2025);
  not csa_tree_add_190_195_groupi_drc_bufs50152(csa_tree_add_190_195_groupi_n_1216 ,csa_tree_add_190_195_groupi_n_1215);
  not csa_tree_add_190_195_groupi_drc_bufs50153(csa_tree_add_190_195_groupi_n_1215 ,csa_tree_add_190_195_groupi_n_2151);
  not csa_tree_add_190_195_groupi_drc_bufs50155(csa_tree_add_190_195_groupi_n_1214 ,csa_tree_add_190_195_groupi_n_1213);
  not csa_tree_add_190_195_groupi_drc_bufs50157(csa_tree_add_190_195_groupi_n_1213 ,csa_tree_add_190_195_groupi_n_2145);
  buf csa_tree_add_190_195_groupi_drc_bufs50159(csa_tree_add_190_195_groupi_n_1678 ,n_47);
  not csa_tree_add_190_195_groupi_drc_bufs50161(csa_tree_add_190_195_groupi_n_1212 ,csa_tree_add_190_195_groupi_n_1211);
  not csa_tree_add_190_195_groupi_drc_bufs50162(csa_tree_add_190_195_groupi_n_1211 ,csa_tree_add_190_195_groupi_n_2224);
  not csa_tree_add_190_195_groupi_drc_bufs50165(csa_tree_add_190_195_groupi_n_1210 ,csa_tree_add_190_195_groupi_n_1209);
  not csa_tree_add_190_195_groupi_drc_bufs50166(csa_tree_add_190_195_groupi_n_1209 ,csa_tree_add_190_195_groupi_n_2186);
  not csa_tree_add_190_195_groupi_drc_bufs50169(csa_tree_add_190_195_groupi_n_1208 ,csa_tree_add_190_195_groupi_n_1207);
  not csa_tree_add_190_195_groupi_drc_bufs50170(csa_tree_add_190_195_groupi_n_1207 ,csa_tree_add_190_195_groupi_n_2183);
  not csa_tree_add_190_195_groupi_drc_bufs50174(csa_tree_add_190_195_groupi_n_2338 ,csa_tree_add_190_195_groupi_n_2072);
  not csa_tree_add_190_195_groupi_drc_bufs50176(csa_tree_add_190_195_groupi_n_1206 ,csa_tree_add_190_195_groupi_n_1205);
  not csa_tree_add_190_195_groupi_drc_bufs50178(csa_tree_add_190_195_groupi_n_1205 ,csa_tree_add_190_195_groupi_n_2028);
  not csa_tree_add_190_195_groupi_drc_bufs50181(csa_tree_add_190_195_groupi_n_1204 ,csa_tree_add_190_195_groupi_n_1203);
  not csa_tree_add_190_195_groupi_drc_bufs50182(csa_tree_add_190_195_groupi_n_1203 ,csa_tree_add_190_195_groupi_n_2069);
  not csa_tree_add_190_195_groupi_drc_bufs50184(csa_tree_add_190_195_groupi_n_1202 ,csa_tree_add_190_195_groupi_n_1201);
  not csa_tree_add_190_195_groupi_drc_bufs50186(csa_tree_add_190_195_groupi_n_1201 ,csa_tree_add_190_195_groupi_n_2021);
  not csa_tree_add_190_195_groupi_drc_bufs50189(csa_tree_add_190_195_groupi_n_1200 ,csa_tree_add_190_195_groupi_n_2341);
  not csa_tree_add_190_195_groupi_drc_bufs50190(csa_tree_add_190_195_groupi_n_2341 ,csa_tree_add_190_195_groupi_n_2018);
  not csa_tree_add_190_195_groupi_drc_bufs50192(csa_tree_add_190_195_groupi_n_1199 ,csa_tree_add_190_195_groupi_n_1198);
  not csa_tree_add_190_195_groupi_drc_bufs50194(csa_tree_add_190_195_groupi_n_1198 ,csa_tree_add_190_195_groupi_n_2014);
  not csa_tree_add_190_195_groupi_drc_bufs50197(csa_tree_add_190_195_groupi_n_1197 ,csa_tree_add_190_195_groupi_n_1196);
  not csa_tree_add_190_195_groupi_drc_bufs50198(csa_tree_add_190_195_groupi_n_1196 ,csa_tree_add_190_195_groupi_n_2167);
  not csa_tree_add_190_195_groupi_drc_bufs50201(csa_tree_add_190_195_groupi_n_1195 ,csa_tree_add_190_195_groupi_n_1194);
  not csa_tree_add_190_195_groupi_drc_bufs50202(csa_tree_add_190_195_groupi_n_1194 ,csa_tree_add_190_195_groupi_n_2096);
  not csa_tree_add_190_195_groupi_drc_bufs50205(csa_tree_add_190_195_groupi_n_1193 ,csa_tree_add_190_195_groupi_n_1192);
  not csa_tree_add_190_195_groupi_drc_bufs50206(csa_tree_add_190_195_groupi_n_1192 ,csa_tree_add_190_195_groupi_n_2071);
  not csa_tree_add_190_195_groupi_drc_bufs50209(csa_tree_add_190_195_groupi_n_1191 ,csa_tree_add_190_195_groupi_n_1190);
  not csa_tree_add_190_195_groupi_drc_bufs50210(csa_tree_add_190_195_groupi_n_1190 ,csa_tree_add_190_195_groupi_n_2010);
  buf csa_tree_add_190_195_groupi_drc_bufs50212(csa_tree_add_190_195_groupi_n_1767 ,n_71);
  buf csa_tree_add_190_195_groupi_drc_bufs50213(csa_tree_add_190_195_groupi_n_1765 ,n_3);
  buf csa_tree_add_190_195_groupi_drc_bufs50214(csa_tree_add_190_195_groupi_n_2085 ,n_131);
  buf csa_tree_add_190_195_groupi_drc_bufs50215(csa_tree_add_190_195_groupi_n_1550 ,n_312);
  buf csa_tree_add_190_195_groupi_drc_bufs50216(csa_tree_add_190_195_groupi_n_1766 ,n_37);
  buf csa_tree_add_190_195_groupi_drc_bufs50217(csa_tree_add_190_195_groupi_n_1763 ,n_161);
  buf csa_tree_add_190_195_groupi_drc_bufs50218(csa_tree_add_190_195_groupi_n_1764 ,n_314);
  buf csa_tree_add_190_195_groupi_drc_bufs50219(csa_tree_add_190_195_groupi_n_1943 ,n_112);
  buf csa_tree_add_190_195_groupi_drc_bufs50220(csa_tree_add_190_195_groupi_n_1942 ,n_95);
  buf csa_tree_add_190_195_groupi_drc_bufs50221(csa_tree_add_190_195_groupi_n_1759 ,n_59);
  buf csa_tree_add_190_195_groupi_drc_bufs50222(csa_tree_add_190_195_groupi_n_1756 ,n_9);
  buf csa_tree_add_190_195_groupi_drc_bufs50223(csa_tree_add_190_195_groupi_n_1755 ,n_8);
  buf csa_tree_add_190_195_groupi_drc_bufs50224(csa_tree_add_190_195_groupi_n_2084 ,n_277);
  buf csa_tree_add_190_195_groupi_drc_bufs50225(csa_tree_add_190_195_groupi_n_1762 ,n_127);
  buf csa_tree_add_190_195_groupi_drc_bufs50226(csa_tree_add_190_195_groupi_n_2083 ,n_260);
  buf csa_tree_add_190_195_groupi_drc_bufs50227(csa_tree_add_190_195_groupi_n_1754 ,n_81);
  buf csa_tree_add_190_195_groupi_drc_bufs50228(csa_tree_add_190_195_groupi_n_2091 ,n_396);
  buf csa_tree_add_190_195_groupi_drc_bufs50229(csa_tree_add_190_195_groupi_n_2086 ,n_379);
  buf csa_tree_add_190_195_groupi_drc_bufs50230(csa_tree_add_190_195_groupi_n_1760 ,n_60);
  buf csa_tree_add_190_195_groupi_drc_bufs50231(csa_tree_add_190_195_groupi_n_2088 ,n_311);
  buf csa_tree_add_190_195_groupi_drc_bufs50232(csa_tree_add_190_195_groupi_n_1758 ,n_43);
  buf csa_tree_add_190_195_groupi_drc_bufs50233(csa_tree_add_190_195_groupi_n_1757 ,n_26);
  buf csa_tree_add_190_195_groupi_drc_bufs50234(csa_tree_add_190_195_groupi_n_2089 ,n_175);
  buf csa_tree_add_190_195_groupi_drc_bufs50235(csa_tree_add_190_195_groupi_n_1761 ,n_94);
  buf csa_tree_add_190_195_groupi_drc_bufs50236(csa_tree_add_190_195_groupi_n_1608 ,n_62);
  buf csa_tree_add_190_195_groupi_drc_bufs50237(csa_tree_add_190_195_groupi_n_1753 ,n_64);
  buf csa_tree_add_190_195_groupi_drc_bufs50238(csa_tree_add_190_195_groupi_n_2090 ,n_328);
  buf csa_tree_add_190_195_groupi_drc_bufs50239(csa_tree_add_190_195_groupi_n_1752 ,n_13);
  buf csa_tree_add_190_195_groupi_drc_bufs50240(csa_tree_add_190_195_groupi_n_2087 ,n_141);
  buf csa_tree_add_190_195_groupi_drc_bufs50241(csa_tree_add_190_195_groupi_n_1944 ,n_129);
  buf csa_tree_add_190_195_groupi_drc_bufs50242(csa_tree_add_190_195_groupi_n_1941 ,n_78);
  buf csa_tree_add_190_195_groupi_drc_bufs50243(csa_tree_add_190_195_groupi_n_2082 ,n_216);
  buf csa_tree_add_190_195_groupi_drc_bufs50244(csa_tree_add_190_195_groupi_n_1609 ,n_283);
  buf csa_tree_add_190_195_groupi_drc_bufs50245(csa_tree_add_190_195_groupi_n_1945 ,n_316);
  buf csa_tree_add_190_195_groupi_drc_bufs50246(csa_tree_add_190_195_groupi_n_1888 ,n_54);
  buf csa_tree_add_190_195_groupi_drc_bufs50247(csa_tree_add_190_195_groupi_n_1887 ,n_20);
  buf csa_tree_add_190_195_groupi_drc_bufs50248(csa_tree_add_190_195_groupi_n_1708 ,n_344);
  buf csa_tree_add_190_195_groupi_drc_bufs50249(csa_tree_add_190_195_groupi_n_1710 ,n_55);
  buf csa_tree_add_190_195_groupi_drc_bufs50250(csa_tree_add_190_195_groupi_n_1709 ,n_4);
  buf csa_tree_add_190_195_groupi_drc_bufs50251(csa_tree_add_190_195_groupi_n_1711 ,n_106);
  buf csa_tree_add_190_195_groupi_drc_bufs50252(csa_tree_add_190_195_groupi_n_1891 ,n_105);
  buf csa_tree_add_190_195_groupi_drc_bufs50253(csa_tree_add_190_195_groupi_n_1892 ,n_122);
  buf csa_tree_add_190_195_groupi_drc_bufs50254(csa_tree_add_190_195_groupi_n_1889 ,n_88);
  buf csa_tree_add_190_195_groupi_drc_bufs50255(csa_tree_add_190_195_groupi_n_1893 ,n_377);
  buf csa_tree_add_190_195_groupi_drc_bufs50256(csa_tree_add_190_195_groupi_n_2155 ,n_301);
  buf csa_tree_add_190_195_groupi_drc_bufs50257(csa_tree_add_190_195_groupi_n_1698 ,n_53);
  buf csa_tree_add_190_195_groupi_drc_bufs50258(csa_tree_add_190_195_groupi_n_1867 ,n_76);
  buf csa_tree_add_190_195_groupi_drc_bufs50259(csa_tree_add_190_195_groupi_n_1871 ,n_315);
  buf csa_tree_add_190_195_groupi_drc_bufs50260(csa_tree_add_190_195_groupi_n_1873 ,n_179);
  buf csa_tree_add_190_195_groupi_drc_bufs50261(csa_tree_add_190_195_groupi_n_1872 ,n_178);
  buf csa_tree_add_190_195_groupi_drc_bufs50262(csa_tree_add_190_195_groupi_n_1869 ,n_280);
  buf csa_tree_add_190_195_groupi_drc_bufs50263(csa_tree_add_190_195_groupi_n_1890 ,n_275);
  buf csa_tree_add_190_195_groupi_drc_bufs50264(csa_tree_add_190_195_groupi_n_1695 ,n_223);
  buf csa_tree_add_190_195_groupi_drc_bufs50265(csa_tree_add_190_195_groupi_n_1870 ,n_110);
  buf csa_tree_add_190_195_groupi_drc_bufs50266(csa_tree_add_190_195_groupi_n_1687 ,n_96);
  buf csa_tree_add_190_195_groupi_drc_bufs50267(csa_tree_add_190_195_groupi_n_1868 ,n_93);
  buf csa_tree_add_190_195_groupi_drc_bufs50268(csa_tree_add_190_195_groupi_n_1586 ,n_23);
  buf csa_tree_add_190_195_groupi_drc_bufs50269(csa_tree_add_190_195_groupi_n_2157 ,n_192);
  buf csa_tree_add_190_195_groupi_drc_bufs50270(csa_tree_add_190_195_groupi_n_2154 ,n_294);
  buf csa_tree_add_190_195_groupi_drc_bufs50271(csa_tree_add_190_195_groupi_n_1865 ,n_400);
  buf csa_tree_add_190_195_groupi_drc_bufs50272(csa_tree_add_190_195_groupi_n_2152 ,n_267);
  buf csa_tree_add_190_195_groupi_drc_bufs50273(csa_tree_add_190_195_groupi_n_1697 ,n_19);
  buf csa_tree_add_190_195_groupi_drc_bufs50274(csa_tree_add_190_195_groupi_n_1696 ,n_2);
  buf csa_tree_add_190_195_groupi_drc_bufs50275(csa_tree_add_190_195_groupi_n_1701 ,n_172);
  buf csa_tree_add_190_195_groupi_drc_bufs50276(csa_tree_add_190_195_groupi_n_1699 ,n_121);
  buf csa_tree_add_190_195_groupi_drc_bufs50277(csa_tree_add_190_195_groupi_n_1864 ,n_213);
  buf csa_tree_add_190_195_groupi_drc_bufs50278(csa_tree_add_190_195_groupi_n_2158 ,n_199);
  buf csa_tree_add_190_195_groupi_drc_bufs50279(csa_tree_add_190_195_groupi_n_1700 ,n_308);
  buf csa_tree_add_190_195_groupi_drc_bufs50280(csa_tree_add_190_195_groupi_n_1693 ,n_109);
  buf csa_tree_add_190_195_groupi_drc_bufs50281(csa_tree_add_190_195_groupi_n_1692 ,n_92);
  buf csa_tree_add_190_195_groupi_drc_bufs50282(csa_tree_add_190_195_groupi_n_2016 ,n_384);
  buf csa_tree_add_190_195_groupi_drc_bufs50283(csa_tree_add_190_195_groupi_n_1859 ,n_30);
  buf csa_tree_add_190_195_groupi_drc_bufs50284(csa_tree_add_190_195_groupi_n_1863 ,n_183);
  buf csa_tree_add_190_195_groupi_drc_bufs50285(csa_tree_add_190_195_groupi_n_2015 ,n_282);
  buf csa_tree_add_190_195_groupi_drc_bufs50286(csa_tree_add_190_195_groupi_n_1861 ,n_115);
  buf csa_tree_add_190_195_groupi_drc_bufs50287(csa_tree_add_190_195_groupi_n_2156 ,n_386);
  buf csa_tree_add_190_195_groupi_drc_bufs50288(csa_tree_add_190_195_groupi_n_1866 ,n_42);
  buf csa_tree_add_190_195_groupi_drc_bufs50289(csa_tree_add_190_195_groupi_n_1686 ,n_11);
  buf csa_tree_add_190_195_groupi_drc_bufs50290(csa_tree_add_190_195_groupi_n_1690 ,n_7);
  buf csa_tree_add_190_195_groupi_drc_bufs50291(csa_tree_add_190_195_groupi_n_1689 ,n_181);
  buf csa_tree_add_190_195_groupi_drc_bufs50292(csa_tree_add_190_195_groupi_n_1862 ,n_319);
  buf csa_tree_add_190_195_groupi_drc_bufs50293(csa_tree_add_190_195_groupi_n_1860 ,n_98);
  buf csa_tree_add_190_195_groupi_drc_bufs50294(csa_tree_add_190_195_groupi_n_1691 ,n_347);
  buf csa_tree_add_190_195_groupi_drc_bufs50295(csa_tree_add_190_195_groupi_n_1585 ,n_18);
  buf csa_tree_add_190_195_groupi_drc_bufs50296(csa_tree_add_190_195_groupi_n_1688 ,n_300);
  buf csa_tree_add_190_195_groupi_drc_bufs50297(csa_tree_add_190_195_groupi_n_2153 ,n_413);
  buf csa_tree_add_190_195_groupi_drc_bufs50298(csa_tree_add_190_195_groupi_n_1970 ,n_128);
  buf csa_tree_add_190_195_groupi_drc_bufs50299(csa_tree_add_190_195_groupi_n_1834 ,n_72);
  buf csa_tree_add_190_195_groupi_drc_bufs50300(csa_tree_add_190_195_groupi_n_1833 ,n_38);
  buf csa_tree_add_190_195_groupi_drc_bufs50301(csa_tree_add_190_195_groupi_n_1971 ,n_298);
  buf csa_tree_add_190_195_groupi_drc_bufs50302(csa_tree_add_190_195_groupi_n_1991 ,n_309);
  buf csa_tree_add_190_195_groupi_drc_bufs50303(csa_tree_add_190_195_groupi_n_1836 ,n_378);
  buf csa_tree_add_190_195_groupi_drc_bufs50304(csa_tree_add_190_195_groupi_n_1835 ,n_123);
  buf csa_tree_add_190_195_groupi_drc_bufs50306(csa_tree_add_190_195_groupi_n_1837 ,n_310);
  buf csa_tree_add_190_195_groupi_drc_bufs50307(csa_tree_add_190_195_groupi_n_2209 ,n_209);
  buf csa_tree_add_190_195_groupi_drc_bufs50308(csa_tree_add_190_195_groupi_n_1993 ,n_190);
  buf csa_tree_add_190_195_groupi_drc_bufs50309(csa_tree_add_190_195_groupi_n_1992 ,n_173);
  buf csa_tree_add_190_195_groupi_drc_bufs50310(csa_tree_add_190_195_groupi_n_1988 ,n_343);
  buf csa_tree_add_190_195_groupi_drc_bufs50311(csa_tree_add_190_195_groupi_n_1966 ,n_77);
  buf csa_tree_add_190_195_groupi_drc_bufs50314(csa_tree_add_190_195_groupi_n_2216 ,n_165);
  buf csa_tree_add_190_195_groupi_drc_bufs50319(csa_tree_add_190_195_groupi_n_1823 ,n_274);
  buf csa_tree_add_190_195_groupi_drc_bufs50321(csa_tree_add_190_195_groupi_n_1965 ,n_246);
  buf csa_tree_add_190_195_groupi_drc_bufs50322(csa_tree_add_190_195_groupi_n_1778 ,n_79);
  buf csa_tree_add_190_195_groupi_drc_bufs50323(csa_tree_add_190_195_groupi_n_1964 ,n_229);
  buf csa_tree_add_190_195_groupi_drc_bufs50324(csa_tree_add_190_195_groupi_n_1987 ,n_224);
  buf csa_tree_add_190_195_groupi_drc_bufs50325(csa_tree_add_190_195_groupi_n_2211 ,n_403);
  buf csa_tree_add_190_195_groupi_drc_bufs50326(csa_tree_add_190_195_groupi_n_2214 ,n_352);
  buf csa_tree_add_190_195_groupi_drc_bufs50327(csa_tree_add_190_195_groupi_n_1990 ,n_139);
  buf csa_tree_add_190_195_groupi_drc_bufs50328(csa_tree_add_190_195_groupi_n_1822 ,n_70);
  buf csa_tree_add_190_195_groupi_drc_bufs50329(csa_tree_add_190_195_groupi_n_1821 ,n_36);
  buf csa_tree_add_190_195_groupi_drc_bufs50330(csa_tree_add_190_195_groupi_n_1968 ,n_111);
  buf csa_tree_add_190_195_groupi_drc_bufs50333(csa_tree_add_190_195_groupi_n_1777 ,n_45);
  buf csa_tree_add_190_195_groupi_drc_bufs50334(csa_tree_add_190_195_groupi_n_1812 ,n_41);
  buf csa_tree_add_190_195_groupi_drc_bufs50335(csa_tree_add_190_195_groupi_n_2116 ,n_214);
  buf csa_tree_add_190_195_groupi_drc_bufs50339(csa_tree_add_190_195_groupi_n_1838 ,n_395);
  buf csa_tree_add_190_195_groupi_drc_bufs50340(csa_tree_add_190_195_groupi_n_2215 ,n_158);
  buf csa_tree_add_190_195_groupi_drc_bufs50341(csa_tree_add_190_195_groupi_n_1967 ,n_281);
  buf csa_tree_add_190_195_groupi_drc_bufs50347(csa_tree_add_190_195_groupi_n_1819 ,n_206);
  buf csa_tree_add_190_195_groupi_drc_bufs50348(csa_tree_add_190_195_groupi_n_1811 ,n_24);
  buf csa_tree_add_190_195_groupi_drc_bufs50349(csa_tree_add_190_195_groupi_n_1818 ,n_177);
  buf csa_tree_add_190_195_groupi_drc_bufs50350(csa_tree_add_190_195_groupi_n_2213 ,n_345);
  buf csa_tree_add_190_195_groupi_drc_bufs50351(csa_tree_add_190_195_groupi_n_1972 ,n_145);
  buf csa_tree_add_190_195_groupi_drc_bufs50352(csa_tree_add_190_195_groupi_n_1951 ,n_132);
  buf csa_tree_add_190_195_groupi_drc_bufs50354(csa_tree_add_190_195_groupi_n_1824 ,n_376);
  buf csa_tree_add_190_195_groupi_drc_bufs50355(csa_tree_add_190_195_groupi_n_1826 ,n_393);
  buf csa_tree_add_190_195_groupi_drc_bufs50356(csa_tree_add_190_195_groupi_n_1820 ,n_342);
  buf csa_tree_add_190_195_groupi_drc_bufs50357(csa_tree_add_190_195_groupi_n_1989 ,n_241);
  buf csa_tree_add_190_195_groupi_drc_bufs50358(csa_tree_add_190_195_groupi_n_1814 ,n_75);
  buf csa_tree_add_190_195_groupi_drc_bufs50359(csa_tree_add_190_195_groupi_n_1776 ,n_28);
  buf csa_tree_add_190_195_groupi_drc_bufs50360(csa_tree_add_190_195_groupi_n_1969 ,n_417);
  buf csa_tree_add_190_195_groupi_drc_bufs50361(csa_tree_add_190_195_groupi_n_1817 ,n_143);
  buf csa_tree_add_190_195_groupi_drc_bufs50362(csa_tree_add_190_195_groupi_n_1780 ,n_130);
  buf csa_tree_add_190_195_groupi_drc_bufs50371(csa_tree_add_190_195_groupi_n_1825 ,n_189);
  buf csa_tree_add_190_195_groupi_drc_bufs50372(csa_tree_add_190_195_groupi_n_1779 ,n_113);
  buf csa_tree_add_190_195_groupi_drc_bufs50373(csa_tree_add_190_195_groupi_n_1949 ,n_251);
  buf csa_tree_add_190_195_groupi_drc_bufs50374(csa_tree_add_190_195_groupi_n_2117 ,n_231);
  buf csa_tree_add_190_195_groupi_drc_bufs50375(csa_tree_add_190_195_groupi_n_2210 ,n_226);
  buf csa_tree_add_190_195_groupi_drc_bufs50376(csa_tree_add_190_195_groupi_n_1813 ,n_58);
  buf csa_tree_add_190_195_groupi_drc_bufs50377(csa_tree_add_190_195_groupi_n_1775 ,n_351);
  buf csa_tree_add_190_195_groupi_drc_bufs50378(csa_tree_add_190_195_groupi_n_2118 ,n_350);
  buf csa_tree_add_190_195_groupi_drc_bufs50379(csa_tree_add_190_195_groupi_n_1950 ,n_285);
  buf csa_tree_add_190_195_groupi_drc_bufs50380(csa_tree_add_190_195_groupi_n_1816 ,n_126);
  buf csa_tree_add_190_195_groupi_drc_bufs50382(csa_tree_add_190_195_groupi_n_2212 ,n_233);
  buf csa_tree_add_190_195_groupi_drc_bufs50383(csa_tree_add_190_195_groupi_n_2119 ,n_146);
  not csa_tree_add_190_195_groupi_drc_bufs50384(csa_tree_add_190_195_groupi_n_1189 ,csa_tree_add_190_195_groupi_n_1187);
  not csa_tree_add_190_195_groupi_drc_bufs50385(csa_tree_add_190_195_groupi_n_1188 ,csa_tree_add_190_195_groupi_n_1187);
  not csa_tree_add_190_195_groupi_drc_bufs50386(csa_tree_add_190_195_groupi_n_1187 ,csa_tree_add_190_195_groupi_n_2173);
  not csa_tree_add_190_195_groupi_drc_bufs50388(csa_tree_add_190_195_groupi_n_1186 ,csa_tree_add_190_195_groupi_n_1184);
  not csa_tree_add_190_195_groupi_drc_bufs50389(csa_tree_add_190_195_groupi_n_1185 ,csa_tree_add_190_195_groupi_n_1184);
  not csa_tree_add_190_195_groupi_drc_bufs50390(csa_tree_add_190_195_groupi_n_1184 ,csa_tree_add_190_195_groupi_n_2169);
  buf csa_tree_add_190_195_groupi_drc_bufs50408(csa_tree_add_190_195_groupi_n_1815 ,n_279);
  not csa_tree_add_190_195_groupi_drc_bufs50428(csa_tree_add_190_195_groupi_n_1183 ,csa_tree_add_190_195_groupi_n_1181);
  not csa_tree_add_190_195_groupi_drc_bufs50429(csa_tree_add_190_195_groupi_n_1182 ,csa_tree_add_190_195_groupi_n_1181);
  not csa_tree_add_190_195_groupi_drc_bufs50430(csa_tree_add_190_195_groupi_n_1181 ,csa_tree_add_190_195_groupi_n_2135);
  not csa_tree_add_190_195_groupi_drc_bufs50444(csa_tree_add_190_195_groupi_n_1180 ,csa_tree_add_190_195_groupi_n_1178);
  not csa_tree_add_190_195_groupi_drc_bufs50445(csa_tree_add_190_195_groupi_n_1179 ,csa_tree_add_190_195_groupi_n_1178);
  not csa_tree_add_190_195_groupi_drc_bufs50446(csa_tree_add_190_195_groupi_n_1178 ,csa_tree_add_190_195_groupi_n_2243);
  not csa_tree_add_190_195_groupi_drc_bufs50448(csa_tree_add_190_195_groupi_n_1177 ,csa_tree_add_190_195_groupi_n_1175);
  not csa_tree_add_190_195_groupi_drc_bufs50449(csa_tree_add_190_195_groupi_n_1176 ,csa_tree_add_190_195_groupi_n_1175);
  not csa_tree_add_190_195_groupi_drc_bufs50450(csa_tree_add_190_195_groupi_n_1175 ,csa_tree_add_190_195_groupi_n_2175);
  not csa_tree_add_190_195_groupi_drc_bufs50452(csa_tree_add_190_195_groupi_n_1174 ,csa_tree_add_190_195_groupi_n_1172);
  not csa_tree_add_190_195_groupi_drc_bufs50453(csa_tree_add_190_195_groupi_n_1173 ,csa_tree_add_190_195_groupi_n_1172);
  not csa_tree_add_190_195_groupi_drc_bufs50454(csa_tree_add_190_195_groupi_n_1172 ,csa_tree_add_190_195_groupi_n_2171);
  buf csa_tree_add_190_195_groupi_drc_bufs50461(csa_tree_add_190_195_groupi_n_1774 ,n_232);
  not csa_tree_add_190_195_groupi_drc_bufs50499(csa_tree_add_190_195_groupi_n_1171 ,csa_tree_add_190_195_groupi_n_1169);
  not csa_tree_add_190_195_groupi_drc_bufs50500(csa_tree_add_190_195_groupi_n_1170 ,csa_tree_add_190_195_groupi_n_1169);
  not csa_tree_add_190_195_groupi_drc_bufs50501(csa_tree_add_190_195_groupi_n_1169 ,csa_tree_add_190_195_groupi_n_2178);
  buf csa_tree_add_190_195_groupi_drc_bufs50503(csa_tree_add_190_195_groupi_n_1948 ,n_234);
  not csa_tree_add_190_195_groupi_drc_bufs50504(csa_tree_add_190_195_groupi_n_1168 ,csa_tree_add_190_195_groupi_n_1166);
  not csa_tree_add_190_195_groupi_drc_bufs50505(csa_tree_add_190_195_groupi_n_1167 ,csa_tree_add_190_195_groupi_n_1166);
  not csa_tree_add_190_195_groupi_drc_bufs50506(csa_tree_add_190_195_groupi_n_1166 ,csa_tree_add_190_195_groupi_n_2148);
  not csa_tree_add_190_195_groupi_drc_bufs50508(csa_tree_add_190_195_groupi_n_1165 ,csa_tree_add_190_195_groupi_n_1163);
  not csa_tree_add_190_195_groupi_drc_bufs50509(csa_tree_add_190_195_groupi_n_1164 ,csa_tree_add_190_195_groupi_n_1163);
  not csa_tree_add_190_195_groupi_drc_bufs50510(csa_tree_add_190_195_groupi_n_1163 ,csa_tree_add_190_195_groupi_n_1919);
  not csa_tree_add_190_195_groupi_drc_bufs50520(csa_tree_add_190_195_groupi_n_1162 ,csa_tree_add_190_195_groupi_n_1160);
  not csa_tree_add_190_195_groupi_drc_bufs50521(csa_tree_add_190_195_groupi_n_1161 ,csa_tree_add_190_195_groupi_n_1160);
  not csa_tree_add_190_195_groupi_drc_bufs50522(csa_tree_add_190_195_groupi_n_1160 ,csa_tree_add_190_195_groupi_n_2139);
  not csa_tree_add_190_195_groupi_drc_bufs50524(csa_tree_add_190_195_groupi_n_1159 ,csa_tree_add_190_195_groupi_n_1157);
  not csa_tree_add_190_195_groupi_drc_bufs50525(csa_tree_add_190_195_groupi_n_1158 ,csa_tree_add_190_195_groupi_n_1157);
  not csa_tree_add_190_195_groupi_drc_bufs50526(csa_tree_add_190_195_groupi_n_1157 ,csa_tree_add_190_195_groupi_n_1771);
  not csa_tree_add_190_195_groupi_drc_bufs50528(csa_tree_add_190_195_groupi_n_1156 ,csa_tree_add_190_195_groupi_n_1154);
  not csa_tree_add_190_195_groupi_drc_bufs50529(csa_tree_add_190_195_groupi_n_1155 ,csa_tree_add_190_195_groupi_n_1154);
  not csa_tree_add_190_195_groupi_drc_bufs50530(csa_tree_add_190_195_groupi_n_1154 ,csa_tree_add_190_195_groupi_n_2137);
  not csa_tree_add_190_195_groupi_drc_bufs50532(csa_tree_add_190_195_groupi_n_1153 ,csa_tree_add_190_195_groupi_n_1151);
  not csa_tree_add_190_195_groupi_drc_bufs50533(csa_tree_add_190_195_groupi_n_1152 ,csa_tree_add_190_195_groupi_n_1151);
  not csa_tree_add_190_195_groupi_drc_bufs50534(csa_tree_add_190_195_groupi_n_1151 ,csa_tree_add_190_195_groupi_n_2137);
  not csa_tree_add_190_195_groupi_drc_bufs50536(csa_tree_add_190_195_groupi_n_1150 ,csa_tree_add_190_195_groupi_n_1148);
  not csa_tree_add_190_195_groupi_drc_bufs50537(csa_tree_add_190_195_groupi_n_1149 ,csa_tree_add_190_195_groupi_n_1148);
  not csa_tree_add_190_195_groupi_drc_bufs50538(csa_tree_add_190_195_groupi_n_1148 ,csa_tree_add_190_195_groupi_n_2135);
  not csa_tree_add_190_195_groupi_drc_bufs50540(csa_tree_add_190_195_groupi_n_1147 ,csa_tree_add_190_195_groupi_n_1145);
  not csa_tree_add_190_195_groupi_drc_bufs50541(csa_tree_add_190_195_groupi_n_1146 ,csa_tree_add_190_195_groupi_n_1145);
  not csa_tree_add_190_195_groupi_drc_bufs50542(csa_tree_add_190_195_groupi_n_1145 ,csa_tree_add_190_195_groupi_n_2129);
  not csa_tree_add_190_195_groupi_drc_bufs50548(csa_tree_add_190_195_groupi_n_1144 ,csa_tree_add_190_195_groupi_n_1142);
  not csa_tree_add_190_195_groupi_drc_bufs50549(csa_tree_add_190_195_groupi_n_1143 ,csa_tree_add_190_195_groupi_n_1142);
  not csa_tree_add_190_195_groupi_drc_bufs50550(csa_tree_add_190_195_groupi_n_1142 ,csa_tree_add_190_195_groupi_n_2219);
  not csa_tree_add_190_195_groupi_drc_bufs50588(csa_tree_add_190_195_groupi_n_1141 ,csa_tree_add_190_195_groupi_n_1139);
  not csa_tree_add_190_195_groupi_drc_bufs50589(csa_tree_add_190_195_groupi_n_1140 ,csa_tree_add_190_195_groupi_n_1139);
  not csa_tree_add_190_195_groupi_drc_bufs50590(csa_tree_add_190_195_groupi_n_1139 ,csa_tree_add_190_195_groupi_n_2175);
  not csa_tree_add_190_195_groupi_drc_bufs50592(csa_tree_add_190_195_groupi_n_1138 ,csa_tree_add_190_195_groupi_n_1136);
  not csa_tree_add_190_195_groupi_drc_bufs50593(csa_tree_add_190_195_groupi_n_1137 ,csa_tree_add_190_195_groupi_n_1136);
  not csa_tree_add_190_195_groupi_drc_bufs50594(csa_tree_add_190_195_groupi_n_1136 ,csa_tree_add_190_195_groupi_n_2173);
  not csa_tree_add_190_195_groupi_drc_bufs50596(csa_tree_add_190_195_groupi_n_1135 ,csa_tree_add_190_195_groupi_n_1133);
  not csa_tree_add_190_195_groupi_drc_bufs50597(csa_tree_add_190_195_groupi_n_1134 ,csa_tree_add_190_195_groupi_n_1133);
  not csa_tree_add_190_195_groupi_drc_bufs50598(csa_tree_add_190_195_groupi_n_1133 ,csa_tree_add_190_195_groupi_n_2171);
  not csa_tree_add_190_195_groupi_drc_bufs50600(csa_tree_add_190_195_groupi_n_1132 ,csa_tree_add_190_195_groupi_n_1130);
  not csa_tree_add_190_195_groupi_drc_bufs50601(csa_tree_add_190_195_groupi_n_1131 ,csa_tree_add_190_195_groupi_n_1130);
  not csa_tree_add_190_195_groupi_drc_bufs50602(csa_tree_add_190_195_groupi_n_1130 ,csa_tree_add_190_195_groupi_n_2169);
  not csa_tree_add_190_195_groupi_drc_bufs50632(csa_tree_add_190_195_groupi_n_1129 ,csa_tree_add_190_195_groupi_n_1127);
  not csa_tree_add_190_195_groupi_drc_bufs50633(csa_tree_add_190_195_groupi_n_1128 ,csa_tree_add_190_195_groupi_n_1127);
  not csa_tree_add_190_195_groupi_drc_bufs50634(csa_tree_add_190_195_groupi_n_1127 ,csa_tree_add_190_195_groupi_n_2125);
  not csa_tree_add_190_195_groupi_drc_bufs50640(csa_tree_add_190_195_groupi_n_1126 ,csa_tree_add_190_195_groupi_n_1124);
  not csa_tree_add_190_195_groupi_drc_bufs50641(csa_tree_add_190_195_groupi_n_1125 ,csa_tree_add_190_195_groupi_n_1124);
  not csa_tree_add_190_195_groupi_drc_bufs50642(csa_tree_add_190_195_groupi_n_1124 ,csa_tree_add_190_195_groupi_n_2044);
  not csa_tree_add_190_195_groupi_drc_bufs50644(csa_tree_add_190_195_groupi_n_1123 ,csa_tree_add_190_195_groupi_n_1121);
  not csa_tree_add_190_195_groupi_drc_bufs50645(csa_tree_add_190_195_groupi_n_1122 ,csa_tree_add_190_195_groupi_n_1121);
  not csa_tree_add_190_195_groupi_drc_bufs50646(csa_tree_add_190_195_groupi_n_1121 ,csa_tree_add_190_195_groupi_n_1947);
  not csa_tree_add_190_195_groupi_drc_bufs50648(csa_tree_add_190_195_groupi_n_1120 ,csa_tree_add_190_195_groupi_n_1118);
  not csa_tree_add_190_195_groupi_drc_bufs50649(csa_tree_add_190_195_groupi_n_1119 ,csa_tree_add_190_195_groupi_n_1118);
  not csa_tree_add_190_195_groupi_drc_bufs50650(csa_tree_add_190_195_groupi_n_1118 ,csa_tree_add_190_195_groupi_n_2034);
  not csa_tree_add_190_195_groupi_drc_bufs50652(csa_tree_add_190_195_groupi_n_1117 ,csa_tree_add_190_195_groupi_n_1115);
  not csa_tree_add_190_195_groupi_drc_bufs50653(csa_tree_add_190_195_groupi_n_1116 ,csa_tree_add_190_195_groupi_n_1115);
  not csa_tree_add_190_195_groupi_drc_bufs50654(csa_tree_add_190_195_groupi_n_1115 ,csa_tree_add_190_195_groupi_n_2032);
  not csa_tree_add_190_195_groupi_drc_bufs50664(csa_tree_add_190_195_groupi_n_1114 ,csa_tree_add_190_195_groupi_n_1112);
  not csa_tree_add_190_195_groupi_drc_bufs50665(csa_tree_add_190_195_groupi_n_1113 ,csa_tree_add_190_195_groupi_n_1112);
  not csa_tree_add_190_195_groupi_drc_bufs50666(csa_tree_add_190_195_groupi_n_1112 ,csa_tree_add_190_195_groupi_n_2139);
  not csa_tree_add_190_195_groupi_drc_bufs50668(csa_tree_add_190_195_groupi_n_1111 ,csa_tree_add_190_195_groupi_n_1109);
  not csa_tree_add_190_195_groupi_drc_bufs50669(csa_tree_add_190_195_groupi_n_1110 ,csa_tree_add_190_195_groupi_n_1109);
  not csa_tree_add_190_195_groupi_drc_bufs50670(csa_tree_add_190_195_groupi_n_1109 ,csa_tree_add_190_195_groupi_n_2221);
  not csa_tree_add_190_195_groupi_drc_bufs50672(csa_tree_add_190_195_groupi_n_1108 ,csa_tree_add_190_195_groupi_n_1106);
  not csa_tree_add_190_195_groupi_drc_bufs50673(csa_tree_add_190_195_groupi_n_1107 ,csa_tree_add_190_195_groupi_n_1106);
  not csa_tree_add_190_195_groupi_drc_bufs50674(csa_tree_add_190_195_groupi_n_1106 ,csa_tree_add_190_195_groupi_n_1771);
  not csa_tree_add_190_195_groupi_drc_bufs50676(csa_tree_add_190_195_groupi_n_1105 ,csa_tree_add_190_195_groupi_n_1103);
  not csa_tree_add_190_195_groupi_drc_bufs50677(csa_tree_add_190_195_groupi_n_1104 ,csa_tree_add_190_195_groupi_n_1103);
  not csa_tree_add_190_195_groupi_drc_bufs50678(csa_tree_add_190_195_groupi_n_1103 ,csa_tree_add_190_195_groupi_n_2129);
  not csa_tree_add_190_195_groupi_drc_bufs50696(csa_tree_add_190_195_groupi_n_1102 ,csa_tree_add_190_195_groupi_n_1100);
  not csa_tree_add_190_195_groupi_drc_bufs50697(csa_tree_add_190_195_groupi_n_1101 ,csa_tree_add_190_195_groupi_n_1100);
  not csa_tree_add_190_195_groupi_drc_bufs50698(csa_tree_add_190_195_groupi_n_1100 ,csa_tree_add_190_195_groupi_n_2239);
  not csa_tree_add_190_195_groupi_drc_bufs50716(csa_tree_add_190_195_groupi_n_1099 ,csa_tree_add_190_195_groupi_n_1097);
  not csa_tree_add_190_195_groupi_drc_bufs50717(csa_tree_add_190_195_groupi_n_1098 ,csa_tree_add_190_195_groupi_n_1097);
  not csa_tree_add_190_195_groupi_drc_bufs50718(csa_tree_add_190_195_groupi_n_1097 ,csa_tree_add_190_195_groupi_n_1986);
  not csa_tree_add_190_195_groupi_drc_bufs50724(csa_tree_add_190_195_groupi_n_1096 ,csa_tree_add_190_195_groupi_n_1094);
  not csa_tree_add_190_195_groupi_drc_bufs50725(csa_tree_add_190_195_groupi_n_1095 ,csa_tree_add_190_195_groupi_n_1094);
  not csa_tree_add_190_195_groupi_drc_bufs50726(csa_tree_add_190_195_groupi_n_1094 ,csa_tree_add_190_195_groupi_n_1980);
  not csa_tree_add_190_195_groupi_drc_bufs50732(csa_tree_add_190_195_groupi_n_1093 ,csa_tree_add_190_195_groupi_n_1091);
  not csa_tree_add_190_195_groupi_drc_bufs50733(csa_tree_add_190_195_groupi_n_1092 ,csa_tree_add_190_195_groupi_n_1091);
  not csa_tree_add_190_195_groupi_drc_bufs50734(csa_tree_add_190_195_groupi_n_1091 ,csa_tree_add_190_195_groupi_n_1953);
  not csa_tree_add_190_195_groupi_drc_bufs50736(csa_tree_add_190_195_groupi_n_1090 ,csa_tree_add_190_195_groupi_n_1088);
  not csa_tree_add_190_195_groupi_drc_bufs50737(csa_tree_add_190_195_groupi_n_1089 ,csa_tree_add_190_195_groupi_n_1088);
  not csa_tree_add_190_195_groupi_drc_bufs50738(csa_tree_add_190_195_groupi_n_1088 ,csa_tree_add_190_195_groupi_n_2112);
  not csa_tree_add_190_195_groupi_drc_bufs50740(csa_tree_add_190_195_groupi_n_1087 ,csa_tree_add_190_195_groupi_n_1085);
  not csa_tree_add_190_195_groupi_drc_bufs50741(csa_tree_add_190_195_groupi_n_1086 ,csa_tree_add_190_195_groupi_n_1085);
  not csa_tree_add_190_195_groupi_drc_bufs50742(csa_tree_add_190_195_groupi_n_1085 ,csa_tree_add_190_195_groupi_n_2109);
  not csa_tree_add_190_195_groupi_drc_bufs50744(csa_tree_add_190_195_groupi_n_1084 ,csa_tree_add_190_195_groupi_n_1082);
  not csa_tree_add_190_195_groupi_drc_bufs50745(csa_tree_add_190_195_groupi_n_1083 ,csa_tree_add_190_195_groupi_n_1082);
  not csa_tree_add_190_195_groupi_drc_bufs50746(csa_tree_add_190_195_groupi_n_1082 ,csa_tree_add_190_195_groupi_n_1794);
  not csa_tree_add_190_195_groupi_drc_bufs50748(csa_tree_add_190_195_groupi_n_1081 ,csa_tree_add_190_195_groupi_n_1079);
  not csa_tree_add_190_195_groupi_drc_bufs50749(csa_tree_add_190_195_groupi_n_1080 ,csa_tree_add_190_195_groupi_n_1079);
  not csa_tree_add_190_195_groupi_drc_bufs50750(csa_tree_add_190_195_groupi_n_1079 ,csa_tree_add_190_195_groupi_n_1786);
  not csa_tree_add_190_195_groupi_drc_bufs50752(csa_tree_add_190_195_groupi_n_1078 ,csa_tree_add_190_195_groupi_n_1076);
  not csa_tree_add_190_195_groupi_drc_bufs50753(csa_tree_add_190_195_groupi_n_1077 ,csa_tree_add_190_195_groupi_n_1076);
  not csa_tree_add_190_195_groupi_drc_bufs50754(csa_tree_add_190_195_groupi_n_1076 ,csa_tree_add_190_195_groupi_n_2180);
  not csa_tree_add_190_195_groupi_drc_bufs50764(csa_tree_add_190_195_groupi_n_1075 ,csa_tree_add_190_195_groupi_n_1073);
  not csa_tree_add_190_195_groupi_drc_bufs50765(csa_tree_add_190_195_groupi_n_1074 ,csa_tree_add_190_195_groupi_n_1073);
  not csa_tree_add_190_195_groupi_drc_bufs50766(csa_tree_add_190_195_groupi_n_1073 ,csa_tree_add_190_195_groupi_n_2038);
  not csa_tree_add_190_195_groupi_drc_bufs50776(csa_tree_add_190_195_groupi_n_1072 ,csa_tree_add_190_195_groupi_n_1070);
  not csa_tree_add_190_195_groupi_drc_bufs50777(csa_tree_add_190_195_groupi_n_1071 ,csa_tree_add_190_195_groupi_n_1070);
  not csa_tree_add_190_195_groupi_drc_bufs50778(csa_tree_add_190_195_groupi_n_1070 ,csa_tree_add_190_195_groupi_n_2160);
  not csa_tree_add_190_195_groupi_drc_bufs50780(csa_tree_add_190_195_groupi_n_1069 ,csa_tree_add_190_195_groupi_n_1067);
  not csa_tree_add_190_195_groupi_drc_bufs50781(csa_tree_add_190_195_groupi_n_1068 ,csa_tree_add_190_195_groupi_n_1067);
  not csa_tree_add_190_195_groupi_drc_bufs50782(csa_tree_add_190_195_groupi_n_1067 ,csa_tree_add_190_195_groupi_n_2046);
  not csa_tree_add_190_195_groupi_drc_bufs50784(csa_tree_add_190_195_groupi_n_1066 ,csa_tree_add_190_195_groupi_n_1064);
  not csa_tree_add_190_195_groupi_drc_bufs50785(csa_tree_add_190_195_groupi_n_1065 ,csa_tree_add_190_195_groupi_n_1064);
  not csa_tree_add_190_195_groupi_drc_bufs50786(csa_tree_add_190_195_groupi_n_1064 ,csa_tree_add_190_195_groupi_n_2046);
  not csa_tree_add_190_195_groupi_drc_bufs50788(csa_tree_add_190_195_groupi_n_1063 ,csa_tree_add_190_195_groupi_n_1061);
  not csa_tree_add_190_195_groupi_drc_bufs50789(csa_tree_add_190_195_groupi_n_1062 ,csa_tree_add_190_195_groupi_n_1061);
  not csa_tree_add_190_195_groupi_drc_bufs50790(csa_tree_add_190_195_groupi_n_1061 ,csa_tree_add_190_195_groupi_n_2036);
  not csa_tree_add_190_195_groupi_drc_bufs50792(csa_tree_add_190_195_groupi_n_1060 ,csa_tree_add_190_195_groupi_n_1058);
  not csa_tree_add_190_195_groupi_drc_bufs50793(csa_tree_add_190_195_groupi_n_1059 ,csa_tree_add_190_195_groupi_n_1058);
  not csa_tree_add_190_195_groupi_drc_bufs50794(csa_tree_add_190_195_groupi_n_1058 ,csa_tree_add_190_195_groupi_n_2036);
  not csa_tree_add_190_195_groupi_drc_bufs50804(csa_tree_add_190_195_groupi_n_1057 ,csa_tree_add_190_195_groupi_n_1055);
  not csa_tree_add_190_195_groupi_drc_bufs50805(csa_tree_add_190_195_groupi_n_1056 ,csa_tree_add_190_195_groupi_n_1055);
  not csa_tree_add_190_195_groupi_drc_bufs50806(csa_tree_add_190_195_groupi_n_1055 ,csa_tree_add_190_195_groupi_n_2034);
  not csa_tree_add_190_195_groupi_drc_bufs50808(csa_tree_add_190_195_groupi_n_1054 ,csa_tree_add_190_195_groupi_n_1052);
  not csa_tree_add_190_195_groupi_drc_bufs50809(csa_tree_add_190_195_groupi_n_1053 ,csa_tree_add_190_195_groupi_n_1052);
  not csa_tree_add_190_195_groupi_drc_bufs50810(csa_tree_add_190_195_groupi_n_1052 ,csa_tree_add_190_195_groupi_n_2032);
  not csa_tree_add_190_195_groupi_drc_bufs50820(csa_tree_add_190_195_groupi_n_1051 ,csa_tree_add_190_195_groupi_n_1049);
  not csa_tree_add_190_195_groupi_drc_bufs50821(csa_tree_add_190_195_groupi_n_1050 ,csa_tree_add_190_195_groupi_n_1049);
  not csa_tree_add_190_195_groupi_drc_bufs50822(csa_tree_add_190_195_groupi_n_1049 ,csa_tree_add_190_195_groupi_n_1926);
  not csa_tree_add_190_195_groupi_drc_bufs50828(csa_tree_add_190_195_groupi_n_1048 ,csa_tree_add_190_195_groupi_n_1046);
  not csa_tree_add_190_195_groupi_drc_bufs50829(csa_tree_add_190_195_groupi_n_1047 ,csa_tree_add_190_195_groupi_n_1046);
  not csa_tree_add_190_195_groupi_drc_bufs50830(csa_tree_add_190_195_groupi_n_1046 ,csa_tree_add_190_195_groupi_n_1913);
  not csa_tree_add_190_195_groupi_drc_bufs50832(csa_tree_add_190_195_groupi_n_1045 ,csa_tree_add_190_195_groupi_n_1043);
  not csa_tree_add_190_195_groupi_drc_bufs50833(csa_tree_add_190_195_groupi_n_1044 ,csa_tree_add_190_195_groupi_n_1043);
  not csa_tree_add_190_195_groupi_drc_bufs50834(csa_tree_add_190_195_groupi_n_1043 ,csa_tree_add_190_195_groupi_n_2143);
  not csa_tree_add_190_195_groupi_drc_bufs50836(csa_tree_add_190_195_groupi_n_1042 ,csa_tree_add_190_195_groupi_n_1040);
  not csa_tree_add_190_195_groupi_drc_bufs50837(csa_tree_add_190_195_groupi_n_1041 ,csa_tree_add_190_195_groupi_n_1040);
  not csa_tree_add_190_195_groupi_drc_bufs50838(csa_tree_add_190_195_groupi_n_1040 ,csa_tree_add_190_195_groupi_n_1769);
  not csa_tree_add_190_195_groupi_drc_bufs50840(csa_tree_add_190_195_groupi_n_1039 ,csa_tree_add_190_195_groupi_n_1037);
  not csa_tree_add_190_195_groupi_drc_bufs50841(csa_tree_add_190_195_groupi_n_1038 ,csa_tree_add_190_195_groupi_n_1037);
  not csa_tree_add_190_195_groupi_drc_bufs50842(csa_tree_add_190_195_groupi_n_1037 ,csa_tree_add_190_195_groupi_n_2141);
  not csa_tree_add_190_195_groupi_drc_bufs50844(csa_tree_add_190_195_groupi_n_1036 ,csa_tree_add_190_195_groupi_n_1034);
  not csa_tree_add_190_195_groupi_drc_bufs50845(csa_tree_add_190_195_groupi_n_1035 ,csa_tree_add_190_195_groupi_n_1034);
  not csa_tree_add_190_195_groupi_drc_bufs50846(csa_tree_add_190_195_groupi_n_1034 ,csa_tree_add_190_195_groupi_n_2141);
  not csa_tree_add_190_195_groupi_drc_bufs50848(csa_tree_add_190_195_groupi_n_1033 ,csa_tree_add_190_195_groupi_n_1031);
  not csa_tree_add_190_195_groupi_drc_bufs50849(csa_tree_add_190_195_groupi_n_1032 ,csa_tree_add_190_195_groupi_n_1031);
  not csa_tree_add_190_195_groupi_drc_bufs50850(csa_tree_add_190_195_groupi_n_1031 ,csa_tree_add_190_195_groupi_n_2225);
  not csa_tree_add_190_195_groupi_drc_bufs50852(csa_tree_add_190_195_groupi_n_1030 ,csa_tree_add_190_195_groupi_n_1028);
  not csa_tree_add_190_195_groupi_drc_bufs50853(csa_tree_add_190_195_groupi_n_1029 ,csa_tree_add_190_195_groupi_n_1028);
  not csa_tree_add_190_195_groupi_drc_bufs50854(csa_tree_add_190_195_groupi_n_1028 ,csa_tree_add_190_195_groupi_n_1875);
  not csa_tree_add_190_195_groupi_drc_bufs50856(csa_tree_add_190_195_groupi_n_1027 ,csa_tree_add_190_195_groupi_n_1025);
  not csa_tree_add_190_195_groupi_drc_bufs50857(csa_tree_add_190_195_groupi_n_1026 ,csa_tree_add_190_195_groupi_n_1025);
  not csa_tree_add_190_195_groupi_drc_bufs50858(csa_tree_add_190_195_groupi_n_1025 ,csa_tree_add_190_195_groupi_n_2131);
  not csa_tree_add_190_195_groupi_drc_bufs50860(csa_tree_add_190_195_groupi_n_1024 ,csa_tree_add_190_195_groupi_n_1022);
  not csa_tree_add_190_195_groupi_drc_bufs50861(csa_tree_add_190_195_groupi_n_1023 ,csa_tree_add_190_195_groupi_n_1022);
  not csa_tree_add_190_195_groupi_drc_bufs50862(csa_tree_add_190_195_groupi_n_1022 ,csa_tree_add_190_195_groupi_n_2127);
  not csa_tree_add_190_195_groupi_drc_bufs50864(csa_tree_add_190_195_groupi_n_1021 ,csa_tree_add_190_195_groupi_n_1019);
  not csa_tree_add_190_195_groupi_drc_bufs50865(csa_tree_add_190_195_groupi_n_1020 ,csa_tree_add_190_195_groupi_n_1019);
  not csa_tree_add_190_195_groupi_drc_bufs50866(csa_tree_add_190_195_groupi_n_1019 ,csa_tree_add_190_195_groupi_n_1879);
  not csa_tree_add_190_195_groupi_drc_bufs50868(csa_tree_add_190_195_groupi_n_1018 ,csa_tree_add_190_195_groupi_n_1016);
  not csa_tree_add_190_195_groupi_drc_bufs50869(csa_tree_add_190_195_groupi_n_1017 ,csa_tree_add_190_195_groupi_n_1016);
  not csa_tree_add_190_195_groupi_drc_bufs50870(csa_tree_add_190_195_groupi_n_1016 ,csa_tree_add_190_195_groupi_n_2133);
  not csa_tree_add_190_195_groupi_drc_bufs50872(csa_tree_add_190_195_groupi_n_1015 ,csa_tree_add_190_195_groupi_n_1013);
  not csa_tree_add_190_195_groupi_drc_bufs50873(csa_tree_add_190_195_groupi_n_1014 ,csa_tree_add_190_195_groupi_n_1013);
  not csa_tree_add_190_195_groupi_drc_bufs50874(csa_tree_add_190_195_groupi_n_1013 ,csa_tree_add_190_195_groupi_n_2133);
  not csa_tree_add_190_195_groupi_drc_bufs50884(csa_tree_add_190_195_groupi_n_1012 ,csa_tree_add_190_195_groupi_n_1010);
  not csa_tree_add_190_195_groupi_drc_bufs50885(csa_tree_add_190_195_groupi_n_1011 ,csa_tree_add_190_195_groupi_n_1010);
  not csa_tree_add_190_195_groupi_drc_bufs50886(csa_tree_add_190_195_groupi_n_1010 ,csa_tree_add_190_195_groupi_n_2245);
  not csa_tree_add_190_195_groupi_drc_bufs50888(csa_tree_add_190_195_groupi_n_1009 ,csa_tree_add_190_195_groupi_n_1007);
  not csa_tree_add_190_195_groupi_drc_bufs50889(csa_tree_add_190_195_groupi_n_1008 ,csa_tree_add_190_195_groupi_n_1007);
  not csa_tree_add_190_195_groupi_drc_bufs50890(csa_tree_add_190_195_groupi_n_1007 ,csa_tree_add_190_195_groupi_n_1732);
  not csa_tree_add_190_195_groupi_drc_bufs50900(csa_tree_add_190_195_groupi_n_1006 ,csa_tree_add_190_195_groupi_n_1004);
  not csa_tree_add_190_195_groupi_drc_bufs50901(csa_tree_add_190_195_groupi_n_1005 ,csa_tree_add_190_195_groupi_n_1004);
  not csa_tree_add_190_195_groupi_drc_bufs50902(csa_tree_add_190_195_groupi_n_1004 ,csa_tree_add_190_195_groupi_n_1737);
  not csa_tree_add_190_195_groupi_drc_bufs50904(csa_tree_add_190_195_groupi_n_1003 ,csa_tree_add_190_195_groupi_n_1001);
  not csa_tree_add_190_195_groupi_drc_bufs50905(csa_tree_add_190_195_groupi_n_1002 ,csa_tree_add_190_195_groupi_n_1001);
  not csa_tree_add_190_195_groupi_drc_bufs50906(csa_tree_add_190_195_groupi_n_1001 ,csa_tree_add_190_195_groupi_n_1740);
  not csa_tree_add_190_195_groupi_drc_bufs50908(csa_tree_add_190_195_groupi_n_1000 ,csa_tree_add_190_195_groupi_n_998);
  not csa_tree_add_190_195_groupi_drc_bufs50909(csa_tree_add_190_195_groupi_n_999 ,csa_tree_add_190_195_groupi_n_998);
  not csa_tree_add_190_195_groupi_drc_bufs50910(csa_tree_add_190_195_groupi_n_998 ,csa_tree_add_190_195_groupi_n_2146);
  not csa_tree_add_190_195_groupi_drc_bufs50912(csa_tree_add_190_195_groupi_n_997 ,csa_tree_add_190_195_groupi_n_995);
  not csa_tree_add_190_195_groupi_drc_bufs50913(csa_tree_add_190_195_groupi_n_996 ,csa_tree_add_190_195_groupi_n_995);
  not csa_tree_add_190_195_groupi_drc_bufs50914(csa_tree_add_190_195_groupi_n_995 ,csa_tree_add_190_195_groupi_n_1858);
  not csa_tree_add_190_195_groupi_drc_bufs50916(csa_tree_add_190_195_groupi_n_994 ,csa_tree_add_190_195_groupi_n_992);
  not csa_tree_add_190_195_groupi_drc_bufs50917(csa_tree_add_190_195_groupi_n_993 ,csa_tree_add_190_195_groupi_n_992);
  not csa_tree_add_190_195_groupi_drc_bufs50918(csa_tree_add_190_195_groupi_n_992 ,csa_tree_add_190_195_groupi_n_1982);
  not csa_tree_add_190_195_groupi_drc_bufs50920(csa_tree_add_190_195_groupi_n_991 ,csa_tree_add_190_195_groupi_n_989);
  not csa_tree_add_190_195_groupi_drc_bufs50921(csa_tree_add_190_195_groupi_n_990 ,csa_tree_add_190_195_groupi_n_989);
  not csa_tree_add_190_195_groupi_drc_bufs50922(csa_tree_add_190_195_groupi_n_989 ,csa_tree_add_190_195_groupi_n_1955);
  not csa_tree_add_190_195_groupi_drc_bufs50924(csa_tree_add_190_195_groupi_n_988 ,csa_tree_add_190_195_groupi_n_986);
  not csa_tree_add_190_195_groupi_drc_bufs50925(csa_tree_add_190_195_groupi_n_987 ,csa_tree_add_190_195_groupi_n_986);
  not csa_tree_add_190_195_groupi_drc_bufs50926(csa_tree_add_190_195_groupi_n_986 ,csa_tree_add_190_195_groupi_n_1980);
  not csa_tree_add_190_195_groupi_drc_bufs50928(csa_tree_add_190_195_groupi_n_985 ,csa_tree_add_190_195_groupi_n_983);
  not csa_tree_add_190_195_groupi_drc_bufs50929(csa_tree_add_190_195_groupi_n_984 ,csa_tree_add_190_195_groupi_n_983);
  not csa_tree_add_190_195_groupi_drc_bufs50930(csa_tree_add_190_195_groupi_n_983 ,csa_tree_add_190_195_groupi_n_1959);
  not csa_tree_add_190_195_groupi_drc_bufs50932(csa_tree_add_190_195_groupi_n_982 ,csa_tree_add_190_195_groupi_n_980);
  not csa_tree_add_190_195_groupi_drc_bufs50933(csa_tree_add_190_195_groupi_n_981 ,csa_tree_add_190_195_groupi_n_980);
  not csa_tree_add_190_195_groupi_drc_bufs50934(csa_tree_add_190_195_groupi_n_980 ,csa_tree_add_190_195_groupi_n_1959);
  not csa_tree_add_190_195_groupi_drc_bufs50936(csa_tree_add_190_195_groupi_n_979 ,csa_tree_add_190_195_groupi_n_977);
  not csa_tree_add_190_195_groupi_drc_bufs50937(csa_tree_add_190_195_groupi_n_978 ,csa_tree_add_190_195_groupi_n_977);
  not csa_tree_add_190_195_groupi_drc_bufs50938(csa_tree_add_190_195_groupi_n_977 ,csa_tree_add_190_195_groupi_n_2410);
  not csa_tree_add_190_195_groupi_drc_bufs50940(csa_tree_add_190_195_groupi_n_976 ,csa_tree_add_190_195_groupi_n_974);
  not csa_tree_add_190_195_groupi_drc_bufs50941(csa_tree_add_190_195_groupi_n_975 ,csa_tree_add_190_195_groupi_n_974);
  not csa_tree_add_190_195_groupi_drc_bufs50942(csa_tree_add_190_195_groupi_n_974 ,csa_tree_add_190_195_groupi_n_2066);
  not csa_tree_add_190_195_groupi_drc_bufs50944(csa_tree_add_190_195_groupi_n_973 ,csa_tree_add_190_195_groupi_n_971);
  not csa_tree_add_190_195_groupi_drc_bufs50945(csa_tree_add_190_195_groupi_n_972 ,csa_tree_add_190_195_groupi_n_971);
  not csa_tree_add_190_195_groupi_drc_bufs50946(csa_tree_add_190_195_groupi_n_971 ,csa_tree_add_190_195_groupi_n_1807);
  not csa_tree_add_190_195_groupi_drc_bufs50948(csa_tree_add_190_195_groupi_n_970 ,csa_tree_add_190_195_groupi_n_968);
  not csa_tree_add_190_195_groupi_drc_bufs50949(csa_tree_add_190_195_groupi_n_969 ,csa_tree_add_190_195_groupi_n_968);
  not csa_tree_add_190_195_groupi_drc_bufs50950(csa_tree_add_190_195_groupi_n_968 ,csa_tree_add_190_195_groupi_n_1803);
  not csa_tree_add_190_195_groupi_drc_bufs50952(csa_tree_add_190_195_groupi_n_967 ,csa_tree_add_190_195_groupi_n_965);
  not csa_tree_add_190_195_groupi_drc_bufs50953(csa_tree_add_190_195_groupi_n_966 ,csa_tree_add_190_195_groupi_n_965);
  not csa_tree_add_190_195_groupi_drc_bufs50954(csa_tree_add_190_195_groupi_n_965 ,csa_tree_add_190_195_groupi_n_1783);
  not csa_tree_add_190_195_groupi_drc_bufs50956(csa_tree_add_190_195_groupi_n_964 ,csa_tree_add_190_195_groupi_n_962);
  not csa_tree_add_190_195_groupi_drc_bufs50957(csa_tree_add_190_195_groupi_n_963 ,csa_tree_add_190_195_groupi_n_962);
  not csa_tree_add_190_195_groupi_drc_bufs50958(csa_tree_add_190_195_groupi_n_962 ,csa_tree_add_190_195_groupi_n_2114);
  not csa_tree_add_190_195_groupi_drc_bufs50960(csa_tree_add_190_195_groupi_n_961 ,csa_tree_add_190_195_groupi_n_959);
  not csa_tree_add_190_195_groupi_drc_bufs50961(csa_tree_add_190_195_groupi_n_960 ,csa_tree_add_190_195_groupi_n_959);
  not csa_tree_add_190_195_groupi_drc_bufs50962(csa_tree_add_190_195_groupi_n_959 ,csa_tree_add_190_195_groupi_n_2105);
  not csa_tree_add_190_195_groupi_drc_bufs50964(csa_tree_add_190_195_groupi_n_958 ,csa_tree_add_190_195_groupi_n_956);
  not csa_tree_add_190_195_groupi_drc_bufs50965(csa_tree_add_190_195_groupi_n_957 ,csa_tree_add_190_195_groupi_n_956);
  not csa_tree_add_190_195_groupi_drc_bufs50966(csa_tree_add_190_195_groupi_n_956 ,csa_tree_add_190_195_groupi_n_1788);
  not csa_tree_add_190_195_groupi_drc_bufs50968(csa_tree_add_190_195_groupi_n_955 ,csa_tree_add_190_195_groupi_n_953);
  not csa_tree_add_190_195_groupi_drc_bufs50969(csa_tree_add_190_195_groupi_n_954 ,csa_tree_add_190_195_groupi_n_953);
  not csa_tree_add_190_195_groupi_drc_bufs50970(csa_tree_add_190_195_groupi_n_953 ,csa_tree_add_190_195_groupi_n_1800);
  not csa_tree_add_190_195_groupi_drc_bufs50972(csa_tree_add_190_195_groupi_n_952 ,csa_tree_add_190_195_groupi_n_950);
  not csa_tree_add_190_195_groupi_drc_bufs50973(csa_tree_add_190_195_groupi_n_951 ,csa_tree_add_190_195_groupi_n_950);
  not csa_tree_add_190_195_groupi_drc_bufs50974(csa_tree_add_190_195_groupi_n_950 ,csa_tree_add_190_195_groupi_n_2048);
  not csa_tree_add_190_195_groupi_drc_bufs50992(csa_tree_add_190_195_groupi_n_949 ,csa_tree_add_190_195_groupi_n_947);
  not csa_tree_add_190_195_groupi_drc_bufs50993(csa_tree_add_190_195_groupi_n_948 ,csa_tree_add_190_195_groupi_n_947);
  not csa_tree_add_190_195_groupi_drc_bufs50994(csa_tree_add_190_195_groupi_n_947 ,csa_tree_add_190_195_groupi_n_2163);
  not csa_tree_add_190_195_groupi_drc_bufs50996(csa_tree_add_190_195_groupi_n_946 ,csa_tree_add_190_195_groupi_n_944);
  not csa_tree_add_190_195_groupi_drc_bufs50997(csa_tree_add_190_195_groupi_n_945 ,csa_tree_add_190_195_groupi_n_944);
  not csa_tree_add_190_195_groupi_drc_bufs50998(csa_tree_add_190_195_groupi_n_944 ,csa_tree_add_190_195_groupi_n_2044);
  not csa_tree_add_190_195_groupi_drc_bufs51000(csa_tree_add_190_195_groupi_n_943 ,csa_tree_add_190_195_groupi_n_941);
  not csa_tree_add_190_195_groupi_drc_bufs51001(csa_tree_add_190_195_groupi_n_942 ,csa_tree_add_190_195_groupi_n_941);
  not csa_tree_add_190_195_groupi_drc_bufs51002(csa_tree_add_190_195_groupi_n_941 ,csa_tree_add_190_195_groupi_n_2038);
  not csa_tree_add_190_195_groupi_drc_bufs51004(csa_tree_add_190_195_groupi_n_940 ,csa_tree_add_190_195_groupi_n_938);
  not csa_tree_add_190_195_groupi_drc_bufs51005(csa_tree_add_190_195_groupi_n_939 ,csa_tree_add_190_195_groupi_n_938);
  not csa_tree_add_190_195_groupi_drc_bufs51006(csa_tree_add_190_195_groupi_n_938 ,csa_tree_add_190_195_groupi_n_2030);
  not csa_tree_add_190_195_groupi_drc_bufs51008(csa_tree_add_190_195_groupi_n_937 ,csa_tree_add_190_195_groupi_n_935);
  not csa_tree_add_190_195_groupi_drc_bufs51009(csa_tree_add_190_195_groupi_n_936 ,csa_tree_add_190_195_groupi_n_935);
  not csa_tree_add_190_195_groupi_drc_bufs51010(csa_tree_add_190_195_groupi_n_935 ,csa_tree_add_190_195_groupi_n_2030);
  not csa_tree_add_190_195_groupi_drc_bufs51012(csa_tree_add_190_195_groupi_n_934 ,csa_tree_add_190_195_groupi_n_932);
  not csa_tree_add_190_195_groupi_drc_bufs51013(csa_tree_add_190_195_groupi_n_933 ,csa_tree_add_190_195_groupi_n_932);
  not csa_tree_add_190_195_groupi_drc_bufs51014(csa_tree_add_190_195_groupi_n_932 ,csa_tree_add_190_195_groupi_n_1947);
  not csa_tree_add_190_195_groupi_drc_bufs51016(csa_tree_add_190_195_groupi_n_931 ,csa_tree_add_190_195_groupi_n_929);
  not csa_tree_add_190_195_groupi_drc_bufs51017(csa_tree_add_190_195_groupi_n_930 ,csa_tree_add_190_195_groupi_n_929);
  not csa_tree_add_190_195_groupi_drc_bufs51018(csa_tree_add_190_195_groupi_n_929 ,csa_tree_add_190_195_groupi_n_2148);
  not csa_tree_add_190_195_groupi_drc_bufs51024(csa_tree_add_190_195_groupi_n_928 ,csa_tree_add_190_195_groupi_n_926);
  not csa_tree_add_190_195_groupi_drc_bufs51025(csa_tree_add_190_195_groupi_n_927 ,csa_tree_add_190_195_groupi_n_926);
  not csa_tree_add_190_195_groupi_drc_bufs51026(csa_tree_add_190_195_groupi_n_926 ,csa_tree_add_190_195_groupi_n_1773);
  not csa_tree_add_190_195_groupi_drc_bufs51028(csa_tree_add_190_195_groupi_n_925 ,csa_tree_add_190_195_groupi_n_923);
  not csa_tree_add_190_195_groupi_drc_bufs51029(csa_tree_add_190_195_groupi_n_924 ,csa_tree_add_190_195_groupi_n_923);
  not csa_tree_add_190_195_groupi_drc_bufs51030(csa_tree_add_190_195_groupi_n_923 ,csa_tree_add_190_195_groupi_n_2143);
  not csa_tree_add_190_195_groupi_drc_bufs51032(csa_tree_add_190_195_groupi_n_922 ,csa_tree_add_190_195_groupi_n_920);
  not csa_tree_add_190_195_groupi_drc_bufs51033(csa_tree_add_190_195_groupi_n_921 ,csa_tree_add_190_195_groupi_n_920);
  not csa_tree_add_190_195_groupi_drc_bufs51034(csa_tree_add_190_195_groupi_n_920 ,csa_tree_add_190_195_groupi_n_1885);
  not csa_tree_add_190_195_groupi_drc_bufs51036(csa_tree_add_190_195_groupi_n_919 ,csa_tree_add_190_195_groupi_n_917);
  not csa_tree_add_190_195_groupi_drc_bufs51037(csa_tree_add_190_195_groupi_n_918 ,csa_tree_add_190_195_groupi_n_917);
  not csa_tree_add_190_195_groupi_drc_bufs51038(csa_tree_add_190_195_groupi_n_917 ,csa_tree_add_190_195_groupi_n_1882);
  not csa_tree_add_190_195_groupi_drc_bufs51040(csa_tree_add_190_195_groupi_n_916 ,csa_tree_add_190_195_groupi_n_914);
  not csa_tree_add_190_195_groupi_drc_bufs51041(csa_tree_add_190_195_groupi_n_915 ,csa_tree_add_190_195_groupi_n_914);
  not csa_tree_add_190_195_groupi_drc_bufs51042(csa_tree_add_190_195_groupi_n_914 ,csa_tree_add_190_195_groupi_n_2131);
  not csa_tree_add_190_195_groupi_drc_bufs51044(csa_tree_add_190_195_groupi_n_913 ,csa_tree_add_190_195_groupi_n_911);
  not csa_tree_add_190_195_groupi_drc_bufs51045(csa_tree_add_190_195_groupi_n_912 ,csa_tree_add_190_195_groupi_n_911);
  not csa_tree_add_190_195_groupi_drc_bufs51046(csa_tree_add_190_195_groupi_n_911 ,csa_tree_add_190_195_groupi_n_2127);
  not csa_tree_add_190_195_groupi_drc_bufs51052(csa_tree_add_190_195_groupi_n_910 ,csa_tree_add_190_195_groupi_n_908);
  not csa_tree_add_190_195_groupi_drc_bufs51053(csa_tree_add_190_195_groupi_n_909 ,csa_tree_add_190_195_groupi_n_908);
  not csa_tree_add_190_195_groupi_drc_bufs51054(csa_tree_add_190_195_groupi_n_908 ,csa_tree_add_190_195_groupi_n_1735);
  not csa_tree_add_190_195_groupi_drc_bufs51056(csa_tree_add_190_195_groupi_n_907 ,csa_tree_add_190_195_groupi_n_905);
  not csa_tree_add_190_195_groupi_drc_bufs51057(csa_tree_add_190_195_groupi_n_906 ,csa_tree_add_190_195_groupi_n_905);
  not csa_tree_add_190_195_groupi_drc_bufs51058(csa_tree_add_190_195_groupi_n_905 ,csa_tree_add_190_195_groupi_n_1721);
  not csa_tree_add_190_195_groupi_drc_bufs51060(csa_tree_add_190_195_groupi_n_904 ,csa_tree_add_190_195_groupi_n_902);
  not csa_tree_add_190_195_groupi_drc_bufs51061(csa_tree_add_190_195_groupi_n_903 ,csa_tree_add_190_195_groupi_n_902);
  not csa_tree_add_190_195_groupi_drc_bufs51062(csa_tree_add_190_195_groupi_n_902 ,csa_tree_add_190_195_groupi_n_1717);
  not csa_tree_add_190_195_groupi_drc_bufs51064(csa_tree_add_190_195_groupi_n_901 ,csa_tree_add_190_195_groupi_n_899);
  not csa_tree_add_190_195_groupi_drc_bufs51065(csa_tree_add_190_195_groupi_n_900 ,csa_tree_add_190_195_groupi_n_899);
  not csa_tree_add_190_195_groupi_drc_bufs51066(csa_tree_add_190_195_groupi_n_899 ,csa_tree_add_190_195_groupi_n_2022);
  not csa_tree_add_190_195_groupi_drc_bufs51068(csa_tree_add_190_195_groupi_n_898 ,csa_tree_add_190_195_groupi_n_896);
  not csa_tree_add_190_195_groupi_drc_bufs51069(csa_tree_add_190_195_groupi_n_897 ,csa_tree_add_190_195_groupi_n_896);
  not csa_tree_add_190_195_groupi_drc_bufs51070(csa_tree_add_190_195_groupi_n_896 ,csa_tree_add_190_195_groupi_n_2024);
  not csa_tree_add_190_195_groupi_drc_bufs51072(csa_tree_add_190_195_groupi_n_895 ,csa_tree_add_190_195_groupi_n_893);
  not csa_tree_add_190_195_groupi_drc_bufs51073(csa_tree_add_190_195_groupi_n_894 ,csa_tree_add_190_195_groupi_n_893);
  not csa_tree_add_190_195_groupi_drc_bufs51074(csa_tree_add_190_195_groupi_n_893 ,csa_tree_add_190_195_groupi_n_2019);
  not csa_tree_add_190_195_groupi_drc_bufs51076(csa_tree_add_190_195_groupi_n_892 ,csa_tree_add_190_195_groupi_n_890);
  not csa_tree_add_190_195_groupi_drc_bufs51077(csa_tree_add_190_195_groupi_n_891 ,csa_tree_add_190_195_groupi_n_890);
  not csa_tree_add_190_195_groupi_drc_bufs51078(csa_tree_add_190_195_groupi_n_890 ,csa_tree_add_190_195_groupi_n_1858);
  not csa_tree_add_190_195_groupi_drc_bufs51080(csa_tree_add_190_195_groupi_n_889 ,csa_tree_add_190_195_groupi_n_887);
  not csa_tree_add_190_195_groupi_drc_bufs51081(csa_tree_add_190_195_groupi_n_888 ,csa_tree_add_190_195_groupi_n_887);
  not csa_tree_add_190_195_groupi_drc_bufs51082(csa_tree_add_190_195_groupi_n_887 ,csa_tree_add_190_195_groupi_n_1984);
  not csa_tree_add_190_195_groupi_drc_bufs51084(csa_tree_add_190_195_groupi_n_886 ,csa_tree_add_190_195_groupi_n_884);
  not csa_tree_add_190_195_groupi_drc_bufs51085(csa_tree_add_190_195_groupi_n_885 ,csa_tree_add_190_195_groupi_n_884);
  not csa_tree_add_190_195_groupi_drc_bufs51086(csa_tree_add_190_195_groupi_n_884 ,csa_tree_add_190_195_groupi_n_1957);
  not csa_tree_add_190_195_groupi_drc_bufs51088(csa_tree_add_190_195_groupi_n_883 ,csa_tree_add_190_195_groupi_n_881);
  not csa_tree_add_190_195_groupi_drc_bufs51089(csa_tree_add_190_195_groupi_n_882 ,csa_tree_add_190_195_groupi_n_881);
  not csa_tree_add_190_195_groupi_drc_bufs51090(csa_tree_add_190_195_groupi_n_881 ,csa_tree_add_190_195_groupi_n_1797);
  not csa_tree_add_190_195_groupi_drc_bufs51092(csa_tree_add_190_195_groupi_n_880 ,csa_tree_add_190_195_groupi_n_878);
  not csa_tree_add_190_195_groupi_drc_bufs51093(csa_tree_add_190_195_groupi_n_879 ,csa_tree_add_190_195_groupi_n_878);
  not csa_tree_add_190_195_groupi_drc_bufs51094(csa_tree_add_190_195_groupi_n_878 ,csa_tree_add_190_195_groupi_n_2066);
  not csa_tree_add_190_195_groupi_drc_bufs51096(csa_tree_add_190_195_groupi_n_877 ,csa_tree_add_190_195_groupi_n_875);
  not csa_tree_add_190_195_groupi_drc_bufs51097(csa_tree_add_190_195_groupi_n_876 ,csa_tree_add_190_195_groupi_n_875);
  not csa_tree_add_190_195_groupi_drc_bufs51098(csa_tree_add_190_195_groupi_n_875 ,csa_tree_add_190_195_groupi_n_1792);
  not csa_tree_add_190_195_groupi_drc_bufs51100(csa_tree_add_190_195_groupi_n_874 ,csa_tree_add_190_195_groupi_n_872);
  not csa_tree_add_190_195_groupi_drc_bufs51101(csa_tree_add_190_195_groupi_n_873 ,csa_tree_add_190_195_groupi_n_872);
  not csa_tree_add_190_195_groupi_drc_bufs51102(csa_tree_add_190_195_groupi_n_872 ,csa_tree_add_190_195_groupi_n_1953);
  not csa_tree_add_190_195_groupi_drc_bufs51104(csa_tree_add_190_195_groupi_n_871 ,csa_tree_add_190_195_groupi_n_869);
  not csa_tree_add_190_195_groupi_drc_bufs51105(csa_tree_add_190_195_groupi_n_870 ,csa_tree_add_190_195_groupi_n_869);
  not csa_tree_add_190_195_groupi_drc_bufs51106(csa_tree_add_190_195_groupi_n_869 ,csa_tree_add_190_195_groupi_n_2048);
  not csa_tree_add_190_195_groupi_drc_bufs51108(csa_tree_add_190_195_groupi_n_868 ,csa_tree_add_190_195_groupi_n_866);
  not csa_tree_add_190_195_groupi_drc_bufs51109(csa_tree_add_190_195_groupi_n_867 ,csa_tree_add_190_195_groupi_n_866);
  not csa_tree_add_190_195_groupi_drc_bufs51110(csa_tree_add_190_195_groupi_n_866 ,csa_tree_add_190_195_groupi_n_1773);
  not csa_tree_add_190_195_groupi_drc_bufs51112(csa_tree_add_190_195_groupi_n_865 ,csa_tree_add_190_195_groupi_n_863);
  not csa_tree_add_190_195_groupi_drc_bufs51113(csa_tree_add_190_195_groupi_n_864 ,csa_tree_add_190_195_groupi_n_863);
  not csa_tree_add_190_195_groupi_drc_bufs51114(csa_tree_add_190_195_groupi_n_863 ,csa_tree_add_190_195_groupi_n_1769);
  not csa_tree_add_190_195_groupi_drc_bufs51116(csa_tree_add_190_195_groupi_n_862 ,csa_tree_add_190_195_groupi_n_860);
  not csa_tree_add_190_195_groupi_drc_bufs51117(csa_tree_add_190_195_groupi_n_861 ,csa_tree_add_190_195_groupi_n_860);
  not csa_tree_add_190_195_groupi_drc_bufs51118(csa_tree_add_190_195_groupi_n_860 ,csa_tree_add_190_195_groupi_n_1727);
  not csa_tree_add_190_195_groupi_drc_bufs51120(csa_tree_add_190_195_groupi_n_859 ,csa_tree_add_190_195_groupi_n_857);
  not csa_tree_add_190_195_groupi_drc_bufs51121(csa_tree_add_190_195_groupi_n_858 ,csa_tree_add_190_195_groupi_n_857);
  not csa_tree_add_190_195_groupi_drc_bufs51122(csa_tree_add_190_195_groupi_n_857 ,csa_tree_add_190_195_groupi_n_1729);
  not csa_tree_add_190_195_groupi_drc_bufs51124(csa_tree_add_190_195_groupi_n_856 ,csa_tree_add_190_195_groupi_n_854);
  not csa_tree_add_190_195_groupi_drc_bufs51125(csa_tree_add_190_195_groupi_n_855 ,csa_tree_add_190_195_groupi_n_854);
  not csa_tree_add_190_195_groupi_drc_bufs51126(csa_tree_add_190_195_groupi_n_854 ,csa_tree_add_190_195_groupi_n_1723);
  not csa_tree_add_190_195_groupi_drc_bufs51128(csa_tree_add_190_195_groupi_n_853 ,csa_tree_add_190_195_groupi_n_851);
  not csa_tree_add_190_195_groupi_drc_bufs51129(csa_tree_add_190_195_groupi_n_852 ,csa_tree_add_190_195_groupi_n_851);
  not csa_tree_add_190_195_groupi_drc_bufs51130(csa_tree_add_190_195_groupi_n_851 ,csa_tree_add_190_195_groupi_n_1939);
  not csa_tree_add_190_195_groupi_drc_bufs51132(csa_tree_add_190_195_groupi_n_850 ,csa_tree_add_190_195_groupi_n_848);
  not csa_tree_add_190_195_groupi_drc_bufs51133(csa_tree_add_190_195_groupi_n_849 ,csa_tree_add_190_195_groupi_n_848);
  not csa_tree_add_190_195_groupi_drc_bufs51134(csa_tree_add_190_195_groupi_n_848 ,csa_tree_add_190_195_groupi_n_2027);
  buf csa_tree_add_190_195_groupi_drc_bufs51136(csa_tree_add_190_195_groupi_n_1933 ,n_21);
  buf csa_tree_add_190_195_groupi_drc_bufs51137(csa_tree_add_190_195_groupi_n_1937 ,n_174);
  not csa_tree_add_190_195_groupi_drc_bufs51138(csa_tree_add_190_195_groupi_n_847 ,csa_tree_add_190_195_groupi_n_845);
  not csa_tree_add_190_195_groupi_drc_bufs51139(csa_tree_add_190_195_groupi_n_846 ,csa_tree_add_190_195_groupi_n_845);
  not csa_tree_add_190_195_groupi_drc_bufs51140(csa_tree_add_190_195_groupi_n_845 ,csa_tree_add_190_195_groupi_n_1986);
  not csa_tree_add_190_195_groupi_drc_bufs51142(csa_tree_add_190_195_groupi_n_844 ,csa_tree_add_190_195_groupi_n_842);
  not csa_tree_add_190_195_groupi_drc_bufs51143(csa_tree_add_190_195_groupi_n_843 ,csa_tree_add_190_195_groupi_n_842);
  not csa_tree_add_190_195_groupi_drc_bufs51144(csa_tree_add_190_195_groupi_n_842 ,csa_tree_add_190_195_groupi_n_1984);
  not csa_tree_add_190_195_groupi_drc_bufs51146(csa_tree_add_190_195_groupi_n_841 ,csa_tree_add_190_195_groupi_n_839);
  not csa_tree_add_190_195_groupi_drc_bufs51147(csa_tree_add_190_195_groupi_n_840 ,csa_tree_add_190_195_groupi_n_839);
  not csa_tree_add_190_195_groupi_drc_bufs51148(csa_tree_add_190_195_groupi_n_839 ,csa_tree_add_190_195_groupi_n_1982);
  not csa_tree_add_190_195_groupi_drc_bufs51150(csa_tree_add_190_195_groupi_n_838 ,csa_tree_add_190_195_groupi_n_836);
  not csa_tree_add_190_195_groupi_drc_bufs51151(csa_tree_add_190_195_groupi_n_837 ,csa_tree_add_190_195_groupi_n_836);
  not csa_tree_add_190_195_groupi_drc_bufs51152(csa_tree_add_190_195_groupi_n_836 ,csa_tree_add_190_195_groupi_n_1957);
  not csa_tree_add_190_195_groupi_drc_bufs51154(csa_tree_add_190_195_groupi_n_835 ,csa_tree_add_190_195_groupi_n_833);
  not csa_tree_add_190_195_groupi_drc_bufs51155(csa_tree_add_190_195_groupi_n_834 ,csa_tree_add_190_195_groupi_n_833);
  not csa_tree_add_190_195_groupi_drc_bufs51156(csa_tree_add_190_195_groupi_n_833 ,csa_tree_add_190_195_groupi_n_1955);
  not csa_tree_add_190_195_groupi_drc_bufs51158(csa_tree_add_190_195_groupi_n_832 ,csa_tree_add_190_195_groupi_n_830);
  not csa_tree_add_190_195_groupi_drc_bufs51159(csa_tree_add_190_195_groupi_n_831 ,csa_tree_add_190_195_groupi_n_830);
  not csa_tree_add_190_195_groupi_drc_bufs51160(csa_tree_add_190_195_groupi_n_830 ,csa_tree_add_190_195_groupi_n_2410);
  not csa_tree_add_190_195_groupi_drc_bufs51162(csa_tree_add_190_195_groupi_n_829 ,csa_tree_add_190_195_groupi_n_827);
  not csa_tree_add_190_195_groupi_drc_bufs51163(csa_tree_add_190_195_groupi_n_828 ,csa_tree_add_190_195_groupi_n_827);
  not csa_tree_add_190_195_groupi_drc_bufs51164(csa_tree_add_190_195_groupi_n_827 ,csa_tree_add_190_195_groupi_n_2411);
  not csa_tree_add_190_195_groupi_drc_bufs51166(csa_tree_add_190_195_groupi_n_826 ,csa_tree_add_190_195_groupi_n_824);
  not csa_tree_add_190_195_groupi_drc_bufs51167(csa_tree_add_190_195_groupi_n_825 ,csa_tree_add_190_195_groupi_n_824);
  not csa_tree_add_190_195_groupi_drc_bufs51168(csa_tree_add_190_195_groupi_n_824 ,csa_tree_add_190_195_groupi_n_2166);
  not csa_tree_add_190_195_groupi_drc_bufs51170(csa_tree_add_190_195_groupi_n_823 ,csa_tree_add_190_195_groupi_n_821);
  not csa_tree_add_190_195_groupi_drc_bufs51171(csa_tree_add_190_195_groupi_n_822 ,csa_tree_add_190_195_groupi_n_821);
  not csa_tree_add_190_195_groupi_drc_bufs51172(csa_tree_add_190_195_groupi_n_821 ,csa_tree_add_190_195_groupi_n_2426);
  buf csa_tree_add_190_195_groupi_drc_bufs51175(csa_tree_add_190_195_groupi_n_1936 ,n_276);
  not csa_tree_add_190_195_groupi_drc_bufs51177(csa_tree_add_190_195_groupi_n_820 ,csa_tree_add_190_195_groupi_n_818);
  not csa_tree_add_190_195_groupi_drc_bufs51178(csa_tree_add_190_195_groupi_n_819 ,csa_tree_add_190_195_groupi_n_818);
  not csa_tree_add_190_195_groupi_drc_bufs51179(csa_tree_add_190_195_groupi_n_818 ,csa_tree_add_190_195_groupi_n_2013);
  not csa_tree_add_190_195_groupi_drc_bufs51181(csa_tree_add_190_195_groupi_n_817 ,csa_tree_add_190_195_groupi_n_815);
  not csa_tree_add_190_195_groupi_drc_bufs51182(csa_tree_add_190_195_groupi_n_816 ,csa_tree_add_190_195_groupi_n_815);
  not csa_tree_add_190_195_groupi_drc_bufs51183(csa_tree_add_190_195_groupi_n_815 ,csa_tree_add_190_195_groupi_n_2011);
  buf csa_tree_add_190_195_groupi_drc_bufs51185(csa_tree_add_190_195_groupi_n_1935 ,n_89);
  buf csa_tree_add_190_195_groupi_drc_bufs51186(csa_tree_add_190_195_groupi_n_2062 ,n_411);
  buf csa_tree_add_190_195_groupi_drc_bufs51187(csa_tree_add_190_195_groupi_n_1747 ,n_84);
  buf csa_tree_add_190_195_groupi_drc_bufs51188(csa_tree_add_190_195_groupi_n_2057 ,n_383);
  buf csa_tree_add_190_195_groupi_drc_bufs51189(csa_tree_add_190_195_groupi_n_1932 ,n_225);
  buf csa_tree_add_190_195_groupi_drc_bufs51190(csa_tree_add_190_195_groupi_n_2051 ,n_349);
  buf csa_tree_add_190_195_groupi_drc_bufs51191(csa_tree_add_190_195_groupi_n_2064 ,n_156);
  buf csa_tree_add_190_195_groupi_drc_bufs51193(csa_tree_add_190_195_groupi_n_1908 ,n_87);
  buf csa_tree_add_190_195_groupi_drc_bufs51194(csa_tree_add_190_195_groupi_n_1909 ,n_291);
  buf csa_tree_add_190_195_groupi_drc_bufs51195(csa_tree_add_190_195_groupi_n_2061 ,n_258);
  buf csa_tree_add_190_195_groupi_drc_bufs51196(csa_tree_add_190_195_groupi_n_2052 ,n_247);
  buf csa_tree_add_190_195_groupi_drc_bufs51197(csa_tree_add_190_195_groupi_n_1749 ,n_91);
  buf csa_tree_add_190_195_groupi_drc_bufs51198(csa_tree_add_190_195_groupi_n_1750 ,n_414);
  buf csa_tree_add_190_195_groupi_drc_bufs51199(csa_tree_add_190_195_groupi_n_2055 ,n_297);
  buf csa_tree_add_190_195_groupi_drc_bufs51200(csa_tree_add_190_195_groupi_n_2063 ,n_292);
  buf csa_tree_add_190_195_groupi_drc_bufs51201(csa_tree_add_190_195_groupi_n_1934 ,n_412);
  buf csa_tree_add_190_195_groupi_drc_bufs51202(csa_tree_add_190_195_groupi_n_1751 ,n_108);
  buf csa_tree_add_190_195_groupi_drc_bufs51204(csa_tree_add_190_195_groupi_n_1748 ,n_322);
  buf csa_tree_add_190_195_groupi_drc_bufs51205(csa_tree_add_190_195_groupi_n_1746 ,n_67);
  buf csa_tree_add_190_195_groupi_drc_bufs51206(csa_tree_add_190_195_groupi_n_2060 ,n_207);
  buf csa_tree_add_190_195_groupi_drc_bufs51207(csa_tree_add_190_195_groupi_n_2059 ,n_196);
  buf csa_tree_add_190_195_groupi_drc_bufs51208(csa_tree_add_190_195_groupi_n_1907 ,n_415);
  buf csa_tree_add_190_195_groupi_drc_bufs51209(csa_tree_add_190_195_groupi_n_2054 ,n_416);
  buf csa_tree_add_190_195_groupi_drc_bufs51210(csa_tree_add_190_195_groupi_n_2049 ,n_212);
  buf csa_tree_add_190_195_groupi_drc_bufs51211(csa_tree_add_190_195_groupi_n_2050 ,n_348);
  buf csa_tree_add_190_195_groupi_drc_bufs51212(csa_tree_add_190_195_groupi_n_1743 ,n_85);
  buf csa_tree_add_190_195_groupi_drc_bufs51213(csa_tree_add_190_195_groupi_n_1744 ,n_136);
  buf csa_tree_add_190_195_groupi_drc_bufs51214(csa_tree_add_190_195_groupi_n_1911 ,n_155);
  buf csa_tree_add_190_195_groupi_drc_bufs51215(csa_tree_add_190_195_groupi_n_1910 ,n_138);
  buf csa_tree_add_190_195_groupi_drc_bufs51219(csa_tree_add_190_195_groupi_n_2058 ,n_195);
  buf csa_tree_add_190_195_groupi_drc_bufs51220(csa_tree_add_190_195_groupi_n_2053 ,n_263);
  buf csa_tree_add_190_195_groupi_drc_bufs51221(csa_tree_add_190_195_groupi_n_1742 ,n_68);
  buf csa_tree_add_190_195_groupi_drc_bufs51222(csa_tree_add_190_195_groupi_n_1702 ,n_222);
  buf csa_tree_add_190_195_groupi_drc_bufs51224(csa_tree_add_190_195_groupi_n_1906 ,n_317);
  buf csa_tree_add_190_195_groupi_drc_bufs51228(csa_tree_add_190_195_groupi_n_2056 ,n_144);
  buf csa_tree_add_190_195_groupi_drc_bufs51229(csa_tree_add_190_195_groupi_n_1706 ,n_307);
  buf csa_tree_add_190_195_groupi_drc_bufs51232(csa_tree_add_190_195_groupi_n_1745 ,n_204);
  buf csa_tree_add_190_195_groupi_drc_bufs51233(csa_tree_add_190_195_groupi_n_1905 ,n_249);
  buf csa_tree_add_190_195_groupi_drc_bufs51234(csa_tree_add_190_195_groupi_n_2040 ,n_404);
  buf csa_tree_add_190_195_groupi_drc_bufs51235(csa_tree_add_190_195_groupi_n_2042 ,n_200);
  buf csa_tree_add_190_195_groupi_drc_bufs51236(csa_tree_add_190_195_groupi_n_1703 ,n_35);
  buf csa_tree_add_190_195_groupi_drc_bufs51237(csa_tree_add_190_195_groupi_n_2041 ,n_353);
  buf csa_tree_add_190_195_groupi_drc_bufs51238(csa_tree_add_190_195_groupi_n_1704 ,n_69);
  buf csa_tree_add_190_195_groupi_drc_bufs51239(csa_tree_add_190_195_groupi_n_2039 ,n_217);
  buf csa_tree_add_190_195_groupi_drc_bufs51240(csa_tree_add_190_195_groupi_n_1904 ,n_334);
  buf csa_tree_add_190_195_groupi_drc_bufs51241(csa_tree_add_190_195_groupi_n_1705 ,n_103);
  buf csa_tree_add_190_195_groupi_drc_bufs51242(csa_tree_add_190_195_groupi_n_1707 ,n_171);
  buf csa_tree_add_190_195_groupi_drc_bufs51243(csa_tree_add_190_195_groupi_n_1999 ,n_327);
  buf csa_tree_add_190_195_groupi_drc_bufs51247(csa_tree_add_190_195_groupi_n_1997 ,n_140);
  buf csa_tree_add_190_195_groupi_drc_bufs51251(csa_tree_add_190_195_groupi_n_1847 ,n_57);
  buf csa_tree_add_190_195_groupi_drc_bufs51252(csa_tree_add_190_195_groupi_n_1995 ,n_259);
  buf csa_tree_add_190_195_groupi_drc_bufs51253(csa_tree_add_190_195_groupi_n_1994 ,n_208);
  buf csa_tree_add_190_195_groupi_drc_bufs51254(csa_tree_add_190_195_groupi_n_1998 ,n_191);
  buf csa_tree_add_190_195_groupi_drc_bufs51256(csa_tree_add_190_195_groupi_n_1996 ,n_293);
  buf csa_tree_add_190_195_groupi_drc_bufs51258(csa_tree_add_190_195_groupi_n_1846 ,n_227);
  buf csa_tree_add_190_195_groupi_drc_bufs51259(csa_tree_add_190_195_groupi_n_1851 ,n_193);
  buf csa_tree_add_190_195_groupi_drc_bufs51260(csa_tree_add_190_195_groupi_n_1674 ,n_286);
  buf csa_tree_add_190_195_groupi_drc_bufs51261(csa_tree_add_190_195_groupi_n_1849 ,n_278);
  buf csa_tree_add_190_195_groupi_drc_bufs51262(csa_tree_add_190_195_groupi_n_1831 ,n_306);
  buf csa_tree_add_190_195_groupi_drc_bufs51264(csa_tree_add_190_195_groupi_n_1840 ,n_288);
  buf csa_tree_add_190_195_groupi_drc_bufs51267(csa_tree_add_190_195_groupi_n_1850 ,n_125);
  buf csa_tree_add_190_195_groupi_drc_bufs51268(csa_tree_add_190_195_groupi_n_1829 ,n_51);
  buf csa_tree_add_190_195_groupi_drc_bufs51270(csa_tree_add_190_195_groupi_n_1845 ,n_431);
  buf csa_tree_add_190_195_groupi_drc_bufs51271(csa_tree_add_190_195_groupi_n_1976 ,n_296);
  buf csa_tree_add_190_195_groupi_drc_bufs51272(csa_tree_add_190_195_groupi_n_1842 ,n_169);
  buf csa_tree_add_190_195_groupi_drc_bufs51274(csa_tree_add_190_195_groupi_n_1843 ,n_390);
  buf csa_tree_add_190_195_groupi_drc_bufs51275(csa_tree_add_190_195_groupi_n_1841 ,n_118);
  buf csa_tree_add_190_195_groupi_drc_bufs51276(csa_tree_add_190_195_groupi_n_1832 ,n_323);
  buf csa_tree_add_190_195_groupi_drc_bufs51277(csa_tree_add_190_195_groupi_n_1830 ,n_289);
  buf csa_tree_add_190_195_groupi_drc_bufs51278(csa_tree_add_190_195_groupi_n_1673 ,n_82);
  buf csa_tree_add_190_195_groupi_drc_bufs51279(csa_tree_add_190_195_groupi_n_1839 ,n_356);
  buf csa_tree_add_190_195_groupi_drc_bufs51281(csa_tree_add_190_195_groupi_n_1675 ,n_133);
  buf csa_tree_add_190_195_groupi_drc_bufs51283(csa_tree_add_190_195_groupi_n_1975 ,n_262);
  buf csa_tree_add_190_195_groupi_drc_bufs51284(csa_tree_add_190_195_groupi_n_1676 ,n_320);
  buf csa_tree_add_190_195_groupi_drc_bufs51285(csa_tree_add_190_195_groupi_n_1848 ,n_74);
  buf csa_tree_add_190_195_groupi_drc_bufs51287(csa_tree_add_190_195_groupi_n_1672 ,n_65);
  buf csa_tree_add_190_195_groupi_drc_bufs51288(csa_tree_add_190_195_groupi_n_1974 ,n_245);
  buf csa_tree_add_190_195_groupi_drc_bufs51290(csa_tree_add_190_195_groupi_n_1844 ,n_203);
  buf csa_tree_add_190_195_groupi_drc_bufs51292(csa_tree_add_190_195_groupi_n_1977 ,n_194);
  buf csa_tree_add_190_195_groupi_drc_bufs51293(csa_tree_add_190_195_groupi_n_1677 ,n_184);
  buf csa_tree_add_190_195_groupi_drc_bufs51294(csa_tree_add_190_195_groupi_n_1963 ,n_147);
  buf csa_tree_add_190_195_groupi_drc_bufs51295(csa_tree_add_190_195_groupi_n_1827 ,n_221);
  buf csa_tree_add_190_195_groupi_drc_bufs51296(csa_tree_add_190_195_groupi_n_1978 ,n_410);
  buf csa_tree_add_190_195_groupi_drc_bufs51297(csa_tree_add_190_195_groupi_n_1960 ,n_215);
  buf csa_tree_add_190_195_groupi_drc_bufs51298(csa_tree_add_190_195_groupi_n_1973 ,n_211);
  buf csa_tree_add_190_195_groupi_drc_bufs51299(csa_tree_add_190_195_groupi_n_1962 ,n_419);
  buf csa_tree_add_190_195_groupi_drc_bufs51300(csa_tree_add_190_195_groupi_n_1828 ,n_408);
  buf csa_tree_add_190_195_groupi_drc_bufs51301(csa_tree_add_190_195_groupi_n_1809 ,n_375);
  buf csa_tree_add_190_195_groupi_drc_bufs51302(csa_tree_add_190_195_groupi_n_1961 ,n_402);
  buf csa_tree_add_190_195_groupi_drc_bufs51303(csa_tree_add_190_195_groupi_n_1808 ,n_273);
  buf csa_tree_add_190_195_groupi_drc_bufs51304(csa_tree_add_190_195_groupi_n_1810 ,n_137);
  buf csa_tree_add_190_195_groupi_drc_bufs51310(csa_tree_add_190_195_groupi_n_1603 ,n_100);
  buf csa_tree_add_190_195_groupi_drc_bufs51311(csa_tree_add_190_195_groupi_n_1607 ,n_321);
  buf csa_tree_add_190_195_groupi_drc_bufs51325(csa_tree_add_190_195_groupi_n_1604 ,n_287);
  buf csa_tree_add_190_195_groupi_drc_bufs51326(csa_tree_add_190_195_groupi_n_1605 ,n_117);
  buf csa_tree_add_190_195_groupi_drc_bufs51347(csa_tree_add_190_195_groupi_n_1602 ,n_49);
  buf csa_tree_add_190_195_groupi_drc_bufs51348(csa_tree_add_190_195_groupi_n_1929 ,n_210);
  buf csa_tree_add_190_195_groupi_drc_bufs51349(csa_tree_add_190_195_groupi_n_1606 ,n_134);
  not csa_tree_add_190_195_groupi_drc_bufs51433(csa_tree_add_190_195_groupi_n_2347 ,csa_tree_add_190_195_groupi_n_2008);
  buf csa_tree_add_190_195_groupi_drc_bufs51472(csa_tree_add_190_195_groupi_n_1921 ,n_220);
  buf csa_tree_add_190_195_groupi_drc_bufs51473(csa_tree_add_190_195_groupi_n_1924 ,n_152);
  not csa_tree_add_190_195_groupi_drc_bufs51512(csa_tree_add_190_195_groupi_n_2344 ,csa_tree_add_190_195_groupi_n_2157);
  buf csa_tree_add_190_195_groupi_drc_bufs51538(csa_tree_add_190_195_groupi_n_1916 ,n_255);
  not csa_tree_add_190_195_groupi_drc_bufs51543(csa_tree_add_190_195_groupi_n_814 ,csa_tree_add_190_195_groupi_n_813);
  not csa_tree_add_190_195_groupi_drc_bufs51545(csa_tree_add_190_195_groupi_n_813 ,csa_tree_add_190_195_groupi_n_1927);
  buf csa_tree_add_190_195_groupi_drc_bufs51568(csa_tree_add_190_195_groupi_n_1931 ,n_380);
  buf csa_tree_add_190_195_groupi_drc_bufs51573(csa_tree_add_190_195_groupi_n_1928 ,n_397);
  not csa_tree_add_190_195_groupi_drc_bufs51604(csa_tree_add_190_195_groupi_n_2386 ,csa_tree_add_190_195_groupi_n_2005);
  buf csa_tree_add_190_195_groupi_drc_bufs51711(csa_tree_add_190_195_groupi_n_1930 ,n_244);
  buf csa_tree_add_190_195_groupi_drc_bufs51712(csa_tree_add_190_195_groupi_n_1923 ,n_305);
  not csa_tree_add_190_195_groupi_drc_bufs51749(csa_tree_add_190_195_groupi_n_2387 ,csa_tree_add_190_195_groupi_n_1815);
  not csa_tree_add_190_195_groupi_drc_bufs51823(csa_tree_add_190_195_groupi_n_812 ,csa_tree_add_190_195_groupi_n_811);
  not csa_tree_add_190_195_groupi_drc_bufs51825(csa_tree_add_190_195_groupi_n_811 ,csa_tree_add_190_195_groupi_n_1914);
  not csa_tree_add_190_195_groupi_drc_bufs51827(csa_tree_add_190_195_groupi_n_810 ,csa_tree_add_190_195_groupi_n_809);
  not csa_tree_add_190_195_groupi_drc_bufs51829(csa_tree_add_190_195_groupi_n_809 ,csa_tree_add_190_195_groupi_n_1714);
  buf csa_tree_add_190_195_groupi_drc_bufs51844(csa_tree_add_190_195_groupi_n_1922 ,n_254);
  buf csa_tree_add_190_195_groupi_drc_bufs51846(csa_tree_add_190_195_groupi_n_1715 ,n_303);
  not csa_tree_add_190_195_groupi_drc_bufs51898(csa_tree_add_190_195_groupi_n_2372 ,csa_tree_add_190_195_groupi_n_2064);
  not csa_tree_add_190_195_groupi_drc_bufs51922(csa_tree_add_190_195_groupi_n_2373 ,csa_tree_add_190_195_groupi_n_2052);
  not csa_tree_add_190_195_groupi_drc_bufs51934(csa_tree_add_190_195_groupi_n_2382 ,csa_tree_add_190_195_groupi_n_1742);
  buf csa_tree_add_190_195_groupi_drc_bufs51948(csa_tree_add_190_195_groupi_n_1920 ,n_153);
  not csa_tree_add_190_195_groupi_drc_bufs51991(csa_tree_add_190_195_groupi_n_2354 ,csa_tree_add_190_195_groupi_n_1837);
  not csa_tree_add_190_195_groupi_drc_bufs52072(csa_tree_add_190_195_groupi_n_2379 ,csa_tree_add_190_195_groupi_n_1816);
  not csa_tree_add_190_195_groupi_drc_bufs52076(csa_tree_add_190_195_groupi_n_2349 ,csa_tree_add_190_195_groupi_n_1813);
  not csa_tree_add_190_195_groupi_drc_bufs52078(csa_tree_add_190_195_groupi_n_808 ,csa_tree_add_190_195_groupi_n_807);
  not csa_tree_add_190_195_groupi_drc_bufs52080(csa_tree_add_190_195_groupi_n_807 ,csa_tree_add_190_195_groupi_n_1801);
  not csa_tree_add_190_195_groupi_drc_bufs52082(csa_tree_add_190_195_groupi_n_806 ,csa_tree_add_190_195_groupi_n_805);
  not csa_tree_add_190_195_groupi_drc_bufs52084(csa_tree_add_190_195_groupi_n_805 ,csa_tree_add_190_195_groupi_n_1795);
  buf csa_tree_add_190_195_groupi_drc_bufs52103(csa_tree_add_190_195_groupi_n_1915 ,n_357);
  not csa_tree_add_190_195_groupi_drc_bufs52104(csa_tree_add_190_195_groupi_n_804 ,csa_tree_add_190_195_groupi_n_803);
  not csa_tree_add_190_195_groupi_drc_bufs52106(csa_tree_add_190_195_groupi_n_803 ,csa_tree_add_190_195_groupi_n_1918);
  not csa_tree_add_190_195_groupi_drc_bufs52114(csa_tree_add_190_195_groupi_n_2370 ,csa_tree_add_190_195_groupi_n_1997);
  not csa_tree_add_190_195_groupi_drc_bufs52126(csa_tree_add_190_195_groupi_n_2343 ,csa_tree_add_190_195_groupi_n_1998);
  not csa_tree_add_190_195_groupi_drc_bufs52144(csa_tree_add_190_195_groupi_n_802 ,csa_tree_add_190_195_groupi_n_801);
  not csa_tree_add_190_195_groupi_drc_bufs52146(csa_tree_add_190_195_groupi_n_801 ,csa_tree_add_190_195_groupi_n_1886);
  not csa_tree_add_190_195_groupi_drc_bufs52148(csa_tree_add_190_195_groupi_n_800 ,csa_tree_add_190_195_groupi_n_799);
  not csa_tree_add_190_195_groupi_drc_bufs52150(csa_tree_add_190_195_groupi_n_799 ,csa_tree_add_190_195_groupi_n_1883);
  not csa_tree_add_190_195_groupi_drc_bufs52160(csa_tree_add_190_195_groupi_n_798 ,csa_tree_add_190_195_groupi_n_797);
  not csa_tree_add_190_195_groupi_drc_bufs52162(csa_tree_add_190_195_groupi_n_797 ,csa_tree_add_190_195_groupi_n_1880);
  not csa_tree_add_190_195_groupi_drc_bufs52239(csa_tree_add_190_195_groupi_n_796 ,csa_tree_add_190_195_groupi_n_795);
  not csa_tree_add_190_195_groupi_drc_bufs52241(csa_tree_add_190_195_groupi_n_795 ,csa_tree_add_190_195_groupi_n_1718);
  not csa_tree_add_190_195_groupi_drc_bufs52271(csa_tree_add_190_195_groupi_n_794 ,csa_tree_add_190_195_groupi_n_793);
  not csa_tree_add_190_195_groupi_drc_bufs52273(csa_tree_add_190_195_groupi_n_793 ,csa_tree_add_190_195_groupi_n_1738);
  not csa_tree_add_190_195_groupi_drc_bufs52283(csa_tree_add_190_195_groupi_n_792 ,csa_tree_add_190_195_groupi_n_791);
  not csa_tree_add_190_195_groupi_drc_bufs52285(csa_tree_add_190_195_groupi_n_791 ,csa_tree_add_190_195_groupi_n_1741);
  buf csa_tree_add_190_195_groupi_drc_bufs52312(csa_tree_add_190_195_groupi_n_1877 ,n_239);
  not csa_tree_add_190_195_groupi_drc_bufs52337(csa_tree_add_190_195_groupi_n_790 ,csa_tree_add_190_195_groupi_n_789);
  not csa_tree_add_190_195_groupi_drc_bufs52339(csa_tree_add_190_195_groupi_n_789 ,csa_tree_add_190_195_groupi_n_1804);
  not csa_tree_add_190_195_groupi_drc_bufs52341(csa_tree_add_190_195_groupi_n_788 ,csa_tree_add_190_195_groupi_n_787);
  not csa_tree_add_190_195_groupi_drc_bufs52343(csa_tree_add_190_195_groupi_n_787 ,csa_tree_add_190_195_groupi_n_1789);
  not csa_tree_add_190_195_groupi_drc_bufs52361(csa_tree_add_190_195_groupi_n_786 ,csa_tree_add_190_195_groupi_n_785);
  not csa_tree_add_190_195_groupi_drc_bufs52363(csa_tree_add_190_195_groupi_n_785 ,csa_tree_add_190_195_groupi_n_1876);
  not csa_tree_add_190_195_groupi_drc_bufs52365(csa_tree_add_190_195_groupi_n_784 ,csa_tree_add_190_195_groupi_n_783);
  not csa_tree_add_190_195_groupi_drc_bufs52367(csa_tree_add_190_195_groupi_n_783 ,csa_tree_add_190_195_groupi_n_1713);
  not csa_tree_add_190_195_groupi_drc_bufs52420(csa_tree_add_190_195_groupi_n_2346 ,csa_tree_add_190_195_groupi_n_1933);
  not csa_tree_add_190_195_groupi_drc_bufs52448(csa_tree_add_190_195_groupi_n_2355 ,csa_tree_add_190_195_groupi_n_1672);
  not csa_tree_add_190_195_groupi_drc_bufs52460(csa_tree_add_190_195_groupi_n_2345 ,csa_tree_add_190_195_groupi_n_1907);
  not csa_tree_add_190_195_groupi_drc_bufs52464(csa_tree_add_190_195_groupi_n_2374 ,csa_tree_add_190_195_groupi_n_1908);
  not csa_tree_add_190_195_groupi_drc_bufs52476(csa_tree_add_190_195_groupi_n_2351 ,csa_tree_add_190_195_groupi_n_1743);
  not csa_tree_add_190_195_groupi_drc_bufs52490(csa_tree_add_190_195_groupi_n_782 ,csa_tree_add_190_195_groupi_n_780);
  not csa_tree_add_190_195_groupi_drc_bufs52491(csa_tree_add_190_195_groupi_n_781 ,csa_tree_add_190_195_groupi_n_780);
  not csa_tree_add_190_195_groupi_drc_bufs52492(csa_tree_add_190_195_groupi_n_780 ,csa_tree_add_190_195_groupi_n_2409);
  not csa_tree_add_190_195_groupi_drc_bufs52498(csa_tree_add_190_195_groupi_n_779 ,csa_tree_add_190_195_groupi_n_778);
  not csa_tree_add_190_195_groupi_drc_bufs52500(csa_tree_add_190_195_groupi_n_778 ,csa_tree_add_190_195_groupi_n_1685);
  not csa_tree_add_190_195_groupi_drc_bufs52502(csa_tree_add_190_195_groupi_n_777 ,csa_tree_add_190_195_groupi_n_776);
  not csa_tree_add_190_195_groupi_drc_bufs52504(csa_tree_add_190_195_groupi_n_776 ,csa_tree_add_190_195_groupi_n_1684);
  not csa_tree_add_190_195_groupi_drc_bufs52506(csa_tree_add_190_195_groupi_n_775 ,csa_tree_add_190_195_groupi_n_774);
  not csa_tree_add_190_195_groupi_drc_bufs52508(csa_tree_add_190_195_groupi_n_774 ,csa_tree_add_190_195_groupi_n_1681);
  not csa_tree_add_190_195_groupi_drc_bufs52510(csa_tree_add_190_195_groupi_n_773 ,csa_tree_add_190_195_groupi_n_772);
  not csa_tree_add_190_195_groupi_drc_bufs52512(csa_tree_add_190_195_groupi_n_772 ,csa_tree_add_190_195_groupi_n_1682);
  not csa_tree_add_190_195_groupi_drc_bufs52521(csa_tree_add_190_195_groupi_n_771 ,csa_tree_add_190_195_groupi_n_769);
  not csa_tree_add_190_195_groupi_drc_bufs52522(csa_tree_add_190_195_groupi_n_770 ,csa_tree_add_190_195_groupi_n_769);
  not csa_tree_add_190_195_groupi_drc_bufs52523(csa_tree_add_190_195_groupi_n_769 ,csa_tree_add_190_195_groupi_n_2408);
  not csa_tree_add_190_195_groupi_drc_bufs52525(csa_tree_add_190_195_groupi_n_768 ,csa_tree_add_190_195_groupi_n_766);
  not csa_tree_add_190_195_groupi_drc_bufs52526(csa_tree_add_190_195_groupi_n_767 ,csa_tree_add_190_195_groupi_n_766);
  not csa_tree_add_190_195_groupi_drc_bufs52527(csa_tree_add_190_195_groupi_n_766 ,csa_tree_add_190_195_groupi_n_2576);
  not csa_tree_add_190_195_groupi_drc_bufs52533(csa_tree_add_190_195_groupi_n_765 ,csa_tree_add_190_195_groupi_n_763);
  not csa_tree_add_190_195_groupi_drc_bufs52534(csa_tree_add_190_195_groupi_n_764 ,csa_tree_add_190_195_groupi_n_763);
  not csa_tree_add_190_195_groupi_drc_bufs52535(csa_tree_add_190_195_groupi_n_763 ,csa_tree_add_190_195_groupi_n_2411);
  not csa_tree_add_190_195_groupi_drc_bufs52537(csa_tree_add_190_195_groupi_n_762 ,csa_tree_add_190_195_groupi_n_761);
  not csa_tree_add_190_195_groupi_drc_bufs52539(csa_tree_add_190_195_groupi_n_761 ,csa_tree_add_190_195_groupi_n_1798);
  not csa_tree_add_190_195_groupi_drc_bufs52541(csa_tree_add_190_195_groupi_n_760 ,csa_tree_add_190_195_groupi_n_759);
  not csa_tree_add_190_195_groupi_drc_bufs52543(csa_tree_add_190_195_groupi_n_759 ,csa_tree_add_190_195_groupi_n_1806);
  not csa_tree_add_190_195_groupi_drc_bufs52549(csa_tree_add_190_195_groupi_n_758 ,csa_tree_add_190_195_groupi_n_757);
  not csa_tree_add_190_195_groupi_drc_bufs52551(csa_tree_add_190_195_groupi_n_757 ,csa_tree_add_190_195_groupi_n_1782);
  not csa_tree_add_190_195_groupi_drc_bufs52565(csa_tree_add_190_195_groupi_n_756 ,csa_tree_add_190_195_groupi_n_755);
  not csa_tree_add_190_195_groupi_drc_bufs52567(csa_tree_add_190_195_groupi_n_755 ,csa_tree_add_190_195_groupi_n_1785);
  not csa_tree_add_190_195_groupi_drc_bufs52583(csa_tree_add_190_195_groupi_n_2377 ,csa_tree_add_190_195_groupi_n_1916);
  not csa_tree_add_190_195_groupi_drc_bufs52589(csa_tree_add_190_195_groupi_n_754 ,csa_tree_add_190_195_groupi_n_1565);
  not csa_tree_add_190_195_groupi_drc_bufs52606(csa_tree_add_190_195_groupi_n_753 ,csa_tree_add_190_195_groupi_n_752);
  not csa_tree_add_190_195_groupi_drc_bufs52608(csa_tree_add_190_195_groupi_n_752 ,csa_tree_add_190_195_groupi_n_1724);
  not csa_tree_add_190_195_groupi_drc_bufs52610(csa_tree_add_190_195_groupi_n_751 ,csa_tree_add_190_195_groupi_n_750);
  not csa_tree_add_190_195_groupi_drc_bufs52612(csa_tree_add_190_195_groupi_n_750 ,csa_tree_add_190_195_groupi_n_1730);
  not csa_tree_add_190_195_groupi_drc_bufs52618(csa_tree_add_190_195_groupi_n_749 ,csa_tree_add_190_195_groupi_n_2342);
  not csa_tree_add_190_195_groupi_drc_bufs52620(csa_tree_add_190_195_groupi_n_2342 ,csa_tree_add_190_195_groupi_n_1720);
  not csa_tree_add_190_195_groupi_drc_bufs52622(csa_tree_add_190_195_groupi_n_748 ,csa_tree_add_190_195_groupi_n_747);
  not csa_tree_add_190_195_groupi_drc_bufs52624(csa_tree_add_190_195_groupi_n_747 ,csa_tree_add_190_195_groupi_n_1734);
  not csa_tree_add_190_195_groupi_drc_bufs52626(csa_tree_add_190_195_groupi_n_746 ,csa_tree_add_190_195_groupi_n_2371);
  not csa_tree_add_190_195_groupi_drc_bufs52628(csa_tree_add_190_195_groupi_n_2371 ,csa_tree_add_190_195_groupi_n_1732);
  not csa_tree_add_190_195_groupi_drc_bufs52634(csa_tree_add_190_195_groupi_n_745 ,csa_tree_add_190_195_groupi_n_743);
  not csa_tree_add_190_195_groupi_drc_bufs52635(csa_tree_add_190_195_groupi_n_744 ,csa_tree_add_190_195_groupi_n_743);
  not csa_tree_add_190_195_groupi_drc_bufs52636(csa_tree_add_190_195_groupi_n_743 ,csa_tree_add_190_195_groupi_n_2415);
  not csa_tree_add_190_195_groupi_drc_bufs52638(csa_tree_add_190_195_groupi_n_742 ,csa_tree_add_190_195_groupi_n_741);
  not csa_tree_add_190_195_groupi_drc_bufs52640(csa_tree_add_190_195_groupi_n_741 ,csa_tree_add_190_195_groupi_n_1791);
  not csa_tree_add_190_195_groupi_drc_bufs52650(csa_tree_add_190_195_groupi_n_740 ,csa_tree_add_190_195_groupi_n_738);
  not csa_tree_add_190_195_groupi_drc_bufs52651(csa_tree_add_190_195_groupi_n_739 ,csa_tree_add_190_195_groupi_n_738);
  not csa_tree_add_190_195_groupi_drc_bufs52652(csa_tree_add_190_195_groupi_n_738 ,csa_tree_add_190_195_groupi_n_2407);
  not csa_tree_add_190_195_groupi_drc_bufs52654(csa_tree_add_190_195_groupi_n_737 ,csa_tree_add_190_195_groupi_n_735);
  not csa_tree_add_190_195_groupi_drc_bufs52655(csa_tree_add_190_195_groupi_n_736 ,csa_tree_add_190_195_groupi_n_735);
  not csa_tree_add_190_195_groupi_drc_bufs52656(csa_tree_add_190_195_groupi_n_735 ,csa_tree_add_190_195_groupi_n_2584);
  not csa_tree_add_190_195_groupi_drc_bufs52658(csa_tree_add_190_195_groupi_n_734 ,csa_tree_add_190_195_groupi_n_732);
  not csa_tree_add_190_195_groupi_drc_bufs52659(csa_tree_add_190_195_groupi_n_733 ,csa_tree_add_190_195_groupi_n_732);
  not csa_tree_add_190_195_groupi_drc_bufs52660(csa_tree_add_190_195_groupi_n_732 ,csa_tree_add_190_195_groupi_n_2417);
  not csa_tree_add_190_195_groupi_drc_bufs52663(csa_tree_add_190_195_groupi_n_731 ,csa_tree_add_190_195_groupi_n_730);
  not csa_tree_add_190_195_groupi_drc_bufs52664(csa_tree_add_190_195_groupi_n_730 ,csa_tree_add_190_195_groupi_n_1545);
  not csa_tree_add_190_195_groupi_drc_bufs52667(csa_tree_add_190_195_groupi_n_729 ,csa_tree_add_190_195_groupi_n_728);
  not csa_tree_add_190_195_groupi_drc_bufs52668(csa_tree_add_190_195_groupi_n_728 ,csa_tree_add_190_195_groupi_n_1549);
  not csa_tree_add_190_195_groupi_drc_bufs52670(csa_tree_add_190_195_groupi_n_727 ,csa_tree_add_190_195_groupi_n_725);
  not csa_tree_add_190_195_groupi_drc_bufs52671(csa_tree_add_190_195_groupi_n_726 ,csa_tree_add_190_195_groupi_n_725);
  not csa_tree_add_190_195_groupi_drc_bufs52672(csa_tree_add_190_195_groupi_n_725 ,csa_tree_add_190_195_groupi_n_2415);
  not csa_tree_add_190_195_groupi_drc_bufs52674(csa_tree_add_190_195_groupi_n_724 ,csa_tree_add_190_195_groupi_n_722);
  not csa_tree_add_190_195_groupi_drc_bufs52675(csa_tree_add_190_195_groupi_n_723 ,csa_tree_add_190_195_groupi_n_722);
  not csa_tree_add_190_195_groupi_drc_bufs52676(csa_tree_add_190_195_groupi_n_722 ,csa_tree_add_190_195_groupi_n_2408);
  not csa_tree_add_190_195_groupi_drc_bufs52678(csa_tree_add_190_195_groupi_n_721 ,csa_tree_add_190_195_groupi_n_719);
  not csa_tree_add_190_195_groupi_drc_bufs52679(csa_tree_add_190_195_groupi_n_720 ,csa_tree_add_190_195_groupi_n_719);
  not csa_tree_add_190_195_groupi_drc_bufs52680(csa_tree_add_190_195_groupi_n_719 ,csa_tree_add_190_195_groupi_n_2588);
  not csa_tree_add_190_195_groupi_drc_bufs52683(csa_tree_add_190_195_groupi_n_718 ,csa_tree_add_190_195_groupi_n_717);
  not csa_tree_add_190_195_groupi_drc_bufs52684(csa_tree_add_190_195_groupi_n_717 ,csa_tree_add_190_195_groupi_n_2426);
  not csa_tree_add_190_195_groupi_drc_bufs52686(csa_tree_add_190_195_groupi_n_716 ,csa_tree_add_190_195_groupi_n_714);
  not csa_tree_add_190_195_groupi_drc_bufs52687(csa_tree_add_190_195_groupi_n_715 ,csa_tree_add_190_195_groupi_n_714);
  not csa_tree_add_190_195_groupi_drc_bufs52688(csa_tree_add_190_195_groupi_n_714 ,csa_tree_add_190_195_groupi_n_2453);
  not csa_tree_add_190_195_groupi_drc_bufs52690(csa_tree_add_190_195_groupi_n_713 ,csa_tree_add_190_195_groupi_n_711);
  not csa_tree_add_190_195_groupi_drc_bufs52691(csa_tree_add_190_195_groupi_n_712 ,csa_tree_add_190_195_groupi_n_711);
  not csa_tree_add_190_195_groupi_drc_bufs52692(csa_tree_add_190_195_groupi_n_711 ,csa_tree_add_190_195_groupi_n_2708);
  not csa_tree_add_190_195_groupi_drc_bufs52695(csa_tree_add_190_195_groupi_n_710 ,csa_tree_add_190_195_groupi_n_709);
  not csa_tree_add_190_195_groupi_drc_bufs52696(csa_tree_add_190_195_groupi_n_709 ,csa_tree_add_190_195_groupi_n_1726);
  not csa_tree_add_190_195_groupi_drc_bufs52698(csa_tree_add_190_195_groupi_n_708 ,csa_tree_add_190_195_groupi_n_706);
  not csa_tree_add_190_195_groupi_drc_bufs52699(csa_tree_add_190_195_groupi_n_707 ,csa_tree_add_190_195_groupi_n_706);
  not csa_tree_add_190_195_groupi_drc_bufs52700(csa_tree_add_190_195_groupi_n_706 ,csa_tree_add_190_195_groupi_n_2424);
  not csa_tree_add_190_195_groupi_drc_bufs52702(csa_tree_add_190_195_groupi_n_705 ,csa_tree_add_190_195_groupi_n_703);
  not csa_tree_add_190_195_groupi_drc_bufs52703(csa_tree_add_190_195_groupi_n_704 ,csa_tree_add_190_195_groupi_n_703);
  not csa_tree_add_190_195_groupi_drc_bufs52704(csa_tree_add_190_195_groupi_n_703 ,csa_tree_add_190_195_groupi_n_2583);
  not csa_tree_add_190_195_groupi_drc_bufs52707(csa_tree_add_190_195_groupi_n_702 ,csa_tree_add_190_195_groupi_n_701);
  not csa_tree_add_190_195_groupi_drc_bufs52708(csa_tree_add_190_195_groupi_n_701 ,csa_tree_add_190_195_groupi_n_1556);
  not csa_tree_add_190_195_groupi_drc_bufs52711(csa_tree_add_190_195_groupi_n_700 ,csa_tree_add_190_195_groupi_n_699);
  not csa_tree_add_190_195_groupi_drc_bufs52712(csa_tree_add_190_195_groupi_n_699 ,csa_tree_add_190_195_groupi_n_1559);
  not csa_tree_add_190_195_groupi_drc_bufs52714(csa_tree_add_190_195_groupi_n_698 ,csa_tree_add_190_195_groupi_n_696);
  not csa_tree_add_190_195_groupi_drc_bufs52715(csa_tree_add_190_195_groupi_n_697 ,csa_tree_add_190_195_groupi_n_696);
  not csa_tree_add_190_195_groupi_drc_bufs52716(csa_tree_add_190_195_groupi_n_696 ,csa_tree_add_190_195_groupi_n_2416);
  not csa_tree_add_190_195_groupi_drc_bufs52718(csa_tree_add_190_195_groupi_n_695 ,csa_tree_add_190_195_groupi_n_693);
  not csa_tree_add_190_195_groupi_drc_bufs52719(csa_tree_add_190_195_groupi_n_694 ,csa_tree_add_190_195_groupi_n_693);
  not csa_tree_add_190_195_groupi_drc_bufs52720(csa_tree_add_190_195_groupi_n_693 ,csa_tree_add_190_195_groupi_n_2581);
  not csa_tree_add_190_195_groupi_drc_bufs52722(csa_tree_add_190_195_groupi_n_692 ,csa_tree_add_190_195_groupi_n_690);
  not csa_tree_add_190_195_groupi_drc_bufs52723(csa_tree_add_190_195_groupi_n_691 ,csa_tree_add_190_195_groupi_n_690);
  not csa_tree_add_190_195_groupi_drc_bufs52724(csa_tree_add_190_195_groupi_n_690 ,csa_tree_add_190_195_groupi_n_2579);
  not csa_tree_add_190_195_groupi_drc_bufs52726(csa_tree_add_190_195_groupi_n_689 ,csa_tree_add_190_195_groupi_n_687);
  not csa_tree_add_190_195_groupi_drc_bufs52727(csa_tree_add_190_195_groupi_n_688 ,csa_tree_add_190_195_groupi_n_687);
  not csa_tree_add_190_195_groupi_drc_bufs52728(csa_tree_add_190_195_groupi_n_687 ,csa_tree_add_190_195_groupi_n_2576);
  not csa_tree_add_190_195_groupi_drc_bufs52730(csa_tree_add_190_195_groupi_n_686 ,csa_tree_add_190_195_groupi_n_684);
  not csa_tree_add_190_195_groupi_drc_bufs52731(csa_tree_add_190_195_groupi_n_685 ,csa_tree_add_190_195_groupi_n_684);
  not csa_tree_add_190_195_groupi_drc_bufs52732(csa_tree_add_190_195_groupi_n_684 ,csa_tree_add_190_195_groupi_n_2586);
  not csa_tree_add_190_195_groupi_drc_bufs52735(csa_tree_add_190_195_groupi_n_683 ,csa_tree_add_190_195_groupi_n_682);
  not csa_tree_add_190_195_groupi_drc_bufs52736(csa_tree_add_190_195_groupi_n_682 ,csa_tree_add_190_195_groupi_n_2432);
  not csa_tree_add_190_195_groupi_drc_bufs52739(csa_tree_add_190_195_groupi_n_681 ,csa_tree_add_190_195_groupi_n_680);
  not csa_tree_add_190_195_groupi_drc_bufs52740(csa_tree_add_190_195_groupi_n_680 ,csa_tree_add_190_195_groupi_n_2594);
  not csa_tree_add_190_195_groupi_drc_bufs52742(csa_tree_add_190_195_groupi_n_679 ,csa_tree_add_190_195_groupi_n_677);
  not csa_tree_add_190_195_groupi_drc_bufs52743(csa_tree_add_190_195_groupi_n_678 ,csa_tree_add_190_195_groupi_n_677);
  not csa_tree_add_190_195_groupi_drc_bufs52744(csa_tree_add_190_195_groupi_n_677 ,csa_tree_add_190_195_groupi_n_2594);
  not csa_tree_add_190_195_groupi_drc_bufs52747(csa_tree_add_190_195_groupi_n_676 ,csa_tree_add_190_195_groupi_n_674);
  not csa_tree_add_190_195_groupi_drc_bufs52748(csa_tree_add_190_195_groupi_n_675 ,csa_tree_add_190_195_groupi_n_674);
  not csa_tree_add_190_195_groupi_drc_bufs52749(csa_tree_add_190_195_groupi_n_674 ,csa_tree_add_190_195_groupi_n_2407);
  not csa_tree_add_190_195_groupi_drc_bufs52751(csa_tree_add_190_195_groupi_n_673 ,csa_tree_add_190_195_groupi_n_671);
  not csa_tree_add_190_195_groupi_drc_bufs52752(csa_tree_add_190_195_groupi_n_672 ,csa_tree_add_190_195_groupi_n_671);
  not csa_tree_add_190_195_groupi_drc_bufs52753(csa_tree_add_190_195_groupi_n_671 ,csa_tree_add_190_195_groupi_n_2432);
  not csa_tree_add_190_195_groupi_drc_bufs52755(csa_tree_add_190_195_groupi_n_670 ,csa_tree_add_190_195_groupi_n_668);
  not csa_tree_add_190_195_groupi_drc_bufs52756(csa_tree_add_190_195_groupi_n_669 ,csa_tree_add_190_195_groupi_n_668);
  not csa_tree_add_190_195_groupi_drc_bufs52757(csa_tree_add_190_195_groupi_n_668 ,csa_tree_add_190_195_groupi_n_2598);
  not csa_tree_add_190_195_groupi_drc_bufs52759(csa_tree_add_190_195_groupi_n_667 ,csa_tree_add_190_195_groupi_n_665);
  not csa_tree_add_190_195_groupi_drc_bufs52760(csa_tree_add_190_195_groupi_n_666 ,csa_tree_add_190_195_groupi_n_665);
  not csa_tree_add_190_195_groupi_drc_bufs52761(csa_tree_add_190_195_groupi_n_665 ,csa_tree_add_190_195_groupi_n_2646);
  not csa_tree_add_190_195_groupi_drc_bufs52763(csa_tree_add_190_195_groupi_n_664 ,csa_tree_add_190_195_groupi_n_662);
  not csa_tree_add_190_195_groupi_drc_bufs52764(csa_tree_add_190_195_groupi_n_663 ,csa_tree_add_190_195_groupi_n_662);
  not csa_tree_add_190_195_groupi_drc_bufs52765(csa_tree_add_190_195_groupi_n_662 ,csa_tree_add_190_195_groupi_n_2644);
  not csa_tree_add_190_195_groupi_drc_bufs52767(csa_tree_add_190_195_groupi_n_661 ,csa_tree_add_190_195_groupi_n_659);
  not csa_tree_add_190_195_groupi_drc_bufs52768(csa_tree_add_190_195_groupi_n_660 ,csa_tree_add_190_195_groupi_n_659);
  not csa_tree_add_190_195_groupi_drc_bufs52769(csa_tree_add_190_195_groupi_n_659 ,csa_tree_add_190_195_groupi_n_2639);
  not csa_tree_add_190_195_groupi_drc_bufs52786(csa_tree_add_190_195_groupi_n_658 ,csa_tree_add_190_195_groupi_n_657);
  not csa_tree_add_190_195_groupi_drc_bufs52788(csa_tree_add_190_195_groupi_n_657 ,csa_tree_add_190_195_groupi_n_1669);
  not csa_tree_add_190_195_groupi_drc_bufs52790(csa_tree_add_190_195_groupi_n_656 ,csa_tree_add_190_195_groupi_n_655);
  not csa_tree_add_190_195_groupi_drc_bufs52792(csa_tree_add_190_195_groupi_n_655 ,csa_tree_add_190_195_groupi_n_1660);
  not csa_tree_add_190_195_groupi_drc_bufs52794(csa_tree_add_190_195_groupi_n_654 ,csa_tree_add_190_195_groupi_n_653);
  not csa_tree_add_190_195_groupi_drc_bufs52796(csa_tree_add_190_195_groupi_n_653 ,csa_tree_add_190_195_groupi_n_1663);
  not csa_tree_add_190_195_groupi_drc_bufs52798(csa_tree_add_190_195_groupi_n_652 ,csa_tree_add_190_195_groupi_n_651);
  not csa_tree_add_190_195_groupi_drc_bufs52800(csa_tree_add_190_195_groupi_n_651 ,csa_tree_add_190_195_groupi_n_1654);
  not csa_tree_add_190_195_groupi_drc_bufs52802(csa_tree_add_190_195_groupi_n_650 ,csa_tree_add_190_195_groupi_n_649);
  not csa_tree_add_190_195_groupi_drc_bufs52804(csa_tree_add_190_195_groupi_n_649 ,csa_tree_add_190_195_groupi_n_1648);
  not csa_tree_add_190_195_groupi_drc_bufs52806(csa_tree_add_190_195_groupi_n_648 ,csa_tree_add_190_195_groupi_n_647);
  not csa_tree_add_190_195_groupi_drc_bufs52808(csa_tree_add_190_195_groupi_n_647 ,csa_tree_add_190_195_groupi_n_1645);
  not csa_tree_add_190_195_groupi_drc_bufs52810(csa_tree_add_190_195_groupi_n_646 ,csa_tree_add_190_195_groupi_n_645);
  not csa_tree_add_190_195_groupi_drc_bufs52812(csa_tree_add_190_195_groupi_n_645 ,csa_tree_add_190_195_groupi_n_1651);
  not csa_tree_add_190_195_groupi_drc_bufs52814(csa_tree_add_190_195_groupi_n_644 ,csa_tree_add_190_195_groupi_n_643);
  not csa_tree_add_190_195_groupi_drc_bufs52816(csa_tree_add_190_195_groupi_n_643 ,csa_tree_add_190_195_groupi_n_1666);
  not csa_tree_add_190_195_groupi_drc_bufs52818(csa_tree_add_190_195_groupi_n_642 ,csa_tree_add_190_195_groupi_n_641);
  not csa_tree_add_190_195_groupi_drc_bufs52820(csa_tree_add_190_195_groupi_n_641 ,csa_tree_add_190_195_groupi_n_1657);
  not csa_tree_add_190_195_groupi_drc_bufs52822(csa_tree_add_190_195_groupi_n_640 ,csa_tree_add_190_195_groupi_n_639);
  not csa_tree_add_190_195_groupi_drc_bufs52824(csa_tree_add_190_195_groupi_n_639 ,csa_tree_add_190_195_groupi_n_1642);
  not csa_tree_add_190_195_groupi_drc_bufs52826(csa_tree_add_190_195_groupi_n_638 ,csa_tree_add_190_195_groupi_n_637);
  not csa_tree_add_190_195_groupi_drc_bufs52828(csa_tree_add_190_195_groupi_n_637 ,csa_tree_add_190_195_groupi_n_1639);
  not csa_tree_add_190_195_groupi_drc_bufs52830(csa_tree_add_190_195_groupi_n_636 ,csa_tree_add_190_195_groupi_n_635);
  not csa_tree_add_190_195_groupi_drc_bufs52832(csa_tree_add_190_195_groupi_n_635 ,csa_tree_add_190_195_groupi_n_1631);
  not csa_tree_add_190_195_groupi_drc_bufs52834(csa_tree_add_190_195_groupi_n_634 ,csa_tree_add_190_195_groupi_n_633);
  not csa_tree_add_190_195_groupi_drc_bufs52836(csa_tree_add_190_195_groupi_n_633 ,csa_tree_add_190_195_groupi_n_1625);
  not csa_tree_add_190_195_groupi_drc_bufs52838(csa_tree_add_190_195_groupi_n_632 ,csa_tree_add_190_195_groupi_n_631);
  not csa_tree_add_190_195_groupi_drc_bufs52840(csa_tree_add_190_195_groupi_n_631 ,csa_tree_add_190_195_groupi_n_1628);
  not csa_tree_add_190_195_groupi_drc_bufs52843(csa_tree_add_190_195_groupi_n_2388 ,csa_tree_add_190_195_groupi_n_629);
  not csa_tree_add_190_195_groupi_drc_bufs52844(csa_tree_add_190_195_groupi_n_630 ,csa_tree_add_190_195_groupi_n_629);
  not csa_tree_add_190_195_groupi_drc_bufs52845(csa_tree_add_190_195_groupi_n_629 ,csa_tree_add_190_195_groupi_n_1634);
  not csa_tree_add_190_195_groupi_drc_bufs53025(csa_tree_add_190_195_groupi_n_628 ,csa_tree_add_190_195_groupi_n_626);
  not csa_tree_add_190_195_groupi_drc_bufs53026(csa_tree_add_190_195_groupi_n_627 ,csa_tree_add_190_195_groupi_n_626);
  not csa_tree_add_190_195_groupi_drc_bufs53027(csa_tree_add_190_195_groupi_n_626 ,csa_tree_add_190_195_groupi_n_2318);
  not csa_tree_add_190_195_groupi_drc_bufs53046(csa_tree_add_190_195_groupi_n_625 ,csa_tree_add_190_195_groupi_n_623);
  not csa_tree_add_190_195_groupi_drc_bufs53047(csa_tree_add_190_195_groupi_n_624 ,csa_tree_add_190_195_groupi_n_623);
  not csa_tree_add_190_195_groupi_drc_bufs53048(csa_tree_add_190_195_groupi_n_623 ,csa_tree_add_190_195_groupi_n_2314);
  not csa_tree_add_190_195_groupi_drc_bufs53050(csa_tree_add_190_195_groupi_n_622 ,csa_tree_add_190_195_groupi_n_620);
  not csa_tree_add_190_195_groupi_drc_bufs53051(csa_tree_add_190_195_groupi_n_621 ,csa_tree_add_190_195_groupi_n_620);
  not csa_tree_add_190_195_groupi_drc_bufs53052(csa_tree_add_190_195_groupi_n_620 ,csa_tree_add_190_195_groupi_n_2327);
  not csa_tree_add_190_195_groupi_drc_bufs53054(csa_tree_add_190_195_groupi_n_619 ,csa_tree_add_190_195_groupi_n_617);
  not csa_tree_add_190_195_groupi_drc_bufs53055(csa_tree_add_190_195_groupi_n_618 ,csa_tree_add_190_195_groupi_n_617);
  not csa_tree_add_190_195_groupi_drc_bufs53056(csa_tree_add_190_195_groupi_n_617 ,csa_tree_add_190_195_groupi_n_2324);
  not csa_tree_add_190_195_groupi_drc_bufs53058(csa_tree_add_190_195_groupi_n_616 ,csa_tree_add_190_195_groupi_n_614);
  not csa_tree_add_190_195_groupi_drc_bufs53059(csa_tree_add_190_195_groupi_n_615 ,csa_tree_add_190_195_groupi_n_614);
  not csa_tree_add_190_195_groupi_drc_bufs53060(csa_tree_add_190_195_groupi_n_614 ,csa_tree_add_190_195_groupi_n_2305);
  not csa_tree_add_190_195_groupi_drc_bufs53062(csa_tree_add_190_195_groupi_n_613 ,csa_tree_add_190_195_groupi_n_611);
  not csa_tree_add_190_195_groupi_drc_bufs53063(csa_tree_add_190_195_groupi_n_612 ,csa_tree_add_190_195_groupi_n_611);
  not csa_tree_add_190_195_groupi_drc_bufs53064(csa_tree_add_190_195_groupi_n_611 ,csa_tree_add_190_195_groupi_n_2321);
  not csa_tree_add_190_195_groupi_drc_bufs53066(csa_tree_add_190_195_groupi_n_610 ,csa_tree_add_190_195_groupi_n_608);
  not csa_tree_add_190_195_groupi_drc_bufs53067(csa_tree_add_190_195_groupi_n_609 ,csa_tree_add_190_195_groupi_n_608);
  not csa_tree_add_190_195_groupi_drc_bufs53068(csa_tree_add_190_195_groupi_n_608 ,csa_tree_add_190_195_groupi_n_2326);
  not csa_tree_add_190_195_groupi_drc_bufs53070(csa_tree_add_190_195_groupi_n_607 ,csa_tree_add_190_195_groupi_n_605);
  not csa_tree_add_190_195_groupi_drc_bufs53071(csa_tree_add_190_195_groupi_n_606 ,csa_tree_add_190_195_groupi_n_605);
  not csa_tree_add_190_195_groupi_drc_bufs53072(csa_tree_add_190_195_groupi_n_605 ,csa_tree_add_190_195_groupi_n_2323);
  not csa_tree_add_190_195_groupi_drc_bufs53074(csa_tree_add_190_195_groupi_n_604 ,csa_tree_add_190_195_groupi_n_602);
  not csa_tree_add_190_195_groupi_drc_bufs53075(csa_tree_add_190_195_groupi_n_603 ,csa_tree_add_190_195_groupi_n_602);
  not csa_tree_add_190_195_groupi_drc_bufs53076(csa_tree_add_190_195_groupi_n_602 ,csa_tree_add_190_195_groupi_n_2320);
  not csa_tree_add_190_195_groupi_drc_bufs53078(csa_tree_add_190_195_groupi_n_601 ,csa_tree_add_190_195_groupi_n_599);
  not csa_tree_add_190_195_groupi_drc_bufs53079(csa_tree_add_190_195_groupi_n_600 ,csa_tree_add_190_195_groupi_n_599);
  not csa_tree_add_190_195_groupi_drc_bufs53080(csa_tree_add_190_195_groupi_n_599 ,csa_tree_add_190_195_groupi_n_2308);
  not csa_tree_add_190_195_groupi_drc_bufs53082(csa_tree_add_190_195_groupi_n_598 ,csa_tree_add_190_195_groupi_n_596);
  not csa_tree_add_190_195_groupi_drc_bufs53083(csa_tree_add_190_195_groupi_n_597 ,csa_tree_add_190_195_groupi_n_596);
  not csa_tree_add_190_195_groupi_drc_bufs53084(csa_tree_add_190_195_groupi_n_596 ,csa_tree_add_190_195_groupi_n_2302);
  not csa_tree_add_190_195_groupi_drc_bufs53097(csa_tree_add_190_195_groupi_n_595 ,csa_tree_add_190_195_groupi_n_593);
  not csa_tree_add_190_195_groupi_drc_bufs53098(csa_tree_add_190_195_groupi_n_594 ,csa_tree_add_190_195_groupi_n_593);
  not csa_tree_add_190_195_groupi_drc_bufs53099(csa_tree_add_190_195_groupi_n_593 ,csa_tree_add_190_195_groupi_n_2300);
  not csa_tree_add_190_195_groupi_drc_bufs53184(csa_tree_add_190_195_groupi_n_592 ,csa_tree_add_190_195_groupi_n_590);
  not csa_tree_add_190_195_groupi_drc_bufs53185(csa_tree_add_190_195_groupi_n_591 ,csa_tree_add_190_195_groupi_n_590);
  not csa_tree_add_190_195_groupi_drc_bufs53186(csa_tree_add_190_195_groupi_n_590 ,csa_tree_add_190_195_groupi_n_2228);
  not csa_tree_add_190_195_groupi_drc_bufs53188(csa_tree_add_190_195_groupi_n_589 ,csa_tree_add_190_195_groupi_n_587);
  not csa_tree_add_190_195_groupi_drc_bufs53189(csa_tree_add_190_195_groupi_n_588 ,csa_tree_add_190_195_groupi_n_587);
  not csa_tree_add_190_195_groupi_drc_bufs53190(csa_tree_add_190_195_groupi_n_587 ,csa_tree_add_190_195_groupi_n_2103);
  not csa_tree_add_190_195_groupi_drc_bufs53192(csa_tree_add_190_195_groupi_n_586 ,csa_tree_add_190_195_groupi_n_584);
  not csa_tree_add_190_195_groupi_drc_bufs53193(csa_tree_add_190_195_groupi_n_585 ,csa_tree_add_190_195_groupi_n_584);
  not csa_tree_add_190_195_groupi_drc_bufs53194(csa_tree_add_190_195_groupi_n_584 ,csa_tree_add_190_195_groupi_n_2318);
  not csa_tree_add_190_195_groupi_drc_bufs53196(csa_tree_add_190_195_groupi_n_583 ,csa_tree_add_190_195_groupi_n_2363);
  not csa_tree_add_190_195_groupi_drc_bufs53198(csa_tree_add_190_195_groupi_n_2363 ,csa_tree_add_190_195_groupi_n_2291);
  not csa_tree_add_190_195_groupi_drc_bufs53200(csa_tree_add_190_195_groupi_n_582 ,csa_tree_add_190_195_groupi_n_580);
  not csa_tree_add_190_195_groupi_drc_bufs53201(csa_tree_add_190_195_groupi_n_581 ,csa_tree_add_190_195_groupi_n_580);
  not csa_tree_add_190_195_groupi_drc_bufs53202(csa_tree_add_190_195_groupi_n_580 ,csa_tree_add_190_195_groupi_n_2314);
  not csa_tree_add_190_195_groupi_drc_bufs53204(csa_tree_add_190_195_groupi_n_579 ,csa_tree_add_190_195_groupi_n_578);
  not csa_tree_add_190_195_groupi_drc_bufs53206(csa_tree_add_190_195_groupi_n_578 ,csa_tree_add_190_195_groupi_n_2231);
  not csa_tree_add_190_195_groupi_drc_bufs53208(csa_tree_add_190_195_groupi_n_577 ,csa_tree_add_190_195_groupi_n_575);
  not csa_tree_add_190_195_groupi_drc_bufs53209(csa_tree_add_190_195_groupi_n_576 ,csa_tree_add_190_195_groupi_n_575);
  not csa_tree_add_190_195_groupi_drc_bufs53210(csa_tree_add_190_195_groupi_n_575 ,csa_tree_add_190_195_groupi_n_2231);
  not csa_tree_add_190_195_groupi_drc_bufs53212(csa_tree_add_190_195_groupi_n_574 ,csa_tree_add_190_195_groupi_n_573);
  not csa_tree_add_190_195_groupi_drc_bufs53214(csa_tree_add_190_195_groupi_n_573 ,csa_tree_add_190_195_groupi_n_2311);
  not csa_tree_add_190_195_groupi_drc_bufs53216(csa_tree_add_190_195_groupi_n_572 ,csa_tree_add_190_195_groupi_n_571);
  not csa_tree_add_190_195_groupi_drc_bufs53218(csa_tree_add_190_195_groupi_n_571 ,csa_tree_add_190_195_groupi_n_2315);
  not csa_tree_add_190_195_groupi_drc_bufs53220(csa_tree_add_190_195_groupi_n_570 ,csa_tree_add_190_195_groupi_n_569);
  not csa_tree_add_190_195_groupi_drc_bufs53222(csa_tree_add_190_195_groupi_n_569 ,csa_tree_add_190_195_groupi_n_2317);
  not csa_tree_add_190_195_groupi_drc_bufs53224(csa_tree_add_190_195_groupi_n_568 ,csa_tree_add_190_195_groupi_n_567);
  not csa_tree_add_190_195_groupi_drc_bufs53226(csa_tree_add_190_195_groupi_n_567 ,csa_tree_add_190_195_groupi_n_2317);
  not csa_tree_add_190_195_groupi_drc_bufs53228(csa_tree_add_190_195_groupi_n_566 ,csa_tree_add_190_195_groupi_n_565);
  not csa_tree_add_190_195_groupi_drc_bufs53230(csa_tree_add_190_195_groupi_n_565 ,csa_tree_add_190_195_groupi_n_2312);
  not csa_tree_add_190_195_groupi_drc_bufs53232(csa_tree_add_190_195_groupi_n_564 ,csa_tree_add_190_195_groupi_n_562);
  not csa_tree_add_190_195_groupi_drc_bufs53233(csa_tree_add_190_195_groupi_n_563 ,csa_tree_add_190_195_groupi_n_562);
  not csa_tree_add_190_195_groupi_drc_bufs53234(csa_tree_add_190_195_groupi_n_562 ,csa_tree_add_190_195_groupi_n_2296);
  not csa_tree_add_190_195_groupi_drc_bufs53236(csa_tree_add_190_195_groupi_n_561 ,csa_tree_add_190_195_groupi_n_559);
  not csa_tree_add_190_195_groupi_drc_bufs53237(csa_tree_add_190_195_groupi_n_560 ,csa_tree_add_190_195_groupi_n_559);
  not csa_tree_add_190_195_groupi_drc_bufs53238(csa_tree_add_190_195_groupi_n_559 ,csa_tree_add_190_195_groupi_n_2233);
  not csa_tree_add_190_195_groupi_drc_bufs53240(csa_tree_add_190_195_groupi_n_558 ,csa_tree_add_190_195_groupi_n_557);
  not csa_tree_add_190_195_groupi_drc_bufs53242(csa_tree_add_190_195_groupi_n_557 ,csa_tree_add_190_195_groupi_n_2230);
  not csa_tree_add_190_195_groupi_drc_bufs53244(csa_tree_add_190_195_groupi_n_556 ,csa_tree_add_190_195_groupi_n_555);
  not csa_tree_add_190_195_groupi_drc_bufs53246(csa_tree_add_190_195_groupi_n_555 ,csa_tree_add_190_195_groupi_n_2324);
  not csa_tree_add_190_195_groupi_drc_bufs53248(csa_tree_add_190_195_groupi_n_554 ,csa_tree_add_190_195_groupi_n_553);
  not csa_tree_add_190_195_groupi_drc_bufs53250(csa_tree_add_190_195_groupi_n_553 ,csa_tree_add_190_195_groupi_n_2327);
  not csa_tree_add_190_195_groupi_drc_bufs53252(csa_tree_add_190_195_groupi_n_552 ,csa_tree_add_190_195_groupi_n_551);
  not csa_tree_add_190_195_groupi_drc_bufs53254(csa_tree_add_190_195_groupi_n_551 ,csa_tree_add_190_195_groupi_n_2305);
  not csa_tree_add_190_195_groupi_drc_bufs53256(csa_tree_add_190_195_groupi_n_550 ,csa_tree_add_190_195_groupi_n_548);
  not csa_tree_add_190_195_groupi_drc_bufs53257(csa_tree_add_190_195_groupi_n_549 ,csa_tree_add_190_195_groupi_n_548);
  not csa_tree_add_190_195_groupi_drc_bufs53258(csa_tree_add_190_195_groupi_n_548 ,csa_tree_add_190_195_groupi_n_2290);
  not csa_tree_add_190_195_groupi_drc_bufs53260(csa_tree_add_190_195_groupi_n_547 ,csa_tree_add_190_195_groupi_n_545);
  not csa_tree_add_190_195_groupi_drc_bufs53261(csa_tree_add_190_195_groupi_n_546 ,csa_tree_add_190_195_groupi_n_545);
  not csa_tree_add_190_195_groupi_drc_bufs53262(csa_tree_add_190_195_groupi_n_545 ,csa_tree_add_190_195_groupi_n_2290);
  not csa_tree_add_190_195_groupi_drc_bufs53264(csa_tree_add_190_195_groupi_n_544 ,csa_tree_add_190_195_groupi_n_542);
  not csa_tree_add_190_195_groupi_drc_bufs53265(csa_tree_add_190_195_groupi_n_543 ,csa_tree_add_190_195_groupi_n_542);
  not csa_tree_add_190_195_groupi_drc_bufs53266(csa_tree_add_190_195_groupi_n_542 ,csa_tree_add_190_195_groupi_n_2284);
  not csa_tree_add_190_195_groupi_drc_bufs53268(csa_tree_add_190_195_groupi_n_541 ,csa_tree_add_190_195_groupi_n_539);
  not csa_tree_add_190_195_groupi_drc_bufs53269(csa_tree_add_190_195_groupi_n_540 ,csa_tree_add_190_195_groupi_n_539);
  not csa_tree_add_190_195_groupi_drc_bufs53270(csa_tree_add_190_195_groupi_n_539 ,csa_tree_add_190_195_groupi_n_2291);
  not csa_tree_add_190_195_groupi_drc_bufs53272(csa_tree_add_190_195_groupi_n_538 ,csa_tree_add_190_195_groupi_n_536);
  not csa_tree_add_190_195_groupi_drc_bufs53273(csa_tree_add_190_195_groupi_n_537 ,csa_tree_add_190_195_groupi_n_536);
  not csa_tree_add_190_195_groupi_drc_bufs53274(csa_tree_add_190_195_groupi_n_536 ,csa_tree_add_190_195_groupi_n_2282);
  not csa_tree_add_190_195_groupi_drc_bufs53276(csa_tree_add_190_195_groupi_n_535 ,csa_tree_add_190_195_groupi_n_534);
  not csa_tree_add_190_195_groupi_drc_bufs53278(csa_tree_add_190_195_groupi_n_534 ,csa_tree_add_190_195_groupi_n_2205);
  not csa_tree_add_190_195_groupi_drc_bufs53280(csa_tree_add_190_195_groupi_n_533 ,csa_tree_add_190_195_groupi_n_532);
  not csa_tree_add_190_195_groupi_drc_bufs53282(csa_tree_add_190_195_groupi_n_532 ,csa_tree_add_190_195_groupi_n_2261);
  not csa_tree_add_190_195_groupi_drc_bufs53284(csa_tree_add_190_195_groupi_n_531 ,csa_tree_add_190_195_groupi_n_530);
  not csa_tree_add_190_195_groupi_drc_bufs53286(csa_tree_add_190_195_groupi_n_530 ,csa_tree_add_190_195_groupi_n_2258);
  not csa_tree_add_190_195_groupi_drc_bufs53288(csa_tree_add_190_195_groupi_n_529 ,csa_tree_add_190_195_groupi_n_527);
  not csa_tree_add_190_195_groupi_drc_bufs53289(csa_tree_add_190_195_groupi_n_528 ,csa_tree_add_190_195_groupi_n_527);
  not csa_tree_add_190_195_groupi_drc_bufs53290(csa_tree_add_190_195_groupi_n_527 ,csa_tree_add_190_195_groupi_n_2285);
  not csa_tree_add_190_195_groupi_drc_bufs53292(csa_tree_add_190_195_groupi_n_526 ,csa_tree_add_190_195_groupi_n_525);
  not csa_tree_add_190_195_groupi_drc_bufs53294(csa_tree_add_190_195_groupi_n_525 ,csa_tree_add_190_195_groupi_n_2269);
  not csa_tree_add_190_195_groupi_drc_bufs53296(csa_tree_add_190_195_groupi_n_524 ,csa_tree_add_190_195_groupi_n_523);
  not csa_tree_add_190_195_groupi_drc_bufs53298(csa_tree_add_190_195_groupi_n_523 ,csa_tree_add_190_195_groupi_n_2273);
  not csa_tree_add_190_195_groupi_drc_bufs53300(csa_tree_add_190_195_groupi_n_522 ,csa_tree_add_190_195_groupi_n_520);
  not csa_tree_add_190_195_groupi_drc_bufs53301(csa_tree_add_190_195_groupi_n_521 ,csa_tree_add_190_195_groupi_n_520);
  not csa_tree_add_190_195_groupi_drc_bufs53302(csa_tree_add_190_195_groupi_n_520 ,csa_tree_add_190_195_groupi_n_2264);
  not csa_tree_add_190_195_groupi_drc_bufs53304(csa_tree_add_190_195_groupi_n_519 ,csa_tree_add_190_195_groupi_n_517);
  not csa_tree_add_190_195_groupi_drc_bufs53305(csa_tree_add_190_195_groupi_n_518 ,csa_tree_add_190_195_groupi_n_517);
  not csa_tree_add_190_195_groupi_drc_bufs53306(csa_tree_add_190_195_groupi_n_517 ,csa_tree_add_190_195_groupi_n_2252);
  not csa_tree_add_190_195_groupi_drc_bufs53308(csa_tree_add_190_195_groupi_n_516 ,csa_tree_add_190_195_groupi_n_515);
  not csa_tree_add_190_195_groupi_drc_bufs53310(csa_tree_add_190_195_groupi_n_515 ,csa_tree_add_190_195_groupi_n_2190);
  not csa_tree_add_190_195_groupi_drc_bufs53312(csa_tree_add_190_195_groupi_n_514 ,csa_tree_add_190_195_groupi_n_513);
  not csa_tree_add_190_195_groupi_drc_bufs53314(csa_tree_add_190_195_groupi_n_513 ,csa_tree_add_190_195_groupi_n_2257);
  not csa_tree_add_190_195_groupi_drc_bufs53316(csa_tree_add_190_195_groupi_n_512 ,csa_tree_add_190_195_groupi_n_511);
  not csa_tree_add_190_195_groupi_drc_bufs53318(csa_tree_add_190_195_groupi_n_511 ,csa_tree_add_190_195_groupi_n_2260);
  not csa_tree_add_190_195_groupi_drc_bufs53320(csa_tree_add_190_195_groupi_n_510 ,csa_tree_add_190_195_groupi_n_509);
  not csa_tree_add_190_195_groupi_drc_bufs53322(csa_tree_add_190_195_groupi_n_509 ,csa_tree_add_190_195_groupi_n_2281);
  not csa_tree_add_190_195_groupi_drc_bufs53324(csa_tree_add_190_195_groupi_n_508 ,csa_tree_add_190_195_groupi_n_507);
  not csa_tree_add_190_195_groupi_drc_bufs53326(csa_tree_add_190_195_groupi_n_507 ,csa_tree_add_190_195_groupi_n_2284);
  not csa_tree_add_190_195_groupi_drc_bufs53328(csa_tree_add_190_195_groupi_n_506 ,csa_tree_add_190_195_groupi_n_505);
  not csa_tree_add_190_195_groupi_drc_bufs53330(csa_tree_add_190_195_groupi_n_505 ,csa_tree_add_190_195_groupi_n_2121);
  not csa_tree_add_190_195_groupi_drc_bufs53332(csa_tree_add_190_195_groupi_n_504 ,csa_tree_add_190_195_groupi_n_503);
  not csa_tree_add_190_195_groupi_drc_bufs53334(csa_tree_add_190_195_groupi_n_503 ,csa_tree_add_190_195_groupi_n_2267);
  not csa_tree_add_190_195_groupi_drc_bufs53336(csa_tree_add_190_195_groupi_n_502 ,csa_tree_add_190_195_groupi_n_500);
  not csa_tree_add_190_195_groupi_drc_bufs53337(csa_tree_add_190_195_groupi_n_501 ,csa_tree_add_190_195_groupi_n_500);
  not csa_tree_add_190_195_groupi_drc_bufs53338(csa_tree_add_190_195_groupi_n_500 ,csa_tree_add_190_195_groupi_n_2266);
  not csa_tree_add_190_195_groupi_drc_bufs53340(csa_tree_add_190_195_groupi_n_499 ,csa_tree_add_190_195_groupi_n_497);
  not csa_tree_add_190_195_groupi_drc_bufs53341(csa_tree_add_190_195_groupi_n_498 ,csa_tree_add_190_195_groupi_n_497);
  not csa_tree_add_190_195_groupi_drc_bufs53342(csa_tree_add_190_195_groupi_n_497 ,csa_tree_add_190_195_groupi_n_2276);
  not csa_tree_add_190_195_groupi_drc_bufs53344(csa_tree_add_190_195_groupi_n_496 ,csa_tree_add_190_195_groupi_n_494);
  not csa_tree_add_190_195_groupi_drc_bufs53345(csa_tree_add_190_195_groupi_n_495 ,csa_tree_add_190_195_groupi_n_494);
  not csa_tree_add_190_195_groupi_drc_bufs53346(csa_tree_add_190_195_groupi_n_494 ,csa_tree_add_190_195_groupi_n_2078);
  not csa_tree_add_190_195_groupi_drc_bufs53348(csa_tree_add_190_195_groupi_n_493 ,csa_tree_add_190_195_groupi_n_492);
  not csa_tree_add_190_195_groupi_drc_bufs53350(csa_tree_add_190_195_groupi_n_492 ,csa_tree_add_190_195_groupi_n_2272);
  not csa_tree_add_190_195_groupi_drc_bufs53352(csa_tree_add_190_195_groupi_n_491 ,csa_tree_add_190_195_groupi_n_489);
  not csa_tree_add_190_195_groupi_drc_bufs53353(csa_tree_add_190_195_groupi_n_490 ,csa_tree_add_190_195_groupi_n_489);
  not csa_tree_add_190_195_groupi_drc_bufs53354(csa_tree_add_190_195_groupi_n_489 ,csa_tree_add_190_195_groupi_n_2077);
  not csa_tree_add_190_195_groupi_drc_bufs53356(csa_tree_add_190_195_groupi_n_488 ,csa_tree_add_190_195_groupi_n_487);
  not csa_tree_add_190_195_groupi_drc_bufs53358(csa_tree_add_190_195_groupi_n_487 ,csa_tree_add_190_195_groupi_n_2102);
  not csa_tree_add_190_195_groupi_drc_bufs53360(csa_tree_add_190_195_groupi_n_486 ,csa_tree_add_190_195_groupi_n_484);
  not csa_tree_add_190_195_groupi_drc_bufs53361(csa_tree_add_190_195_groupi_n_485 ,csa_tree_add_190_195_groupi_n_484);
  not csa_tree_add_190_195_groupi_drc_bufs53362(csa_tree_add_190_195_groupi_n_484 ,csa_tree_add_190_195_groupi_n_2227);
  not csa_tree_add_190_195_groupi_drc_bufs53364(csa_tree_add_190_195_groupi_n_483 ,csa_tree_add_190_195_groupi_n_481);
  not csa_tree_add_190_195_groupi_drc_bufs53365(csa_tree_add_190_195_groupi_n_482 ,csa_tree_add_190_195_groupi_n_481);
  not csa_tree_add_190_195_groupi_drc_bufs53366(csa_tree_add_190_195_groupi_n_481 ,csa_tree_add_190_195_groupi_n_2311);
  not csa_tree_add_190_195_groupi_drc_bufs53368(csa_tree_add_190_195_groupi_n_480 ,csa_tree_add_190_195_groupi_n_478);
  not csa_tree_add_190_195_groupi_drc_bufs53369(csa_tree_add_190_195_groupi_n_479 ,csa_tree_add_190_195_groupi_n_478);
  not csa_tree_add_190_195_groupi_drc_bufs53370(csa_tree_add_190_195_groupi_n_478 ,csa_tree_add_190_195_groupi_n_2236);
  not csa_tree_add_190_195_groupi_drc_bufs53372(csa_tree_add_190_195_groupi_n_477 ,csa_tree_add_190_195_groupi_n_476);
  not csa_tree_add_190_195_groupi_drc_bufs53374(csa_tree_add_190_195_groupi_n_476 ,csa_tree_add_190_195_groupi_n_2202);
  not csa_tree_add_190_195_groupi_drc_bufs53376(csa_tree_add_190_195_groupi_n_475 ,csa_tree_add_190_195_groupi_n_474);
  not csa_tree_add_190_195_groupi_drc_bufs53378(csa_tree_add_190_195_groupi_n_474 ,csa_tree_add_190_195_groupi_n_2208);
  not csa_tree_add_190_195_groupi_drc_bufs53380(csa_tree_add_190_195_groupi_n_473 ,csa_tree_add_190_195_groupi_n_471);
  not csa_tree_add_190_195_groupi_drc_bufs53381(csa_tree_add_190_195_groupi_n_472 ,csa_tree_add_190_195_groupi_n_471);
  not csa_tree_add_190_195_groupi_drc_bufs53382(csa_tree_add_190_195_groupi_n_471 ,csa_tree_add_190_195_groupi_n_2257);
  not csa_tree_add_190_195_groupi_drc_bufs53384(csa_tree_add_190_195_groupi_n_470 ,csa_tree_add_190_195_groupi_n_2329);
  not csa_tree_add_190_195_groupi_drc_bufs53386(csa_tree_add_190_195_groupi_n_2329 ,csa_tree_add_190_195_groupi_n_2258);
  not csa_tree_add_190_195_groupi_drc_bufs53388(csa_tree_add_190_195_groupi_n_469 ,csa_tree_add_190_195_groupi_n_467);
  not csa_tree_add_190_195_groupi_drc_bufs53389(csa_tree_add_190_195_groupi_n_468 ,csa_tree_add_190_195_groupi_n_467);
  not csa_tree_add_190_195_groupi_drc_bufs53390(csa_tree_add_190_195_groupi_n_467 ,csa_tree_add_190_195_groupi_n_2306);
  not csa_tree_add_190_195_groupi_drc_bufs53392(csa_tree_add_190_195_groupi_n_466 ,csa_tree_add_190_195_groupi_n_2331);
  not csa_tree_add_190_195_groupi_drc_bufs53394(csa_tree_add_190_195_groupi_n_2331 ,csa_tree_add_190_195_groupi_n_2282);
  not csa_tree_add_190_195_groupi_drc_bufs53396(csa_tree_add_190_195_groupi_n_465 ,csa_tree_add_190_195_groupi_n_2334);
  not csa_tree_add_190_195_groupi_drc_bufs53398(csa_tree_add_190_195_groupi_n_2334 ,csa_tree_add_190_195_groupi_n_2255);
  not csa_tree_add_190_195_groupi_drc_bufs53400(csa_tree_add_190_195_groupi_n_464 ,csa_tree_add_190_195_groupi_n_2333);
  not csa_tree_add_190_195_groupi_drc_bufs53402(csa_tree_add_190_195_groupi_n_2333 ,csa_tree_add_190_195_groupi_n_2208);
  not csa_tree_add_190_195_groupi_drc_bufs53404(csa_tree_add_190_195_groupi_n_463 ,csa_tree_add_190_195_groupi_n_462);
  not csa_tree_add_190_195_groupi_drc_bufs53406(csa_tree_add_190_195_groupi_n_462 ,csa_tree_add_190_195_groupi_n_2326);
  not csa_tree_add_190_195_groupi_drc_bufs53408(csa_tree_add_190_195_groupi_n_461 ,csa_tree_add_190_195_groupi_n_460);
  not csa_tree_add_190_195_groupi_drc_bufs53410(csa_tree_add_190_195_groupi_n_460 ,csa_tree_add_190_195_groupi_n_2279);
  not csa_tree_add_190_195_groupi_drc_bufs53412(csa_tree_add_190_195_groupi_n_459 ,csa_tree_add_190_195_groupi_n_2359);
  not csa_tree_add_190_195_groupi_drc_bufs53414(csa_tree_add_190_195_groupi_n_2359 ,csa_tree_add_190_195_groupi_n_2261);
  not csa_tree_add_190_195_groupi_drc_bufs53416(csa_tree_add_190_195_groupi_n_458 ,csa_tree_add_190_195_groupi_n_2364);
  not csa_tree_add_190_195_groupi_drc_bufs53418(csa_tree_add_190_195_groupi_n_2364 ,csa_tree_add_190_195_groupi_n_2272);
  not csa_tree_add_190_195_groupi_drc_bufs53420(csa_tree_add_190_195_groupi_n_457 ,csa_tree_add_190_195_groupi_n_455);
  not csa_tree_add_190_195_groupi_drc_bufs53421(csa_tree_add_190_195_groupi_n_456 ,csa_tree_add_190_195_groupi_n_455);
  not csa_tree_add_190_195_groupi_drc_bufs53422(csa_tree_add_190_195_groupi_n_455 ,csa_tree_add_190_195_groupi_n_2234);
  not csa_tree_add_190_195_groupi_drc_bufs53424(csa_tree_add_190_195_groupi_n_454 ,csa_tree_add_190_195_groupi_n_2330);
  not csa_tree_add_190_195_groupi_drc_bufs53426(csa_tree_add_190_195_groupi_n_2330 ,csa_tree_add_190_195_groupi_n_2285);
  not csa_tree_add_190_195_groupi_drc_bufs53428(csa_tree_add_190_195_groupi_n_453 ,csa_tree_add_190_195_groupi_n_452);
  not csa_tree_add_190_195_groupi_drc_bufs53430(csa_tree_add_190_195_groupi_n_452 ,csa_tree_add_190_195_groupi_n_2306);
  not csa_tree_add_190_195_groupi_drc_bufs53432(csa_tree_add_190_195_groupi_n_451 ,csa_tree_add_190_195_groupi_n_450);
  not csa_tree_add_190_195_groupi_drc_bufs53434(csa_tree_add_190_195_groupi_n_450 ,csa_tree_add_190_195_groupi_n_2315);
  not csa_tree_add_190_195_groupi_drc_bufs53436(csa_tree_add_190_195_groupi_n_449 ,csa_tree_add_190_195_groupi_n_447);
  not csa_tree_add_190_195_groupi_drc_bufs53437(csa_tree_add_190_195_groupi_n_448 ,csa_tree_add_190_195_groupi_n_447);
  not csa_tree_add_190_195_groupi_drc_bufs53438(csa_tree_add_190_195_groupi_n_447 ,csa_tree_add_190_195_groupi_n_2205);
  not csa_tree_add_190_195_groupi_drc_bufs53440(csa_tree_add_190_195_groupi_n_446 ,csa_tree_add_190_195_groupi_n_444);
  not csa_tree_add_190_195_groupi_drc_bufs53441(csa_tree_add_190_195_groupi_n_445 ,csa_tree_add_190_195_groupi_n_444);
  not csa_tree_add_190_195_groupi_drc_bufs53442(csa_tree_add_190_195_groupi_n_444 ,csa_tree_add_190_195_groupi_n_2309);
  not csa_tree_add_190_195_groupi_drc_bufs53444(csa_tree_add_190_195_groupi_n_443 ,csa_tree_add_190_195_groupi_n_441);
  not csa_tree_add_190_195_groupi_drc_bufs53445(csa_tree_add_190_195_groupi_n_442 ,csa_tree_add_190_195_groupi_n_441);
  not csa_tree_add_190_195_groupi_drc_bufs53446(csa_tree_add_190_195_groupi_n_441 ,csa_tree_add_190_195_groupi_n_2303);
  not csa_tree_add_190_195_groupi_drc_bufs53448(csa_tree_add_190_195_groupi_n_440 ,csa_tree_add_190_195_groupi_n_438);
  not csa_tree_add_190_195_groupi_drc_bufs53449(csa_tree_add_190_195_groupi_n_439 ,csa_tree_add_190_195_groupi_n_438);
  not csa_tree_add_190_195_groupi_drc_bufs53450(csa_tree_add_190_195_groupi_n_438 ,csa_tree_add_190_195_groupi_n_2299);
  not csa_tree_add_190_195_groupi_drc_bufs53452(csa_tree_add_190_195_groupi_n_437 ,csa_tree_add_190_195_groupi_n_2335);
  not csa_tree_add_190_195_groupi_drc_bufs53454(csa_tree_add_190_195_groupi_n_2335 ,csa_tree_add_190_195_groupi_n_2122);
  not csa_tree_add_190_195_groupi_drc_bufs53456(csa_tree_add_190_195_groupi_n_436 ,csa_tree_add_190_195_groupi_n_2366);
  not csa_tree_add_190_195_groupi_drc_bufs53458(csa_tree_add_190_195_groupi_n_2366 ,csa_tree_add_190_195_groupi_n_2251);
  not csa_tree_add_190_195_groupi_drc_bufs53460(csa_tree_add_190_195_groupi_n_435 ,csa_tree_add_190_195_groupi_n_433);
  not csa_tree_add_190_195_groupi_drc_bufs53461(csa_tree_add_190_195_groupi_n_434 ,csa_tree_add_190_195_groupi_n_433);
  not csa_tree_add_190_195_groupi_drc_bufs53462(csa_tree_add_190_195_groupi_n_433 ,csa_tree_add_190_195_groupi_n_2321);
  not csa_tree_add_190_195_groupi_drc_bufs53464(csa_tree_add_190_195_groupi_n_432 ,csa_tree_add_190_195_groupi_n_430);
  not csa_tree_add_190_195_groupi_drc_bufs53465(csa_tree_add_190_195_groupi_n_431 ,csa_tree_add_190_195_groupi_n_430);
  not csa_tree_add_190_195_groupi_drc_bufs53466(csa_tree_add_190_195_groupi_n_430 ,csa_tree_add_190_195_groupi_n_2297);
  not csa_tree_add_190_195_groupi_drc_bufs53468(csa_tree_add_190_195_groupi_n_429 ,csa_tree_add_190_195_groupi_n_427);
  not csa_tree_add_190_195_groupi_drc_bufs53469(csa_tree_add_190_195_groupi_n_428 ,csa_tree_add_190_195_groupi_n_427);
  not csa_tree_add_190_195_groupi_drc_bufs53470(csa_tree_add_190_195_groupi_n_427 ,csa_tree_add_190_195_groupi_n_2275);
  not csa_tree_add_190_195_groupi_drc_bufs53472(csa_tree_add_190_195_groupi_n_426 ,csa_tree_add_190_195_groupi_n_424);
  not csa_tree_add_190_195_groupi_drc_bufs53473(csa_tree_add_190_195_groupi_n_425 ,csa_tree_add_190_195_groupi_n_424);
  not csa_tree_add_190_195_groupi_drc_bufs53474(csa_tree_add_190_195_groupi_n_424 ,csa_tree_add_190_195_groupi_n_2323);
  not csa_tree_add_190_195_groupi_drc_bufs53476(csa_tree_add_190_195_groupi_n_423 ,csa_tree_add_190_195_groupi_n_421);
  not csa_tree_add_190_195_groupi_drc_bufs53477(csa_tree_add_190_195_groupi_n_422 ,csa_tree_add_190_195_groupi_n_421);
  not csa_tree_add_190_195_groupi_drc_bufs53478(csa_tree_add_190_195_groupi_n_421 ,csa_tree_add_190_195_groupi_n_2201);
  not csa_tree_add_190_195_groupi_drc_bufs53480(csa_tree_add_190_195_groupi_n_420 ,csa_tree_add_190_195_groupi_n_2339);
  not csa_tree_add_190_195_groupi_drc_bufs53482(csa_tree_add_190_195_groupi_n_2339 ,csa_tree_add_190_195_groupi_n_2278);
  not csa_tree_add_190_195_groupi_drc_bufs53484(csa_tree_add_190_195_groupi_n_419 ,csa_tree_add_190_195_groupi_n_418);
  not csa_tree_add_190_195_groupi_drc_bufs53486(csa_tree_add_190_195_groupi_n_418 ,csa_tree_add_190_195_groupi_n_2270);
  not csa_tree_add_190_195_groupi_drc_bufs53488(csa_tree_add_190_195_groupi_n_417 ,csa_tree_add_190_195_groupi_n_415);
  not csa_tree_add_190_195_groupi_drc_bufs53489(csa_tree_add_190_195_groupi_n_416 ,csa_tree_add_190_195_groupi_n_415);
  not csa_tree_add_190_195_groupi_drc_bufs53490(csa_tree_add_190_195_groupi_n_415 ,csa_tree_add_190_195_groupi_n_2204);
  not csa_tree_add_190_195_groupi_drc_bufs53493(csa_tree_add_190_195_groupi_n_414 ,csa_tree_add_190_195_groupi_n_413);
  not csa_tree_add_190_195_groupi_drc_bufs53494(csa_tree_add_190_195_groupi_n_413 ,csa_tree_add_190_195_groupi_n_2294);
  not csa_tree_add_190_195_groupi_drc_bufs53496(csa_tree_add_190_195_groupi_n_412 ,csa_tree_add_190_195_groupi_n_410);
  not csa_tree_add_190_195_groupi_drc_bufs53497(csa_tree_add_190_195_groupi_n_411 ,csa_tree_add_190_195_groupi_n_410);
  not csa_tree_add_190_195_groupi_drc_bufs53498(csa_tree_add_190_195_groupi_n_410 ,csa_tree_add_190_195_groupi_n_2293);
  not csa_tree_add_190_195_groupi_drc_bufs53501(csa_tree_add_190_195_groupi_n_409 ,csa_tree_add_190_195_groupi_n_408);
  not csa_tree_add_190_195_groupi_drc_bufs53502(csa_tree_add_190_195_groupi_n_408 ,csa_tree_add_190_195_groupi_n_2181);
  not csa_tree_add_190_195_groupi_drc_bufs53505(csa_tree_add_190_195_groupi_n_407 ,csa_tree_add_190_195_groupi_n_406);
  not csa_tree_add_190_195_groupi_drc_bufs53506(csa_tree_add_190_195_groupi_n_406 ,csa_tree_add_190_195_groupi_n_2177);
  not csa_tree_add_190_195_groupi_drc_bufs53509(csa_tree_add_190_195_groupi_n_405 ,csa_tree_add_190_195_groupi_n_404);
  not csa_tree_add_190_195_groupi_drc_bufs53510(csa_tree_add_190_195_groupi_n_404 ,csa_tree_add_190_195_groupi_n_2161);
  not csa_tree_add_190_195_groupi_drc_bufs53513(csa_tree_add_190_195_groupi_n_403 ,csa_tree_add_190_195_groupi_n_402);
  not csa_tree_add_190_195_groupi_drc_bufs53514(csa_tree_add_190_195_groupi_n_402 ,csa_tree_add_190_195_groupi_n_2297);
  not csa_tree_add_190_195_groupi_drc_bufs53517(csa_tree_add_190_195_groupi_n_401 ,csa_tree_add_190_195_groupi_n_400);
  not csa_tree_add_190_195_groupi_drc_bufs53518(csa_tree_add_190_195_groupi_n_400 ,csa_tree_add_190_195_groupi_n_2296);
  not csa_tree_add_190_195_groupi_drc_bufs53520(csa_tree_add_190_195_groupi_n_399 ,csa_tree_add_190_195_groupi_n_397);
  not csa_tree_add_190_195_groupi_drc_bufs53521(csa_tree_add_190_195_groupi_n_398 ,csa_tree_add_190_195_groupi_n_397);
  not csa_tree_add_190_195_groupi_drc_bufs53522(csa_tree_add_190_195_groupi_n_397 ,csa_tree_add_190_195_groupi_n_2312);
  not csa_tree_add_190_195_groupi_drc_bufs53525(csa_tree_add_190_195_groupi_n_396 ,csa_tree_add_190_195_groupi_n_395);
  not csa_tree_add_190_195_groupi_drc_bufs53526(csa_tree_add_190_195_groupi_n_395 ,csa_tree_add_190_195_groupi_n_2108);
  not csa_tree_add_190_195_groupi_drc_bufs53528(csa_tree_add_190_195_groupi_n_394 ,csa_tree_add_190_195_groupi_n_392);
  not csa_tree_add_190_195_groupi_drc_bufs53529(csa_tree_add_190_195_groupi_n_393 ,csa_tree_add_190_195_groupi_n_392);
  not csa_tree_add_190_195_groupi_drc_bufs53530(csa_tree_add_190_195_groupi_n_392 ,csa_tree_add_190_195_groupi_n_2237);
  not csa_tree_add_190_195_groupi_drc_bufs53533(csa_tree_add_190_195_groupi_n_391 ,csa_tree_add_190_195_groupi_n_390);
  not csa_tree_add_190_195_groupi_drc_bufs53534(csa_tree_add_190_195_groupi_n_390 ,csa_tree_add_190_195_groupi_n_2151);
  not csa_tree_add_190_195_groupi_drc_bufs53537(csa_tree_add_190_195_groupi_n_389 ,csa_tree_add_190_195_groupi_n_388);
  not csa_tree_add_190_195_groupi_drc_bufs53538(csa_tree_add_190_195_groupi_n_388 ,csa_tree_add_190_195_groupi_n_2111);
  not csa_tree_add_190_195_groupi_drc_bufs53540(csa_tree_add_190_195_groupi_n_387 ,csa_tree_add_190_195_groupi_n_385);
  not csa_tree_add_190_195_groupi_drc_bufs53541(csa_tree_add_190_195_groupi_n_386 ,csa_tree_add_190_195_groupi_n_385);
  not csa_tree_add_190_195_groupi_drc_bufs53542(csa_tree_add_190_195_groupi_n_385 ,csa_tree_add_190_195_groupi_n_2106);
  not csa_tree_add_190_195_groupi_drc_bufs53545(csa_tree_add_190_195_groupi_n_384 ,csa_tree_add_190_195_groupi_n_383);
  not csa_tree_add_190_195_groupi_drc_bufs53546(csa_tree_add_190_195_groupi_n_383 ,csa_tree_add_190_195_groupi_n_2236);
  not csa_tree_add_190_195_groupi_drc_bufs53549(csa_tree_add_190_195_groupi_n_382 ,csa_tree_add_190_195_groupi_n_381);
  not csa_tree_add_190_195_groupi_drc_bufs53550(csa_tree_add_190_195_groupi_n_381 ,csa_tree_add_190_195_groupi_n_2233);
  not csa_tree_add_190_195_groupi_drc_bufs53553(csa_tree_add_190_195_groupi_n_380 ,csa_tree_add_190_195_groupi_n_379);
  not csa_tree_add_190_195_groupi_drc_bufs53554(csa_tree_add_190_195_groupi_n_379 ,csa_tree_add_190_195_groupi_n_2115);
  not csa_tree_add_190_195_groupi_drc_bufs53556(csa_tree_add_190_195_groupi_n_378 ,csa_tree_add_190_195_groupi_n_376);
  not csa_tree_add_190_195_groupi_drc_bufs53557(csa_tree_add_190_195_groupi_n_377 ,csa_tree_add_190_195_groupi_n_376);
  not csa_tree_add_190_195_groupi_drc_bufs53558(csa_tree_add_190_195_groupi_n_376 ,csa_tree_add_190_195_groupi_n_2150);
  not csa_tree_add_190_195_groupi_drc_bufs53561(csa_tree_add_190_195_groupi_n_375 ,csa_tree_add_190_195_groupi_n_374);
  not csa_tree_add_190_195_groupi_drc_bufs53562(csa_tree_add_190_195_groupi_n_374 ,csa_tree_add_190_195_groupi_n_2281);
  not csa_tree_add_190_195_groupi_drc_bufs53565(csa_tree_add_190_195_groupi_n_373 ,csa_tree_add_190_195_groupi_n_372);
  not csa_tree_add_190_195_groupi_drc_bufs53566(csa_tree_add_190_195_groupi_n_372 ,csa_tree_add_190_195_groupi_n_2269);
  not csa_tree_add_190_195_groupi_drc_bufs53568(csa_tree_add_190_195_groupi_n_371 ,csa_tree_add_190_195_groupi_n_369);
  not csa_tree_add_190_195_groupi_drc_bufs53569(csa_tree_add_190_195_groupi_n_370 ,csa_tree_add_190_195_groupi_n_369);
  not csa_tree_add_190_195_groupi_drc_bufs53570(csa_tree_add_190_195_groupi_n_369 ,csa_tree_add_190_195_groupi_n_2273);
  not csa_tree_add_190_195_groupi_drc_bufs53573(csa_tree_add_190_195_groupi_n_368 ,csa_tree_add_190_195_groupi_n_367);
  not csa_tree_add_190_195_groupi_drc_bufs53574(csa_tree_add_190_195_groupi_n_367 ,csa_tree_add_190_195_groupi_n_2186);
  not csa_tree_add_190_195_groupi_drc_bufs53577(csa_tree_add_190_195_groupi_n_366 ,csa_tree_add_190_195_groupi_n_365);
  not csa_tree_add_190_195_groupi_drc_bufs53578(csa_tree_add_190_195_groupi_n_365 ,csa_tree_add_190_195_groupi_n_2207);
  not csa_tree_add_190_195_groupi_drc_bufs53581(csa_tree_add_190_195_groupi_n_364 ,csa_tree_add_190_195_groupi_n_363);
  not csa_tree_add_190_195_groupi_drc_bufs53582(csa_tree_add_190_195_groupi_n_363 ,csa_tree_add_190_195_groupi_n_2074);
  not csa_tree_add_190_195_groupi_drc_bufs53585(csa_tree_add_190_195_groupi_n_362 ,csa_tree_add_190_195_groupi_n_361);
  not csa_tree_add_190_195_groupi_drc_bufs53586(csa_tree_add_190_195_groupi_n_361 ,csa_tree_add_190_195_groupi_n_2254);
  not csa_tree_add_190_195_groupi_drc_bufs53589(csa_tree_add_190_195_groupi_n_360 ,csa_tree_add_190_195_groupi_n_359);
  not csa_tree_add_190_195_groupi_drc_bufs53590(csa_tree_add_190_195_groupi_n_359 ,csa_tree_add_190_195_groupi_n_2249);
  not csa_tree_add_190_195_groupi_drc_bufs53593(csa_tree_add_190_195_groupi_n_358 ,csa_tree_add_190_195_groupi_n_357);
  not csa_tree_add_190_195_groupi_drc_bufs53594(csa_tree_add_190_195_groupi_n_357 ,csa_tree_add_190_195_groupi_n_2308);
  not csa_tree_add_190_195_groupi_drc_bufs53596(csa_tree_add_190_195_groupi_n_356 ,csa_tree_add_190_195_groupi_n_354);
  not csa_tree_add_190_195_groupi_drc_bufs53597(csa_tree_add_190_195_groupi_n_355 ,csa_tree_add_190_195_groupi_n_354);
  not csa_tree_add_190_195_groupi_drc_bufs53598(csa_tree_add_190_195_groupi_n_354 ,csa_tree_add_190_195_groupi_n_2072);
  not csa_tree_add_190_195_groupi_drc_bufs53601(csa_tree_add_190_195_groupi_n_353 ,csa_tree_add_190_195_groupi_n_352);
  not csa_tree_add_190_195_groupi_drc_bufs53602(csa_tree_add_190_195_groupi_n_352 ,csa_tree_add_190_195_groupi_n_2099);
  not csa_tree_add_190_195_groupi_drc_bufs53604(csa_tree_add_190_195_groupi_n_351 ,csa_tree_add_190_195_groupi_n_349);
  not csa_tree_add_190_195_groupi_drc_bufs53605(csa_tree_add_190_195_groupi_n_350 ,csa_tree_add_190_195_groupi_n_349);
  not csa_tree_add_190_195_groupi_drc_bufs53606(csa_tree_add_190_195_groupi_n_349 ,csa_tree_add_190_195_groupi_n_2093);
  not csa_tree_add_190_195_groupi_drc_bufs53608(csa_tree_add_190_195_groupi_n_348 ,csa_tree_add_190_195_groupi_n_346);
  not csa_tree_add_190_195_groupi_drc_bufs53609(csa_tree_add_190_195_groupi_n_347 ,csa_tree_add_190_195_groupi_n_346);
  not csa_tree_add_190_195_groupi_drc_bufs53610(csa_tree_add_190_195_groupi_n_346 ,csa_tree_add_190_195_groupi_n_2195);
  not csa_tree_add_190_195_groupi_drc_bufs53613(csa_tree_add_190_195_groupi_n_345 ,csa_tree_add_190_195_groupi_n_344);
  not csa_tree_add_190_195_groupi_drc_bufs53614(csa_tree_add_190_195_groupi_n_344 ,csa_tree_add_190_195_groupi_n_2300);
  not csa_tree_add_190_195_groupi_drc_bufs53616(csa_tree_add_190_195_groupi_n_343 ,csa_tree_add_190_195_groupi_n_341);
  not csa_tree_add_190_195_groupi_drc_bufs53617(csa_tree_add_190_195_groupi_n_342 ,csa_tree_add_190_195_groupi_n_341);
  not csa_tree_add_190_195_groupi_drc_bufs53618(csa_tree_add_190_195_groupi_n_341 ,csa_tree_add_190_195_groupi_n_2320);
  not csa_tree_add_190_195_groupi_drc_bufs53621(csa_tree_add_190_195_groupi_n_340 ,csa_tree_add_190_195_groupi_n_339);
  not csa_tree_add_190_195_groupi_drc_bufs53622(csa_tree_add_190_195_groupi_n_339 ,csa_tree_add_190_195_groupi_n_2187);
  not csa_tree_add_190_195_groupi_drc_bufs53625(csa_tree_add_190_195_groupi_n_338 ,csa_tree_add_190_195_groupi_n_337);
  not csa_tree_add_190_195_groupi_drc_bufs53626(csa_tree_add_190_195_groupi_n_337 ,csa_tree_add_190_195_groupi_n_2249);
  not csa_tree_add_190_195_groupi_drc_bufs53629(csa_tree_add_190_195_groupi_n_336 ,csa_tree_add_190_195_groupi_n_335);
  not csa_tree_add_190_195_groupi_drc_bufs53630(csa_tree_add_190_195_groupi_n_335 ,csa_tree_add_190_195_groupi_n_2184);
  not csa_tree_add_190_195_groupi_drc_bufs53633(csa_tree_add_190_195_groupi_n_334 ,csa_tree_add_190_195_groupi_n_333);
  not csa_tree_add_190_195_groupi_drc_bufs53634(csa_tree_add_190_195_groupi_n_333 ,csa_tree_add_190_195_groupi_n_2094);
  not csa_tree_add_190_195_groupi_drc_bufs53637(csa_tree_add_190_195_groupi_n_332 ,csa_tree_add_190_195_groupi_n_331);
  not csa_tree_add_190_195_groupi_drc_bufs53638(csa_tree_add_190_195_groupi_n_331 ,csa_tree_add_190_195_groupi_n_2266);
  not csa_tree_add_190_195_groupi_drc_bufs53641(csa_tree_add_190_195_groupi_n_330 ,csa_tree_add_190_195_groupi_n_329);
  not csa_tree_add_190_195_groupi_drc_bufs53642(csa_tree_add_190_195_groupi_n_329 ,csa_tree_add_190_195_groupi_n_2276);
  not csa_tree_add_190_195_groupi_drc_bufs53645(csa_tree_add_190_195_groupi_n_328 ,csa_tree_add_190_195_groupi_n_327);
  not csa_tree_add_190_195_groupi_drc_bufs53646(csa_tree_add_190_195_groupi_n_327 ,csa_tree_add_190_195_groupi_n_2190);
  not csa_tree_add_190_195_groupi_drc_bufs53648(csa_tree_add_190_195_groupi_n_326 ,csa_tree_add_190_195_groupi_n_324);
  not csa_tree_add_190_195_groupi_drc_bufs53649(csa_tree_add_190_195_groupi_n_325 ,csa_tree_add_190_195_groupi_n_324);
  not csa_tree_add_190_195_groupi_drc_bufs53650(csa_tree_add_190_195_groupi_n_324 ,csa_tree_add_190_195_groupi_n_2184);
  not csa_tree_add_190_195_groupi_drc_bufs53653(csa_tree_add_190_195_groupi_n_323 ,csa_tree_add_190_195_groupi_n_322);
  not csa_tree_add_190_195_groupi_drc_bufs53654(csa_tree_add_190_195_groupi_n_322 ,csa_tree_add_190_195_groupi_n_2263);
  not csa_tree_add_190_195_groupi_drc_bufs53657(csa_tree_add_190_195_groupi_n_321 ,csa_tree_add_190_195_groupi_n_320);
  not csa_tree_add_190_195_groupi_drc_bufs53658(csa_tree_add_190_195_groupi_n_320 ,csa_tree_add_190_195_groupi_n_2264);
  not csa_tree_add_190_195_groupi_drc_bufs53661(csa_tree_add_190_195_groupi_n_319 ,csa_tree_add_190_195_groupi_n_318);
  not csa_tree_add_190_195_groupi_drc_bufs53662(csa_tree_add_190_195_groupi_n_318 ,csa_tree_add_190_195_groupi_n_2248);
  not csa_tree_add_190_195_groupi_drc_bufs53665(csa_tree_add_190_195_groupi_n_317 ,csa_tree_add_190_195_groupi_n_316);
  not csa_tree_add_190_195_groupi_drc_bufs53666(csa_tree_add_190_195_groupi_n_316 ,csa_tree_add_190_195_groupi_n_2193);
  not csa_tree_add_190_195_groupi_drc_bufs53669(csa_tree_add_190_195_groupi_n_315 ,csa_tree_add_190_195_groupi_n_314);
  not csa_tree_add_190_195_groupi_drc_bufs53670(csa_tree_add_190_195_groupi_n_314 ,csa_tree_add_190_195_groupi_n_2069);
  not csa_tree_add_190_195_groupi_drc_bufs53672(csa_tree_add_190_195_groupi_n_313 ,csa_tree_add_190_195_groupi_n_311);
  not csa_tree_add_190_195_groupi_drc_bufs53673(csa_tree_add_190_195_groupi_n_312 ,csa_tree_add_190_195_groupi_n_311);
  not csa_tree_add_190_195_groupi_drc_bufs53674(csa_tree_add_190_195_groupi_n_311 ,csa_tree_add_190_195_groupi_n_2275);
  not csa_tree_add_190_195_groupi_drc_bufs53676(csa_tree_add_190_195_groupi_n_310 ,csa_tree_add_190_195_groupi_n_308);
  not csa_tree_add_190_195_groupi_drc_bufs53677(csa_tree_add_190_195_groupi_n_309 ,csa_tree_add_190_195_groupi_n_308);
  not csa_tree_add_190_195_groupi_drc_bufs53678(csa_tree_add_190_195_groupi_n_308 ,csa_tree_add_190_195_groupi_n_2183);
  not csa_tree_add_190_195_groupi_drc_bufs53681(csa_tree_add_190_195_groupi_n_307 ,csa_tree_add_190_195_groupi_n_306);
  not csa_tree_add_190_195_groupi_drc_bufs53682(csa_tree_add_190_195_groupi_n_306 ,csa_tree_add_190_195_groupi_n_2302);
  not csa_tree_add_190_195_groupi_drc_bufs53684(csa_tree_add_190_195_groupi_n_305 ,csa_tree_add_190_195_groupi_n_303);
  not csa_tree_add_190_195_groupi_drc_bufs53685(csa_tree_add_190_195_groupi_n_304 ,csa_tree_add_190_195_groupi_n_303);
  not csa_tree_add_190_195_groupi_drc_bufs53686(csa_tree_add_190_195_groupi_n_303 ,csa_tree_add_190_195_groupi_n_2202);
  not csa_tree_add_190_195_groupi_drc_bufs53688(csa_tree_add_190_195_groupi_n_302 ,csa_tree_add_190_195_groupi_n_2332);
  not csa_tree_add_190_195_groupi_drc_bufs53690(csa_tree_add_190_195_groupi_n_2332 ,csa_tree_add_190_195_groupi_n_2267);
  not csa_tree_add_190_195_groupi_drc_bufs53693(csa_tree_add_190_195_groupi_n_301 ,csa_tree_add_190_195_groupi_n_300);
  not csa_tree_add_190_195_groupi_drc_bufs53694(csa_tree_add_190_195_groupi_n_300 ,csa_tree_add_190_195_groupi_n_2255);
  not csa_tree_add_190_195_groupi_drc_bufs53697(csa_tree_add_190_195_groupi_n_299 ,csa_tree_add_190_195_groupi_n_298);
  not csa_tree_add_190_195_groupi_drc_bufs53698(csa_tree_add_190_195_groupi_n_298 ,csa_tree_add_190_195_groupi_n_2252);
  not csa_tree_add_190_195_groupi_drc_bufs53701(csa_tree_add_190_195_groupi_n_297 ,csa_tree_add_190_195_groupi_n_296);
  not csa_tree_add_190_195_groupi_drc_bufs53702(csa_tree_add_190_195_groupi_n_296 ,csa_tree_add_190_195_groupi_n_2279);
  not csa_tree_add_190_195_groupi_drc_bufs53705(csa_tree_add_190_195_groupi_n_295 ,csa_tree_add_190_195_groupi_n_294);
  not csa_tree_add_190_195_groupi_drc_bufs53706(csa_tree_add_190_195_groupi_n_294 ,csa_tree_add_190_195_groupi_n_2309);
  not csa_tree_add_190_195_groupi_drc_bufs53709(csa_tree_add_190_195_groupi_n_293 ,csa_tree_add_190_195_groupi_n_292);
  not csa_tree_add_190_195_groupi_drc_bufs53710(csa_tree_add_190_195_groupi_n_292 ,csa_tree_add_190_195_groupi_n_2278);
  not csa_tree_add_190_195_groupi_drc_bufs53713(csa_tree_add_190_195_groupi_n_291 ,csa_tree_add_190_195_groupi_n_290);
  not csa_tree_add_190_195_groupi_drc_bufs53714(csa_tree_add_190_195_groupi_n_290 ,csa_tree_add_190_195_groupi_n_2195);
  not csa_tree_add_190_195_groupi_drc_bufs53717(csa_tree_add_190_195_groupi_n_289 ,csa_tree_add_190_195_groupi_n_288);
  not csa_tree_add_190_195_groupi_drc_bufs53718(csa_tree_add_190_195_groupi_n_288 ,csa_tree_add_190_195_groupi_n_2251);
  not csa_tree_add_190_195_groupi_drc_bufs53720(csa_tree_add_190_195_groupi_n_287 ,csa_tree_add_190_195_groupi_n_285);
  not csa_tree_add_190_195_groupi_drc_bufs53721(csa_tree_add_190_195_groupi_n_286 ,csa_tree_add_190_195_groupi_n_285);
  not csa_tree_add_190_195_groupi_drc_bufs53722(csa_tree_add_190_195_groupi_n_285 ,csa_tree_add_190_195_groupi_n_2254);
  not csa_tree_add_190_195_groupi_drc_bufs53724(csa_tree_add_190_195_groupi_n_284 ,csa_tree_add_190_195_groupi_n_282);
  not csa_tree_add_190_195_groupi_drc_bufs53725(csa_tree_add_190_195_groupi_n_283 ,csa_tree_add_190_195_groupi_n_282);
  not csa_tree_add_190_195_groupi_drc_bufs53726(csa_tree_add_190_195_groupi_n_282 ,csa_tree_add_190_195_groupi_n_1940);
  not csa_tree_add_190_195_groupi_drc_bufs53729(csa_tree_add_190_195_groupi_n_281 ,csa_tree_add_190_195_groupi_n_280);
  not csa_tree_add_190_195_groupi_drc_bufs53730(csa_tree_add_190_195_groupi_n_280 ,csa_tree_add_190_195_groupi_n_2303);
  not csa_tree_add_190_195_groupi_drc_bufs53733(csa_tree_add_190_195_groupi_n_279 ,csa_tree_add_190_195_groupi_n_278);
  not csa_tree_add_190_195_groupi_drc_bufs53734(csa_tree_add_190_195_groupi_n_278 ,csa_tree_add_190_195_groupi_n_2288);
  not csa_tree_add_190_195_groupi_drc_bufs53736(csa_tree_add_190_195_groupi_n_277 ,csa_tree_add_190_195_groupi_n_275);
  not csa_tree_add_190_195_groupi_drc_bufs53737(csa_tree_add_190_195_groupi_n_276 ,csa_tree_add_190_195_groupi_n_275);
  not csa_tree_add_190_195_groupi_drc_bufs53738(csa_tree_add_190_195_groupi_n_275 ,csa_tree_add_190_195_groupi_n_2068);
  not csa_tree_add_190_195_groupi_drc_bufs53740(csa_tree_add_190_195_groupi_n_274 ,csa_tree_add_190_195_groupi_n_272);
  not csa_tree_add_190_195_groupi_drc_bufs53741(csa_tree_add_190_195_groupi_n_273 ,csa_tree_add_190_195_groupi_n_272);
  not csa_tree_add_190_195_groupi_drc_bufs53742(csa_tree_add_190_195_groupi_n_272 ,csa_tree_add_190_195_groupi_n_2299);
  not csa_tree_add_190_195_groupi_drc_bufs53744(csa_tree_add_190_195_groupi_n_271 ,csa_tree_add_190_195_groupi_n_269);
  not csa_tree_add_190_195_groupi_drc_bufs53745(csa_tree_add_190_195_groupi_n_270 ,csa_tree_add_190_195_groupi_n_269);
  not csa_tree_add_190_195_groupi_drc_bufs53746(csa_tree_add_190_195_groupi_n_269 ,csa_tree_add_190_195_groupi_n_2198);
  not csa_tree_add_190_195_groupi_drc_bufs53749(csa_tree_add_190_195_groupi_n_268 ,csa_tree_add_190_195_groupi_n_267);
  not csa_tree_add_190_195_groupi_drc_bufs53750(csa_tree_add_190_195_groupi_n_267 ,csa_tree_add_190_195_groupi_n_2196);
  not csa_tree_add_190_195_groupi_drc_bufs53753(csa_tree_add_190_195_groupi_n_266 ,csa_tree_add_190_195_groupi_n_265);
  not csa_tree_add_190_195_groupi_drc_bufs53754(csa_tree_add_190_195_groupi_n_265 ,csa_tree_add_190_195_groupi_n_2097);
  not csa_tree_add_190_195_groupi_drc_bufs53757(csa_tree_add_190_195_groupi_n_264 ,csa_tree_add_190_195_groupi_n_263);
  not csa_tree_add_190_195_groupi_drc_bufs53758(csa_tree_add_190_195_groupi_n_263 ,csa_tree_add_190_195_groupi_n_2080);
  not csa_tree_add_190_195_groupi_drc_bufs53760(csa_tree_add_190_195_groupi_n_262 ,csa_tree_add_190_195_groupi_n_260);
  not csa_tree_add_190_195_groupi_drc_bufs53761(csa_tree_add_190_195_groupi_n_261 ,csa_tree_add_190_195_groupi_n_260);
  not csa_tree_add_190_195_groupi_drc_bufs53762(csa_tree_add_190_195_groupi_n_260 ,csa_tree_add_190_195_groupi_n_2192);
  not csa_tree_add_190_195_groupi_drc_bufs53765(csa_tree_add_190_195_groupi_n_259 ,csa_tree_add_190_195_groupi_n_258);
  not csa_tree_add_190_195_groupi_drc_bufs53766(csa_tree_add_190_195_groupi_n_258 ,csa_tree_add_190_195_groupi_n_2100);
  not csa_tree_add_190_195_groupi_drc_bufs53768(csa_tree_add_190_195_groupi_n_257 ,csa_tree_add_190_195_groupi_n_255);
  not csa_tree_add_190_195_groupi_drc_bufs53769(csa_tree_add_190_195_groupi_n_256 ,csa_tree_add_190_195_groupi_n_255);
  not csa_tree_add_190_195_groupi_drc_bufs53770(csa_tree_add_190_195_groupi_n_255 ,csa_tree_add_190_195_groupi_n_2222);
  not csa_tree_add_190_195_groupi_drc_bufs53773(csa_tree_add_190_195_groupi_n_254 ,csa_tree_add_190_195_groupi_n_2369);
  not csa_tree_add_190_195_groupi_drc_bufs53774(csa_tree_add_190_195_groupi_n_2369 ,csa_tree_add_190_195_groupi_n_2218);
  not csa_tree_add_190_195_groupi_drc_bufs53776(csa_tree_add_190_195_groupi_n_253 ,csa_tree_add_190_195_groupi_n_251);
  not csa_tree_add_190_195_groupi_drc_bufs53777(csa_tree_add_190_195_groupi_n_252 ,csa_tree_add_190_195_groupi_n_251);
  not csa_tree_add_190_195_groupi_drc_bufs53778(csa_tree_add_190_195_groupi_n_251 ,csa_tree_add_190_195_groupi_n_2124);
  not csa_tree_add_190_195_groupi_drc_bufs53781(csa_tree_add_190_195_groupi_n_250 ,csa_tree_add_190_195_groupi_n_249);
  not csa_tree_add_190_195_groupi_drc_bufs53782(csa_tree_add_190_195_groupi_n_249 ,csa_tree_add_190_195_groupi_n_2288);
  not csa_tree_add_190_195_groupi_drc_bufs53785(csa_tree_add_190_195_groupi_n_248 ,csa_tree_add_190_195_groupi_n_2336);
  not csa_tree_add_190_195_groupi_drc_bufs53786(csa_tree_add_190_195_groupi_n_2336 ,csa_tree_add_190_195_groupi_n_2081);
  not csa_tree_add_190_195_groupi_drc_bufs53789(csa_tree_add_190_195_groupi_n_247 ,csa_tree_add_190_195_groupi_n_2328);
  not csa_tree_add_190_195_groupi_drc_bufs53790(csa_tree_add_190_195_groupi_n_2328 ,csa_tree_add_190_195_groupi_n_2270);
  not csa_tree_add_190_195_groupi_drc_bufs53793(csa_tree_add_190_195_groupi_n_246 ,csa_tree_add_190_195_groupi_n_245);
  not csa_tree_add_190_195_groupi_drc_bufs53794(csa_tree_add_190_195_groupi_n_245 ,csa_tree_add_190_195_groupi_n_2260);
  not csa_tree_add_190_195_groupi_drc_bufs53796(csa_tree_add_190_195_groupi_n_244 ,csa_tree_add_190_195_groupi_n_242);
  not csa_tree_add_190_195_groupi_drc_bufs53797(csa_tree_add_190_195_groupi_n_243 ,csa_tree_add_190_195_groupi_n_242);
  not csa_tree_add_190_195_groupi_drc_bufs53798(csa_tree_add_190_195_groupi_n_242 ,csa_tree_add_190_195_groupi_n_2018);
  not csa_tree_add_190_195_groupi_drc_bufs53800(csa_tree_add_190_195_groupi_n_241 ,csa_tree_add_190_195_groupi_n_239);
  not csa_tree_add_190_195_groupi_drc_bufs53801(csa_tree_add_190_195_groupi_n_240 ,csa_tree_add_190_195_groupi_n_239);
  not csa_tree_add_190_195_groupi_drc_bufs53802(csa_tree_add_190_195_groupi_n_239 ,csa_tree_add_190_195_groupi_n_2198);
  not csa_tree_add_190_195_groupi_drc_bufs53804(csa_tree_add_190_195_groupi_n_238 ,csa_tree_add_190_195_groupi_n_236);
  not csa_tree_add_190_195_groupi_drc_bufs53805(csa_tree_add_190_195_groupi_n_237 ,csa_tree_add_190_195_groupi_n_236);
  not csa_tree_add_190_195_groupi_drc_bufs53806(csa_tree_add_190_195_groupi_n_236 ,csa_tree_add_190_195_groupi_n_2096);
  not csa_tree_add_190_195_groupi_drc_bufs53809(csa_tree_add_190_195_groupi_n_235 ,csa_tree_add_190_195_groupi_n_2367);
  not csa_tree_add_190_195_groupi_drc_bufs53810(csa_tree_add_190_195_groupi_n_2367 ,csa_tree_add_190_195_groupi_n_2187);
  not csa_tree_add_190_195_groupi_drc_bufs53812(csa_tree_add_190_195_groupi_n_234 ,csa_tree_add_190_195_groupi_n_232);
  not csa_tree_add_190_195_groupi_drc_bufs53813(csa_tree_add_190_195_groupi_n_233 ,csa_tree_add_190_195_groupi_n_232);
  not csa_tree_add_190_195_groupi_drc_bufs53814(csa_tree_add_190_195_groupi_n_232 ,csa_tree_add_190_195_groupi_n_2071);
  not csa_tree_add_190_195_groupi_drc_bufs53817(csa_tree_add_190_195_groupi_n_231 ,csa_tree_add_190_195_groupi_n_2368);
  not csa_tree_add_190_195_groupi_drc_bufs53818(csa_tree_add_190_195_groupi_n_2368 ,csa_tree_add_190_195_groupi_n_2287);
  not csa_tree_add_190_195_groupi_drc_bufs53821(csa_tree_add_190_195_groupi_n_230 ,csa_tree_add_190_195_groupi_n_2362);
  not csa_tree_add_190_195_groupi_drc_bufs53822(csa_tree_add_190_195_groupi_n_2362 ,csa_tree_add_190_195_groupi_n_2199);
  not csa_tree_add_190_195_groupi_drc_bufs53825(csa_tree_add_190_195_groupi_n_229 ,csa_tree_add_190_195_groupi_n_2340);
  not csa_tree_add_190_195_groupi_drc_bufs53826(csa_tree_add_190_195_groupi_n_2340 ,csa_tree_add_190_195_groupi_n_2075);
  not csa_tree_add_190_195_groupi_drc_bufs53829(csa_tree_add_190_195_groupi_n_228 ,csa_tree_add_190_195_groupi_n_2361);
  not csa_tree_add_190_195_groupi_drc_bufs53830(csa_tree_add_190_195_groupi_n_2361 ,csa_tree_add_190_195_groupi_n_2192);
  not csa_tree_add_190_195_groupi_drc_bufs53832(csa_tree_add_190_195_groupi_n_227 ,csa_tree_add_190_195_groupi_n_225);
  not csa_tree_add_190_195_groupi_drc_bufs53833(csa_tree_add_190_195_groupi_n_226 ,csa_tree_add_190_195_groupi_n_225);
  not csa_tree_add_190_195_groupi_drc_bufs53834(csa_tree_add_190_195_groupi_n_225 ,csa_tree_add_190_195_groupi_n_2025);
  not csa_tree_add_190_195_groupi_drc_bufs53837(csa_tree_add_190_195_groupi_n_224 ,csa_tree_add_190_195_groupi_n_2360);
  not csa_tree_add_190_195_groupi_drc_bufs53838(csa_tree_add_190_195_groupi_n_2360 ,csa_tree_add_190_195_groupi_n_2263);
  not csa_tree_add_190_195_groupi_drc_bufs53841(csa_tree_add_190_195_groupi_n_223 ,csa_tree_add_190_195_groupi_n_2365);
  not csa_tree_add_190_195_groupi_drc_bufs53842(csa_tree_add_190_195_groupi_n_2365 ,csa_tree_add_190_195_groupi_n_2189);
  not csa_tree_add_190_195_groupi_drc_bufs53844(csa_tree_add_190_195_groupi_n_222 ,csa_tree_add_190_195_groupi_n_220);
  not csa_tree_add_190_195_groupi_drc_bufs53845(csa_tree_add_190_195_groupi_n_221 ,csa_tree_add_190_195_groupi_n_220);
  not csa_tree_add_190_195_groupi_drc_bufs53846(csa_tree_add_190_195_groupi_n_220 ,csa_tree_add_190_195_groupi_n_2240);
  not csa_tree_add_190_195_groupi_drc_bufs53848(csa_tree_add_190_195_groupi_n_219 ,csa_tree_add_190_195_groupi_n_217);
  not csa_tree_add_190_195_groupi_drc_bufs53849(csa_tree_add_190_195_groupi_n_218 ,csa_tree_add_190_195_groupi_n_217);
  not csa_tree_add_190_195_groupi_drc_bufs53850(csa_tree_add_190_195_groupi_n_217 ,csa_tree_add_190_195_groupi_n_2242);
  not csa_tree_add_190_195_groupi_drc_bufs53852(csa_tree_add_190_195_groupi_n_216 ,csa_tree_add_190_195_groupi_n_214);
  not csa_tree_add_190_195_groupi_drc_bufs53853(csa_tree_add_190_195_groupi_n_215 ,csa_tree_add_190_195_groupi_n_214);
  not csa_tree_add_190_195_groupi_drc_bufs53854(csa_tree_add_190_195_groupi_n_214 ,csa_tree_add_190_195_groupi_n_2246);
  not csa_tree_add_190_195_groupi_drc_bufs53856(csa_tree_add_190_195_groupi_n_213 ,csa_tree_add_190_195_groupi_n_211);
  not csa_tree_add_190_195_groupi_drc_bufs53857(csa_tree_add_190_195_groupi_n_212 ,csa_tree_add_190_195_groupi_n_211);
  not csa_tree_add_190_195_groupi_drc_bufs53858(csa_tree_add_190_195_groupi_n_211 ,csa_tree_add_190_195_groupi_n_2224);
  not csa_tree_add_190_195_groupi_drc_bufs53860(csa_tree_add_190_195_groupi_n_210 ,csa_tree_add_190_195_groupi_n_208);
  not csa_tree_add_190_195_groupi_drc_bufs53861(csa_tree_add_190_195_groupi_n_209 ,csa_tree_add_190_195_groupi_n_208);
  not csa_tree_add_190_195_groupi_drc_bufs53862(csa_tree_add_190_195_groupi_n_208 ,csa_tree_add_190_195_groupi_n_2167);
  not csa_tree_add_190_195_groupi_drc_bufs53864(csa_tree_add_190_195_groupi_n_207 ,csa_tree_add_190_195_groupi_n_205);
  not csa_tree_add_190_195_groupi_drc_bufs53865(csa_tree_add_190_195_groupi_n_206 ,csa_tree_add_190_195_groupi_n_205);
  not csa_tree_add_190_195_groupi_drc_bufs53866(csa_tree_add_190_195_groupi_n_205 ,csa_tree_add_190_195_groupi_n_2164);
  not csa_tree_add_190_195_groupi_drc_bufs53868(csa_tree_add_190_195_groupi_n_204 ,csa_tree_add_190_195_groupi_n_203);
  not csa_tree_add_190_195_groupi_drc_bufs53870(csa_tree_add_190_195_groupi_n_203 ,csa_tree_add_190_195_groupi_n_2010);
  not csa_tree_add_190_195_groupi_drc_bufs53872(csa_tree_add_190_195_groupi_n_202 ,csa_tree_add_190_195_groupi_n_200);
  not csa_tree_add_190_195_groupi_drc_bufs53873(csa_tree_add_190_195_groupi_n_201 ,csa_tree_add_190_195_groupi_n_200);
  not csa_tree_add_190_195_groupi_drc_bufs53874(csa_tree_add_190_195_groupi_n_200 ,csa_tree_add_190_195_groupi_n_2145);
  not csa_tree_add_190_195_groupi_drc_bufs53876(csa_tree_add_190_195_groupi_n_199 ,csa_tree_add_190_195_groupi_n_197);
  not csa_tree_add_190_195_groupi_drc_bufs53877(csa_tree_add_190_195_groupi_n_198 ,csa_tree_add_190_195_groupi_n_197);
  not csa_tree_add_190_195_groupi_drc_bufs53878(csa_tree_add_190_195_groupi_n_197 ,csa_tree_add_190_195_groupi_n_2014);
  not csa_tree_add_190_195_groupi_drc_bufs53880(csa_tree_add_190_195_groupi_n_196 ,csa_tree_add_190_195_groupi_n_195);
  not csa_tree_add_190_195_groupi_drc_bufs53882(csa_tree_add_190_195_groupi_n_195 ,csa_tree_add_190_195_groupi_n_2021);
  not csa_tree_add_190_195_groupi_drc_bufs53884(csa_tree_add_190_195_groupi_n_194 ,csa_tree_add_190_195_groupi_n_192);
  not csa_tree_add_190_195_groupi_drc_bufs53885(csa_tree_add_190_195_groupi_n_193 ,csa_tree_add_190_195_groupi_n_192);
  not csa_tree_add_190_195_groupi_drc_bufs53886(csa_tree_add_190_195_groupi_n_192 ,csa_tree_add_190_195_groupi_n_2028);
  not csa_tree_add_190_195_groupi_drc_bufs53888(csa_tree_add_190_195_groupi_n_191 ,csa_tree_add_190_195_groupi_n_189);
  not csa_tree_add_190_195_groupi_drc_bufs53889(csa_tree_add_190_195_groupi_n_190 ,csa_tree_add_190_195_groupi_n_189);
  not csa_tree_add_190_195_groupi_drc_bufs53890(csa_tree_add_190_195_groupi_n_189 ,csa_tree_add_190_195_groupi_n_2248);
  not csa_tree_add_190_195_groupi_drc_bufs53892(csa_tree_add_190_195_groupi_n_188 ,csa_tree_add_190_195_groupi_n_187);
  not csa_tree_add_190_195_groupi_drc_bufs53894(csa_tree_add_190_195_groupi_n_187 ,csa_tree_add_190_195_groupi_n_2287);
  xor csa_tree_add_190_195_groupi_g2(csa_tree_add_190_195_groupi_n_186 ,csa_tree_add_190_195_groupi_n_12590 ,csa_tree_add_190_195_groupi_n_12542);
  xor csa_tree_add_190_195_groupi_g53896(csa_tree_add_190_195_groupi_n_185 ,csa_tree_add_190_195_groupi_n_12585 ,csa_tree_add_190_195_groupi_n_12562);
  xor csa_tree_add_190_195_groupi_g53897(csa_tree_add_190_195_groupi_n_184 ,csa_tree_add_190_195_groupi_n_12560 ,csa_tree_add_190_195_groupi_n_12503);
  xor csa_tree_add_190_195_groupi_g53898(csa_tree_add_190_195_groupi_n_183 ,csa_tree_add_190_195_groupi_n_12531 ,csa_tree_add_190_195_groupi_n_12525);
  xor csa_tree_add_190_195_groupi_g53899(csa_tree_add_190_195_groupi_n_182 ,csa_tree_add_190_195_groupi_n_12486 ,csa_tree_add_190_195_groupi_n_12500);
  xor csa_tree_add_190_195_groupi_g53900(out1[10] ,csa_tree_add_190_195_groupi_n_12490 ,csa_tree_add_190_195_groupi_n_12449);
  xor csa_tree_add_190_195_groupi_g53901(csa_tree_add_190_195_groupi_n_180 ,csa_tree_add_190_195_groupi_n_12454 ,csa_tree_add_190_195_groupi_n_12457);
  xor csa_tree_add_190_195_groupi_g53902(out1[9] ,csa_tree_add_190_195_groupi_n_12429 ,csa_tree_add_190_195_groupi_n_12416);
  xor csa_tree_add_190_195_groupi_g53903(out1[8] ,csa_tree_add_190_195_groupi_n_12353 ,csa_tree_add_190_195_groupi_n_12333);
  xor csa_tree_add_190_195_groupi_g53904(csa_tree_add_190_195_groupi_n_177 ,csa_tree_add_190_195_groupi_n_12300 ,csa_tree_add_190_195_groupi_n_12273);
  xor csa_tree_add_190_195_groupi_g53905(csa_tree_add_190_195_groupi_n_176 ,csa_tree_add_190_195_groupi_n_12219 ,csa_tree_add_190_195_groupi_n_12164);
  xor csa_tree_add_190_195_groupi_g53906(csa_tree_add_190_195_groupi_n_175 ,csa_tree_add_190_195_groupi_n_11998 ,csa_tree_add_190_195_groupi_n_12081);
  xor csa_tree_add_190_195_groupi_g53907(csa_tree_add_190_195_groupi_n_174 ,csa_tree_add_190_195_groupi_n_12006 ,csa_tree_add_190_195_groupi_n_12091);
  xor csa_tree_add_190_195_groupi_g53908(csa_tree_add_190_195_groupi_n_173 ,csa_tree_add_190_195_groupi_n_11827 ,csa_tree_add_190_195_groupi_n_11648);
  xor csa_tree_add_190_195_groupi_g53909(csa_tree_add_190_195_groupi_n_172 ,csa_tree_add_190_195_groupi_n_11824 ,csa_tree_add_190_195_groupi_n_11638);
  xor csa_tree_add_190_195_groupi_g53910(csa_tree_add_190_195_groupi_n_171 ,csa_tree_add_190_195_groupi_n_11450 ,csa_tree_add_190_195_groupi_n_11718);
  xor csa_tree_add_190_195_groupi_g53911(csa_tree_add_190_195_groupi_n_170 ,csa_tree_add_190_195_groupi_n_11596 ,csa_tree_add_190_195_groupi_n_11726);
  xor csa_tree_add_190_195_groupi_g53912(csa_tree_add_190_195_groupi_n_169 ,csa_tree_add_190_195_groupi_n_11477 ,csa_tree_add_190_195_groupi_n_11611);
  xor csa_tree_add_190_195_groupi_g53913(csa_tree_add_190_195_groupi_n_168 ,csa_tree_add_190_195_groupi_n_11473 ,csa_tree_add_190_195_groupi_n_11479);
  xor csa_tree_add_190_195_groupi_g53914(csa_tree_add_190_195_groupi_n_167 ,csa_tree_add_190_195_groupi_n_11471 ,csa_tree_add_190_195_groupi_n_11356);
  xor csa_tree_add_190_195_groupi_g53915(csa_tree_add_190_195_groupi_n_166 ,csa_tree_add_190_195_groupi_n_11247 ,csa_tree_add_190_195_groupi_n_11466);
  xor csa_tree_add_190_195_groupi_g53916(csa_tree_add_190_195_groupi_n_165 ,csa_tree_add_190_195_groupi_n_11073 ,csa_tree_add_190_195_groupi_n_11338);
  xor csa_tree_add_190_195_groupi_g53917(csa_tree_add_190_195_groupi_n_164 ,csa_tree_add_190_195_groupi_n_11042 ,csa_tree_add_190_195_groupi_n_11264);
  xor csa_tree_add_190_195_groupi_g53918(csa_tree_add_190_195_groupi_n_163 ,csa_tree_add_190_195_groupi_n_11182 ,csa_tree_add_190_195_groupi_n_11358);
  xor csa_tree_add_190_195_groupi_g53919(csa_tree_add_190_195_groupi_n_162 ,csa_tree_add_190_195_groupi_n_11175 ,csa_tree_add_190_195_groupi_n_11484);
  xor csa_tree_add_190_195_groupi_g53920(csa_tree_add_190_195_groupi_n_161 ,csa_tree_add_190_195_groupi_n_11171 ,csa_tree_add_190_195_groupi_n_11189);
  xor csa_tree_add_190_195_groupi_g53921(csa_tree_add_190_195_groupi_n_160 ,csa_tree_add_190_195_groupi_n_10962 ,csa_tree_add_190_195_groupi_n_11083);
  xor csa_tree_add_190_195_groupi_g53922(csa_tree_add_190_195_groupi_n_159 ,csa_tree_add_190_195_groupi_n_10983 ,csa_tree_add_190_195_groupi_n_11198);
  xor csa_tree_add_190_195_groupi_g53923(csa_tree_add_190_195_groupi_n_158 ,csa_tree_add_190_195_groupi_n_10978 ,csa_tree_add_190_195_groupi_n_11342);
  xor csa_tree_add_190_195_groupi_g53924(csa_tree_add_190_195_groupi_n_157 ,csa_tree_add_190_195_groupi_n_10975 ,csa_tree_add_190_195_groupi_n_11360);
  xor csa_tree_add_190_195_groupi_g53925(csa_tree_add_190_195_groupi_n_156 ,csa_tree_add_190_195_groupi_n_10766 ,csa_tree_add_190_195_groupi_n_10971);
  xor csa_tree_add_190_195_groupi_g53926(csa_tree_add_190_195_groupi_n_155 ,csa_tree_add_190_195_groupi_n_10196 ,csa_tree_add_190_195_groupi_n_10796);
  xor csa_tree_add_190_195_groupi_g53927(csa_tree_add_190_195_groupi_n_154 ,csa_tree_add_190_195_groupi_n_10458 ,csa_tree_add_190_195_groupi_n_10783);
  xor csa_tree_add_190_195_groupi_g53928(csa_tree_add_190_195_groupi_n_153 ,csa_tree_add_190_195_groupi_n_10778 ,csa_tree_add_190_195_groupi_n_11201);
  xor csa_tree_add_190_195_groupi_g53929(csa_tree_add_190_195_groupi_n_152 ,csa_tree_add_190_195_groupi_n_9952 ,csa_tree_add_190_195_groupi_n_10698);
  xor csa_tree_add_190_195_groupi_g53930(csa_tree_add_190_195_groupi_n_151 ,csa_tree_add_190_195_groupi_n_10696 ,csa_tree_add_190_195_groupi_n_10815);
  xor csa_tree_add_190_195_groupi_g53931(csa_tree_add_190_195_groupi_n_150 ,csa_tree_add_190_195_groupi_n_10577 ,csa_tree_add_190_195_groupi_n_10812);
  xor csa_tree_add_190_195_groupi_g53932(csa_tree_add_190_195_groupi_n_149 ,csa_tree_add_190_195_groupi_n_9913 ,csa_tree_add_190_195_groupi_n_10353);
  xor csa_tree_add_190_195_groupi_g53933(csa_tree_add_190_195_groupi_n_148 ,csa_tree_add_190_195_groupi_n_10352 ,csa_tree_add_190_195_groupi_n_10371);
  xor csa_tree_add_190_195_groupi_g53934(csa_tree_add_190_195_groupi_n_147 ,csa_tree_add_190_195_groupi_n_10052 ,csa_tree_add_190_195_groupi_n_10336);
  xor csa_tree_add_190_195_groupi_g53935(csa_tree_add_190_195_groupi_n_146 ,csa_tree_add_190_195_groupi_n_9628 ,csa_tree_add_190_195_groupi_n_10227);
  xor csa_tree_add_190_195_groupi_g53936(csa_tree_add_190_195_groupi_n_145 ,csa_tree_add_190_195_groupi_n_9922 ,csa_tree_add_190_195_groupi_n_10224);
  xor csa_tree_add_190_195_groupi_g53937(csa_tree_add_190_195_groupi_n_144 ,csa_tree_add_190_195_groupi_n_10085 ,csa_tree_add_190_195_groupi_n_10367);
  xor csa_tree_add_190_195_groupi_g53938(csa_tree_add_190_195_groupi_n_143 ,csa_tree_add_190_195_groupi_n_10084 ,csa_tree_add_190_195_groupi_n_8251);
  xor csa_tree_add_190_195_groupi_g53939(csa_tree_add_190_195_groupi_n_142 ,csa_tree_add_190_195_groupi_n_9317 ,csa_tree_add_190_195_groupi_n_10081);
  xor csa_tree_add_190_195_groupi_g53940(csa_tree_add_190_195_groupi_n_141 ,csa_tree_add_190_195_groupi_n_7350 ,csa_tree_add_190_195_groupi_n_10076);
  xor csa_tree_add_190_195_groupi_g53941(csa_tree_add_190_195_groupi_n_140 ,csa_tree_add_190_195_groupi_n_10075 ,csa_tree_add_190_195_groupi_n_10384);
  xor csa_tree_add_190_195_groupi_g53942(csa_tree_add_190_195_groupi_n_139 ,csa_tree_add_190_195_groupi_n_10073 ,csa_tree_add_190_195_groupi_n_10361);
  xor csa_tree_add_190_195_groupi_g53943(csa_tree_add_190_195_groupi_n_138 ,csa_tree_add_190_195_groupi_n_10072 ,csa_tree_add_190_195_groupi_n_9839);
  xor csa_tree_add_190_195_groupi_g53944(csa_tree_add_190_195_groupi_n_137 ,csa_tree_add_190_195_groupi_n_10070 ,csa_tree_add_190_195_groupi_n_10368);
  xor csa_tree_add_190_195_groupi_g53945(csa_tree_add_190_195_groupi_n_136 ,csa_tree_add_190_195_groupi_n_7162 ,csa_tree_add_190_195_groupi_n_9956);
  xor csa_tree_add_190_195_groupi_g53946(csa_tree_add_190_195_groupi_n_135 ,csa_tree_add_190_195_groupi_n_9797 ,csa_tree_add_190_195_groupi_n_10107);
  xor csa_tree_add_190_195_groupi_g53947(csa_tree_add_190_195_groupi_n_134 ,csa_tree_add_190_195_groupi_n_9779 ,csa_tree_add_190_195_groupi_n_10223);
  xor csa_tree_add_190_195_groupi_g53948(csa_tree_add_190_195_groupi_n_133 ,csa_tree_add_190_195_groupi_n_9007 ,csa_tree_add_190_195_groupi_n_9668);
  xor csa_tree_add_190_195_groupi_g53949(csa_tree_add_190_195_groupi_n_132 ,csa_tree_add_190_195_groupi_n_6909 ,csa_tree_add_190_195_groupi_n_9653);
  xor csa_tree_add_190_195_groupi_g53950(csa_tree_add_190_195_groupi_n_131 ,csa_tree_add_190_195_groupi_n_6956 ,csa_tree_add_190_195_groupi_n_9467);
  xor csa_tree_add_190_195_groupi_g53951(csa_tree_add_190_195_groupi_n_130 ,csa_tree_add_190_195_groupi_n_8820 ,csa_tree_add_190_195_groupi_n_9361);
  xor csa_tree_add_190_195_groupi_g53952(csa_tree_add_190_195_groupi_n_129 ,csa_tree_add_190_195_groupi_n_8614 ,csa_tree_add_190_195_groupi_n_9353);
  xor csa_tree_add_190_195_groupi_g53953(csa_tree_add_190_195_groupi_n_128 ,csa_tree_add_190_195_groupi_n_6955 ,csa_tree_add_190_195_groupi_n_9198);
  xor csa_tree_add_190_195_groupi_g53954(csa_tree_add_190_195_groupi_n_127 ,csa_tree_add_190_195_groupi_n_9197 ,csa_tree_add_190_195_groupi_n_9546);
  xor csa_tree_add_190_195_groupi_g53955(csa_tree_add_190_195_groupi_n_126 ,csa_tree_add_190_195_groupi_n_7368 ,csa_tree_add_190_195_groupi_n_9189);
  xor csa_tree_add_190_195_groupi_g53956(csa_tree_add_190_195_groupi_n_125 ,csa_tree_add_190_195_groupi_n_7338 ,csa_tree_add_190_195_groupi_n_9051);
  xor csa_tree_add_190_195_groupi_g53957(csa_tree_add_190_195_groupi_n_124 ,csa_tree_add_190_195_groupi_n_8653 ,csa_tree_add_190_195_groupi_n_9046);
  xor csa_tree_add_190_195_groupi_g53958(csa_tree_add_190_195_groupi_n_123 ,csa_tree_add_190_195_groupi_n_8685 ,csa_tree_add_190_195_groupi_n_8868);
  xor csa_tree_add_190_195_groupi_g53959(csa_tree_add_190_195_groupi_n_122 ,csa_tree_add_190_195_groupi_n_7629 ,csa_tree_add_190_195_groupi_n_8857);
  xor csa_tree_add_190_195_groupi_g53960(csa_tree_add_190_195_groupi_n_121 ,csa_tree_add_190_195_groupi_n_7981 ,csa_tree_add_190_195_groupi_n_8717);
  xor csa_tree_add_190_195_groupi_g53961(csa_tree_add_190_195_groupi_n_120 ,csa_tree_add_190_195_groupi_n_8716 ,csa_tree_add_190_195_groupi_n_6621);
  xor csa_tree_add_190_195_groupi_g53962(csa_tree_add_190_195_groupi_n_119 ,csa_tree_add_190_195_groupi_n_8534 ,csa_tree_add_190_195_groupi_n_8584);
  xor csa_tree_add_190_195_groupi_g53963(csa_tree_add_190_195_groupi_n_118 ,csa_tree_add_190_195_groupi_n_8373 ,csa_tree_add_190_195_groupi_n_8532);
  xor csa_tree_add_190_195_groupi_g53964(csa_tree_add_190_195_groupi_n_117 ,csa_tree_add_190_195_groupi_n_8510 ,csa_tree_add_190_195_groupi_n_8886);
  xor csa_tree_add_190_195_groupi_g53965(csa_tree_add_190_195_groupi_n_116 ,csa_tree_add_190_195_groupi_n_7993 ,csa_tree_add_190_195_groupi_n_8393);
  xor csa_tree_add_190_195_groupi_g53966(csa_tree_add_190_195_groupi_n_115 ,csa_tree_add_190_195_groupi_n_4789 ,csa_tree_add_190_195_groupi_n_8379);
  and csa_tree_add_190_195_groupi_g53967(csa_tree_add_190_195_groupi_n_114 ,csa_tree_add_190_195_groupi_n_5983 ,csa_tree_add_190_195_groupi_n_8234);
  xor csa_tree_add_190_195_groupi_g53968(csa_tree_add_190_195_groupi_n_113 ,csa_tree_add_190_195_groupi_n_7330 ,csa_tree_add_190_195_groupi_n_8225);
  xor csa_tree_add_190_195_groupi_g53969(csa_tree_add_190_195_groupi_n_112 ,csa_tree_add_190_195_groupi_n_8209 ,csa_tree_add_190_195_groupi_n_7941);
  xor csa_tree_add_190_195_groupi_g53970(csa_tree_add_190_195_groupi_n_111 ,csa_tree_add_190_195_groupi_n_8208 ,csa_tree_add_190_195_groupi_n_8553);
  xor csa_tree_add_190_195_groupi_g53971(csa_tree_add_190_195_groupi_n_110 ,csa_tree_add_190_195_groupi_n_8048 ,csa_tree_add_190_195_groupi_n_8911);
  xor csa_tree_add_190_195_groupi_g53972(csa_tree_add_190_195_groupi_n_109 ,csa_tree_add_190_195_groupi_n_8039 ,csa_tree_add_190_195_groupi_n_6703);
  xor csa_tree_add_190_195_groupi_g53973(csa_tree_add_190_195_groupi_n_108 ,csa_tree_add_190_195_groupi_n_7151 ,csa_tree_add_190_195_groupi_n_7854);
  xor csa_tree_add_190_195_groupi_g53974(csa_tree_add_190_195_groupi_n_107 ,csa_tree_add_190_195_groupi_n_7853 ,csa_tree_add_190_195_groupi_n_7063);
  xor csa_tree_add_190_195_groupi_g53975(csa_tree_add_190_195_groupi_n_106 ,csa_tree_add_190_195_groupi_n_4765 ,csa_tree_add_190_195_groupi_n_7431);
  xor csa_tree_add_190_195_groupi_g53976(csa_tree_add_190_195_groupi_n_105 ,csa_tree_add_190_195_groupi_n_7422 ,csa_tree_add_190_195_groupi_n_8271);
  xor csa_tree_add_190_195_groupi_g53977(csa_tree_add_190_195_groupi_n_104 ,csa_tree_add_190_195_groupi_n_7416 ,csa_tree_add_190_195_groupi_n_1678);
  xor csa_tree_add_190_195_groupi_g53978(csa_tree_add_190_195_groupi_n_103 ,csa_tree_add_190_195_groupi_n_7387 ,csa_tree_add_190_195_groupi_n_8267);
  xor csa_tree_add_190_195_groupi_g53979(csa_tree_add_190_195_groupi_n_102 ,csa_tree_add_190_195_groupi_n_6267 ,csa_tree_add_190_195_groupi_n_7223);
  xor csa_tree_add_190_195_groupi_g53980(csa_tree_add_190_195_groupi_n_101 ,csa_tree_add_190_195_groupi_n_4568 ,csa_tree_add_190_195_groupi_n_86);
  xor csa_tree_add_190_195_groupi_g53981(csa_tree_add_190_195_groupi_n_100 ,csa_tree_add_190_195_groupi_n_7003 ,csa_tree_add_190_195_groupi_n_1775);
  xor csa_tree_add_190_195_groupi_g53982(csa_tree_add_190_195_groupi_n_99 ,csa_tree_add_190_195_groupi_n_6919 ,csa_tree_add_190_195_groupi_n_8511);
  xor csa_tree_add_190_195_groupi_g53983(csa_tree_add_190_195_groupi_n_98 ,csa_tree_add_190_195_groupi_n_5031 ,csa_tree_add_190_195_groupi_n_6586);
  xor csa_tree_add_190_195_groupi_g53984(csa_tree_add_190_195_groupi_n_97 ,csa_tree_add_190_195_groupi_n_6579 ,csa_tree_add_190_195_groupi_n_70);
  and csa_tree_add_190_195_groupi_g53985(csa_tree_add_190_195_groupi_n_96 ,csa_tree_add_190_195_groupi_n_2398 ,csa_tree_add_190_195_groupi_n_5546);
  and csa_tree_add_190_195_groupi_g53986(csa_tree_add_190_195_groupi_n_95 ,csa_tree_add_190_195_groupi_n_2397 ,csa_tree_add_190_195_groupi_n_5541);
  and csa_tree_add_190_195_groupi_g53987(csa_tree_add_190_195_groupi_n_94 ,csa_tree_add_190_195_groupi_n_2403 ,csa_tree_add_190_195_groupi_n_5411);
  and csa_tree_add_190_195_groupi_g53988(csa_tree_add_190_195_groupi_n_93 ,csa_tree_add_190_195_groupi_n_2396 ,csa_tree_add_190_195_groupi_n_5322);
  and csa_tree_add_190_195_groupi_g53989(csa_tree_add_190_195_groupi_n_92 ,csa_tree_add_190_195_groupi_n_2399 ,csa_tree_add_190_195_groupi_n_5269);
  and csa_tree_add_190_195_groupi_g53990(csa_tree_add_190_195_groupi_n_91 ,csa_tree_add_190_195_groupi_n_2404 ,csa_tree_add_190_195_groupi_n_5252);
  and csa_tree_add_190_195_groupi_g53991(csa_tree_add_190_195_groupi_n_90 ,csa_tree_add_190_195_groupi_n_2401 ,csa_tree_add_190_195_groupi_n_5244);
  xor csa_tree_add_190_195_groupi_g53992(csa_tree_add_190_195_groupi_n_89 ,csa_tree_add_190_195_groupi_n_5173 ,csa_tree_add_190_195_groupi_n_6708);
  xor csa_tree_add_190_195_groupi_g53993(csa_tree_add_190_195_groupi_n_88 ,csa_tree_add_190_195_groupi_n_5159 ,csa_tree_add_190_195_groupi_n_3201);
  xor csa_tree_add_190_195_groupi_g53994(csa_tree_add_190_195_groupi_n_87 ,csa_tree_add_190_195_groupi_n_5131 ,csa_tree_add_190_195_groupi_n_5874);
  xor csa_tree_add_190_195_groupi_g53995(csa_tree_add_190_195_groupi_n_86 ,csa_tree_add_190_195_groupi_n_4832 ,csa_tree_add_190_195_groupi_n_6087);
  xor csa_tree_add_190_195_groupi_g53996(csa_tree_add_190_195_groupi_n_85 ,csa_tree_add_190_195_groupi_n_4814 ,csa_tree_add_190_195_groupi_n_3804);
  xor csa_tree_add_190_195_groupi_g53997(csa_tree_add_190_195_groupi_n_84 ,csa_tree_add_190_195_groupi_n_5986 ,csa_tree_add_190_195_groupi_n_3200);
  xor csa_tree_add_190_195_groupi_g53998(csa_tree_add_190_195_groupi_n_83 ,csa_tree_add_190_195_groupi_n_264 ,csa_tree_add_190_195_groupi_n_2388);
  xor csa_tree_add_190_195_groupi_g53999(csa_tree_add_190_195_groupi_n_82 ,csa_tree_add_190_195_groupi_n_1715 ,csa_tree_add_190_195_groupi_n_1542);
  xor csa_tree_add_190_195_groupi_g54000(csa_tree_add_190_195_groupi_n_81 ,csa_tree_add_190_195_groupi_n_4014 ,csa_tree_add_190_195_groupi_n_717);
  xor csa_tree_add_190_195_groupi_g54001(csa_tree_add_190_195_groupi_n_80 ,csa_tree_add_190_195_groupi_n_4051 ,csa_tree_add_190_195_groupi_n_578);
  xor csa_tree_add_190_195_groupi_g54002(csa_tree_add_190_195_groupi_n_79 ,csa_tree_add_190_195_groupi_n_5513 ,csa_tree_add_190_195_groupi_n_573);
  xor csa_tree_add_190_195_groupi_g54003(csa_tree_add_190_195_groupi_n_78 ,csa_tree_add_190_195_groupi_n_6038 ,csa_tree_add_190_195_groupi_n_571);
  xor csa_tree_add_190_195_groupi_g54004(csa_tree_add_190_195_groupi_n_77 ,csa_tree_add_190_195_groupi_n_3743 ,csa_tree_add_190_195_groupi_n_569);
  xor csa_tree_add_190_195_groupi_g54005(csa_tree_add_190_195_groupi_n_76 ,csa_tree_add_190_195_groupi_n_3980 ,csa_tree_add_190_195_groupi_n_567);
  xor csa_tree_add_190_195_groupi_g54006(csa_tree_add_190_195_groupi_n_75 ,csa_tree_add_190_195_groupi_n_4069 ,csa_tree_add_190_195_groupi_n_565);
  xor csa_tree_add_190_195_groupi_g54007(csa_tree_add_190_195_groupi_n_74 ,csa_tree_add_190_195_groupi_n_6066 ,csa_tree_add_190_195_groupi_n_557);
  xor csa_tree_add_190_195_groupi_g54008(csa_tree_add_190_195_groupi_n_73 ,csa_tree_add_190_195_groupi_n_6022 ,csa_tree_add_190_195_groupi_n_555);
  xor csa_tree_add_190_195_groupi_g54009(csa_tree_add_190_195_groupi_n_72 ,csa_tree_add_190_195_groupi_n_7919 ,csa_tree_add_190_195_groupi_n_553);
  xor csa_tree_add_190_195_groupi_g54010(csa_tree_add_190_195_groupi_n_71 ,csa_tree_add_190_195_groupi_n_4111 ,csa_tree_add_190_195_groupi_n_551);
  xor csa_tree_add_190_195_groupi_g54011(csa_tree_add_190_195_groupi_n_70 ,csa_tree_add_190_195_groupi_n_3914 ,csa_tree_add_190_195_groupi_n_534);
  xor csa_tree_add_190_195_groupi_g54012(csa_tree_add_190_195_groupi_n_69 ,csa_tree_add_190_195_groupi_n_514 ,csa_tree_add_190_195_groupi_n_532);
  and csa_tree_add_190_195_groupi_g54013(csa_tree_add_190_195_groupi_n_68 ,csa_tree_add_190_195_groupi_n_530 ,csa_tree_add_190_195_groupi_n_245);
  and csa_tree_add_190_195_groupi_g54014(csa_tree_add_190_195_groupi_n_67 ,csa_tree_add_190_195_groupi_n_525 ,csa_tree_add_190_195_groupi_n_460);
  xor csa_tree_add_190_195_groupi_g54015(csa_tree_add_190_195_groupi_n_66 ,csa_tree_add_190_195_groupi_n_3905 ,csa_tree_add_190_195_groupi_n_523);
  xor csa_tree_add_190_195_groupi_g54016(csa_tree_add_190_195_groupi_n_65 ,csa_tree_add_190_195_groupi_n_4130 ,csa_tree_add_190_195_groupi_n_515);
  xor csa_tree_add_190_195_groupi_g54017(csa_tree_add_190_195_groupi_n_64 ,csa_tree_add_190_195_groupi_n_4027 ,csa_tree_add_190_195_groupi_n_513);
  xor csa_tree_add_190_195_groupi_g54018(csa_tree_add_190_195_groupi_n_63 ,csa_tree_add_190_195_groupi_n_826 ,csa_tree_add_190_195_groupi_n_511);
  and csa_tree_add_190_195_groupi_g54019(csa_tree_add_190_195_groupi_n_62 ,csa_tree_add_190_195_groupi_n_509 ,csa_tree_add_190_195_groupi_n_249);
  xor csa_tree_add_190_195_groupi_g54020(csa_tree_add_190_195_groupi_n_61 ,csa_tree_add_190_195_groupi_n_82 ,csa_tree_add_190_195_groupi_n_507);
  xnor csa_tree_add_190_195_groupi_g54021(csa_tree_add_190_195_groupi_n_60 ,csa_tree_add_190_195_groupi_n_4847 ,csa_tree_add_190_195_groupi_n_505);
  xor csa_tree_add_190_195_groupi_g54022(csa_tree_add_190_195_groupi_n_59 ,csa_tree_add_190_195_groupi_n_3850 ,csa_tree_add_190_195_groupi_n_503);
  xor csa_tree_add_190_195_groupi_g54023(csa_tree_add_190_195_groupi_n_58 ,csa_tree_add_190_195_groupi_n_4122 ,csa_tree_add_190_195_groupi_n_492);
  xor csa_tree_add_190_195_groupi_g54024(csa_tree_add_190_195_groupi_n_57 ,csa_tree_add_190_195_groupi_n_5582 ,csa_tree_add_190_195_groupi_n_487);
  xor csa_tree_add_190_195_groupi_g54025(csa_tree_add_190_195_groupi_n_56 ,csa_tree_add_190_195_groupi_n_3791 ,csa_tree_add_190_195_groupi_n_476);
  xor csa_tree_add_190_195_groupi_g54026(csa_tree_add_190_195_groupi_n_55 ,csa_tree_add_190_195_groupi_n_3757 ,csa_tree_add_190_195_groupi_n_474);
  xor csa_tree_add_190_195_groupi_g54027(csa_tree_add_190_195_groupi_n_54 ,csa_tree_add_190_195_groupi_n_3880 ,csa_tree_add_190_195_groupi_n_462);
  xor csa_tree_add_190_195_groupi_g54028(csa_tree_add_190_195_groupi_n_53 ,csa_tree_add_190_195_groupi_n_3837 ,csa_tree_add_190_195_groupi_n_452);
  xor csa_tree_add_190_195_groupi_g54029(csa_tree_add_190_195_groupi_n_52 ,csa_tree_add_190_195_groupi_n_4091 ,csa_tree_add_190_195_groupi_n_450);
  and csa_tree_add_190_195_groupi_g54030(csa_tree_add_190_195_groupi_n_51 ,csa_tree_add_190_195_groupi_n_329 ,csa_tree_add_190_195_groupi_n_418);
  xor csa_tree_add_190_195_groupi_g54031(csa_tree_add_190_195_groupi_n_50 ,csa_tree_add_190_195_groupi_n_4060 ,csa_tree_add_190_195_groupi_n_413);
  xor csa_tree_add_190_195_groupi_g54032(csa_tree_add_190_195_groupi_n_49 ,csa_tree_add_190_195_groupi_n_40 ,csa_tree_add_190_195_groupi_n_408);
  xor csa_tree_add_190_195_groupi_g54033(csa_tree_add_190_195_groupi_n_48 ,csa_tree_add_190_195_groupi_n_3944 ,csa_tree_add_190_195_groupi_n_406);
  xor csa_tree_add_190_195_groupi_g54034(csa_tree_add_190_195_groupi_n_47 ,csa_tree_add_190_195_groupi_n_885 ,csa_tree_add_190_195_groupi_n_404);
  xor csa_tree_add_190_195_groupi_g54035(csa_tree_add_190_195_groupi_n_46 ,csa_tree_add_190_195_groupi_n_7031 ,csa_tree_add_190_195_groupi_n_402);
  xor csa_tree_add_190_195_groupi_g54036(csa_tree_add_190_195_groupi_n_45 ,csa_tree_add_190_195_groupi_n_235 ,csa_tree_add_190_195_groupi_n_400);
  xor csa_tree_add_190_195_groupi_g54037(csa_tree_add_190_195_groupi_n_44 ,csa_tree_add_190_195_groupi_n_621 ,csa_tree_add_190_195_groupi_n_395);
  xor csa_tree_add_190_195_groupi_g54038(csa_tree_add_190_195_groupi_n_43 ,csa_tree_add_190_195_groupi_n_6689 ,csa_tree_add_190_195_groupi_n_390);
  xor csa_tree_add_190_195_groupi_g54039(csa_tree_add_190_195_groupi_n_42 ,csa_tree_add_190_195_groupi_n_3938 ,csa_tree_add_190_195_groupi_n_388);
  xor csa_tree_add_190_195_groupi_g54040(csa_tree_add_190_195_groupi_n_41 ,csa_tree_add_190_195_groupi_n_4572 ,csa_tree_add_190_195_groupi_n_383);
  xor csa_tree_add_190_195_groupi_g54041(csa_tree_add_190_195_groupi_n_40 ,csa_tree_add_190_195_groupi_n_268 ,csa_tree_add_190_195_groupi_n_381);
  xor csa_tree_add_190_195_groupi_g54042(csa_tree_add_190_195_groupi_n_39 ,csa_tree_add_190_195_groupi_n_377 ,csa_tree_add_190_195_groupi_n_379);
  xor csa_tree_add_190_195_groupi_g54043(csa_tree_add_190_195_groupi_n_38 ,csa_tree_add_190_195_groupi_n_3824 ,csa_tree_add_190_195_groupi_n_374);
  xor csa_tree_add_190_195_groupi_g54044(csa_tree_add_190_195_groupi_n_37 ,csa_tree_add_190_195_groupi_n_3903 ,csa_tree_add_190_195_groupi_n_372);
  xor csa_tree_add_190_195_groupi_g54045(csa_tree_add_190_195_groupi_n_36 ,csa_tree_add_190_195_groupi_n_6589 ,csa_tree_add_190_195_groupi_n_367);
  xor csa_tree_add_190_195_groupi_g54046(csa_tree_add_190_195_groupi_n_35 ,csa_tree_add_190_195_groupi_n_5179 ,csa_tree_add_190_195_groupi_n_365);
  xor csa_tree_add_190_195_groupi_g54047(csa_tree_add_190_195_groupi_n_34 ,csa_tree_add_190_195_groupi_n_853 ,csa_tree_add_190_195_groupi_n_363);
  xor csa_tree_add_190_195_groupi_g54048(csa_tree_add_190_195_groupi_n_33 ,csa_tree_add_190_195_groupi_n_237 ,csa_tree_add_190_195_groupi_n_361);
  xor csa_tree_add_190_195_groupi_g54049(csa_tree_add_190_195_groupi_n_32 ,csa_tree_add_190_195_groupi_n_3802 ,csa_tree_add_190_195_groupi_n_359);
  xor csa_tree_add_190_195_groupi_g54050(csa_tree_add_190_195_groupi_n_31 ,csa_tree_add_190_195_groupi_n_4003 ,csa_tree_add_190_195_groupi_n_357);
  xor csa_tree_add_190_195_groupi_g54051(csa_tree_add_190_195_groupi_n_30 ,csa_tree_add_190_195_groupi_n_6029 ,csa_tree_add_190_195_groupi_n_352);
  xor csa_tree_add_190_195_groupi_g54052(csa_tree_add_190_195_groupi_n_29 ,csa_tree_add_190_195_groupi_n_4009 ,csa_tree_add_190_195_groupi_n_344);
  xor csa_tree_add_190_195_groupi_g54053(csa_tree_add_190_195_groupi_n_28 ,csa_tree_add_190_195_groupi_n_3764 ,csa_tree_add_190_195_groupi_n_339);
  xor csa_tree_add_190_195_groupi_g54054(csa_tree_add_190_195_groupi_n_27 ,csa_tree_add_190_195_groupi_n_4099 ,csa_tree_add_190_195_groupi_n_337);
  xor csa_tree_add_190_195_groupi_g54055(csa_tree_add_190_195_groupi_n_26 ,csa_tree_add_190_195_groupi_n_4078 ,csa_tree_add_190_195_groupi_n_335);
  xor csa_tree_add_190_195_groupi_g54056(csa_tree_add_190_195_groupi_n_25 ,csa_tree_add_190_195_groupi_n_8274 ,csa_tree_add_190_195_groupi_n_333);
  xor csa_tree_add_190_195_groupi_g54057(csa_tree_add_190_195_groupi_n_24 ,csa_tree_add_190_195_groupi_n_4021 ,csa_tree_add_190_195_groupi_n_331);
  xor csa_tree_add_190_195_groupi_g54058(csa_tree_add_190_195_groupi_n_23 ,csa_tree_add_190_195_groupi_n_5978 ,csa_tree_add_190_195_groupi_n_327);
  xor csa_tree_add_190_195_groupi_g54059(csa_tree_add_190_195_groupi_n_22 ,csa_tree_add_190_195_groupi_n_7201 ,csa_tree_add_190_195_groupi_n_322);
  xor csa_tree_add_190_195_groupi_g54060(csa_tree_add_190_195_groupi_n_21 ,csa_tree_add_190_195_groupi_n_6011 ,csa_tree_add_190_195_groupi_n_320);
  xor csa_tree_add_190_195_groupi_g54061(csa_tree_add_190_195_groupi_n_20 ,csa_tree_add_190_195_groupi_n_3970 ,csa_tree_add_190_195_groupi_n_318);
  xnor csa_tree_add_190_195_groupi_g54062(csa_tree_add_190_195_groupi_n_19 ,csa_tree_add_190_195_groupi_n_5602 ,csa_tree_add_190_195_groupi_n_316);
  xor csa_tree_add_190_195_groupi_g54063(csa_tree_add_190_195_groupi_n_18 ,csa_tree_add_190_195_groupi_n_3891 ,csa_tree_add_190_195_groupi_n_314);
  xor csa_tree_add_190_195_groupi_g54064(csa_tree_add_190_195_groupi_n_17 ,csa_tree_add_190_195_groupi_n_3844 ,csa_tree_add_190_195_groupi_n_306);
  xor csa_tree_add_190_195_groupi_g54065(csa_tree_add_190_195_groupi_n_16 ,csa_tree_add_190_195_groupi_n_3788 ,csa_tree_add_190_195_groupi_n_300);
  xor csa_tree_add_190_195_groupi_g54066(csa_tree_add_190_195_groupi_n_15 ,csa_tree_add_190_195_groupi_n_270 ,csa_tree_add_190_195_groupi_n_298);
  xor csa_tree_add_190_195_groupi_g54067(csa_tree_add_190_195_groupi_n_14 ,csa_tree_add_190_195_groupi_n_4097 ,csa_tree_add_190_195_groupi_n_296);
  xor csa_tree_add_190_195_groupi_g54068(csa_tree_add_190_195_groupi_n_13 ,csa_tree_add_190_195_groupi_n_7467 ,csa_tree_add_190_195_groupi_n_294);
  xor csa_tree_add_190_195_groupi_g54069(csa_tree_add_190_195_groupi_n_12 ,csa_tree_add_190_195_groupi_n_256 ,csa_tree_add_190_195_groupi_n_292);
  xor csa_tree_add_190_195_groupi_g54070(csa_tree_add_190_195_groupi_n_11 ,csa_tree_add_190_195_groupi_n_3760 ,csa_tree_add_190_195_groupi_n_290);
  xor csa_tree_add_190_195_groupi_g54071(csa_tree_add_190_195_groupi_n_10 ,csa_tree_add_190_195_groupi_n_4049 ,csa_tree_add_190_195_groupi_n_288);
  xor csa_tree_add_190_195_groupi_g54072(csa_tree_add_190_195_groupi_n_9 ,csa_tree_add_190_195_groupi_n_3762 ,csa_tree_add_190_195_groupi_n_280);
  xor csa_tree_add_190_195_groupi_g54073(csa_tree_add_190_195_groupi_n_8 ,csa_tree_add_190_195_groupi_n_4110 ,csa_tree_add_190_195_groupi_n_278);
  xor csa_tree_add_190_195_groupi_g54074(csa_tree_add_190_195_groupi_n_7 ,csa_tree_add_190_195_groupi_n_4028 ,csa_tree_add_190_195_groupi_n_267);
  xor csa_tree_add_190_195_groupi_g54075(csa_tree_add_190_195_groupi_n_6 ,csa_tree_add_190_195_groupi_n_3972 ,csa_tree_add_190_195_groupi_n_265);
  xor csa_tree_add_190_195_groupi_g54076(csa_tree_add_190_195_groupi_n_5 ,csa_tree_add_190_195_groupi_n_4573 ,csa_tree_add_190_195_groupi_n_263);
  xor csa_tree_add_190_195_groupi_g54077(csa_tree_add_190_195_groupi_n_4 ,csa_tree_add_190_195_groupi_n_6611 ,csa_tree_add_190_195_groupi_n_258);
  xor csa_tree_add_190_195_groupi_g54078(csa_tree_add_190_195_groupi_n_3 ,csa_tree_add_190_195_groupi_n_203 ,csa_tree_add_190_195_groupi_n_1624);
  xor csa_tree_add_190_195_groupi_g54079(csa_tree_add_190_195_groupi_n_2 ,csa_tree_add_190_195_groupi_n_195 ,csa_tree_add_190_195_groupi_n_1643);
  xor csa_tree_add_190_195_groupi_g54080(csa_tree_add_190_195_groupi_n_1 ,csa_tree_add_190_195_groupi_n_187 ,csa_tree_add_190_195_groupi_n_1214);
  xor csa_tree_add_190_195_groupi_g54081(csa_tree_add_190_195_groupi_n_0 ,csa_tree_add_190_195_groupi_n_2338 ,in56[4]);
  xnor inc_add_191_21_g197(out2[16] ,inc_add_191_21_n_66 ,out1[28]);
  xnor inc_add_191_21_g198(out2[15] ,inc_add_191_21_n_62 ,out1[27]);
  or inc_add_191_21_g199(inc_add_191_21_n_66 ,inc_add_191_21_n_7 ,inc_add_191_21_n_61);
  xnor inc_add_191_21_g200(out2[14] ,inc_add_191_21_n_57 ,out1[26]);
  xnor inc_add_191_21_g201(out2[13] ,inc_add_191_21_n_56 ,out1[25]);
  xnor inc_add_191_21_g202(out2[11] ,inc_add_191_21_n_55 ,out1[23]);
  or inc_add_191_21_g203(inc_add_191_21_n_62 ,inc_add_191_21_n_7 ,inc_add_191_21_n_57);
  or inc_add_191_21_g204(inc_add_191_21_n_61 ,inc_add_191_21_n_16 ,inc_add_191_21_n_57);
  xor inc_add_191_21_g205(out2[12] ,inc_add_191_21_n_51 ,out1[24]);
  xor inc_add_191_21_g206(out2[10] ,inc_add_191_21_n_49 ,out1[22]);
  xnor inc_add_191_21_g207(out2[9] ,inc_add_191_21_n_53 ,out1[21]);
  or inc_add_191_21_g208(inc_add_191_21_n_57 ,inc_add_191_21_n_26 ,inc_add_191_21_n_52);
  or inc_add_191_21_g209(inc_add_191_21_n_56 ,inc_add_191_21_n_8 ,inc_add_191_21_n_52);
  or inc_add_191_21_g210(inc_add_191_21_n_55 ,inc_add_191_21_n_17 ,inc_add_191_21_n_50);
  xnor inc_add_191_21_g211(out2[8] ,inc_add_191_21_n_47 ,out1[20]);
  or inc_add_191_21_g212(inc_add_191_21_n_53 ,inc_add_191_21_n_14 ,inc_add_191_21_n_47);
  not inc_add_191_21_g213(inc_add_191_21_n_52 ,inc_add_191_21_n_51);
  and inc_add_191_21_g214(inc_add_191_21_n_51 ,inc_add_191_21_n_34 ,inc_add_191_21_n_46);
  not inc_add_191_21_g215(inc_add_191_21_n_50 ,inc_add_191_21_n_49);
  and inc_add_191_21_g216(inc_add_191_21_n_49 ,inc_add_191_21_n_24 ,inc_add_191_21_n_46);
  xnor inc_add_191_21_g217(out2[7] ,inc_add_191_21_n_43 ,out1[19]);
  not inc_add_191_21_g218(inc_add_191_21_n_46 ,inc_add_191_21_n_47);
  or inc_add_191_21_g219(inc_add_191_21_n_47 ,inc_add_191_21_n_2 ,inc_add_191_21_n_42);
  xnor inc_add_191_21_g220(out2[6] ,inc_add_191_21_n_38 ,inc_add_191_21_n_15);
  xnor inc_add_191_21_g221(out2[5] ,inc_add_191_21_n_40 ,out1[17]);
  or inc_add_191_21_g222(inc_add_191_21_n_43 ,inc_add_191_21_n_2 ,inc_add_191_21_n_39);
  or inc_add_191_21_g223(inc_add_191_21_n_42 ,inc_add_191_21_n_13 ,inc_add_191_21_n_39);
  xnor inc_add_191_21_g224(out2[4] ,inc_add_191_21_n_37 ,inc_add_191_21_n_5);
  or inc_add_191_21_g225(inc_add_191_21_n_40 ,inc_add_191_21_n_6 ,inc_add_191_21_n_37);
  not inc_add_191_21_g226(inc_add_191_21_n_39 ,inc_add_191_21_n_38);
  and inc_add_191_21_g227(inc_add_191_21_n_38 ,inc_add_191_21_n_22 ,inc_add_191_21_n_36);
  not inc_add_191_21_g229(inc_add_191_21_n_37 ,inc_add_191_21_n_36);
  and inc_add_191_21_g230(inc_add_191_21_n_36 ,out1[15] ,inc_add_191_21_n_33);
  xnor inc_add_191_21_g231(out2[2] ,inc_add_191_21_n_29 ,out1[14]);
  nor inc_add_191_21_g232(inc_add_191_21_n_34 ,inc_add_191_21_n_17 ,inc_add_191_21_n_28);
  and inc_add_191_21_g234(inc_add_191_21_n_33 ,out1[14] ,inc_add_191_21_n_30);
  nor inc_add_191_21_g235(inc_add_191_21_n_32 ,inc_add_191_21_n_30 ,inc_add_191_21_n_31);
  nor inc_add_191_21_g236(inc_add_191_21_n_31 ,out1[13] ,inc_add_191_21_n_21);
  not inc_add_191_21_g237(inc_add_191_21_n_30 ,inc_add_191_21_n_29);
  or inc_add_191_21_g238(inc_add_191_21_n_29 ,inc_add_191_21_n_19 ,inc_add_191_21_n_20);
  or inc_add_191_21_g239(inc_add_191_21_n_28 ,inc_add_191_21_n_12 ,inc_add_191_21_n_23);
  nor inc_add_191_21_g240(inc_add_191_21_n_27 ,inc_add_191_21_n_21 ,inc_add_191_21_n_25);
  or inc_add_191_21_g241(inc_add_191_21_n_26 ,inc_add_191_21_n_9 ,inc_add_191_21_n_8);
  nor inc_add_191_21_g242(inc_add_191_21_n_25 ,out1[12] ,in62);
  not inc_add_191_21_g243(inc_add_191_21_n_24 ,inc_add_191_21_n_23);
  or inc_add_191_21_g244(inc_add_191_21_n_23 ,inc_add_191_21_n_10 ,inc_add_191_21_n_14);
  and inc_add_191_21_g245(inc_add_191_21_n_22 ,out1[17] ,inc_add_191_21_n_5);
  not inc_add_191_21_g246(inc_add_191_21_n_21 ,inc_add_191_21_n_20);
  or inc_add_191_21_g247(inc_add_191_21_n_20 ,inc_add_191_21_n_18 ,inc_add_191_21_n_11);
  not inc_add_191_21_g248(inc_add_191_21_n_19 ,out1[13]);
  not inc_add_191_21_g249(inc_add_191_21_n_18 ,out1[12]);
  not inc_add_191_21_g250(inc_add_191_21_n_17 ,out1[22]);
  not inc_add_191_21_g251(inc_add_191_21_n_16 ,out1[27]);
  not inc_add_191_21_g252(inc_add_191_21_n_15 ,out1[18]);
  not inc_add_191_21_g253(inc_add_191_21_n_14 ,out1[20]);
  not inc_add_191_21_g254(inc_add_191_21_n_13 ,out1[19]);
  not inc_add_191_21_g255(inc_add_191_21_n_12 ,out1[23]);
  not inc_add_191_21_g256(inc_add_191_21_n_11 ,in62);
  not inc_add_191_21_g258(inc_add_191_21_n_10 ,out1[21]);
  not inc_add_191_21_g259(inc_add_191_21_n_9 ,out1[25]);
  not inc_add_191_21_g260(inc_add_191_21_n_8 ,out1[24]);
  not inc_add_191_21_g261(inc_add_191_21_n_7 ,out1[26]);
  not inc_add_191_21_drc_bufs(inc_add_191_21_n_5 ,inc_add_191_21_n_6);
  not inc_add_191_21_drc_bufs263(inc_add_191_21_n_6 ,out1[16]);
  buf inc_add_191_21_drc_bufs265(out2[1] ,inc_add_191_21_n_32);
  buf inc_add_191_21_drc_bufs266(out2[0] ,inc_add_191_21_n_27);
  not inc_add_191_21_drc_bufs268(inc_add_191_21_n_2 ,inc_add_191_21_n_1);
  not inc_add_191_21_drc_bufs269(inc_add_191_21_n_1 ,inc_add_191_21_n_15);
  xor inc_add_191_21_g2(out2[3] ,inc_add_191_21_n_33 ,out1[15]);
  buf g54082(csa_tree_add_190_195_groupi_n_4834 ,csa_tree_add_190_195_groupi_n_4171);
endmodule
