module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, out1, out2);
  input [12:0] in1, in35, in39;
  input [6:0] in2, in21, in26, in42;
  input in3, in5, in6, in7, in8, in9, in10, in11, in12, in14, in15, in16, in17, in18, in19, in20, in22, in27, in30, in31, in32, in33, in34, in36, in37, in38, in40;
  input [3:0] in4, in23;
  input [5:0] in13;
  input [8:0] in24, in28, in29;
  input [2:0] in25, in41;
  output [12:0] out1, out2;
  wire [12:0] in1, in35, in39;
  wire [6:0] in2, in21, in26, in42;
  wire in3, in5, in6, in7, in8, in9, in10, in11, in12, in14, in15, in16, in17, in18, in19, in20, in22, in27, in30, in31, in32, in33, in34, in36, in37, in38, in40;
  wire [3:0] in4, in23;
  wire [5:0] in13;
  wire [8:0] in24, in28, in29;
  wire [2:0] in25, in41;
  wire [12:0] out1, out2;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__139, w__140, w__141, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__157, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__171, w__172, w__173, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__665, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__680;
  wire w__681, w__682, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__697, w__698, w__699, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__714, w__715, w__716, w__717, w__718, w__719, w__720;
  wire w__721, w__722, w__723, w__724, w__725, w__726, w__727, w__728;
  wire w__729, w__730, w__731, w__732, w__733, w__734, w__735, w__736;
  wire w__737, w__738, w__739, w__740, w__741, w__742, w__743, w__744;
  wire w__745, w__746, w__747, w__748, w__749, w__750, w__751, w__752;
  wire w__753, w__754, w__755, w__756, w__757, w__758, w__759, w__760;
  wire w__761, w__762, w__763, w__764, w__765, w__766, w__767, w__768;
  wire w__769, w__770, w__771, w__772, w__773, w__774, w__775, w__776;
  wire w__777, w__778, w__779, w__780, w__781, w__782, w__783, w__784;
  wire w__785, w__786, w__787, w__788, w__789, w__790, w__791, w__792;
  wire w__793, w__794, w__795, w__796, w__797, w__798, w__799, w__800;
  wire w__801, w__802, w__803, w__804, w__805, w__806, w__807, w__808;
  wire w__809, w__810, w__811, w__812, w__813, w__814, w__815, w__816;
  wire w__817, w__818, w__819, w__820, w__821, w__822, w__823, w__824;
  wire w__825, w__826, w__827, w__828, w__829, w__830, w__831, w__832;
  wire w__833, w__834, w__835, w__836, w__837, w__838, w__839, w__840;
  wire w__841, w__842, w__843, w__844, w__845, w__846, w__847, w__848;
  wire w__849, w__850, w__851, w__852, w__853, w__854, w__855, w__856;
  wire w__857, w__858, w__859, w__860, w__861, w__862, w__863, w__864;
  wire w__865, w__866, w__867, w__868, w__869, w__870, w__871, w__872;
  wire w__873, w__874, w__875, w__876, w__877, w__878, w__879, w__880;
  wire w__881, w__882, w__883, w__884, w__885, w__886, w__887, w__888;
  wire w__889, w__890, w__891, w__892, w__893, w__894, w__895, w__896;
  wire w__897, w__898, w__899, w__900, w__901, w__902, w__903, w__904;
  wire w__905, w__906, w__907, w__908, w__909, w__910, w__911, w__912;
  wire w__913, w__914, w__915, w__916, w__917, w__918, w__919, w__920;
  wire w__921, w__922, w__923, w__924, w__925, w__926, w__927, w__928;
  wire w__929, w__930, w__931, w__932, w__933, w__934, w__935, w__936;
  wire w__937, w__938, w__939, w__940, w__941, w__942, w__943, w__944;
  wire w__945, w__946, w__947, w__948, w__949, w__950, w__951, w__952;
  wire w__953, w__954, w__955, w__956, w__957, w__958, w__959, w__960;
  wire w__961, w__962, w__963, w__964, w__965, w__966, w__967, w__968;
  wire w__969, w__970, w__971, w__972, w__973, w__974, w__975, w__976;
  wire w__977, w__978, w__979, w__980, w__981, w__982, w__983, w__984;
  wire w__985, w__986, w__987, w__988, w__989, w__990, w__991, w__992;
  wire w__993, w__994, w__995, w__996, w__997, w__998, w__999, w__1000;
  wire w__1001, w__1002, w__1003, w__1004, w__1005, w__1006, w__1007, w__1008;
  wire w__1009, w__1010, w__1011, w__1012, w__1013, w__1014, w__1015, w__1016;
  wire w__1017, w__1018, w__1019, w__1020, w__1021, w__1022, w__1023, w__1024;
  wire w__1025, w__1026, w__1027, w__1028, w__1029, w__1030, w__1031, w__1032;
  wire w__1033, w__1034, w__1035, w__1036, w__1037, w__1038, w__1039, w__1040;
  wire w__1041, w__1042, w__1043, w__1044, w__1045, w__1046, w__1047, w__1048;
  wire w__1049, w__1050, w__1051, w__1052, w__1053, w__1054, w__1055, w__1056;
  wire w__1057, w__1058, w__1059, w__1060, w__1061, w__1062, w__1063, w__1064;
  wire w__1065, w__1066, w__1067, w__1068, w__1069, w__1070, w__1071, w__1072;
  wire w__1073, w__1074, w__1075, w__1076, w__1077, w__1078, w__1079, w__1080;
  wire w__1081, w__1082, w__1083, w__1084, w__1085, w__1086, w__1087, w__1088;
  wire w__1089, w__1090, w__1091, w__1092, w__1093, w__1094, w__1095, w__1096;
  wire w__1097, w__1098, w__1099, w__1100, w__1101, w__1102, w__1103, w__1104;
  wire w__1105, w__1106, w__1107, w__1108, w__1109, w__1110, w__1111, w__1112;
  wire w__1113, w__1114, w__1115, w__1116, w__1117, w__1118, w__1119, w__1120;
  wire w__1121, w__1122, w__1123, w__1124, w__1125, w__1126, w__1127, w__1128;
  wire w__1129, w__1130, w__1131, w__1132, w__1133, w__1134, w__1135, w__1136;
  wire w__1137, w__1138, w__1139, w__1140, w__1141, w__1142, w__1143, w__1144;
  wire w__1145, w__1146, w__1147, w__1148, w__1149, w__1150, w__1151, w__1152;
  wire w__1153, w__1154, w__1155, w__1156, w__1157, w__1158, w__1159, w__1160;
  wire w__1161, w__1162, w__1163, w__1164, w__1165, w__1166, w__1167, w__1168;
  wire w__1169, w__1170, w__1171, w__1172, w__1173, w__1174, w__1175, w__1176;
  wire w__1177, w__1178, w__1179, w__1180, w__1181, w__1182, w__1183, w__1184;
  wire w__1185, w__1186, w__1187, w__1188, w__1189, w__1190, w__1191, w__1192;
  wire w__1193, w__1194, w__1195, w__1196, w__1197, w__1198, w__1199, w__1200;
  wire w__1201, w__1202, w__1203, w__1204, w__1205, w__1206, w__1207, w__1208;
  wire w__1209, w__1210, w__1211, w__1212, w__1213, w__1214, w__1215, w__1216;
  wire w__1217, w__1218, w__1219, w__1220, w__1221, w__1222, w__1223, w__1224;
  wire w__1225, w__1226, w__1227, w__1228, w__1229, w__1230, w__1231, w__1232;
  wire w__1233, w__1234, w__1235, w__1236, w__1237, w__1238, w__1239, w__1240;
  wire w__1241, w__1242, w__1243, w__1244, w__1245, w__1246, w__1247, w__1248;
  wire w__1249, w__1250, w__1251, w__1252, w__1253, w__1254, w__1255, w__1256;
  wire w__1257, w__1258, w__1259, w__1260, w__1261, w__1262, w__1263, w__1264;
  wire w__1265, w__1266, w__1267, w__1268, w__1269, w__1270, w__1271, w__1272;
  wire w__1273, w__1274, w__1275, w__1276, w__1277, w__1278, w__1279, w__1280;
  wire w__1281, w__1282, w__1283, w__1284, w__1285, w__1286, w__1287, w__1288;
  wire w__1289, w__1290, w__1291, w__1292, w__1293, w__1294, w__1295, w__1296;
  wire w__1297, w__1298, w__1299, w__1300, w__1301, w__1302, w__1303, w__1304;
  wire w__1305, w__1306, w__1307, w__1308, w__1309, w__1310, w__1311, w__1312;
  wire w__1313, w__1314, w__1315, w__1316, w__1317, w__1318, w__1319, w__1320;
  wire w__1321, w__1322, w__1323, w__1324, w__1325, w__1326, w__1327, w__1328;
  wire w__1329, w__1330, w__1331, w__1332, w__1333, w__1334, w__1335, w__1336;
  wire w__1337, w__1338, w__1339, w__1340, w__1341, w__1342, w__1343, w__1344;
  wire w__1345, w__1346, w__1347, w__1348, w__1349, w__1350, w__1351, w__1352;
  wire w__1353, w__1354, w__1355, w__1356, w__1357, w__1358, w__1359, w__1360;
  wire w__1361, w__1362, w__1363, w__1364, w__1365, w__1366, w__1367, w__1368;
  wire w__1369, w__1370, w__1371, w__1372, w__1373, w__1374, w__1375, w__1376;
  wire w__1377, w__1378, w__1379, w__1380, w__1381, w__1382, w__1383, w__1384;
  wire w__1385, w__1386, w__1387, w__1388, w__1389, w__1390, w__1391, w__1392;
  wire w__1393, w__1394, w__1395, w__1396, w__1397, w__1398, w__1399, w__1400;
  wire w__1401, w__1402, w__1403, w__1404, w__1405, w__1406, w__1407, w__1408;
  wire w__1409, w__1410, w__1411, w__1412, w__1413, w__1414, w__1415, w__1416;
  wire w__1417, w__1418, w__1419, w__1420, w__1421, w__1422, w__1423, w__1424;
  wire w__1425, w__1426, w__1427, w__1428, w__1429, w__1430, w__1431, w__1432;
  wire w__1433, w__1434, w__1435, w__1436, w__1437, w__1438, w__1439, w__1440;
  wire w__1441, w__1442, w__1443, w__1444, w__1445, w__1446, w__1447, w__1448;
  wire w__1449, w__1450, w__1451, w__1452, w__1453, w__1454, w__1455, w__1456;
  wire w__1457, w__1458, w__1459, w__1460, w__1461, w__1462, w__1463, w__1464;
  wire w__1465, w__1466, w__1467, w__1468, w__1469, w__1470, w__1471, w__1472;
  wire w__1473, w__1474, w__1475, w__1476, w__1477, w__1478, w__1479, w__1480;
  wire w__1481, w__1482, w__1483, w__1484, w__1485, w__1486, w__1487, w__1488;
  wire w__1489, w__1490, w__1491, w__1492, w__1493, w__1494, w__1495, w__1496;
  wire w__1497, w__1498, w__1499, w__1500, w__1501, w__1502, w__1503, w__1504;
  wire w__1505, w__1506, w__1507, w__1508, w__1509, w__1510, w__1511, w__1512;
  wire w__1513, w__1514, w__1515, w__1516, w__1517, w__1518, w__1519, w__1520;
  wire w__1521, w__1522, w__1523, w__1524, w__1525, w__1526, w__1527, w__1528;
  wire w__1529, w__1530, w__1531, w__1532, w__1533, w__1534, w__1535, w__1536;
  wire w__1537, w__1538, w__1539, w__1540, w__1541, w__1542, w__1543, w__1544;
  wire w__1545, w__1546, w__1547, w__1548, w__1549, w__1550, w__1551, w__1552;
  wire w__1553, w__1554, w__1555, w__1556, w__1557, w__1558, w__1559, w__1560;
  wire w__1561, w__1562, w__1563, w__1564, w__1565, w__1566, w__1567, w__1568;
  wire w__1569, w__1570, w__1571, w__1572, w__1573, w__1574, w__1575, w__1576;
  wire w__1577, w__1578, w__1579, w__1580, w__1581, w__1582, w__1583, w__1584;
  wire w__1585, w__1586, w__1587, w__1588, w__1589, w__1590, w__1591, w__1592;
  wire w__1593, w__1594, w__1595, w__1596, w__1597, w__1598, w__1599, w__1600;
  wire w__1601, w__1602, w__1603, w__1604, w__1605, w__1606, w__1607, w__1608;
  wire w__1609, w__1610, w__1611, w__1612, w__1613, w__1614, w__1615, w__1616;
  wire w__1617, w__1618, w__1619, w__1620, w__1621, w__1622, w__1623, w__1624;
  wire w__1625, w__1626, w__1627, w__1628, w__1629, w__1630, w__1631, w__1632;
  wire w__1633, w__1634, w__1635, w__1636, w__1637, w__1638, w__1639, w__1640;
  wire w__1641, w__1642, w__1643, w__1644, w__1645, w__1646, w__1647, w__1648;
  wire w__1649, w__1650, w__1651, w__1652, w__1653, w__1654, w__1655, w__1656;
  wire w__1657, w__1658, w__1659, w__1660, w__1661, w__1662, w__1663, w__1664;
  wire w__1665, w__1666, w__1667, w__1668, w__1669, w__1670, w__1671, w__1672;
  wire w__1673, w__1674, w__1675, w__1676, w__1677, w__1678, w__1679, w__1680;
  wire w__1681, w__1682, w__1683, w__1684, w__1685, w__1686, w__1687, w__1688;
  wire w__1689, w__1690, w__1691, w__1692, w__1693, w__1694, w__1695, w__1696;
  wire w__1697, w__1698, w__1699, w__1700, w__1701, w__1702, w__1703, w__1704;
  wire w__1705, w__1706, w__1707, w__1708, w__1709, w__1710, w__1711, w__1712;
  wire w__1713, w__1714, w__1715, w__1716, w__1717, w__1718, w__1719, w__1720;
  wire w__1721, w__1722, w__1723, w__1724, w__1725, w__1726, w__1727, w__1728;
  wire w__1729, w__1730, w__1731, w__1732, w__1733, w__1734, w__1735, w__1736;
  wire w__1737, w__1738, w__1739, w__1740, w__1741, w__1742, w__1743, w__1744;
  wire w__1745, w__1746, w__1747, w__1748, w__1749, w__1750, w__1751, w__1752;
  wire w__1753, w__1754, w__1755, w__1756, w__1757, w__1758, w__1759, w__1760;
  wire w__1761, w__1762, w__1763, w__1764, w__1765, w__1766, w__1767, w__1768;
  wire w__1769, w__1770, w__1771, w__1772, w__1773, w__1774, w__1775, w__1776;
  wire w__1777, w__1778, w__1779, w__1780, w__1781, w__1782, w__1783, w__1784;
  wire w__1785, w__1786, w__1787, w__1788, w__1789, w__1790, w__1791, w__1792;
  wire w__1793, w__1794, w__1795, w__1796, w__1797, w__1798, w__1799, w__1800;
  wire w__1801, w__1802, w__1803, w__1804, w__1805, w__1806, w__1807, w__1808;
  wire w__1809, w__1810, w__1811, w__1812, w__1813, w__1814, w__1815, w__1816;
  wire w__1817, w__1818, w__1819, w__1820, w__1821, w__1822, w__1823, w__1824;
  wire w__1825, w__1826, w__1827, w__1828, w__1829, w__1830, w__1831, w__1832;
  wire w__1833, w__1834, w__1835, w__1836, w__1837, w__1838, w__1839, w__1840;
  wire w__1841, w__1842, w__1843, w__1844, w__1845, w__1846, w__1847, w__1848;
  wire w__1849, w__1850, w__1851, w__1852, w__1853, w__1854, w__1855, w__1856;
  wire w__1857, w__1858, w__1859, w__1860, w__1861, w__1862, w__1863, w__1864;
  wire w__1865, w__1866, w__1867, w__1868, w__1869, w__1870, w__1871, w__1872;
  wire w__1873, w__1874, w__1875, w__1876, w__1877, w__1878, w__1879, w__1880;
  wire w__1881, w__1882, w__1883, w__1884, w__1885, w__1886, w__1887, w__1888;
  wire w__1889, w__1890, w__1891, w__1892, w__1893, w__1894, w__1895, w__1896;
  wire w__1897, w__1898, w__1899, w__1900, w__1901, w__1902, w__1903, w__1904;
  wire w__1905, w__1906, w__1907, w__1908, w__1909, w__1910, w__1911, w__1912;
  wire w__1913, w__1914, w__1915, w__1916, w__1917, w__1918, w__1919, w__1920;
  wire w__1921, w__1922, w__1923, w__1924, w__1925, w__1926, w__1927, w__1928;
  wire w__1929, w__1930, w__1931, w__1932, w__1933, w__1934, w__1935, w__1936;
  wire w__1937, w__1938, w__1939, w__1940, w__1941, w__1942, w__1943, w__1944;
  wire w__1945, w__1946, w__1947, w__1948, w__1949, w__1950, w__1951, w__1952;
  wire w__1953, w__1954, w__1955, w__1956, w__1957, w__1958, w__1959, w__1960;
  wire w__1961, w__1962, w__1963, w__1964, w__1965, w__1966, w__1967, w__1968;
  wire w__1969, w__1970, w__1971, w__1972, w__1973, w__1974, w__1975, w__1976;
  wire w__1977, w__1978, w__1979, w__1980, w__1981, w__1982, w__1983, w__1984;
  wire w__1985, w__1986, w__1987, w__1988, w__1989, w__1990, w__1991, w__1992;
  wire w__1993, w__1994, w__1995, w__1996, w__1997, w__1998, w__1999, w__2000;
  wire w__2001, w__2002, w__2003, w__2004, w__2005, w__2006, w__2007, w__2008;
  wire w__2009, w__2010, w__2011, w__2012, w__2013, w__2014, w__2015, w__2016;
  wire w__2017, w__2018, w__2019, w__2020, w__2021, w__2022, w__2023, w__2024;
  wire w__2025, w__2026, w__2027, w__2028, w__2029, w__2030, w__2031, w__2032;
  wire w__2033, w__2034, w__2035, w__2036, w__2037, w__2038, w__2039, w__2040;
  wire w__2041, w__2042, w__2043, w__2044, w__2045, w__2046, w__2047, w__2048;
  wire w__2049, w__2050, w__2051, w__2052, w__2053, w__2054, w__2055, w__2056;
  wire w__2057, w__2058, w__2059, w__2060, w__2061, w__2062, w__2063, w__2064;
  wire w__2065, w__2066, w__2067, w__2068, w__2069, w__2070, w__2071, w__2072;
  wire w__2073, w__2074, w__2075, w__2076, w__2077, w__2078, w__2079, w__2080;
  wire w__2081, w__2082, w__2083, w__2084, w__2085, w__2086, w__2087, w__2088;
  wire w__2089, w__2090, w__2091, w__2092, w__2093, w__2094, w__2095, w__2096;
  wire w__2097, w__2098, w__2099, w__2100, w__2101, w__2102, w__2103, w__2104;
  wire w__2105, w__2106, w__2107, w__2108, w__2109, w__2110, w__2111, w__2112;
  wire w__2113, w__2114, w__2115, w__2116, w__2117, w__2118, w__2119, w__2120;
  wire w__2121, w__2122, w__2123, w__2124, w__2125, w__2126, w__2127, w__2128;
  wire w__2129, w__2130, w__2131, w__2132, w__2133, w__2134, w__2135, w__2136;
  wire w__2137, w__2138, w__2139, w__2140, w__2141, w__2142, w__2143, w__2144;
  wire w__2145, w__2146, w__2147, w__2148, w__2149, w__2150, w__2151, w__2152;
  wire w__2153, w__2154, w__2155, w__2156, w__2157, w__2158, w__2159, w__2160;
  wire w__2161, w__2162, w__2163, w__2164, w__2165, w__2166, w__2167, w__2168;
  wire w__2169, w__2170, w__2171, w__2172, w__2173, w__2174, w__2175, w__2176;
  wire w__2177, w__2178, w__2179, w__2180, w__2181, w__2182, w__2183, w__2184;
  wire w__2185, w__2186, w__2187, w__2188, w__2189, w__2190, w__2191, w__2192;
  wire w__2193, w__2194, w__2195, w__2196, w__2197, w__2198, w__2199, w__2200;
  wire w__2201, w__2202, w__2203, w__2204, w__2205, w__2206, w__2207, w__2208;
  wire w__2209, w__2210, w__2211, w__2212, w__2213, w__2214, w__2215, w__2216;
  wire w__2217, w__2218, w__2219, w__2220, w__2221, w__2222, w__2223, w__2224;
  wire w__2225, w__2226, w__2227, w__2228, w__2229, w__2230, w__2231, w__2232;
  wire w__2233, w__2234, w__2235, w__2236, w__2237, w__2238, w__2239, w__2240;
  wire w__2241, w__2242, w__2243, w__2244, w__2245, w__2246, w__2247, w__2248;
  wire w__2249, w__2250, w__2251, w__2252, w__2253, w__2254, w__2255, w__2256;
  wire w__2257, w__2258, w__2259, w__2260, w__2261, w__2262, w__2263, w__2264;
  wire w__2265, w__2266, w__2267, w__2268, w__2269, w__2270, w__2271, w__2272;
  wire w__2273, w__2274, w__2275, w__2276, w__2277, w__2278, w__2279, w__2280;
  wire w__2281, w__2282, w__2283, w__2284, w__2285, w__2286, w__2287, w__2288;
  wire w__2289, w__2290, w__2291, w__2292, w__2293, w__2294, w__2295, w__2296;
  wire w__2297, w__2298, w__2299, w__2300, w__2301, w__2302, w__2303, w__2304;
  wire w__2305, w__2306, w__2307, w__2308, w__2309, w__2310, w__2311, w__2312;
  wire w__2313, w__2314, w__2315, w__2316, w__2317, w__2318, w__2319, w__2320;
  wire w__2321, w__2322, w__2323, w__2324, w__2325, w__2326, w__2327, w__2328;
  wire w__2329, w__2330, w__2331, w__2332, w__2333, w__2334, w__2335, w__2336;
  wire w__2337, w__2338, w__2339, w__2340, w__2341, w__2342, w__2343, w__2344;
  wire w__2345, w__2346, w__2347, w__2348, w__2349, w__2350, w__2351, w__2352;
  wire w__2353, w__2354, w__2355, w__2356, w__2357, w__2358, w__2359, w__2360;
  wire w__2361, w__2362, w__2363, w__2364, w__2365, w__2366, w__2367, w__2368;
  wire w__2369, w__2370, w__2371, w__2372, w__2373, w__2374, w__2375, w__2376;
  wire w__2377, w__2378, w__2379, w__2380, w__2381, w__2382, w__2383, w__2384;
  wire w__2385, w__2386, w__2387, w__2388, w__2389, w__2390, w__2391, w__2392;
  wire w__2393, w__2394, w__2395, w__2396, w__2397, w__2398, w__2399, w__2400;
  wire w__2401, w__2402, w__2403, w__2404, w__2405, w__2406, w__2407, w__2408;
  wire w__2409, w__2410, w__2411, w__2412, w__2413, w__2414, w__2415, w__2416;
  wire w__2417, w__2418, w__2419, w__2420, w__2421, w__2422, w__2423, w__2424;
  wire w__2425, w__2426, w__2427, w__2428, w__2429, w__2430, w__2431, w__2432;
  wire w__2433, w__2434, w__2435, w__2436, w__2437, w__2438, w__2439, w__2440;
  wire w__2441, w__2442, w__2443, w__2444, w__2445, w__2446, w__2447, w__2448;
  wire w__2449, w__2450, w__2451, w__2452, w__2453, w__2454, w__2455, w__2456;
  wire w__2457, w__2458, w__2459, w__2460, w__2461, w__2462, w__2463, w__2464;
  wire w__2465, w__2466, w__2467, w__2468, w__2469, w__2470, w__2471, w__2472;
  wire w__2473, w__2474, w__2475, w__2476, w__2477, w__2478, w__2479, w__2480;
  wire w__2481, w__2482, w__2483, w__2484, w__2485, w__2486, w__2487, w__2488;
  wire w__2489, w__2490, w__2491, w__2492, w__2493, w__2494, w__2495, w__2496;
  wire w__2497, w__2498, w__2499, w__2500, w__2501, w__2502, w__2503, w__2504;
  wire w__2505, w__2506, w__2507, w__2508, w__2509, w__2510, w__2511, w__2512;
  wire w__2513, w__2514, w__2515, w__2516, w__2517, w__2518, w__2519, w__2520;
  wire w__2521, w__2522, w__2523, w__2524, w__2525, w__2526, w__2527, w__2528;
  wire w__2529, w__2530, w__2531, w__2532, w__2533, w__2534, w__2535, w__2536;
  wire w__2537, w__2538, w__2539, w__2540, w__2541, w__2542, w__2543, w__2544;
  wire w__2545, w__2546, w__2547, w__2548, w__2549, w__2550, w__2551, w__2552;
  wire w__2553, w__2554, w__2555, w__2556, w__2557, w__2558, w__2559, w__2560;
  wire w__2561, w__2562, w__2563, w__2564, w__2565, w__2566, w__2567, w__2568;
  wire w__2569, w__2570, w__2571, w__2572, w__2573, w__2574, w__2575, w__2576;
  wire w__2577, w__2578, w__2579, w__2580, w__2581, w__2582, w__2583, w__2584;
  wire w__2585, w__2586, w__2587, w__2588, w__2589, w__2590, w__2591, w__2592;
  wire w__2593, w__2594, w__2595, w__2596, w__2597, w__2598, w__2599, w__2600;
  wire w__2601, w__2602, w__2603, w__2604, w__2605, w__2606, w__2607, w__2608;
  wire w__2609, w__2610, w__2611, w__2612, w__2613, w__2614, w__2615, w__2616;
  wire w__2617, w__2618, w__2619, w__2620, w__2621, w__2622, w__2623, w__2624;
  wire w__2625, w__2626, w__2627, w__2628, w__2629, w__2630, w__2631, w__2632;
  wire w__2633, w__2634, w__2635, w__2636, w__2637, w__2638, w__2639, w__2640;
  wire w__2641, w__2642, w__2643, w__2644, w__2645, w__2646, w__2647, w__2648;
  wire w__2649, w__2650, w__2651, w__2652, w__2653, w__2654, w__2655, w__2656;
  wire w__2657, w__2658, w__2659, w__2660, w__2661, w__2662, w__2663, w__2664;
  wire w__2665, w__2666, w__2667, w__2668, w__2669, w__2670, w__2671, w__2672;
  wire w__2673, w__2674, w__2675, w__2676, w__2677, w__2678, w__2679, w__2680;
  wire w__2681, w__2682, w__2683, w__2684, w__2685, w__2686, w__2687, w__2688;
  wire w__2689, w__2690, w__2691, w__2692, w__2693, w__2694, w__2695, w__2696;
  wire w__2697, w__2698, w__2699, w__2700, w__2701, w__2702, w__2703, w__2704;
  wire w__2705, w__2706, w__2707, w__2708, w__2709, w__2710, w__2711, w__2712;
  wire w__2713, w__2714, w__2715, w__2716, w__2717, w__2718, w__2719, w__2720;
  wire w__2721, w__2722, w__2723, w__2724, w__2725, w__2726, w__2727, w__2728;
  wire w__2729, w__2730, w__2731, w__2732, w__2733, w__2734, w__2735, w__2736;
  wire w__2737, w__2738, w__2739, w__2740, w__2741, w__2742, w__2743, w__2744;
  wire w__2745, w__2746, w__2747, w__2748, w__2749, w__2750, w__2751, w__2752;
  wire w__2753, w__2754, w__2755, w__2756, w__2757, w__2758, w__2759, w__2760;
  wire w__2761, w__2762, w__2763, w__2764, w__2765, w__2766, w__2767, w__2768;
  wire w__2769, w__2770, w__2771, w__2772, w__2773, w__2774, w__2775, w__2776;
  wire w__2777, w__2778, w__2779, w__2780, w__2781, w__2782, w__2783, w__2784;
  wire w__2785, w__2786, w__2787, w__2788, w__2789, w__2790, w__2791, w__2792;
  wire w__2793, w__2794, w__2795, w__2796, w__2797, w__2798, w__2799, w__2800;
  wire w__2801, w__2802, w__2803, w__2804, w__2805, w__2806, w__2807, w__2808;
  wire w__2809, w__2810, w__2811, w__2812, w__2813, w__2814, w__2815, w__2816;
  wire w__2817, w__2818, w__2819, w__2820, w__2821, w__2822, w__2823, w__2824;
  wire w__2825, w__2826, w__2827, w__2828, w__2829, w__2830, w__2831, w__2832;
  wire w__2833, w__2834, w__2835, w__2836, w__2837, w__2838, w__2839, w__2840;
  wire w__2841, w__2842, w__2843, w__2844, w__2845, w__2846, w__2847, w__2848;
  wire w__2849, w__2850, w__2851, w__2852, w__2853, w__2854, w__2855, w__2856;
  wire w__2857, w__2858, w__2859, w__2860, w__2861, w__2862, w__2863, w__2864;
  wire w__2865, w__2866, w__2867, w__2868, w__2869, w__2870, w__2871, w__2872;
  wire w__2873, w__2874, w__2875, w__2876, w__2877, w__2878, w__2879, w__2880;
  wire w__2881, w__2882, w__2883, w__2884, w__2885, w__2886, w__2887, w__2888;
  wire w__2889, w__2890, w__2891, w__2892, w__2893, w__2894, w__2895, w__2896;
  wire w__2897, w__2898, w__2899, w__2900, w__2901, w__2902, w__2903, w__2904;
  wire w__2905, w__2906, w__2907, w__2908, w__2909, w__2910, w__2911, w__2912;
  wire w__2913, w__2914, w__2915, w__2916, w__2917, w__2918, w__2919, w__2920;
  wire w__2921, w__2922, w__2923, w__2924, w__2925, w__2926, w__2927, w__2928;
  wire w__2929, w__2930, w__2931, w__2932, w__2933, w__2934, w__2935, w__2936;
  wire w__2937, w__2938, w__2939, w__2940, w__2941, w__2942, w__2943, w__2944;
  wire w__2945, w__2946, w__2947, w__2948, w__2949, w__2950, w__2951, w__2952;
  wire w__2953, w__2954, w__2955, w__2956, w__2957, w__2958, w__2959, w__2960;
  wire w__2961, w__2962, w__2963, w__2964, w__2965, w__2966, w__2967, w__2968;
  wire w__2969, w__2970, w__2971, w__2972, w__2973, w__2974, w__2975, w__2976;
  wire w__2977, w__2978, w__2979, w__2980, w__2981, w__2982, w__2983, w__2984;
  wire w__2985, w__2986, w__2987, w__2988, w__2989, w__2990, w__2991, w__2992;
  wire w__2993, w__2994, w__2995, w__2996, w__2997, w__2998, w__2999, w__3000;
  wire w__3001, w__3002, w__3003, w__3004, w__3005, w__3006, w__3007, w__3008;
  wire w__3009, w__3010, w__3011, w__3012, w__3013, w__3014, w__3015, w__3016;
  wire w__3017, w__3018, w__3019, w__3020, w__3021, w__3022, w__3023, w__3024;
  wire w__3025, w__3026, w__3027, w__3028, w__3029, w__3030, w__3031, w__3032;
  wire w__3033, w__3034, w__3035, w__3036, w__3037, w__3038, w__3039, w__3040;
  wire w__3041, w__3042, w__3043, w__3044, w__3045, w__3046, w__3047, w__3048;
  wire w__3049, w__3050, w__3051, w__3052, w__3053, w__3054, w__3055, w__3056;
  wire w__3057, w__3058, w__3059, w__3060, w__3061, w__3062, w__3063, w__3064;
  wire w__3065, w__3066, w__3067, w__3068, w__3069, w__3070, w__3071, w__3072;
  wire w__3073, w__3074, w__3075, w__3076, w__3077, w__3078, w__3079, w__3080;
  wire w__3081, w__3082, w__3083, w__3084, w__3085, w__3086, w__3087, w__3088;
  wire w__3089, w__3090, w__3091, w__3092, w__3093, w__3094, w__3095, w__3096;
  wire w__3097, w__3098, w__3099, w__3100, w__3101, w__3102, w__3103, w__3104;
  wire w__3105, w__3106, w__3107, w__3108, w__3109, w__3110, w__3111, w__3112;
  wire w__3113, w__3114, w__3115, w__3116, w__3117, w__3118, w__3119, w__3120;
  wire w__3121, w__3122, w__3123, w__3124, w__3125, w__3126, w__3127, w__3128;
  wire w__3129, w__3130, w__3131, w__3132, w__3133, w__3134;
  not g__1(w__2081 ,in31);
  not g__2(w__2080 ,in9);
  xor g__3(w__2079 ,in2[6] ,in3);
  xor g__4(w__2078 ,in2[4] ,in3);
  xor g__5(w__2077 ,in2[2] ,in3);
  xor g__6(w__2076 ,in2[0] ,in3);
  xor g__7(w__2075 ,in2[5] ,in3);
  xor g__8(w__2074 ,in2[1] ,in3);
  xor g__9(w__2073 ,in2[3] ,in3);
  buf g__10(w__2397 ,w__2079);
  buf g__11(w__2394 ,w__2073);
  buf g__12(w__2392 ,w__2074);
  buf g__13(w__2396 ,w__2075);
  buf g__14(w__2391 ,w__2076);
  buf g__15(w__2393 ,w__2077);
  buf g__16(w__2395 ,w__2078);
  or g__17(w__2212 ,w__1835 ,w__2067);
  or g__18(w__2217 ,w__1880 ,w__2072);
  or g__19(w__2216 ,w__1878 ,w__2071);
  or g__20(w__2215 ,w__1877 ,w__2070);
  or g__21(w__2214 ,w__1876 ,w__2069);
  or g__22(w__2213 ,w__1836 ,w__2068);
  or g__23(w__2110 ,w__2059 ,w__2038);
  or g__24(w__2205 ,w__1826 ,w__2060);
  or g__25(w__2210 ,w__1833 ,w__2065);
  or g__26(w__2209 ,w__1832 ,w__2064);
  or g__27(w__2208 ,w__1831 ,w__2063);
  or g__28(w__2207 ,w__1829 ,w__2062);
  or g__29(w__2206 ,w__2061 ,w__2028);
  or g__30(w__2211 ,w__1834 ,w__2066);
  or g__31(w__2118 ,w__2048 ,w__2045);
  or g__32(w__2109 ,w__2058 ,w__2057);
  or g__33(w__2115 ,w__2055 ,w__2054);
  or g__34(w__2114 ,w__2047 ,w__2044);
  or g__35(w__2072 ,w__1705 ,w__2053);
  or g__36(w__2120 ,w__2049 ,w__2040);
  or g__37(w__2071 ,w__1725 ,w__2051);
  or g__38(w__2070 ,w__1723 ,w__2046);
  or g__39(w__2113 ,w__2039 ,w__2037);
  or g__40(w__2069 ,w__1722 ,w__2043);
  or g__41(w__2068 ,w__1980 ,w__2042);
  or g__42(w__2067 ,w__1976 ,w__2041);
  or g__43(w__2066 ,w__1972 ,w__2019);
  or g__44(w__2065 ,w__1968 ,w__2036);
  or g__45(w__2064 ,w__1965 ,w__2034);
  or g__46(w__2112 ,w__2033 ,w__2031);
  or g__47(w__2063 ,w__1963 ,w__2032);
  or g__48(w__2121 ,w__2052 ,w__2050);
  or g__49(w__2062 ,w__1961 ,w__2030);
  or g__50(w__2117 ,w__2035 ,w__2027);
  or g__51(w__2111 ,w__2026 ,w__2024);
  or g__52(w__2061 ,w__1702 ,w__2029);
  or g__53(w__2060 ,w__1954 ,w__2025);
  or g__54(w__2119 ,w__2023 ,w__2056);
  or g__55(w__2116 ,w__2022 ,w__2021);
  or g__56(w__2059 ,w__1733 ,w__2020);
  or g__57(w__2058 ,w__1948 ,w__1998);
  or g__58(w__2057 ,w__1990 ,w__2135);
  or g__59(w__2056 ,w__1991 ,w__2018);
  or g__60(w__2055 ,w__1947 ,w__1989);
  or g__61(w__2054 ,w__2016 ,w__2141);
  or g__62(w__2053 ,w__1946 ,w__2015);
  or g__63(w__2052 ,w__1926 ,w__1995);
  or g__64(w__2051 ,w__1945 ,w__2014);
  or g__65(w__2050 ,w__1974 ,w__2147);
  or g__66(w__2049 ,w__1939 ,w__1964);
  or g__67(w__2048 ,w__1941 ,w__2009);
  or g__68(w__2047 ,w__1943 ,w__2012);
  or g__69(w__2046 ,w__1944 ,w__2013);
  or g__70(w__2045 ,w__1979 ,w__2144);
  or g__71(w__2044 ,w__1982 ,w__1988);
  or g__72(w__2043 ,w__1942 ,w__2011);
  or g__73(w__2042 ,w__2010 ,w__1978);
  or g__74(w__2041 ,w__2007 ,w__1975);
  or g__75(w__2040 ,w__2008 ,w__1985);
  or g__76(w__2039 ,w__1937 ,w__1971);
  or g__77(w__2038 ,w__1419 ,w__1981);
  or g__78(w__2037 ,w__2005 ,w__2139);
  or g__79(w__2036 ,w__2004 ,w__1966);
  or g__80(w__2035 ,w__1919 ,w__2000);
  or g__81(w__2034 ,w__2003 ,w__1983);
  or g__82(w__2033 ,w__1950 ,w__2002);
  or g__83(w__2032 ,w__2001 ,w__1962);
  or g__84(w__2031 ,w__1960 ,w__1987);
  or g__85(w__2030 ,w__1999 ,w__1958);
  or g__86(w__2029 ,w__2017 ,w__1956);
  or g__87(w__2028 ,w__1871 ,w__1955);
  or g__88(w__2027 ,w__1957 ,w__2143);
  or g__89(w__2026 ,w__1927 ,w__1967);
  or g__90(w__2025 ,w__1997 ,w__1959);
  or g__91(w__2136 ,w__1419 ,w__1969);
  or g__92(w__2024 ,w__1996 ,w__1986);
  or g__93(w__2023 ,w__1924 ,w__1993);
  or g__94(w__2022 ,w__1925 ,w__1973);
  or g__95(w__2021 ,w__1992 ,w__1984);
  or g__96(w__2020 ,w__1994 ,w__1977);
  or g__97(w__2019 ,w__2006 ,w__1970);
  and g__98(w__2017 ,w__2304 ,w__1599);
  and g__99(w__2016 ,w__2276 ,w__1596);
  and g__100(w__2015 ,w__2315 ,w__1429);
  and g__101(w__2014 ,w__2314 ,w__1522);
  and g__102(w__2013 ,w__2313 ,w__1445);
  and g__103(w__2012 ,w__2275 ,w__1441);
  and g__104(w__2011 ,w__2312 ,w__1521);
  and g__105(w__2010 ,w__2311 ,w__1483);
  and g__106(w__2009 ,w__2279 ,w__1546);
  and g__107(w__2008 ,w__2281 ,w__1443);
  and g__108(w__2007 ,w__2310 ,w__1483);
  and g__109(w__2006 ,w__2309 ,w__1429);
  and g__110(w__2005 ,w__2274 ,w__1545);
  and g__111(w__2004 ,w__2308 ,w__1445);
  and g__112(w__2003 ,w__2307 ,w__1598);
  and g__113(w__2002 ,w__2273 ,w__1455);
  and g__114(w__2001 ,w__2306 ,w__1521);
  and g__115(w__2000 ,w__2278 ,w__1455);
  and g__116(w__1999 ,w__2305 ,w__1482);
  and g__117(w__1998 ,w__2270 ,w__1441);
  and g__118(w__1997 ,w__2303 ,w__1522);
  and g__119(w__1996 ,w__2272 ,w__1443);
  and g__120(w__1995 ,w__2282 ,w__1595);
  and g__121(w__1994 ,w__2271 ,w__1545);
  and g__122(w__1993 ,w__2280 ,w__1454);
  and g__123(w__1992 ,w__2277 ,w__1546);
  and g__124(w__1991 ,w__2313 ,w__1590);
  and g__125(w__2198 ,in42[0] ,w__1552);
  and g__126(w__1990 ,w__2303 ,w__1439);
  and g__127(w__2199 ,in42[1] ,w__1549);
  and g__128(w__1989 ,w__2309 ,w__1543);
  and g__129(w__2200 ,in42[2] ,w__1551);
  and g__130(w__2204 ,in42[6] ,w__1537);
  and g__131(w__2203 ,in42[5] ,w__1536);
  and g__132(w__2202 ,in42[4] ,w__1552);
  and g__133(w__2201 ,in42[3] ,w__1551);
  or g__134(w__2141 ,w__1837 ,w__1930);
  or g__135(w__2135 ,w__1882 ,w__1922);
  or g__136(w__2018 ,w__1881 ,w__1921);
  and g__137(w__1983 ,in28[4] ,w__1524);
  and g__138(w__1982 ,w__2308 ,w__1427);
  or g__139(w__1981 ,w__1910 ,w__1949);
  or g__140(w__1980 ,w__1856 ,w__1940);
  and g__141(w__1979 ,w__2312 ,w__1542);
  and g__142(w__1978 ,in28[8] ,w__1525);
  and g__143(w__1977 ,w__2304 ,w__1452);
  or g__144(w__1976 ,w__1854 ,w__1938);
  and g__145(w__1975 ,in28[7] ,w__1525);
  and g__146(w__1974 ,w__2315 ,w__1452);
  and g__147(w__1973 ,w__2310 ,w__1439);
  or g__148(w__1972 ,w__1853 ,w__1936);
  and g__149(w__1971 ,w__2307 ,w__1427);
  and g__150(w__1970 ,in28[6] ,w__1537);
  or g__151(w__1969 ,w__1733 ,w__1912);
  or g__152(w__1968 ,w__1851 ,w__1935);
  and g__153(w__1967 ,w__2305 ,w__1589);
  and g__154(w__1966 ,in28[5] ,w__1524);
  or g__155(w__1965 ,w__1849 ,w__1934);
  and g__156(w__1964 ,w__2314 ,w__1542);
  or g__157(w__1963 ,w__1848 ,w__1933);
  and g__158(w__1962 ,in28[3] ,w__1548);
  or g__159(w__1961 ,w__1847 ,w__1951);
  and g__160(w__1960 ,w__2306 ,w__1451);
  and g__161(w__1959 ,in28[0] ,w__1548);
  and g__162(w__1958 ,in28[2] ,w__1549);
  and g__163(w__1957 ,w__2311 ,w__1543);
  and g__164(w__1956 ,in28[1] ,w__1536);
  or g__165(w__1955 ,w__1827 ,w__1929);
  or g__166(w__1954 ,w__1842 ,w__1928);
  or g__167(w__1988 ,w__1875 ,w__1917);
  or g__168(w__1987 ,w__1828 ,w__1913);
  or g__169(w__2139 ,w__1873 ,w__1915);
  or g__170(w__1986 ,w__1869 ,w__1918);
  or g__171(w__1985 ,w__1830 ,w__1914);
  or g__172(w__2147 ,w__1872 ,w__1920);
  or g__173(w__1984 ,w__1892 ,w__1923);
  or g__174(w__2144 ,w__1874 ,w__1916);
  or g__175(w__2143 ,w__1870 ,w__1911);
  and g__176(w__1951 ,w__2272 ,w__1587);
  and g__177(w__1950 ,w__1640 ,w__1605);
  and g__178(w__1949 ,w__1628 ,w__1423);
  and g__179(w__1948 ,w__1655 ,w__1528);
  and g__180(w__1947 ,w__1619 ,w__1501);
  and g__181(w__1946 ,w__2282 ,w__1460);
  and g__182(w__1945 ,w__2281 ,w__1540);
  and g__183(w__1944 ,w__2280 ,w__1437);
  and g__184(w__1943 ,w__1637 ,w__1527);
  and g__185(w__1942 ,w__2279 ,w__1539);
  and g__186(w__1941 ,w__1646 ,w__1469);
  and g__187(w__1940 ,w__2278 ,w__1458);
  and g__188(w__1939 ,w__1649 ,w__1469);
  and g__189(w__1938 ,w__2277 ,w__1458);
  and g__190(w__1937 ,w__1643 ,w__1423);
  and g__191(w__1936 ,w__2276 ,w__1460);
  and g__192(w__1935 ,w__2275 ,w__1437);
  and g__193(w__1934 ,w__2274 ,w__1586);
  and g__194(w__1933 ,w__2273 ,w__1539);
  and g__195(w__1953 ,w__1695 ,w__1908);
  and g__196(w__1952 ,w__1693 ,w__1909);
  or g__197(w__1930 ,w__1859 ,w__1901);
  and g__198(w__1929 ,w__2271 ,w__1457);
  and g__199(w__1928 ,w__2270 ,w__1540);
  and g__200(w__1927 ,w__1634 ,w__1501);
  and g__201(w__1926 ,w__1631 ,w__1604);
  and g__202(w__1925 ,w__1622 ,w__1527);
  and g__203(w__1924 ,w__1625 ,w__1468);
  or g__204(w__1923 ,w__1817 ,w__1903);
  or g__205(w__1922 ,w__1816 ,w__1904);
  or g__206(w__1921 ,w__1814 ,w__1902);
  or g__207(w__1920 ,w__1818 ,w__1905);
  and g__208(w__1919 ,w__1652 ,w__1528);
  or g__209(w__1918 ,w__1794 ,w__1894);
  or g__210(w__1917 ,w__1807 ,w__1900);
  or g__211(w__1916 ,w__1804 ,w__1898);
  or g__212(w__1915 ,w__1802 ,w__1899);
  or g__213(w__1914 ,w__1843 ,w__1895);
  or g__214(w__1913 ,w__1844 ,w__1897);
  or g__215(w__1912 ,w__1868 ,w__1910);
  or g__216(w__1911 ,w__1795 ,w__1896);
  and g__217(w__1932 ,in11 ,w__1908);
  and g__218(w__1931 ,in19 ,w__1909);
  or g__219(w__1907 ,w__1786 ,w__2126);
  or g__220(w__1906 ,w__1784 ,w__2127);
  and g__221(w__1905 ,w__2269 ,w__1593);
  and g__222(w__1904 ,w__2257 ,w__1421);
  and g__223(w__1903 ,w__2264 ,w__1510);
  and g__224(w__1902 ,w__2267 ,w__1471);
  and g__225(w__1901 ,w__2263 ,w__1509);
  and g__226(w__1900 ,w__2262 ,w__1489);
  and g__227(w__1899 ,w__2261 ,w__1489);
  and g__228(w__1898 ,w__2266 ,w__1421);
  and g__229(w__1897 ,w__2260 ,w__1471);
  and g__230(w__1896 ,w__2265 ,w__1592);
  and g__231(w__1895 ,w__2268 ,w__1509);
  and g__232(w__1894 ,w__2259 ,w__1488);
  or g__233(w__1893 ,w__1783 ,w__2128);
  or g__234(w__1892 ,w__1704 ,w__1864);
  or g__235(w__1891 ,w__1780 ,w__2132);
  or g__236(w__1890 ,w__1793 ,w__2131);
  or g__237(w__1889 ,w__1785 ,w__2130);
  or g__238(w__1888 ,w__1782 ,w__2129);
  and g__239(w__1910 ,w__2258 ,w__1510);
  and g__240(w__1909 ,w__1687 ,w__1866);
  and g__241(w__1908 ,w__1696 ,w__1868);
  or g__242(w__1885 ,w__1819 ,w__2125);
  or g__243(w__1884 ,w__1820 ,w__2124);
  or g__244(w__1883 ,w__1778 ,w__1825);
  or g__245(w__2158 ,w__1792 ,w__2122);
  or g__246(w__1882 ,w__1726 ,w__1863);
  or g__247(w__1881 ,w__1712 ,w__1862);
  or g__248(w__1880 ,w__1815 ,w__1861);
  or g__249(w__1879 ,w__1779 ,w__2133);
  or g__250(w__1878 ,w__1812 ,w__1860);
  or g__251(w__1877 ,w__1811 ,w__1858);
  or g__252(w__2170 ,w__1781 ,w__2134);
  or g__253(w__1876 ,w__1810 ,w__1857);
  or g__254(w__1875 ,w__1720 ,w__1855);
  or g__255(w__1874 ,w__1728 ,w__1852);
  or g__256(w__1873 ,w__1754 ,w__1850);
  or g__257(w__1872 ,w__1709 ,w__1846);
  or g__258(w__1871 ,w__1797 ,w__1845);
  or g__259(w__1870 ,w__1740 ,w__1841);
  or g__260(w__1869 ,w__1710 ,w__1867);
  or g__261(w__2123 ,w__1734 ,w__1838);
  and g__262(w__1887 ,in10 ,w__1868);
  and g__263(w__1886 ,in18 ,w__1865);
  and g__264(w__1867 ,w__2367 ,w__1611);
  nor g__265(w__1866 ,in17 ,w__1822);
  nor g__266(w__1865 ,in17 ,w__1822);
  and g__267(w__1864 ,w__2372 ,w__1495);
  and g__268(w__1863 ,w__2365 ,w__1513);
  and g__269(w__1862 ,w__2375 ,w__1493);
  and g__270(w__1861 ,w__2269 ,w__1581);
  and g__271(w__1860 ,w__2268 ,w__1449);
  and g__272(w__1859 ,w__2371 ,w__1512);
  and g__273(w__1858 ,w__2267 ,w__1516);
  and g__274(w__1857 ,w__2266 ,w__1433);
  and g__275(w__1856 ,w__2265 ,w__1515);
  and g__276(w__1855 ,w__2370 ,w__1480);
  and g__277(w__1854 ,w__2264 ,w__1474);
  and g__278(w__1853 ,w__2263 ,w__1474);
  and g__279(w__1852 ,w__2374 ,w__1480);
  and g__280(w__1851 ,w__2262 ,w__1449);
  and g__281(w__1850 ,w__2369 ,w__1495);
  and g__282(w__1849 ,w__2261 ,w__1433);
  and g__283(w__1848 ,w__2260 ,w__1580);
  and g__284(w__1847 ,w__2259 ,w__1515);
  and g__285(w__1846 ,w__2377 ,w__1493);
  and g__286(w__1845 ,w__2258 ,w__1473);
  and g__287(w__1844 ,w__2368 ,w__1610);
  and g__288(w__1843 ,w__2376 ,w__1512);
  and g__289(w__1842 ,w__2257 ,w__1516);
  and g__290(w__1841 ,w__2373 ,w__1479);
  and g__291(w__1868 ,w__1688 ,w__1823);
  or g__292(w__1838 ,w__1566 ,w__1790);
  or g__293(w__1837 ,w__1703 ,w__1813);
  or g__294(w__1836 ,w__1730 ,w__1809);
  or g__295(w__1835 ,w__1718 ,w__1808);
  or g__296(w__1834 ,w__1724 ,w__1806);
  or g__297(w__1833 ,w__1713 ,w__1805);
  or g__298(w__1832 ,w__1711 ,w__1803);
  or g__299(w__1831 ,w__1739 ,w__1801);
  or g__300(w__1830 ,w__1708 ,w__1800);
  or g__301(w__1829 ,w__1706 ,w__1799);
  or g__302(w__1828 ,w__1715 ,w__1798);
  and g__303(w__1827 ,in17 ,w__1821);
  or g__304(w__1826 ,w__1701 ,w__1796);
  or g__305(w__1825 ,w__1734 ,w__1790);
  and g__306(w__1840 ,w__2366 ,w__1513);
  or g__307(w__2134 ,w__1657 ,w__1771);
  or g__308(w__2133 ,w__1657 ,w__1770);
  or g__309(w__2132 ,w__1732 ,w__1773);
  or g__310(w__2131 ,w__1732 ,w__1769);
  or g__311(w__2130 ,w__1719 ,w__1768);
  or g__312(w__2129 ,w__1698 ,w__1766);
  or g__313(w__2128 ,w__1741 ,w__1765);
  or g__314(w__2127 ,w__1721 ,w__1764);
  or g__315(w__2126 ,w__1714 ,w__1763);
  or g__316(w__2125 ,w__1700 ,w__1762);
  or g__317(w__2124 ,w__1742 ,w__1761);
  or g__318(w__2122 ,w__1753 ,w__1767);
  and g__319(w__1839 ,in8 ,w__1823);
  not g__320(w__1822 ,w__1821);
  and g__321(w__1820 ,w__1633 ,w__1565);
  and g__322(w__1819 ,w__1639 ,w__1578);
  and g__323(w__1818 ,w__2256 ,w__1602);
  and g__324(w__1817 ,w__2251 ,w__1447);
  and g__325(w__1816 ,w__2244 ,w__1519);
  and g__326(w__1815 ,w__2256 ,w__1608);
  and g__327(w__1814 ,w__2254 ,w__1431);
  and g__328(w__1813 ,w__2250 ,w__1518);
  and g__329(w__1812 ,w__2255 ,w__1499);
  and g__330(w__1811 ,w__2254 ,w__1534);
  and g__331(w__1810 ,w__2253 ,w__1497);
  and g__332(w__1809 ,w__2252 ,w__1533);
  and g__333(w__1808 ,w__2251 ,w__1466);
  and g__334(w__1807 ,w__2249 ,w__1477);
  and g__335(w__1806 ,w__2250 ,w__1466);
  and g__336(w__1805 ,w__2249 ,w__1499);
  and g__337(w__1804 ,w__2253 ,w__1477);
  and g__338(w__1803 ,w__2248 ,w__1497);
  and g__339(w__1802 ,w__2248 ,w__1447);
  and g__340(w__1801 ,w__2247 ,w__1607);
  and g__341(w__1800 ,w__2255 ,w__1431);
  and g__342(w__1799 ,w__2246 ,w__1533);
  and g__343(w__1798 ,w__2247 ,w__1601);
  and g__344(w__1797 ,w__2245 ,w__1465);
  and g__345(w__1796 ,w__2244 ,w__1534);
  and g__346(w__1795 ,w__2252 ,w__1518);
  and g__347(w__1794 ,w__2246 ,w__1476);
  and g__348(w__2149 ,w__1674 ,w__1568);
  and g__349(w__1793 ,w__1645 ,w__1562);
  and g__350(w__1792 ,w__1654 ,w__1575);
  and g__351(w__1791 ,w__1680 ,w__1565);
  and g__352(w__2155 ,w__1664 ,w__1569);
  and g__353(w__2153 ,w__1666 ,w__1577);
  and g__354(w__2151 ,w__1679 ,w__1578);
  and g__355(w__1824 ,w__2245 ,w__1519);
  and g__356(w__1823 ,w__1694 ,w__1716);
  and g__357(w__1821 ,w__1690 ,w__1699);
  and g__358(w__2150 ,w__1677 ,w__1566);
  and g__359(w__1787 ,w__1672 ,w__1575);
  and g__360(w__1786 ,w__1642 ,w__1572);
  and g__361(w__1785 ,w__1651 ,w__1562);
  and g__362(w__1784 ,w__1636 ,w__1574);
  and g__363(w__2154 ,w__1662 ,w__1571);
  and g__364(w__2152 ,w__1668 ,w__1574);
  and g__365(w__1783 ,w__1618 ,w__1569);
  and g__366(w__1782 ,w__1621 ,w__1563);
  and g__367(w__2156 ,w__1670 ,w__1568);
  and g__368(w__1781 ,w__1630 ,w__1563);
  and g__369(w__1780 ,w__1624 ,w__1577);
  and g__370(w__1779 ,w__1648 ,w__1572);
  and g__371(w__1778 ,w__1627 ,w__1571);
  or g__372(w__2438 ,w__2439 ,w__1743);
  or g__373(w__2437 ,w__1735 ,w__1744);
  or g__374(w__2436 ,w__1736 ,w__1748);
  or g__375(w__1777 ,w__1752 ,w__1751);
  or g__376(w__1776 ,w__1729 ,w__1745);
  or g__377(w__1775 ,w__1727 ,w__1750);
  or g__378(w__1774 ,w__1707 ,w__1746);
  or g__379(w__2235 ,w__1738 ,w__1749);
  and g__380(w__1773 ,in39[10] ,w__1584);
  or g__381(w__1772 ,w__1717 ,w__1747);
  and g__382(w__1771 ,in39[12] ,w__1435);
  and g__383(w__1770 ,in39[11] ,w__1531);
  and g__384(w__1769 ,in39[9] ,w__1425);
  and g__385(w__1768 ,in39[8] ,w__1530);
  and g__386(w__1767 ,in39[0] ,w__1463);
  and g__387(w__1766 ,in39[7] ,w__1463);
  and g__388(w__1765 ,in39[6] ,w__1435);
  and g__389(w__1764 ,in39[5] ,w__1425);
  and g__390(w__1763 ,in39[4] ,w__1583);
  and g__391(w__1762 ,in39[3] ,w__1530);
  and g__392(w__1761 ,in39[2] ,w__1462);
  and g__393(w__1790 ,in39[1] ,w__1531);
  and g__394(w__1789 ,in16 ,w__1697);
  and g__395(w__1788 ,in7 ,w__1737);
  not g__396(w__1758 ,w__1755);
  not g__397(w__1757 ,w__1755);
  not g__398(w__1756 ,w__1755);
  and g__399(w__1754 ,in5 ,w__2222);
  and g__400(w__1753 ,in37 ,w__1672);
  and g__401(w__1752 ,in29[5] ,w__1675);
  and g__402(w__2405 ,w__1622 ,w__1556);
  and g__403(w__2400 ,w__1634 ,w__1557);
  and g__404(w__1751 ,in28[5] ,w__1557);
  and g__405(w__1750 ,in28[2] ,w__1486);
  and g__406(w__1749 ,in28[0] ,w__1504);
  and g__407(w__1748 ,in28[6] ,w__1506);
  and g__408(w__2407 ,w__1646 ,w__1556);
  and g__409(w__2403 ,w__1637 ,w__1503);
  and g__410(w__1747 ,in28[3] ,w__1485);
  and g__411(w__2399 ,w__1628 ,w__1503);
  and g__412(w__1746 ,in28[1] ,w__1486);
  and g__413(w__2404 ,w__1619 ,w__1559);
  and g__414(w__1745 ,in28[4] ,w__1613);
  and g__415(w__2398 ,w__1655 ,w__1559);
  and g__416(w__2401 ,w__1640 ,w__1560);
  and g__417(w__2409 ,w__1649 ,w__1560);
  and g__418(w__1744 ,in28[7] ,w__1491);
  and g__419(w__2402 ,w__1643 ,w__1507);
  and g__420(w__2410 ,w__1631 ,w__1504);
  and g__421(w__2406 ,w__1652 ,w__1506);
  and g__422(w__1743 ,in28[8] ,w__1507);
  and g__423(w__2408 ,w__1625 ,w__1491);
  and g__424(w__1742 ,in37 ,w__1677);
  and g__425(w__1741 ,in37 ,w__1662);
  and g__426(w__1740 ,in5 ,w__2239);
  and g__427(w__1739 ,in14 ,w__2221);
  and g__428(w__1738 ,in29[0] ,w__1682);
  nor g__429(w__1737 ,in5 ,in6);
  and g__430(w__1736 ,in29[6] ,w__1554);
  and g__431(w__1735 ,in29[7] ,w__1660);
  and g__432(w__2439 ,in29[8] ,w__1675);
  and g__433(w__1760 ,in6 ,w__1686);
  and g__434(w__1759 ,in15 ,w__1691);
  or g__435(w__1755 ,w__1689 ,in37);
  and g__436(w__1730 ,in14 ,w__2239);
  and g__437(w__1729 ,in29[4] ,w__1554);
  and g__438(w__1728 ,in5 ,w__2240);
  and g__439(w__1727 ,in29[2] ,w__1659);
  and g__440(w__1726 ,in5 ,w__2218);
  and g__441(w__1725 ,in14 ,w__2242);
  and g__442(w__1724 ,in14 ,w__2237);
  and g__443(w__1723 ,in14 ,w__2241);
  and g__444(w__1722 ,in14 ,w__2240);
  and g__445(w__1721 ,in37 ,w__1666);
  and g__446(w__1720 ,in5 ,w__2236);
  and g__447(w__1719 ,in37 ,w__1670);
  and g__448(w__1718 ,in14 ,w__2238);
  and g__449(w__1717 ,in29[3] ,w__1659);
  nor g__450(w__1716 ,in5 ,in6);
  and g__451(w__1715 ,in5 ,w__2221);
  and g__452(w__1714 ,in37 ,w__1668);
  and g__453(w__1713 ,in14 ,w__2236);
  and g__454(w__1712 ,in5 ,w__2241);
  and g__455(w__1711 ,in14 ,w__2222);
  and g__456(w__1710 ,in5 ,w__2220);
  and g__457(w__1709 ,in5 ,w__2243);
  and g__458(w__1708 ,in5 ,w__2242);
  and g__459(w__1707 ,in29[1] ,w__1660);
  and g__460(w__1706 ,in14 ,w__2220);
  and g__461(w__1705 ,in14 ,w__2243);
  and g__462(w__1704 ,in5 ,w__2238);
  and g__463(w__1703 ,in5 ,w__2237);
  and g__464(w__1702 ,in14 ,w__2219);
  and g__465(w__1701 ,in14 ,w__2218);
  and g__466(w__1700 ,in37 ,w__1679);
  nor g__467(w__1699 ,in14 ,in15);
  and g__468(w__1698 ,in37 ,w__1664);
  nor g__469(w__1697 ,in14 ,in15);
  and g__470(w__1734 ,in37 ,w__1674);
  and g__471(w__1733 ,in5 ,w__2219);
  and g__472(w__1732 ,in37 ,w__1680);
  and g__473(w__1731 ,w__1692 ,w__1689);
  not g__474(w__1696 ,in10);
  not g__475(w__1695 ,in11);
  not g__476(w__1694 ,in7);
  not g__477(w__1693 ,in19);
  not g__478(w__1692 ,in37);
  not g__479(w__1691 ,in14);
  not g__480(w__1690 ,in16);
  not g__481(w__1689 ,in38);
  not g__482(w__1688 ,in8);
  not g__483(w__1687 ,in18);
  not g__484(w__1686 ,in5);
  not g__485(w__1685 ,in30);
  not g__486(w__1684 ,in30);
  not g__487(w__1683 ,w__1681);
  not g__488(w__1682 ,w__1681);
  not g__489(w__1681 ,in30);
  not g__490(w__1679 ,w__1678);
  not g__491(w__1678 ,w__2332);
  not g__492(w__1677 ,w__1676);
  not g__493(w__1676 ,w__2331);
  not g__494(w__1675 ,w__1681);
  not g__495(w__1674 ,w__1673);
  not g__496(w__1673 ,w__2330);
  not g__497(w__1672 ,w__1671);
  not g__498(w__1671 ,w__2316);
  not g__499(w__1670 ,w__1669);
  not g__500(w__1669 ,w__2337);
  not g__501(w__1668 ,w__1667);
  not g__502(w__1667 ,w__2333);
  not g__503(w__1666 ,w__1665);
  not g__504(w__1665 ,w__2334);
  not g__505(w__1664 ,w__1663);
  not g__506(w__1663 ,w__2336);
  not g__507(w__1662 ,w__1661);
  not g__508(w__1661 ,w__2335);
  not g__509(w__1660 ,w__1658);
  not g__510(w__1659 ,w__1658);
  not g__511(w__1658 ,w__1683);
  not g__512(w__1657 ,w__1656);
  not g__513(w__1656 ,w__1732);
  not g__514(w__1655 ,w__1653);
  not g__515(w__1654 ,w__1653);
  not g__516(w__1653 ,w__2411);
  not g__517(w__1652 ,w__1650);
  not g__518(w__1651 ,w__1650);
  not g__519(w__1650 ,w__2419);
  not g__520(w__1649 ,w__1647);
  not g__521(w__1648 ,w__1647);
  not g__522(w__1647 ,w__2422);
  not g__523(w__1646 ,w__1644);
  not g__524(w__1645 ,w__1644);
  not g__525(w__1644 ,w__2420);
  not g__526(w__1643 ,w__1641);
  not g__527(w__1642 ,w__1641);
  not g__528(w__1641 ,w__2415);
  not g__529(w__1640 ,w__1638);
  not g__530(w__1639 ,w__1638);
  not g__531(w__1638 ,w__2414);
  not g__532(w__1637 ,w__1635);
  not g__533(w__1636 ,w__1635);
  not g__534(w__1635 ,w__2416);
  not g__535(w__1634 ,w__1632);
  not g__536(w__1633 ,w__1632);
  not g__537(w__1632 ,w__2413);
  not g__538(w__1631 ,w__1629);
  not g__539(w__1630 ,w__1629);
  not g__540(w__1629 ,w__2423);
  not g__541(w__1628 ,w__1626);
  not g__542(w__1627 ,w__1626);
  not g__543(w__1626 ,w__2412);
  not g__544(w__1625 ,w__1623);
  not g__545(w__1624 ,w__1623);
  not g__546(w__1623 ,w__2421);
  not g__547(w__1622 ,w__1620);
  not g__548(w__1621 ,w__1620);
  not g__549(w__1620 ,w__2418);
  not g__550(w__1619 ,w__1617);
  not g__551(w__1618 ,w__1617);
  not g__552(w__1617 ,w__2417);
  buf g__553(w__2140 ,w__1988);
  buf g__554(w__2145 ,w__2018);
  buf g__555(w__2138 ,w__1987);
  buf g__556(w__2137 ,w__1986);
  buf g__557(w__2146 ,w__1985);
  buf g__558(w__2142 ,w__1984);
  buf g__559(w__2163 ,w__1906);
  buf g__560(w__2161 ,w__1885);
  buf g__561(w__2165 ,w__1888);
  buf g__562(w__2160 ,w__1884);
  buf g__563(w__2159 ,w__1883);
  buf g__564(w__2169 ,w__1879);
  buf g__565(w__2168 ,w__1891);
  buf g__566(w__2167 ,w__1890);
  buf g__567(w__2166 ,w__1889);
  buf g__568(w__2164 ,w__1893);
  buf g__569(w__2162 ,w__1907);
  buf g__570(w__2434 ,w__1776);
  buf g__571(w__2435 ,w__1777);
  buf g__572(w__2433 ,w__1772);
  buf g__573(w__2432 ,w__1775);
  buf g__574(w__2431 ,w__1774);
  buf g__575(w__2157 ,w__1791);
  buf g__576(w__2148 ,w__1787);
  not g__577(w__1616 ,w__1615);
  not g__578(w__1615 ,w__1952);
  not g__579(w__1614 ,w__1612);
  not g__580(w__1613 ,w__1612);
  not g__581(w__1612 ,w__1685);
  not g__582(w__1611 ,w__1609);
  not g__583(w__1610 ,w__1609);
  not g__584(w__1609 ,w__1788);
  not g__585(w__1608 ,w__1606);
  not g__586(w__1607 ,w__1606);
  not g__587(w__1606 ,w__1759);
  not g__588(w__1605 ,w__1603);
  not g__589(w__1604 ,w__1603);
  not g__590(w__1603 ,w__1887);
  not g__591(w__1602 ,w__1600);
  not g__592(w__1601 ,w__1600);
  not g__593(w__1600 ,w__1760);
  not g__594(w__1599 ,w__1597);
  not g__595(w__1598 ,w__1597);
  not g__596(w__1597 ,w__1931);
  not g__597(w__1596 ,w__1594);
  not g__598(w__1595 ,w__1594);
  not g__599(w__1594 ,w__1932);
  not g__600(w__1593 ,w__1591);
  not g__601(w__1592 ,w__1591);
  not g__602(w__1591 ,w__1839);
  not g__603(w__1590 ,w__1588);
  not g__604(w__1589 ,w__1588);
  not g__605(w__1588 ,w__1953);
  not g__606(w__1587 ,w__1585);
  not g__607(w__1586 ,w__1585);
  not g__608(w__1585 ,w__1886);
  not g__609(w__1584 ,w__1582);
  not g__610(w__1583 ,w__1582);
  not g__611(w__1582 ,w__1731);
  not g__612(w__1581 ,w__1579);
  not g__613(w__1580 ,w__1579);
  not g__614(w__1579 ,w__1789);
  buf g__615(w__1680 ,w__2338);
  not g__616(w__1578 ,w__1576);
  not g__617(w__1577 ,w__1576);
  not g__618(w__1576 ,w__1758);
  not g__619(w__1575 ,w__1573);
  not g__620(w__1574 ,w__1573);
  not g__621(w__1573 ,w__1757);
  not g__622(w__1572 ,w__1570);
  not g__623(w__1571 ,w__1570);
  not g__624(w__1570 ,w__1756);
  not g__625(w__1569 ,w__1567);
  not g__626(w__1568 ,w__1567);
  not g__627(w__1567 ,w__1757);
  not g__628(w__1566 ,w__1564);
  not g__629(w__1565 ,w__1564);
  not g__630(w__1564 ,w__1756);
  not g__631(w__1563 ,w__1561);
  not g__632(w__1562 ,w__1561);
  not g__633(w__1561 ,w__1758);
  not g__634(w__1560 ,w__1558);
  not g__635(w__1559 ,w__1558);
  not g__636(w__1558 ,w__1684);
  not g__637(w__1557 ,w__1555);
  not g__638(w__1556 ,w__1555);
  not g__639(w__1555 ,w__1684);
  not g__640(w__1554 ,w__1553);
  not g__641(w__1553 ,w__1682);
  not g__642(w__1552 ,w__1550);
  not g__643(w__1551 ,w__1550);
  not g__644(w__1550 ,w__1952);
  not g__645(w__1549 ,w__1547);
  not g__646(w__1548 ,w__1547);
  not g__647(w__1547 ,w__1616);
  not g__648(w__1546 ,w__1544);
  not g__649(w__1545 ,w__1544);
  not g__650(w__1544 ,w__1932);
  not g__651(w__1543 ,w__1541);
  not g__652(w__1542 ,w__1541);
  not g__653(w__1541 ,w__1953);
  not g__654(w__1540 ,w__1538);
  not g__655(w__1539 ,w__1538);
  not g__656(w__1538 ,w__1886);
  not g__657(w__1537 ,w__1535);
  not g__658(w__1536 ,w__1535);
  not g__659(w__1535 ,w__1616);
  not g__660(w__1534 ,w__1532);
  not g__661(w__1533 ,w__1532);
  not g__662(w__1532 ,w__1759);
  not g__663(w__1531 ,w__1529);
  not g__664(w__1530 ,w__1529);
  not g__665(w__1529 ,w__1731);
  not g__666(w__1528 ,w__1526);
  not g__667(w__1527 ,w__1526);
  not g__668(w__1526 ,w__1887);
  not g__669(w__1525 ,w__1523);
  not g__670(w__1524 ,w__1523);
  not g__671(w__1523 ,w__1952);
  not g__672(w__1522 ,w__1520);
  not g__673(w__1521 ,w__1520);
  not g__674(w__1520 ,w__1931);
  not g__675(w__1519 ,w__1517);
  not g__676(w__1518 ,w__1517);
  not g__677(w__1517 ,w__1760);
  not g__678(w__1516 ,w__1514);
  not g__679(w__1515 ,w__1514);
  not g__680(w__1514 ,w__1789);
  not g__681(w__1513 ,w__1511);
  not g__682(w__1512 ,w__1511);
  not g__683(w__1511 ,w__1788);
  not g__684(w__1510 ,w__1508);
  not g__685(w__1509 ,w__1508);
  not g__686(w__1508 ,w__1839);
  not g__687(w__1507 ,w__1505);
  not g__688(w__1506 ,w__1505);
  not g__689(w__1505 ,w__1685);
  not g__690(w__1504 ,w__1502);
  not g__691(w__1503 ,w__1502);
  not g__692(w__1502 ,w__1614);
  not g__693(w__1501 ,w__1500);
  not g__694(w__1500 ,w__1605);
  not g__695(w__1499 ,w__1498);
  not g__696(w__1498 ,w__1607);
  not g__697(w__1497 ,w__1496);
  not g__698(w__1496 ,w__1608);
  not g__699(w__1495 ,w__1494);
  not g__700(w__1494 ,w__1610);
  not g__701(w__1493 ,w__1492);
  not g__702(w__1492 ,w__1611);
  not g__703(w__1491 ,w__1490);
  not g__704(w__1490 ,w__1613);
  not g__705(w__1489 ,w__1487);
  not g__706(w__1488 ,w__1487);
  not g__707(w__1487 ,w__1839);
  not g__708(w__1486 ,w__1484);
  not g__709(w__1485 ,w__1484);
  not g__710(w__1484 ,w__1685);
  not g__711(w__1483 ,w__1481);
  not g__712(w__1482 ,w__1481);
  not g__713(w__1481 ,w__1931);
  not g__714(w__1480 ,w__1478);
  not g__715(w__1479 ,w__1478);
  not g__716(w__1478 ,w__1788);
  not g__717(w__1477 ,w__1475);
  not g__718(w__1476 ,w__1475);
  not g__719(w__1475 ,w__1760);
  not g__720(w__1474 ,w__1472);
  not g__721(w__1473 ,w__1472);
  not g__722(w__1472 ,w__1789);
  not g__723(w__1471 ,w__1470);
  not g__724(w__1470 ,w__1593);
  not g__725(w__1469 ,w__1467);
  not g__726(w__1468 ,w__1467);
  not g__727(w__1467 ,w__1887);
  not g__728(w__1466 ,w__1464);
  not g__729(w__1465 ,w__1464);
  not g__730(w__1464 ,w__1759);
  not g__731(w__1463 ,w__1461);
  not g__732(w__1462 ,w__1461);
  not g__733(w__1461 ,w__1731);
  not g__734(w__1460 ,w__1459);
  not g__735(w__1459 ,w__1586);
  not g__736(w__1458 ,w__1456);
  not g__737(w__1457 ,w__1456);
  not g__738(w__1456 ,w__1886);
  not g__739(w__1455 ,w__1453);
  not g__740(w__1454 ,w__1453);
  not g__741(w__1453 ,w__1932);
  not g__742(w__1452 ,w__1450);
  not g__743(w__1451 ,w__1450);
  not g__744(w__1450 ,w__1953);
  not g__745(w__1449 ,w__1448);
  not g__746(w__1448 ,w__1580);
  not g__747(w__1447 ,w__1446);
  not g__748(w__1446 ,w__1601);
  not g__749(w__1445 ,w__1444);
  not g__750(w__1444 ,w__1599);
  not g__751(w__1443 ,w__1442);
  not g__752(w__1442 ,w__1596);
  not g__753(w__1441 ,w__1440);
  not g__754(w__1440 ,w__1595);
  not g__755(w__1439 ,w__1438);
  not g__756(w__1438 ,w__1589);
  not g__757(w__1437 ,w__1436);
  not g__758(w__1436 ,w__1587);
  not g__759(w__1435 ,w__1434);
  not g__760(w__1434 ,w__1583);
  not g__761(w__1433 ,w__1432);
  not g__762(w__1432 ,w__1581);
  not g__763(w__1431 ,w__1430);
  not g__764(w__1430 ,w__1602);
  not g__765(w__1429 ,w__1428);
  not g__766(w__1428 ,w__1598);
  not g__767(w__1427 ,w__1426);
  not g__768(w__1426 ,w__1590);
  not g__769(w__1425 ,w__1424);
  not g__770(w__1424 ,w__1584);
  not g__771(w__1423 ,w__1422);
  not g__772(w__1422 ,w__1604);
  not g__773(w__1421 ,w__1420);
  not g__774(w__1420 ,w__1592);
  or g__775(w__1419 ,w__1824 ,w__1840);
  xor g__776(w__1418 ,in21[6] ,in22);
  xor g__777(w__1417 ,in21[4] ,in22);
  xor g__778(w__1416 ,in21[2] ,in22);
  xor g__779(w__1415 ,in21[0] ,in22);
  xor g__780(w__1414 ,in21[5] ,in22);
  xor g__781(w__1413 ,in21[1] ,in22);
  xor g__782(w__1412 ,in21[3] ,in22);
  buf g__783(w__2302 ,w__1418);
  buf g__784(w__2299 ,w__1412);
  buf g__785(w__2297 ,w__1413);
  buf g__786(w__2301 ,w__1414);
  buf g__787(w__2296 ,w__1415);
  buf g__788(w__2298 ,w__1416);
  buf g__789(w__2300 ,w__1417);
  xor g__790(w__2430 ,in26[6] ,in27);
  xor g__791(w__2428 ,in26[4] ,in27);
  xor g__792(w__2426 ,in26[2] ,in27);
  xor g__793(w__1411 ,in26[0] ,in27);
  xor g__794(w__2429 ,in26[5] ,in27);
  xor g__795(w__1410 ,in26[1] ,in27);
  xor g__796(w__2427 ,in26[3] ,in27);
  buf g__797(w__2424 ,w__1411);
  buf g__798(w__2425 ,w__1410);
  buf g__799(w__2588 ,w__2484);
  buf g__800(w__2587 ,w__2471);
  buf g__801(w__2586 ,w__2485);
  buf g__802(w__2585 ,w__2472);
  buf g__803(w__2584 ,w__2486);
  buf g__804(w__2583 ,w__2473);
  buf g__805(w__2582 ,w__2487);
  buf g__806(w__2581 ,w__2474);
  buf g__807(w__2580 ,w__2488);
  buf g__808(w__2579 ,w__2475);
  buf g__809(w__2578 ,w__2489);
  buf g__810(w__2577 ,w__2476);
  buf g__811(w__2576 ,w__2490);
  buf g__812(w__2575 ,w__2477);
  buf g__813(w__2574 ,w__2491);
  buf g__814(w__2573 ,w__2478);
  buf g__815(w__2572 ,w__2492);
  buf g__816(w__2571 ,w__2479);
  buf g__817(w__2570 ,w__2493);
  buf g__818(w__2569 ,w__2494);
  buf g__819(w__2568 ,w__2481);
  buf g__820(w__2567 ,w__2495);
  buf g__821(w__2566 ,w__2496);
  buf g__822(w__2565 ,w__2480);
  buf g__823(w__2564 ,w__2482);
  buf g__824(w__2563 ,w__2483);
  or g__825(w__2197 ,w__2507 ,w__2551);
  or g__826(w__2562 ,w__2509 ,w__2546);
  or g__827(w__2561 ,w__2536 ,w__2548);
  or g__828(w__2560 ,w__2508 ,w__2547);
  or g__829(w__2559 ,w__2504 ,w__2543);
  or g__830(w__2558 ,w__2505 ,w__2545);
  or g__831(w__2185 ,w__2506 ,w__2550);
  or g__832(w__2557 ,w__2537 ,w__2544);
  or g__833(w__2556 ,w__2501 ,w__2540);
  or g__834(w__2555 ,w__2500 ,w__2538);
  or g__835(w__2554 ,w__2502 ,w__2541);
  or g__836(w__2553 ,w__2499 ,w__2539);
  or g__837(w__2552 ,w__2503 ,w__2542);
  and g__838(w__2551 ,w__2587 ,w__2465);
  and g__839(w__2550 ,w__2563 ,w__2463);
  and g__840(w__2548 ,w__2575 ,w__2462);
  and g__841(w__2547 ,w__2573 ,w__2441);
  and g__842(w__2546 ,w__2581 ,w__2448);
  and g__843(w__2545 ,w__2571 ,w__2443);
  and g__844(w__2544 ,w__2585 ,w__2448);
  and g__845(w__2543 ,w__2579 ,w__2447);
  and g__846(w__2542 ,w__2565 ,w__2443);
  and g__847(w__2541 ,w__2568 ,w__2445);
  and g__848(w__2540 ,w__2583 ,w__2447);
  and g__849(w__2539 ,w__2564 ,w__2445);
  and g__850(w__2538 ,w__2577 ,w__2441);
  and g__851(w__2537 ,w__2453 ,w__2586);
  and g__852(w__2536 ,w__2456 ,w__2576);
  and g__853(w__2509 ,w__2457 ,w__2582);
  and g__854(w__2508 ,w__2454 ,w__2574);
  and g__855(w__2507 ,w__2457 ,w__2588);
  and g__856(w__2506 ,w__2460 ,w__2566);
  and g__857(w__2505 ,w__2459 ,w__2572);
  and g__858(w__2504 ,w__2451 ,w__2580);
  and g__859(w__2503 ,w__2454 ,w__2570);
  and g__860(w__2502 ,w__2450 ,w__2569);
  and g__861(w__2501 ,w__2459 ,w__2584);
  and g__862(w__2500 ,w__2451 ,w__2578);
  and g__863(w__2499 ,w__2460 ,w__2567);
  not g__864(w__2498 ,w__2470);
  not g__865(w__2497 ,w__2470);
  not g__866(w__2470 ,w__2468);
  not g__867(w__2469 ,w__2468);
  not g__868(w__2468 ,w__2467);
  not g__869(w__2467 ,w__2081);
  buf g__870(w__2188 ,w__2552);
  buf g__871(w__2186 ,w__2553);
  buf g__872(w__2187 ,w__2554);
  buf g__873(w__2192 ,w__2555);
  buf g__874(w__2195 ,w__2556);
  buf g__875(w__2196 ,w__2557);
  buf g__876(w__2191 ,w__2561);
  buf g__877(w__2193 ,w__2559);
  buf g__878(w__2190 ,w__2560);
  buf g__879(w__2189 ,w__2558);
  buf g__880(w__2194 ,w__2562);
  not g__881(w__2466 ,w__2464);
  not g__882(w__2465 ,w__2464);
  not g__883(w__2464 ,w__2469);
  not g__884(w__2463 ,w__2461);
  not g__885(w__2462 ,w__2461);
  not g__886(w__2461 ,w__2469);
  not g__887(w__2460 ,w__2458);
  not g__888(w__2459 ,w__2458);
  not g__889(w__2458 ,w__2497);
  not g__890(w__2457 ,w__2455);
  not g__891(w__2456 ,w__2455);
  not g__892(w__2455 ,w__2498);
  not g__893(w__2454 ,w__2452);
  not g__894(w__2453 ,w__2452);
  not g__895(w__2452 ,w__2498);
  not g__896(w__2451 ,w__2449);
  not g__897(w__2450 ,w__2449);
  not g__898(w__2449 ,w__2497);
  not g__899(w__2448 ,w__2446);
  not g__900(w__2447 ,w__2446);
  not g__901(w__2446 ,w__2466);
  not g__902(w__2445 ,w__2444);
  not g__903(w__2444 ,w__2462);
  not g__904(w__2443 ,w__2442);
  not g__905(w__2442 ,w__2463);
  not g__906(w__2441 ,w__2440);
  not g__907(w__2440 ,w__2465);
  buf g__908(w__2761 ,w__2223);
  buf g__909(w__2760 ,w__2230);
  buf g__910(w__2759 ,w__2224);
  buf g__911(w__2758 ,w__2225);
  buf g__912(w__2757 ,w__2226);
  buf g__913(w__2756 ,w__2227);
  buf g__914(w__2755 ,w__2228);
  buf g__915(w__2754 ,w__2229);
  buf g__916(w__2753 ,w__2231);
  buf g__917(w__2752 ,w__2232);
  buf g__918(w__2751 ,w__2233);
  buf g__919(w__2750 ,w__2234);
  buf g__920(w__2749 ,w__2235);
  or g__921(w__2364 ,w__2716 ,w__2737);
  or g__922(w__2363 ,w__2719 ,w__2742);
  or g__923(w__2359 ,w__2721 ,w__2745);
  or g__924(w__2353 ,w__2720 ,w__2744);
  or g__925(w__2358 ,w__2717 ,w__2735);
  or g__926(w__2352 ,w__2718 ,w__2743);
  or g__927(w__2354 ,w__2709 ,w__2747);
  or g__928(w__2357 ,w__2714 ,w__2739);
  or g__929(w__2748 ,w__2710 ,w__2746);
  or g__930(w__2360 ,w__2712 ,w__2736);
  or g__931(w__2356 ,w__2713 ,w__2738);
  or g__932(w__2355 ,w__2711 ,w__2741);
  or g__933(w__2361 ,w__2715 ,w__2740);
  or g__934(w__2747 ,w__2667 ,w__2733);
  or g__935(w__2746 ,w__2649 ,w__2730);
  or g__936(w__2745 ,w__2665 ,w__2731);
  or g__937(w__2744 ,w__2664 ,w__2732);
  or g__938(w__2743 ,w__2660 ,w__2729);
  or g__939(w__2742 ,w__2653 ,w__2725);
  or g__940(w__2741 ,w__2642 ,w__2723);
  or g__941(w__2740 ,w__2652 ,w__2726);
  or g__942(w__2739 ,w__2651 ,w__2727);
  or g__943(w__2738 ,w__2647 ,w__2724);
  or g__944(w__2737 ,w__2659 ,w__2734);
  or g__945(w__2736 ,w__2643 ,w__2728);
  or g__946(w__2735 ,w__2656 ,w__2722);
  nor g__947(w__2734 ,w__2674 ,w__2698);
  nor g__948(w__2733 ,w__2672 ,w__2708);
  nor g__949(w__2732 ,w__2678 ,w__2706);
  nor g__950(w__2731 ,w__2693 ,w__2702);
  nor g__951(w__2730 ,w__2692 ,w__2705);
  nor g__952(w__2729 ,w__2676 ,w__2707);
  nor g__953(w__2728 ,w__2677 ,w__2696);
  nor g__954(w__2727 ,w__2694 ,w__2703);
  nor g__955(w__2726 ,w__2671 ,w__2701);
  nor g__956(w__2725 ,w__2673 ,w__2700);
  nor g__957(w__2724 ,w__2670 ,w__2699);
  nor g__958(w__2723 ,w__2669 ,w__2697);
  nor g__959(w__2722 ,w__2675 ,w__2704);
  and g__960(w__2721 ,w__2418 ,w__2622);
  and g__961(w__2720 ,w__2412 ,w__2602);
  and g__962(w__2719 ,w__2422 ,w__2611);
  and g__963(w__2718 ,w__2411 ,w__2595);
  and g__964(w__2717 ,w__2417 ,w__2612);
  and g__965(w__2716 ,w__2423 ,w__2593);
  and g__966(w__2715 ,w__2420 ,w__2593);
  and g__967(w__2714 ,w__2416 ,w__2602);
  and g__968(w__2713 ,w__2415 ,w__2595);
  and g__969(w__2712 ,w__2419 ,w__2623);
  and g__970(w__2711 ,w__2414 ,w__2612);
  and g__971(w__2710 ,w__2421 ,w__2592);
  and g__972(w__2709 ,w__2413 ,w__2611);
  or g__973(w__2708 ,w__2666 ,w__2625);
  or g__974(w__2707 ,w__2657 ,w__2590);
  or g__975(w__2706 ,w__2663 ,w__2614);
  or g__976(w__2705 ,w__2658 ,w__2597);
  or g__977(w__2704 ,w__2654 ,w__2615);
  or g__978(w__2703 ,w__2650 ,w__2600);
  or g__979(w__2702 ,w__2646 ,w__2600);
  or g__980(w__2701 ,w__2648 ,w__2590);
  or g__981(w__2700 ,w__2644 ,w__2597);
  or g__982(w__2699 ,w__2645 ,w__2626);
  or g__983(w__2698 ,w__2655 ,w__2615);
  or g__984(w__2697 ,w__2661 ,w__2599);
  or g__985(w__2696 ,w__2668 ,w__2614);
  nor g__986(w__2694 ,w__2606 ,w__2760);
  nor g__987(w__2693 ,w__2604 ,w__2755);
  nor g__988(w__2692 ,w__2628 ,w__2758);
  nor g__989(w__2678 ,w__2604 ,w__2750);
  nor g__990(w__2677 ,w__2609 ,w__2756);
  nor g__991(w__2676 ,w__2629 ,w__2749);
  nor g__992(w__2675 ,w__2617 ,w__2754);
  nor g__993(w__2674 ,w__2618 ,w__2761);
  nor g__994(w__2673 ,w__2609 ,w__2759);
  nor g__995(w__2672 ,w__2617 ,w__2751);
  nor g__996(w__2671 ,w__2618 ,w__2757);
  nor g__997(w__2670 ,w__2607 ,w__2753);
  nor g__998(w__2669 ,w__2607 ,w__2752);
  nor g__999(w__2668 ,w__2632 ,in35[8]);
  and g__1000(w__2667 ,in32 ,w__2367);
  nor g__1001(w__2666 ,w__2631 ,in35[2]);
  and g__1002(w__2665 ,in32 ,w__2372);
  and g__1003(w__2664 ,in32 ,w__2366);
  nor g__1004(w__2663 ,w__2636 ,in35[1]);
  and g__1005(w__2695 ,in33 ,w__2641);
  nor g__1006(w__2661 ,w__2620 ,in35[3]);
  and g__1007(w__2660 ,in32 ,w__2365);
  and g__1008(w__2659 ,in32 ,w__2377);
  nor g__1009(w__2658 ,w__2631 ,in35[10]);
  nor g__1010(w__2657 ,w__2634 ,in35[0]);
  and g__1011(w__2656 ,in32 ,w__2371);
  nor g__1012(w__2655 ,w__2620 ,in35[12]);
  nor g__1013(w__2654 ,w__2636 ,in35[6]);
  and g__1014(w__2653 ,in32 ,w__2376);
  and g__1015(w__2652 ,in32 ,w__2374);
  and g__1016(w__2651 ,in32 ,w__2370);
  nor g__1017(w__2650 ,w__2632 ,in35[5]);
  and g__1018(w__2649 ,in32 ,w__2375);
  nor g__1019(w__2648 ,w__2635 ,in35[9]);
  and g__1020(w__2647 ,in32 ,w__2369);
  nor g__1021(w__2646 ,w__2640 ,in35[7]);
  nor g__1022(w__2645 ,w__2635 ,in35[4]);
  nor g__1023(w__2644 ,w__2634 ,in35[11]);
  and g__1024(w__2643 ,in32 ,w__2373);
  and g__1025(w__2642 ,in32 ,w__2368);
  or g__1026(w__2662 ,in32 ,in33);
  not g__1027(w__2641 ,in32);
  not g__1028(w__2640 ,w__2638);
  not g__1029(w__2639 ,w__2638);
  not g__1030(w__2638 ,in34);
  not g__1031(w__2637 ,in34);
  not g__1032(w__2636 ,w__2638);
  not g__1033(w__2635 ,w__2633);
  not g__1034(w__2634 ,w__2633);
  not g__1035(w__2633 ,w__2639);
  not g__1036(w__2632 ,w__2630);
  not g__1037(w__2631 ,w__2630);
  not g__1038(w__2630 ,w__2639);
  buf g__1039(w__2362 ,w__2748);
  not g__1040(w__2629 ,w__2627);
  not g__1041(w__2628 ,w__2627);
  not g__1042(w__2627 ,w__2637);
  not g__1043(w__2626 ,w__2624);
  not g__1044(w__2625 ,w__2624);
  not g__1045(w__2624 ,w__2662);
  not g__1046(w__2623 ,w__2621);
  not g__1047(w__2622 ,w__2621);
  not g__1048(w__2621 ,w__2695);
  not g__1049(w__2620 ,w__2619);
  not g__1050(w__2619 ,w__2640);
  not g__1051(w__2618 ,w__2616);
  not g__1052(w__2617 ,w__2616);
  not g__1053(w__2616 ,w__2637);
  not g__1054(w__2615 ,w__2613);
  not g__1055(w__2614 ,w__2613);
  not g__1056(w__2613 ,w__2662);
  not g__1057(w__2612 ,w__2610);
  not g__1058(w__2611 ,w__2610);
  not g__1059(w__2610 ,w__2695);
  not g__1060(w__2609 ,w__2608);
  not g__1061(w__2608 ,w__2628);
  not g__1062(w__2607 ,w__2605);
  not g__1063(w__2606 ,w__2605);
  not g__1064(w__2605 ,w__2637);
  not g__1065(w__2604 ,w__2603);
  not g__1066(w__2603 ,w__2629);
  not g__1067(w__2602 ,w__2601);
  not g__1068(w__2601 ,w__2623);
  not g__1069(w__2600 ,w__2598);
  not g__1070(w__2599 ,w__2598);
  not g__1071(w__2598 ,w__2662);
  not g__1072(w__2597 ,w__2596);
  not g__1073(w__2596 ,w__2625);
  not g__1074(w__2595 ,w__2594);
  not g__1075(w__2594 ,w__2622);
  not g__1076(w__2593 ,w__2591);
  not g__1077(w__2592 ,w__2591);
  not g__1078(w__2591 ,w__2695);
  not g__1079(w__2590 ,w__2589);
  not g__1080(w__2589 ,w__2626);
  buf g__1081(w__2793 ,w__2317);
  buf g__1082(w__2792 ,w__2318);
  buf g__1083(w__2791 ,w__2320);
  buf g__1084(w__2790 ,w__2326);
  buf g__1085(w__2789 ,w__2328);
  buf g__1086(w__2788 ,w__2321);
  buf g__1087(w__2787 ,w__2325);
  buf g__1088(w__2786 ,w__2329);
  buf g__1089(w__2785 ,w__2319);
  buf g__1090(w__2784 ,w__2322);
  buf g__1091(w__2783 ,w__2324);
  buf g__1092(w__2782 ,w__2327);
  buf g__1093(w__2781 ,w__2323);
  not g__1094(w__2780 ,in33);
  not g__1095(w__2779 ,in32);
  and g__1096(w__2351 ,w__2793 ,w__2766);
  and g__1097(w__2350 ,w__2792 ,w__2765);
  and g__1098(w__2347 ,w__2788 ,w__2766);
  and g__1099(w__2342 ,w__2790 ,w__2764);
  and g__1100(w__2341 ,w__2782 ,w__2763);
  and g__1101(w__2340 ,w__2789 ,w__2776);
  and g__1102(w__2343 ,w__2787 ,w__2762);
  and g__1103(w__2346 ,w__2784 ,w__2764);
  and g__1104(w__2778 ,w__2786 ,w__2762);
  and g__1105(w__2345 ,w__2781 ,w__2763);
  and g__1106(w__2348 ,w__2791 ,w__2765);
  and g__1107(w__2344 ,w__2783 ,w__2774);
  and g__1108(w__2777 ,w__2785 ,w__2775);
  and g__1109(w__2776 ,in34 ,w__2771);
  and g__1110(w__2775 ,in34 ,w__2772);
  and g__1111(w__2774 ,in34 ,w__2767);
  and g__1112(w__2773 ,w__2779 ,w__2780);
  buf g__1113(w__2349 ,w__2777);
  buf g__1114(w__2339 ,w__2778);
  not g__1115(w__2772 ,w__2770);
  not g__1116(w__2771 ,w__2770);
  not g__1117(w__2770 ,w__2773);
  not g__1118(w__2769 ,w__2768);
  not g__1119(w__2768 ,w__2773);
  not g__1120(w__2767 ,w__2768);
  and g__1121(w__2766 ,in34 ,w__2769);
  and g__1122(w__2765 ,in34 ,w__2772);
  and g__1123(w__2764 ,in34 ,w__2769);
  and g__1124(w__2763 ,in34 ,w__2771);
  and g__1125(w__2762 ,in34 ,w__2767);
  buf g__1126(w__2927 ,w__2521);
  buf g__1127(w__2926 ,w__2522);
  buf g__1128(w__2925 ,w__2533);
  buf g__1129(w__2924 ,w__2535);
  buf g__1130(w__2923 ,w__2520);
  buf g__1131(w__2922 ,w__2534);
  buf g__1132(w__2921 ,w__2523);
  buf g__1133(w__2920 ,w__2510);
  buf g__1134(w__2919 ,w__2524);
  buf g__1135(w__2918 ,w__2511);
  buf g__1136(w__2917 ,w__2525);
  buf g__1137(w__2916 ,w__2512);
  buf g__1138(w__2915 ,w__2526);
  buf g__1139(w__2914 ,w__2513);
  buf g__1140(w__2913 ,w__2527);
  buf g__1141(w__2912 ,w__2514);
  buf g__1142(w__2911 ,w__2528);
  buf g__1143(w__2910 ,w__2515);
  buf g__1144(w__2909 ,w__2529);
  buf g__1145(w__2908 ,w__2516);
  buf g__1146(w__2907 ,w__2530);
  buf g__1147(w__2906 ,w__2517);
  buf g__1148(w__2905 ,w__2531);
  buf g__1149(w__2904 ,w__2518);
  buf g__1150(w__2903 ,w__2532);
  buf g__1151(w__2902 ,w__2519);
  or g__1152(w__2184 ,w__2872 ,w__2889);
  or g__1153(w__2901 ,w__2874 ,w__2885);
  or g__1154(w__2900 ,w__2875 ,w__2887);
  or g__1155(w__2899 ,w__2873 ,w__2886);
  or g__1156(w__2898 ,w__2869 ,w__2882);
  or g__1157(w__2897 ,w__2870 ,w__2884);
  or g__1158(w__2896 ,w__2871 ,w__2888);
  or g__1159(w__2895 ,w__2876 ,w__2883);
  or g__1160(w__2894 ,w__2866 ,w__2879);
  or g__1161(w__2893 ,w__2865 ,w__2877);
  or g__1162(w__2892 ,w__2867 ,w__2880);
  or g__1163(w__2891 ,w__2864 ,w__2878);
  or g__1164(w__2890 ,w__2868 ,w__2881);
  and g__1165(w__2889 ,w__2920 ,w__2855);
  and g__1166(w__2887 ,w__2908 ,w__2852);
  and g__1167(w__2886 ,w__2906 ,w__2795);
  and g__1168(w__2885 ,w__2914 ,w__2815);
  and g__1169(w__2884 ,w__2904 ,w__2797);
  and g__1170(w__2883 ,w__2918 ,w__2815);
  and g__1171(w__2882 ,w__2912 ,w__2814);
  and g__1172(w__2881 ,w__2902 ,w__2797);
  and g__1173(w__2880 ,w__2923 ,w__2799);
  and g__1174(w__2879 ,w__2916 ,w__2814);
  and g__1175(w__2878 ,w__2927 ,w__2799);
  and g__1176(w__2877 ,w__2910 ,w__2795);
  and g__1177(w__2876 ,w__2820 ,w__2919);
  and g__1178(w__2875 ,w__2823 ,w__2909);
  and g__1179(w__2874 ,w__2824 ,w__2915);
  and g__1180(w__2873 ,w__2821 ,w__2907);
  and g__1181(w__2872 ,w__2824 ,w__2921);
  and g__1182(w__2870 ,w__2849 ,w__2905);
  and g__1183(w__2869 ,w__2818 ,w__2913);
  and g__1184(w__2868 ,w__2821 ,w__2903);
  and g__1185(w__2867 ,w__2817 ,w__2925);
  and g__1186(w__2866 ,w__2849 ,w__2917);
  and g__1187(w__2865 ,w__2818 ,w__2911);
  and g__1188(w__2864 ,w__2850 ,w__2922);
  not g__1189(w__2863 ,w__2860);
  not g__1190(w__2861 ,w__2860);
  not g__1191(w__2860 ,w__2858);
  not g__1192(w__2859 ,w__2858);
  not g__1193(w__2858 ,w__2857);
  not g__1194(w__2857 ,w__2081);
  buf g__1195(w__2175 ,w__2890);
  buf g__1196(w__2173 ,w__2891);
  buf g__1197(w__2174 ,w__2892);
  buf g__1198(w__2179 ,w__2893);
  buf g__1199(w__2182 ,w__2894);
  buf g__1200(w__2177 ,w__2899);
  buf g__1201(w__2178 ,w__2900);
  buf g__1202(w__2176 ,w__2897);
  buf g__1203(w__2180 ,w__2898);
  buf g__1204(w__2181 ,w__2901);
  buf g__1205(w__2172 ,w__2896);
  buf g__1206(w__2183 ,w__2895);
  not g__1207(w__2856 ,w__2854);
  not g__1208(w__2855 ,w__2854);
  not g__1209(w__2854 ,w__2859);
  not g__1210(w__2853 ,w__2851);
  not g__1211(w__2852 ,w__2851);
  not g__1212(w__2851 ,w__2859);
  not g__1213(w__2850 ,w__2825);
  not g__1214(w__2849 ,w__2825);
  not g__1215(w__2825 ,w__2861);
  not g__1216(w__2824 ,w__2822);
  not g__1217(w__2823 ,w__2822);
  not g__1218(w__2822 ,w__2863);
  not g__1219(w__2821 ,w__2819);
  not g__1220(w__2820 ,w__2819);
  not g__1221(w__2819 ,w__2863);
  not g__1222(w__2818 ,w__2816);
  not g__1223(w__2817 ,w__2816);
  not g__1224(w__2816 ,w__2861);
  not g__1225(w__2815 ,w__2813);
  not g__1226(w__2814 ,w__2813);
  not g__1227(w__2813 ,w__2856);
  not g__1228(w__2799 ,w__2798);
  not g__1229(w__2798 ,w__2852);
  not g__1230(w__2797 ,w__2796);
  not g__1231(w__2796 ,w__2853);
  not g__1232(w__2795 ,w__2794);
  not g__1233(w__2794 ,w__2855);
  buf g__1234(w__2934 ,w__2205);
  not g__1235(w__2933 ,w__2549);
  or g__1236(w__2932 ,w__2930 ,w__2931);
  nor g__1237(w__2931 ,w__2933 ,w__2929);
  and g__1238(w__2930 ,w__2929 ,w__2934);
  not g__1239(w__2929 ,w__2928);
  not g__1240(w__2928 ,w__2081);
  buf g__1241(w__2171 ,w__2932);
  buf g__1242(w__3030 ,w__2688);
  buf g__1243(w__3029 ,w__2800);
  buf g__1244(w__3028 ,w__2679);
  buf g__1245(w__3027 ,w__2801);
  buf g__1246(w__3026 ,w__2680);
  buf g__1247(w__3025 ,w__2802);
  buf g__1248(w__3024 ,w__2681);
  buf g__1249(w__3023 ,w__2803);
  buf g__1250(w__3022 ,w__2682);
  buf g__1251(w__3021 ,w__2804);
  buf g__1252(w__3020 ,w__2683);
  buf g__1253(w__3019 ,w__2805);
  buf g__1254(w__3018 ,w__2684);
  buf g__1255(w__3017 ,w__2806);
  buf g__1256(w__3016 ,w__2685);
  buf g__1257(w__3015 ,w__2807);
  buf g__1258(w__3014 ,w__2686);
  buf g__1259(w__3013 ,w__2808);
  buf g__1260(w__3012 ,w__2687);
  buf g__1261(w__3011 ,w__2809);
  buf g__1262(w__3010 ,w__2691);
  buf g__1263(w__3009 ,w__2810);
  buf g__1264(w__3008 ,w__2689);
  buf g__1265(w__3007 ,w__2811);
  buf g__1266(w__3006 ,w__2690);
  buf g__1267(w__3005 ,w__2812);
  or g__1268(w__2108 ,w__2976 ,w__2993);
  or g__1269(w__3004 ,w__2978 ,w__2989);
  or g__1270(w__3003 ,w__2979 ,w__2991);
  or g__1271(w__3002 ,w__2977 ,w__2990);
  or g__1272(w__3001 ,w__2973 ,w__2986);
  or g__1273(w__3000 ,w__2974 ,w__2988);
  or g__1274(w__2096 ,w__2975 ,w__2992);
  or g__1275(w__2999 ,w__2980 ,w__2987);
  or g__1276(w__2998 ,w__2970 ,w__2983);
  or g__1277(w__2997 ,w__2969 ,w__2981);
  or g__1278(w__2996 ,w__2971 ,w__2984);
  or g__1279(w__2995 ,w__2968 ,w__2982);
  or g__1280(w__2994 ,w__2972 ,w__2985);
  and g__1281(w__2993 ,w__3028 ,w__2960);
  and g__1282(w__2992 ,w__3010 ,w__2958);
  and g__1283(w__2991 ,w__3016 ,w__2957);
  and g__1284(w__2990 ,w__3014 ,w__2936);
  and g__1285(w__2989 ,w__3022 ,w__2943);
  and g__1286(w__2988 ,w__3012 ,w__2938);
  and g__1287(w__2987 ,w__3026 ,w__2943);
  and g__1288(w__2986 ,w__3020 ,w__2942);
  and g__1289(w__2985 ,w__3030 ,w__2938);
  and g__1290(w__2984 ,w__3008 ,w__2940);
  and g__1291(w__2983 ,w__3024 ,w__2942);
  and g__1292(w__2982 ,w__3006 ,w__2940);
  and g__1293(w__2981 ,w__3018 ,w__2936);
  and g__1294(w__2980 ,w__2948 ,w__3027);
  and g__1295(w__2979 ,w__2951 ,w__3017);
  and g__1296(w__2978 ,w__2952 ,w__3023);
  and g__1297(w__2977 ,w__2949 ,w__3015);
  and g__1298(w__2976 ,w__2952 ,w__3029);
  and g__1299(w__2975 ,w__2955 ,w__3005);
  and g__1300(w__2974 ,w__2954 ,w__3013);
  and g__1301(w__2973 ,w__2946 ,w__3021);
  and g__1302(w__2972 ,w__2949 ,w__3011);
  and g__1303(w__2971 ,w__2945 ,w__3009);
  and g__1304(w__2970 ,w__2954 ,w__3025);
  and g__1305(w__2969 ,w__2946 ,w__3019);
  and g__1306(w__2968 ,w__2955 ,w__3007);
  not g__1307(w__2967 ,w__2965);
  not g__1308(w__2966 ,w__2965);
  not g__1309(w__2965 ,w__2963);
  not g__1310(w__2964 ,w__2963);
  not g__1311(w__2963 ,w__2962);
  not g__1312(w__2962 ,w__2080);
  buf g__1313(w__2099 ,w__2994);
  buf g__1314(w__2097 ,w__2995);
  buf g__1315(w__2098 ,w__2996);
  buf g__1316(w__2103 ,w__2997);
  buf g__1317(w__2106 ,w__2998);
  buf g__1318(w__2107 ,w__2999);
  buf g__1319(w__2102 ,w__3003);
  buf g__1320(w__2104 ,w__3001);
  buf g__1321(w__2101 ,w__3002);
  buf g__1322(w__2100 ,w__3000);
  buf g__1323(w__2105 ,w__3004);
  not g__1324(w__2961 ,w__2959);
  not g__1325(w__2960 ,w__2959);
  not g__1326(w__2959 ,w__2964);
  not g__1327(w__2958 ,w__2956);
  not g__1328(w__2957 ,w__2956);
  not g__1329(w__2956 ,w__2964);
  not g__1330(w__2955 ,w__2953);
  not g__1331(w__2954 ,w__2953);
  not g__1332(w__2953 ,w__2966);
  not g__1333(w__2952 ,w__2950);
  not g__1334(w__2951 ,w__2950);
  not g__1335(w__2950 ,w__2967);
  not g__1336(w__2949 ,w__2947);
  not g__1337(w__2948 ,w__2947);
  not g__1338(w__2947 ,w__2967);
  not g__1339(w__2946 ,w__2944);
  not g__1340(w__2945 ,w__2944);
  not g__1341(w__2944 ,w__2966);
  not g__1342(w__2943 ,w__2941);
  not g__1343(w__2942 ,w__2941);
  not g__1344(w__2941 ,w__2961);
  not g__1345(w__2940 ,w__2939);
  not g__1346(w__2939 ,w__2957);
  not g__1347(w__2938 ,w__2937);
  not g__1348(w__2937 ,w__2958);
  not g__1349(w__2936 ,w__2935);
  not g__1350(w__2935 ,w__2960);
  buf g__1351(w__3127 ,w__2838);
  buf g__1352(w__3126 ,w__2826);
  buf g__1353(w__3125 ,w__2839);
  buf g__1354(w__3124 ,w__2827);
  buf g__1355(w__3123 ,w__2840);
  buf g__1356(w__3122 ,w__2828);
  buf g__1357(w__3121 ,w__2841);
  buf g__1358(w__3120 ,w__2829);
  buf g__1359(w__3119 ,w__2842);
  buf g__1360(w__3118 ,w__2830);
  buf g__1361(w__3117 ,w__2843);
  buf g__1362(w__3116 ,w__2831);
  buf g__1363(w__3115 ,w__2844);
  buf g__1364(w__3114 ,w__2845);
  buf g__1365(w__3113 ,w__2833);
  buf g__1366(w__3112 ,w__2846);
  buf g__1367(w__3111 ,w__2834);
  buf g__1368(w__3110 ,w__2847);
  buf g__1369(w__3109 ,w__2848);
  buf g__1370(w__3108 ,w__2836);
  buf g__1371(w__3107 ,w__2149);
  buf g__1372(w__3106 ,w__2158);
  buf g__1373(w__3105 ,w__2109);
  buf g__1374(w__3104 ,w__2837);
  buf g__1375(w__3103 ,w__2832);
  buf g__1376(w__3102 ,w__2835);
  or g__1377(w__2095 ,w__3072 ,w__3089);
  or g__1378(w__3101 ,w__3074 ,w__3085);
  or g__1379(w__3100 ,w__3075 ,w__3087);
  or g__1380(w__3099 ,w__3073 ,w__3086);
  or g__1381(w__3098 ,w__3069 ,w__3082);
  or g__1382(w__3097 ,w__3070 ,w__3084);
  or g__1383(w__3096 ,w__3071 ,w__3088);
  or g__1384(w__3095 ,w__3076 ,w__3083);
  or g__1385(w__3094 ,w__3066 ,w__3079);
  or g__1386(w__3093 ,w__3065 ,w__3077);
  or g__1387(w__3092 ,w__3067 ,w__3080);
  or g__1388(w__3091 ,w__3064 ,w__3078);
  or g__1389(w__3090 ,w__3068 ,w__3081);
  and g__1390(w__3089 ,w__3126 ,w__3056);
  and g__1391(w__3088 ,w__3104 ,w__3054);
  and g__1392(w__3087 ,w__3103 ,w__3053);
  and g__1393(w__3086 ,w__3113 ,w__3032);
  and g__1394(w__3085 ,w__3120 ,w__3039);
  and g__1395(w__3084 ,w__3111 ,w__3034);
  and g__1396(w__3083 ,w__3124 ,w__3039);
  and g__1397(w__3082 ,w__3118 ,w__3038);
  and g__1398(w__3081 ,w__3102 ,w__3034);
  and g__1399(w__3080 ,w__3108 ,w__3036);
  and g__1400(w__3079 ,w__3122 ,w__3038);
  and g__1401(w__3078 ,w__3106 ,w__3036);
  and g__1402(w__3077 ,w__3116 ,w__3032);
  and g__1403(w__3076 ,w__3044 ,w__3125);
  and g__1404(w__3075 ,w__3047 ,w__3115);
  and g__1405(w__3074 ,w__3048 ,w__3121);
  and g__1406(w__3073 ,w__3045 ,w__3114);
  and g__1407(w__3072 ,w__3048 ,w__3127);
  and g__1408(w__3071 ,w__3051 ,w__3105);
  and g__1409(w__3070 ,w__3050 ,w__3112);
  and g__1410(w__3069 ,w__3042 ,w__3119);
  and g__1411(w__3068 ,w__3045 ,w__3110);
  and g__1412(w__3067 ,w__3041 ,w__3109);
  and g__1413(w__3066 ,w__3050 ,w__3123);
  and g__1414(w__3065 ,w__3042 ,w__3117);
  and g__1415(w__3064 ,w__3051 ,w__3107);
  not g__1416(w__3063 ,w__3061);
  not g__1417(w__3062 ,w__3061);
  not g__1418(w__3061 ,w__3059);
  not g__1419(w__3060 ,w__3059);
  not g__1420(w__3059 ,w__3058);
  not g__1421(w__3058 ,w__2080);
  buf g__1422(w__2086 ,w__3090);
  buf g__1423(w__2084 ,w__3091);
  buf g__1424(w__2085 ,w__3092);
  buf g__1425(w__2090 ,w__3093);
  buf g__1426(w__2093 ,w__3094);
  buf g__1427(w__2088 ,w__3099);
  buf g__1428(w__2089 ,w__3100);
  buf g__1429(w__2087 ,w__3097);
  buf g__1430(w__2091 ,w__3098);
  buf g__1431(w__2092 ,w__3101);
  buf g__1432(w__2083 ,w__3096);
  buf g__1433(w__2094 ,w__3095);
  not g__1434(w__3057 ,w__3055);
  not g__1435(w__3056 ,w__3055);
  not g__1436(w__3055 ,w__3060);
  not g__1437(w__3054 ,w__3052);
  not g__1438(w__3053 ,w__3052);
  not g__1439(w__3052 ,w__3060);
  not g__1440(w__3051 ,w__3049);
  not g__1441(w__3050 ,w__3049);
  not g__1442(w__3049 ,w__3062);
  not g__1443(w__3048 ,w__3046);
  not g__1444(w__3047 ,w__3046);
  not g__1445(w__3046 ,w__3063);
  not g__1446(w__3045 ,w__3043);
  not g__1447(w__3044 ,w__3043);
  not g__1448(w__3043 ,w__3063);
  not g__1449(w__3042 ,w__3040);
  not g__1450(w__3041 ,w__3040);
  not g__1451(w__3040 ,w__3062);
  not g__1452(w__3039 ,w__3037);
  not g__1453(w__3038 ,w__3037);
  not g__1454(w__3037 ,w__3057);
  not g__1455(w__3036 ,w__3035);
  not g__1456(w__3035 ,w__3053);
  not g__1457(w__3034 ,w__3033);
  not g__1458(w__3033 ,w__3054);
  not g__1459(w__3032 ,w__3031);
  not g__1460(w__3031 ,w__3056);
  buf g__1461(w__3134 ,w__2122);
  not g__1462(w__3133 ,w__2862);
  or g__1463(w__3132 ,w__3130 ,w__3131);
  nor g__1464(w__3131 ,w__3133 ,w__3129);
  and g__1465(w__3130 ,w__3129 ,w__3134);
  not g__1466(w__3129 ,w__3128);
  not g__1467(w__3128 ,w__2080);
  buf g__1468(w__2082 ,w__3132);
  xnor g__1469(w__2377 ,w__48 ,w__2390);
  or g__1470(w__48 ,w__19 ,w__47);
  or g__1471(w__47 ,w__14 ,w__46);
  or g__1472(w__46 ,w__20 ,w__45);
  or g__1473(w__45 ,w__16 ,w__44);
  or g__1474(w__44 ,w__17 ,w__43);
  or g__1475(w__43 ,w__13 ,w__42);
  or g__1476(w__42 ,w__18 ,w__41);
  and g__1477(w__2369 ,w__41 ,w__40);
  or g__1478(w__41 ,w__15 ,w__39);
  or g__1479(w__40 ,w__2 ,w__38);
  not g__1480(w__39 ,w__38);
  or g__1481(w__38 ,w__26 ,w__37);
  xnor g__1482(w__2368 ,w__36 ,w__30);
  and g__1483(w__37 ,w__24 ,w__36);
  or g__1484(w__36 ,w__25 ,w__35);
  xnor g__1485(w__2367 ,w__34 ,w__32);
  and g__1486(w__35 ,w__23 ,w__34);
  xor g__1487(w__2366 ,w__22 ,w__31);
  or g__1488(w__34 ,w__29 ,w__33);
  nor g__1489(w__33 ,w__22 ,w__27);
  and g__1490(w__2365 ,w__22 ,w__28);
  xnor g__1491(w__32 ,w__5 ,in4[2]);
  xnor g__1492(w__31 ,w__10 ,in4[1]);
  xnor g__1493(w__30 ,w__8 ,in4[3]);
  and g__1494(w__29 ,w__10 ,in4[1]);
  or g__1495(w__28 ,w__1 ,in4[0]);
  nor g__1496(w__27 ,w__11 ,in4[1]);
  and g__1497(w__26 ,w__7 ,in4[3]);
  and g__1498(w__25 ,w__4 ,in4[2]);
  or g__1499(w__24 ,w__8 ,in4[3]);
  or g__1500(w__23 ,w__5 ,in4[2]);
  or g__1501(w__22 ,w__12 ,w__21);
  not g__1502(w__21 ,in4[0]);
  not g__1503(w__11 ,w__9);
  not g__1504(w__10 ,w__9);
  not g__1505(w__9 ,w__2379);
  not g__1506(w__8 ,w__6);
  not g__1507(w__7 ,w__6);
  not g__1508(w__6 ,w__2381);
  not g__1509(w__5 ,w__3);
  not g__1510(w__4 ,w__3);
  not g__1511(w__3 ,w__2380);
  not g__1512(w__18 ,w__2383);
  not g__1513(w__2 ,w__15);
  not g__1514(w__15 ,w__2382);
  not g__1515(w__16 ,w__2386);
  not g__1516(w__17 ,w__2385);
  not g__1517(w__14 ,w__2388);
  not g__1518(w__19 ,w__2389);
  not g__1519(w__20 ,w__2387);
  not g__1520(w__13 ,w__2384);
  not g__1521(w__1 ,w__12);
  not g__1522(w__12 ,w__2378);
  xor g__1523(w__2370 ,w__41 ,w__18);
  xor g__1524(w__2373 ,w__44 ,w__16);
  xor g__1525(w__2372 ,w__43 ,w__17);
  xor g__1526(w__2375 ,w__46 ,w__14);
  xor g__1527(w__2376 ,w__47 ,w__19);
  xor g__1528(w__2374 ,w__45 ,w__20);
  xor g__1529(w__2371 ,w__42 ,w__13);
  xnor g__1530(w__2243 ,w__108 ,w__2390);
  or g__1531(w__108 ,w__68 ,w__107);
  or g__1532(w__107 ,w__69 ,w__106);
  or g__1533(w__106 ,w__70 ,w__105);
  or g__1534(w__105 ,w__72 ,w__104);
  or g__1535(w__104 ,w__66 ,w__103);
  and g__1536(w__2237 ,w__103 ,w__102);
  or g__1537(w__103 ,w__67 ,w__101);
  or g__1538(w__102 ,w__50 ,w__100);
  not g__1539(w__101 ,w__100);
  or g__1540(w__100 ,w__85 ,w__99);
  xnor g__1541(w__2236 ,w__98 ,w__90);
  and g__1542(w__99 ,w__75 ,w__98);
  or g__1543(w__98 ,w__83 ,w__97);
  xnor g__1544(w__2222 ,w__96 ,w__89);
  and g__1545(w__97 ,w__77 ,w__96);
  or g__1546(w__96 ,w__81 ,w__95);
  xnor g__1547(w__2221 ,w__94 ,w__88);
  and g__1548(w__95 ,w__84 ,w__94);
  or g__1549(w__94 ,w__76 ,w__93);
  xnor g__1550(w__2220 ,w__92 ,w__87);
  and g__1551(w__93 ,w__74 ,w__92);
  xor g__1552(w__2219 ,w__79 ,w__86);
  or g__1553(w__92 ,w__78 ,w__91);
  nor g__1554(w__91 ,w__79 ,w__80);
  and g__1555(w__2218 ,w__79 ,w__82);
  xnor g__1556(w__90 ,w__56 ,in13[5]);
  xnor g__1557(w__89 ,w__53 ,in13[4]);
  xnor g__1558(w__88 ,w__62 ,in13[3]);
  xnor g__1559(w__87 ,w__59 ,in13[2]);
  xnor g__1560(w__86 ,w__64 ,in13[1]);
  and g__1561(w__85 ,in13[5] ,w__55);
  or g__1562(w__84 ,in13[3] ,w__61);
  and g__1563(w__83 ,in13[4] ,w__52);
  or g__1564(w__82 ,in13[0] ,w__49);
  and g__1565(w__81 ,in13[3] ,w__62);
  nor g__1566(w__80 ,in13[1] ,w__65);
  and g__1567(w__78 ,in13[1] ,w__64);
  or g__1568(w__77 ,in13[4] ,w__53);
  and g__1569(w__76 ,in13[2] ,w__58);
  or g__1570(w__75 ,in13[5] ,w__56);
  or g__1571(w__74 ,in13[2] ,w__59);
  or g__1572(w__79 ,w__73 ,w__71);
  not g__1573(w__73 ,in13[0]);
  not g__1574(w__65 ,w__63);
  not g__1575(w__64 ,w__63);
  not g__1576(w__63 ,w__2379);
  not g__1577(w__62 ,w__60);
  not g__1578(w__61 ,w__60);
  not g__1579(w__60 ,w__2381);
  not g__1580(w__59 ,w__57);
  not g__1581(w__58 ,w__57);
  not g__1582(w__57 ,w__2380);
  not g__1583(w__56 ,w__54);
  not g__1584(w__55 ,w__54);
  not g__1585(w__54 ,w__2383);
  not g__1586(w__53 ,w__51);
  not g__1587(w__52 ,w__51);
  not g__1588(w__51 ,w__2382);
  not g__1589(w__66 ,w__2385);
  not g__1590(w__72 ,w__2386);
  not g__1591(w__70 ,w__2387);
  not g__1592(w__68 ,w__2389);
  not g__1593(w__69 ,w__2388);
  not g__1594(w__50 ,w__67);
  not g__1595(w__67 ,w__2384);
  not g__1596(w__49 ,w__71);
  not g__1597(w__71 ,w__2378);
  xor g__1598(w__2238 ,w__103 ,w__66);
  xor g__1599(w__2239 ,w__104 ,w__72);
  xor g__1600(w__2240 ,w__105 ,w__70);
  xor g__1601(w__2242 ,w__107 ,w__68);
  xor g__1602(w__2241 ,w__106 ,w__69);
  xnor g__1603(w__2256 ,w__168 ,w__2295);
  or g__1604(w__168 ,w__128 ,w__167);
  or g__1605(w__167 ,w__129 ,w__166);
  or g__1606(w__166 ,w__130 ,w__165);
  or g__1607(w__165 ,w__132 ,w__164);
  or g__1608(w__164 ,w__126 ,w__163);
  and g__1609(w__2250 ,w__163 ,w__162);
  or g__1610(w__163 ,w__127 ,w__161);
  or g__1611(w__162 ,w__110 ,w__160);
  not g__1612(w__161 ,w__160);
  or g__1613(w__160 ,w__145 ,w__159);
  xnor g__1614(w__2249 ,w__158 ,w__150);
  and g__1615(w__159 ,w__135 ,w__158);
  or g__1616(w__158 ,w__143 ,w__157);
  xnor g__1617(w__2248 ,w__156 ,w__149);
  and g__1618(w__157 ,w__137 ,w__156);
  or g__1619(w__156 ,w__141 ,w__155);
  xnor g__1620(w__2247 ,w__154 ,w__148);
  and g__1621(w__155 ,w__144 ,w__154);
  or g__1622(w__154 ,w__136 ,w__153);
  xnor g__1623(w__2246 ,w__152 ,w__147);
  and g__1624(w__153 ,w__134 ,w__152);
  xor g__1625(w__2245 ,w__139 ,w__146);
  or g__1626(w__152 ,w__138 ,w__151);
  nor g__1627(w__151 ,w__139 ,w__140);
  and g__1628(w__2244 ,w__139 ,w__142);
  xnor g__1629(w__150 ,w__116 ,in13[5]);
  xnor g__1630(w__149 ,w__113 ,in13[4]);
  xnor g__1631(w__148 ,w__122 ,in13[3]);
  xnor g__1632(w__147 ,w__119 ,in13[2]);
  xnor g__1633(w__146 ,w__124 ,in13[1]);
  and g__1634(w__145 ,in13[5] ,w__115);
  or g__1635(w__144 ,in13[3] ,w__121);
  and g__1636(w__143 ,in13[4] ,w__112);
  or g__1637(w__142 ,in13[0] ,w__109);
  and g__1638(w__141 ,in13[3] ,w__122);
  nor g__1639(w__140 ,in13[1] ,w__125);
  and g__1640(w__138 ,in13[1] ,w__124);
  or g__1641(w__137 ,in13[4] ,w__113);
  and g__1642(w__136 ,in13[2] ,w__118);
  or g__1643(w__135 ,in13[5] ,w__116);
  or g__1644(w__134 ,in13[2] ,w__119);
  or g__1645(w__139 ,w__133 ,w__131);
  not g__1646(w__133 ,in13[0]);
  not g__1647(w__125 ,w__123);
  not g__1648(w__124 ,w__123);
  not g__1649(w__123 ,w__2284);
  not g__1650(w__122 ,w__120);
  not g__1651(w__121 ,w__120);
  not g__1652(w__120 ,w__2286);
  not g__1653(w__119 ,w__117);
  not g__1654(w__118 ,w__117);
  not g__1655(w__117 ,w__2285);
  not g__1656(w__116 ,w__114);
  not g__1657(w__115 ,w__114);
  not g__1658(w__114 ,w__2288);
  not g__1659(w__113 ,w__111);
  not g__1660(w__112 ,w__111);
  not g__1661(w__111 ,w__2287);
  not g__1662(w__126 ,w__2290);
  not g__1663(w__132 ,w__2291);
  not g__1664(w__130 ,w__2292);
  not g__1665(w__128 ,w__2294);
  not g__1666(w__129 ,w__2293);
  not g__1667(w__110 ,w__127);
  not g__1668(w__127 ,w__2289);
  not g__1669(w__109 ,w__131);
  not g__1670(w__131 ,w__2283);
  xor g__1671(w__2251 ,w__163 ,w__126);
  xor g__1672(w__2252 ,w__164 ,w__132);
  xor g__1673(w__2253 ,w__165 ,w__130);
  xor g__1674(w__2255 ,w__167 ,w__128);
  xor g__1675(w__2254 ,w__166 ,w__129);
  xnor g__1676(w__2269 ,w__210 ,w__2295);
  or g__1677(w__210 ,w__183 ,w__209);
  or g__1678(w__209 ,w__180 ,w__208);
  or g__1679(w__208 ,w__184 ,w__207);
  or g__1680(w__207 ,w__181 ,w__206);
  or g__1681(w__206 ,w__182 ,w__205);
  or g__1682(w__205 ,w__179 ,w__204);
  or g__1683(w__204 ,w__177 ,w__203);
  or g__1684(w__203 ,w__185 ,w__201);
  and g__1685(w__2260 ,w__201 ,w__202);
  or g__1686(w__202 ,w__170 ,w__199);
  or g__1687(w__201 ,w__178 ,w__200);
  not g__1688(w__200 ,w__199);
  or g__1689(w__199 ,w__193 ,w__198);
  xnor g__1690(w__2259 ,w__197 ,w__194);
  and g__1691(w__198 ,w__189 ,w__197);
  xor g__1692(w__2258 ,w__190 ,w__195);
  or g__1693(w__197 ,w__188 ,w__196);
  nor g__1694(w__196 ,w__190 ,w__191);
  and g__1695(w__2257 ,w__190 ,w__192);
  xnor g__1696(w__195 ,w__175 ,in41[1]);
  xnor g__1697(w__194 ,w__173 ,in41[2]);
  and g__1698(w__193 ,w__172 ,in41[2]);
  or g__1699(w__192 ,w__169 ,in41[0]);
  nor g__1700(w__191 ,w__176 ,in41[1]);
  or g__1701(w__190 ,w__186 ,w__187);
  or g__1702(w__189 ,w__173 ,in41[2]);
  and g__1703(w__188 ,w__175 ,in41[1]);
  not g__1704(w__187 ,in41[0]);
  not g__1705(w__176 ,w__174);
  not g__1706(w__175 ,w__174);
  not g__1707(w__174 ,w__2284);
  not g__1708(w__173 ,w__171);
  not g__1709(w__172 ,w__171);
  not g__1710(w__171 ,w__2285);
  not g__1711(w__170 ,w__178);
  not g__1712(w__178 ,w__2286);
  not g__1713(w__177 ,w__2288);
  not g__1714(w__185 ,w__2287);
  not g__1715(w__181 ,w__2291);
  not g__1716(w__182 ,w__2290);
  not g__1717(w__183 ,w__2294);
  not g__1718(w__180 ,w__2293);
  not g__1719(w__184 ,w__2292);
  not g__1720(w__179 ,w__2289);
  not g__1721(w__169 ,w__186);
  not g__1722(w__186 ,w__2283);
  xor g__1723(w__2262 ,w__203 ,w__177);
  xor g__1724(w__2261 ,w__201 ,w__185);
  xor g__1725(w__2265 ,w__206 ,w__181);
  xor g__1726(w__2264 ,w__205 ,w__182);
  xor g__1727(w__2268 ,w__209 ,w__183);
  xor g__1728(w__2267 ,w__208 ,w__180);
  xor g__1729(w__2266 ,w__207 ,w__184);
  xor g__1730(w__2263 ,w__204 ,w__179);
  xnor g__1731(w__258 ,w__254 ,in24[8]);
  and g__1732(w__257 ,in24[8] ,w__253);
  and g__1733(w__256 ,w__255 ,w__254);
  or g__1734(w__255 ,in24[7] ,w__250);
  not g__1735(w__253 ,w__254);
  or g__1736(w__254 ,w__212 ,w__251);
  and g__1737(w__252 ,w__251 ,w__249);
  not g__1738(w__250 ,w__251);
  or g__1739(w__251 ,w__211 ,w__248);
  or g__1740(w__249 ,in24[6] ,w__247);
  not g__1741(w__248 ,w__247);
  or g__1742(w__247 ,w__218 ,w__245);
  xnor g__1743(w__246 ,w__244 ,w__229);
  and g__1744(w__245 ,w__225 ,w__244);
  or g__1745(w__244 ,w__224 ,w__242);
  xnor g__1746(w__243 ,w__241 ,w__228);
  and g__1747(w__242 ,w__222 ,w__241);
  or g__1748(w__241 ,w__221 ,w__239);
  xnor g__1749(w__240 ,w__238 ,w__227);
  and g__1750(w__239 ,w__226 ,w__238);
  or g__1751(w__238 ,w__216 ,w__236);
  xnor g__1752(w__237 ,w__234 ,w__231);
  and g__1753(w__236 ,w__215 ,w__234);
  xor g__1754(w__235 ,w__220 ,w__230);
  or g__1755(w__234 ,w__217 ,w__233);
  nor g__1756(w__233 ,w__220 ,w__223);
  and g__1757(w__232 ,w__220 ,w__219);
  xnor g__1758(w__231 ,in13[2] ,in24[2]);
  xnor g__1759(w__230 ,in13[1] ,in24[1]);
  xnor g__1760(w__229 ,in13[5] ,in24[5]);
  xnor g__1761(w__228 ,in13[4] ,in24[4]);
  xnor g__1762(w__227 ,in13[3] ,in24[3]);
  or g__1763(w__226 ,in13[3] ,in24[3]);
  or g__1764(w__225 ,in13[5] ,in24[5]);
  and g__1765(w__224 ,in13[4] ,in24[4]);
  nor g__1766(w__223 ,in13[1] ,in24[1]);
  or g__1767(w__222 ,in13[4] ,in24[4]);
  and g__1768(w__221 ,in13[3] ,in24[3]);
  or g__1769(w__219 ,in13[0] ,in24[0]);
  and g__1770(w__218 ,in13[5] ,in24[5]);
  and g__1771(w__217 ,in13[1] ,in24[1]);
  and g__1772(w__216 ,in13[2] ,in24[2]);
  or g__1773(w__215 ,in13[2] ,in24[2]);
  or g__1774(w__220 ,w__213 ,w__214);
  not g__1775(w__214 ,in24[0]);
  not g__1776(w__213 ,in13[0]);
  not g__1777(w__212 ,in24[7]);
  not g__1778(w__211 ,in24[6]);
  buf g__1779(w__2338 ,w__257);
  buf g__1780(w__2334 ,w__246);
  buf g__1781(w__2331 ,w__237);
  buf g__1782(w__2333 ,w__243);
  buf g__1783(w__2332 ,w__240);
  buf g__1784(w__2330 ,w__235);
  buf g__1785(w__2337 ,w__258);
  buf g__1786(w__2336 ,w__256);
  buf g__1787(w__2316 ,w__232);
  buf g__1788(w__2335 ,w__252);
  xnor g__1789(w__2315 ,w__356 ,w__331);
  or g__1790(w__356 ,w__313 ,w__355);
  xnor g__1791(w__2314 ,w__354 ,w__334);
  and g__1792(w__355 ,w__303 ,w__354);
  or g__1793(w__354 ,w__300 ,w__353);
  xnor g__1794(w__2313 ,w__352 ,w__333);
  and g__1795(w__353 ,w__315 ,w__352);
  or g__1796(w__352 ,w__316 ,w__351);
  xnor g__1797(w__2312 ,w__350 ,w__332);
  and g__1798(w__351 ,w__319 ,w__350);
  or g__1799(w__350 ,w__302 ,w__349);
  xnor g__1800(w__2311 ,w__348 ,w__327);
  and g__1801(w__349 ,w__320 ,w__348);
  or g__1802(w__348 ,w__318 ,w__347);
  xnor g__1803(w__2310 ,w__346 ,w__326);
  and g__1804(w__347 ,w__311 ,w__346);
  or g__1805(w__346 ,w__314 ,w__345);
  xnor g__1806(w__2309 ,w__344 ,w__325);
  and g__1807(w__345 ,w__299 ,w__344);
  or g__1808(w__344 ,w__306 ,w__343);
  xnor g__1809(w__2308 ,w__342 ,w__324);
  and g__1810(w__343 ,w__309 ,w__342);
  or g__1811(w__342 ,w__301 ,w__341);
  xnor g__1812(w__2307 ,w__340 ,w__330);
  and g__1813(w__341 ,w__305 ,w__340);
  or g__1814(w__340 ,w__308 ,w__339);
  xnor g__1815(w__2306 ,w__338 ,w__329);
  and g__1816(w__339 ,w__321 ,w__338);
  or g__1817(w__338 ,w__304 ,w__337);
  xnor g__1818(w__2305 ,w__336 ,w__323);
  and g__1819(w__337 ,w__322 ,w__336);
  xor g__1820(w__2304 ,w__310 ,w__328);
  or g__1821(w__336 ,w__317 ,w__335);
  and g__1822(w__2303 ,w__310 ,w__307);
  nor g__1823(w__335 ,w__310 ,w__312);
  xnor g__1824(w__334 ,w__264 ,in1[11]);
  xnor g__1825(w__333 ,w__261 ,in1[10]);
  xnor g__1826(w__332 ,w__266 ,in1[9]);
  xnor g__1827(w__331 ,w__268 ,in1[12]);
  xnor g__1828(w__330 ,w__281 ,in1[4]);
  xnor g__1829(w__329 ,w__290 ,in1[3]);
  xnor g__1830(w__328 ,w__286 ,in1[1]);
  xnor g__1831(w__327 ,w__284 ,in1[8]);
  xnor g__1832(w__326 ,w__272 ,in1[7]);
  xnor g__1833(w__325 ,w__275 ,in1[6]);
  xnor g__1834(w__324 ,w__278 ,in1[5]);
  xnor g__1835(w__323 ,w__293 ,in1[2]);
  or g__1836(w__322 ,in1[2] ,w__292);
  or g__1837(w__321 ,in1[3] ,w__289);
  or g__1838(w__320 ,in1[8] ,w__283);
  or g__1839(w__319 ,in1[9] ,w__261);
  and g__1840(w__318 ,in1[7] ,w__271);
  and g__1841(w__317 ,in1[1] ,w__286);
  and g__1842(w__316 ,in1[9] ,w__264);
  or g__1843(w__315 ,in1[10] ,w__266);
  and g__1844(w__314 ,in1[6] ,w__274);
  and g__1845(w__313 ,in1[11] ,w__268);
  nor g__1846(w__312 ,in1[1] ,w__287);
  or g__1847(w__311 ,in1[7] ,w__272);
  or g__1848(w__309 ,in1[5] ,w__277);
  and g__1849(w__308 ,in1[3] ,w__290);
  or g__1850(w__307 ,in1[0] ,w__269);
  and g__1851(w__306 ,in1[5] ,w__278);
  or g__1852(w__305 ,in1[4] ,w__280);
  and g__1853(w__304 ,in1[2] ,w__293);
  or g__1854(w__303 ,in1[11] ,w__260);
  and g__1855(w__302 ,in1[8] ,w__284);
  and g__1856(w__301 ,in1[4] ,w__281);
  and g__1857(w__300 ,in1[10] ,w__263);
  or g__1858(w__299 ,in1[6] ,w__275);
  or g__1859(w__310 ,w__298 ,w__297);
  not g__1860(w__298 ,in1[0]);
  not g__1861(w__296 ,w__294);
  not g__1862(w__295 ,w__294);
  not g__1863(w__294 ,w__2338);
  not g__1864(w__293 ,w__291);
  not g__1865(w__292 ,w__291);
  not g__1866(w__291 ,w__2331);
  not g__1867(w__290 ,w__288);
  not g__1868(w__289 ,w__288);
  not g__1869(w__288 ,w__2332);
  not g__1870(w__287 ,w__285);
  not g__1871(w__286 ,w__285);
  not g__1872(w__285 ,w__2330);
  not g__1873(w__284 ,w__282);
  not g__1874(w__283 ,w__282);
  not g__1875(w__282 ,w__2337);
  not g__1876(w__281 ,w__279);
  not g__1877(w__280 ,w__279);
  not g__1878(w__279 ,w__2333);
  not g__1879(w__278 ,w__276);
  not g__1880(w__277 ,w__276);
  not g__1881(w__276 ,w__2334);
  not g__1882(w__275 ,w__273);
  not g__1883(w__274 ,w__273);
  not g__1884(w__273 ,w__2335);
  not g__1885(w__272 ,w__270);
  not g__1886(w__271 ,w__270);
  not g__1887(w__270 ,w__2336);
  not g__1888(w__269 ,w__297);
  not g__1889(w__297 ,w__2316);
  not g__1890(w__268 ,w__267);
  not g__1891(w__267 ,w__296);
  not g__1892(w__266 ,w__265);
  not g__1893(w__265 ,w__295);
  not g__1894(w__264 ,w__262);
  not g__1895(w__263 ,w__262);
  not g__1896(w__262 ,w__296);
  not g__1897(w__261 ,w__259);
  not g__1898(w__260 ,w__259);
  not g__1899(w__259 ,w__295);
  xnor g__1900(w__430 ,w__429 ,w__388);
  or g__1901(w__429 ,w__358 ,w__427);
  xnor g__1902(w__428 ,w__426 ,w__393);
  and g__1903(w__427 ,w__360 ,w__426);
  or g__1904(w__426 ,w__375 ,w__424);
  xnor g__1905(w__425 ,w__423 ,w__392);
  and g__1906(w__424 ,w__376 ,w__423);
  or g__1907(w__423 ,w__374 ,w__421);
  xnor g__1908(w__422 ,w__420 ,w__391);
  and g__1909(w__421 ,w__377 ,w__420);
  or g__1910(w__420 ,w__368 ,w__418);
  xnor g__1911(w__419 ,w__417 ,w__390);
  and g__1912(w__418 ,w__366 ,w__417);
  or g__1913(w__417 ,w__370 ,w__415);
  xnor g__1914(w__416 ,w__414 ,w__389);
  and g__1915(w__415 ,w__378 ,w__414);
  or g__1916(w__414 ,w__371 ,w__412);
  xnor g__1917(w__413 ,w__411 ,w__384);
  and g__1918(w__412 ,w__357 ,w__411);
  or g__1919(w__411 ,w__361 ,w__409);
  xnor g__1920(w__410 ,w__408 ,w__383);
  and g__1921(w__409 ,w__373 ,w__408);
  or g__1922(w__408 ,w__379 ,w__406);
  xnor g__1923(w__407 ,w__405 ,w__382);
  and g__1924(w__406 ,w__363 ,w__405);
  or g__1925(w__405 ,w__367 ,w__403);
  xnor g__1926(w__404 ,w__402 ,w__387);
  and g__1927(w__403 ,w__364 ,w__402);
  or g__1928(w__402 ,w__369 ,w__400);
  xnor g__1929(w__401 ,w__399 ,w__381);
  and g__1930(w__400 ,w__362 ,w__399);
  or g__1931(w__399 ,w__365 ,w__397);
  xnor g__1932(w__398 ,w__395 ,w__386);
  and g__1933(w__397 ,w__372 ,w__395);
  xnor g__1934(w__396 ,w__385 ,in22);
  or g__1935(w__395 ,w__359 ,w__394);
  and g__1936(w__394 ,in1[0] ,w__380);
  xnor g__1937(w__393 ,in1[11] ,in22);
  xnor g__1938(w__392 ,in1[10] ,in22);
  xnor g__1939(w__391 ,in1[9] ,in22);
  xnor g__1940(w__390 ,in1[8] ,in22);
  xnor g__1941(w__389 ,in1[7] ,in22);
  xnor g__1942(w__388 ,in1[12] ,in22);
  xnor g__1943(w__387 ,w__2299 ,in1[3]);
  xnor g__1944(w__386 ,w__2297 ,in1[1]);
  xnor g__1945(w__385 ,w__2296 ,in1[0]);
  xnor g__1946(w__384 ,w__2302 ,in1[6]);
  xnor g__1947(w__383 ,w__2301 ,in1[5]);
  xnor g__1948(w__382 ,w__2300 ,in1[4]);
  xnor g__1949(w__381 ,w__2298 ,in1[2]);
  or g__1950(w__380 ,w__2296 ,in22);
  and g__1951(w__379 ,in1[4] ,w__2300);
  or g__1952(w__378 ,in1[7] ,in22);
  or g__1953(w__377 ,in1[9] ,in22);
  or g__1954(w__376 ,in1[10] ,in22);
  and g__1955(w__375 ,in1[10] ,in22);
  and g__1956(w__374 ,in1[9] ,in22);
  or g__1957(w__373 ,in1[5] ,w__2301);
  or g__1958(w__372 ,in1[1] ,w__2297);
  and g__1959(w__371 ,in1[6] ,w__2302);
  and g__1960(w__370 ,in1[7] ,in22);
  and g__1961(w__369 ,in1[2] ,w__2298);
  and g__1962(w__368 ,in1[8] ,in22);
  and g__1963(w__367 ,in1[3] ,w__2299);
  or g__1964(w__366 ,in1[8] ,in22);
  and g__1965(w__365 ,in1[1] ,w__2297);
  or g__1966(w__364 ,in1[3] ,w__2299);
  or g__1967(w__363 ,in1[4] ,w__2300);
  or g__1968(w__362 ,in1[2] ,w__2298);
  and g__1969(w__361 ,in1[5] ,w__2301);
  or g__1970(w__360 ,in1[11] ,in22);
  and g__1971(w__359 ,w__2296 ,in22);
  and g__1972(w__358 ,in1[11] ,in22);
  or g__1973(w__357 ,in1[6] ,w__2302);
  buf g__1974(w__2295 ,w__430);
  buf g__1975(w__2294 ,w__428);
  buf g__1976(w__2284 ,w__398);
  buf g__1977(w__2285 ,w__401);
  buf g__1978(w__2286 ,w__404);
  buf g__1979(w__2287 ,w__407);
  buf g__1980(w__2292 ,w__422);
  buf g__1981(w__2289 ,w__413);
  buf g__1982(w__2290 ,w__416);
  buf g__1983(w__2291 ,w__419);
  buf g__1984(w__2288 ,w__410);
  buf g__1985(w__2293 ,w__425);
  buf g__1986(w__2283 ,w__396);
  xnor g__1987(w__504 ,w__503 ,w__462);
  or g__1988(w__503 ,w__432 ,w__501);
  xnor g__1989(w__502 ,w__500 ,w__467);
  and g__1990(w__501 ,w__434 ,w__500);
  or g__1991(w__500 ,w__449 ,w__498);
  xnor g__1992(w__499 ,w__497 ,w__466);
  and g__1993(w__498 ,w__450 ,w__497);
  or g__1994(w__497 ,w__448 ,w__495);
  xnor g__1995(w__496 ,w__494 ,w__465);
  and g__1996(w__495 ,w__451 ,w__494);
  or g__1997(w__494 ,w__442 ,w__492);
  xnor g__1998(w__493 ,w__491 ,w__464);
  and g__1999(w__492 ,w__440 ,w__491);
  or g__2000(w__491 ,w__444 ,w__489);
  xnor g__2001(w__490 ,w__488 ,w__463);
  and g__2002(w__489 ,w__452 ,w__488);
  or g__2003(w__488 ,w__445 ,w__486);
  xnor g__2004(w__487 ,w__485 ,w__458);
  and g__2005(w__486 ,w__431 ,w__485);
  or g__2006(w__485 ,w__435 ,w__483);
  xnor g__2007(w__484 ,w__482 ,w__457);
  and g__2008(w__483 ,w__447 ,w__482);
  or g__2009(w__482 ,w__453 ,w__480);
  xnor g__2010(w__481 ,w__479 ,w__456);
  and g__2011(w__480 ,w__437 ,w__479);
  or g__2012(w__479 ,w__441 ,w__477);
  xnor g__2013(w__478 ,w__476 ,w__461);
  and g__2014(w__477 ,w__438 ,w__476);
  or g__2015(w__476 ,w__443 ,w__474);
  xnor g__2016(w__475 ,w__473 ,w__455);
  and g__2017(w__474 ,w__436 ,w__473);
  or g__2018(w__473 ,w__439 ,w__471);
  xnor g__2019(w__472 ,w__469 ,w__460);
  and g__2020(w__471 ,w__446 ,w__469);
  xnor g__2021(w__470 ,w__459 ,in3);
  or g__2022(w__469 ,w__433 ,w__468);
  and g__2023(w__468 ,in1[0] ,w__454);
  xnor g__2024(w__467 ,in1[11] ,in3);
  xnor g__2025(w__466 ,in1[10] ,in3);
  xnor g__2026(w__465 ,in1[9] ,in3);
  xnor g__2027(w__464 ,in1[8] ,in3);
  xnor g__2028(w__463 ,in1[7] ,in3);
  xnor g__2029(w__462 ,in1[12] ,in3);
  xnor g__2030(w__461 ,w__2394 ,in1[3]);
  xnor g__2031(w__460 ,w__2392 ,in1[1]);
  xnor g__2032(w__459 ,w__2391 ,in1[0]);
  xnor g__2033(w__458 ,w__2397 ,in1[6]);
  xnor g__2034(w__457 ,w__2396 ,in1[5]);
  xnor g__2035(w__456 ,w__2395 ,in1[4]);
  xnor g__2036(w__455 ,w__2393 ,in1[2]);
  or g__2037(w__454 ,w__2391 ,in3);
  and g__2038(w__453 ,in1[4] ,w__2395);
  or g__2039(w__452 ,in1[7] ,in3);
  or g__2040(w__451 ,in1[9] ,in3);
  or g__2041(w__450 ,in1[10] ,in3);
  and g__2042(w__449 ,in1[10] ,in3);
  and g__2043(w__448 ,in1[9] ,in3);
  or g__2044(w__447 ,in1[5] ,w__2396);
  or g__2045(w__446 ,in1[1] ,w__2392);
  and g__2046(w__445 ,in1[6] ,w__2397);
  and g__2047(w__444 ,in1[7] ,in3);
  and g__2048(w__443 ,in1[2] ,w__2393);
  and g__2049(w__442 ,in1[8] ,in3);
  and g__2050(w__441 ,in1[3] ,w__2394);
  or g__2051(w__440 ,in1[8] ,in3);
  and g__2052(w__439 ,in1[1] ,w__2392);
  or g__2053(w__438 ,in1[3] ,w__2394);
  or g__2054(w__437 ,in1[4] ,w__2395);
  or g__2055(w__436 ,in1[2] ,w__2393);
  and g__2056(w__435 ,in1[5] ,w__2396);
  or g__2057(w__434 ,in1[11] ,in3);
  and g__2058(w__433 ,w__2391 ,in3);
  and g__2059(w__432 ,in1[11] ,in3);
  or g__2060(w__431 ,in1[6] ,w__2397);
  buf g__2061(w__2390 ,w__504);
  buf g__2062(w__2389 ,w__502);
  buf g__2063(w__2379 ,w__472);
  buf g__2064(w__2380 ,w__475);
  buf g__2065(w__2381 ,w__478);
  buf g__2066(w__2382 ,w__481);
  buf g__2067(w__2387 ,w__496);
  buf g__2068(w__2384 ,w__487);
  buf g__2069(w__2385 ,w__490);
  buf g__2070(w__2386 ,w__493);
  buf g__2071(w__2383 ,w__484);
  buf g__2072(w__2388 ,w__499);
  buf g__2073(w__2378 ,w__470);
  xnor g__2074(w__2423 ,w__550 ,w__614);
  nor g__2075(w__614 ,w__537 ,w__613);
  xnor g__2076(w__2422 ,w__612 ,w__542);
  nor g__2077(w__613 ,w__538 ,w__612);
  and g__2078(w__612 ,w__533 ,w__611);
  xnor g__2079(w__2421 ,w__610 ,w__552);
  or g__2080(w__611 ,w__534 ,w__610);
  and g__2081(w__610 ,w__536 ,w__609);
  xnor g__2082(w__2420 ,w__608 ,w__551);
  or g__2083(w__609 ,w__535 ,w__608);
  and g__2084(w__608 ,w__555 ,w__607);
  or g__2085(w__607 ,w__554 ,w__606);
  and g__2086(w__606 ,w__559 ,w__605);
  or g__2087(w__605 ,w__565 ,w__604);
  and g__2088(w__604 ,w__564 ,w__603);
  or g__2089(w__603 ,w__566 ,w__602);
  and g__2090(w__602 ,w__563 ,w__601);
  xnor g__2091(w__2416 ,w__599 ,w__572);
  or g__2092(w__601 ,w__561 ,w__600);
  not g__2093(w__600 ,w__599);
  or g__2094(w__599 ,w__560 ,w__598);
  xnor g__2095(w__2415 ,w__597 ,w__573);
  and g__2096(w__598 ,w__567 ,w__597);
  or g__2097(w__597 ,w__583 ,w__596);
  xnor g__2098(w__2414 ,w__595 ,w__584);
  nor g__2099(w__596 ,w__582 ,w__595);
  and g__2100(w__595 ,w__588 ,w__594);
  xnor g__2101(w__2413 ,w__592 ,w__589);
  or g__2102(w__594 ,w__587 ,w__593);
  xnor g__2103(w__2412 ,w__581 ,w__590);
  not g__2104(w__593 ,w__592);
  or g__2105(w__592 ,w__586 ,w__591);
  nor g__2106(w__591 ,w__581 ,w__585);
  xnor g__2107(w__590 ,w__531 ,w__576);
  xnor g__2108(w__589 ,w__571 ,w__580);
  xor g__2109(w__2411 ,w__578 ,w__2424);
  or g__2110(w__588 ,w__570 ,w__579);
  nor g__2111(w__587 ,w__571 ,w__580);
  nor g__2112(w__586 ,w__531 ,w__577);
  and g__2113(w__585 ,w__531 ,w__577);
  xnor g__2114(w__584 ,w__544 ,w__568);
  nor g__2115(w__583 ,w__544 ,w__569);
  and g__2116(w__582 ,w__544 ,w__569);
  and g__2117(w__581 ,w__532 ,w__562);
  not g__2118(w__579 ,w__580);
  xnor g__2119(w__580 ,w__541 ,w__2426);
  xnor g__2120(w__578 ,w__549 ,in27);
  not g__2121(w__577 ,w__576);
  xnor g__2122(w__576 ,w__543 ,w__2425);
  xnor g__2123(w__575 ,w__528 ,w__557);
  xnor g__2124(w__574 ,w__530 ,w__547);
  xnor g__2125(w__573 ,w__527 ,w__546);
  xnor g__2126(w__572 ,w__529 ,w__548);
  not g__2127(w__570 ,w__571);
  not g__2128(w__569 ,w__568);
  or g__2129(w__567 ,w__526 ,w__545);
  and g__2130(w__566 ,w__530 ,w__547);
  and g__2131(w__565 ,w__528 ,w__557);
  or g__2132(w__564 ,w__530 ,w__547);
  or g__2133(w__571 ,w__524 ,w__553);
  or g__2134(w__568 ,w__539 ,w__556);
  or g__2135(w__563 ,w__529 ,w__548);
  or g__2136(w__562 ,w__522 ,w__549);
  and g__2137(w__561 ,w__529 ,w__548);
  nor g__2138(w__560 ,w__527 ,w__546);
  or g__2139(w__559 ,w__528 ,w__557);
  xnor g__2140(w__558 ,w__540 ,in1[8]);
  and g__2141(w__556 ,w__2426 ,w__523);
  or g__2142(w__555 ,in1[8] ,w__540);
  and g__2143(w__554 ,in1[8] ,w__540);
  and g__2144(w__553 ,in25[1] ,w__525);
  xnor g__2145(w__552 ,in1[10] ,in1[9]);
  xnor g__2146(w__551 ,in1[9] ,in1[8]);
  xnor g__2147(w__550 ,in1[12] ,in1[11]);
  xnor g__2148(w__557 ,in1[7] ,in27);
  not g__2149(w__545 ,w__546);
  xnor g__2150(w__543 ,in25[1] ,in1[1]);
  xnor g__2151(w__542 ,in1[11] ,in1[10]);
  xnor g__2152(w__541 ,in25[2] ,in1[2]);
  xnor g__2153(w__549 ,in25[0] ,in1[0]);
  xnor g__2154(w__548 ,w__2429 ,in1[5]);
  xnor g__2155(w__547 ,w__2430 ,in1[6]);
  xnor g__2156(w__546 ,w__2428 ,in1[4]);
  xnor g__2157(w__544 ,w__2427 ,in1[3]);
  and g__2158(w__539 ,in25[2] ,in1[2]);
  nor g__2159(w__538 ,w__507 ,in1[10]);
  nor g__2160(w__537 ,w__505 ,in1[11]);
  or g__2161(w__536 ,w__515 ,in1[9]);
  nor g__2162(w__535 ,w__506 ,in1[8]);
  nor g__2163(w__534 ,w__505 ,in1[9]);
  or g__2164(w__533 ,w__506 ,in1[10]);
  or g__2165(w__532 ,w__517 ,w__516);
  and g__2166(w__540 ,in27 ,w__514);
  not g__2167(w__526 ,w__527);
  or g__2168(w__525 ,in1[1] ,w__2425);
  and g__2169(w__524 ,in1[1] ,w__2425);
  or g__2170(w__523 ,in25[2] ,in1[2]);
  nor g__2171(w__522 ,w__2424 ,in27);
  or g__2172(w__531 ,w__519 ,w__509);
  or g__2173(w__530 ,w__518 ,w__508);
  or g__2174(w__529 ,w__513 ,w__510);
  or g__2175(w__528 ,w__521 ,w__512);
  or g__2176(w__527 ,w__520 ,w__511);
  not g__2177(w__521 ,in1[6]);
  not g__2178(w__520 ,in1[3]);
  not g__2179(w__519 ,in25[0]);
  not g__2180(w__518 ,in1[5]);
  not g__2181(w__517 ,w__2424);
  not g__2182(w__516 ,in27);
  not g__2183(w__515 ,in1[8]);
  not g__2184(w__514 ,in1[7]);
  not g__2185(w__513 ,in1[4]);
  not g__2186(w__512 ,w__2430);
  not g__2187(w__511 ,w__2427);
  not g__2188(w__510 ,w__2428);
  not g__2189(w__509 ,in1[0]);
  not g__2190(w__508 ,w__2429);
  not g__2191(w__507 ,in1[11]);
  not g__2192(w__506 ,in1[9]);
  not g__2193(w__505 ,in1[10]);
  xor g__2194(w__2419 ,w__606 ,w__558);
  xor g__2195(w__2418 ,w__604 ,w__575);
  xor g__2196(w__2417 ,w__602 ,w__574);
  xnor g__2197(w__2324 ,w__637 ,w__2403);
  xnor g__2198(w__2325 ,w__636 ,w__2402);
  xnor g__2199(w__2326 ,w__635 ,w__2401);
  xnor g__2200(w__2327 ,w__634 ,w__2400);
  xnor g__2201(w__2328 ,w__633 ,w__2399);
  or g__2202(w__2230 ,w__627 ,w__638);
  or g__2203(w__2232 ,w__632 ,w__641);
  or g__2204(w__2323 ,w__628 ,w__642);
  or g__2205(w__2233 ,w__625 ,w__640);
  or g__2206(w__2231 ,w__623 ,w__639);
  xor g__2207(w__2319 ,w__616 ,w__2408);
  and g__2208(w__642 ,w__2403 ,w__630);
  and g__2209(w__641 ,w__2400 ,w__631);
  and g__2210(w__640 ,w__2399 ,w__626);
  and g__2211(w__639 ,w__2401 ,w__629);
  xor g__2212(w__2229 ,w__2436 ,w__2404);
  xor g__2213(w__2318 ,w__619 ,w__2409);
  xor g__2214(w__2329 ,w__2398 ,in13[0]);
  and g__2215(w__638 ,w__2402 ,w__624);
  xor g__2216(w__2317 ,w__619 ,w__2410);
  xor g__2217(w__2322 ,w__2437 ,w__2405);
  xor g__2218(w__2321 ,w__2438 ,w__2406);
  xor g__2219(w__2320 ,w__621 ,w__2407);
  xnor g__2220(w__637 ,w__2435 ,in13[5]);
  xnor g__2221(w__636 ,w__2434 ,in13[4]);
  xnor g__2222(w__635 ,w__2433 ,in13[3]);
  xnor g__2223(w__634 ,w__2432 ,in13[2]);
  xnor g__2224(w__633 ,w__2431 ,in13[1]);
  and g__2225(w__632 ,in13[2] ,w__2432);
  or g__2226(w__631 ,in13[2] ,w__2432);
  or g__2227(w__630 ,in13[5] ,w__2435);
  or g__2228(w__629 ,in13[3] ,w__2433);
  and g__2229(w__628 ,in13[5] ,w__2435);
  and g__2230(w__2224 ,w__618 ,w__2408);
  and g__2231(w__2226 ,w__2438 ,w__2406);
  and g__2232(w__2223 ,w__616 ,w__2409);
  and g__2233(w__627 ,in13[4] ,w__2434);
  or g__2234(w__626 ,in13[1] ,w__2431);
  and g__2235(w__625 ,in13[1] ,w__2431);
  or g__2236(w__624 ,in13[4] ,w__2434);
  and g__2237(w__623 ,in13[3] ,w__2433);
  and g__2238(w__2225 ,w__618 ,w__2407);
  and g__2239(w__2228 ,w__2436 ,w__2404);
  and g__2240(w__2227 ,w__2437 ,w__2405);
  and g__2241(w__2234 ,in13[0] ,w__2398);
  not g__2242(w__622 ,w__620);
  not g__2243(w__621 ,w__620);
  not g__2244(w__620 ,w__2439);
  not g__2245(w__619 ,w__617);
  not g__2246(w__618 ,w__617);
  not g__2247(w__617 ,w__622);
  not g__2248(w__616 ,w__615);
  not g__2249(w__615 ,w__621);
  xnor g__2250(w__2282 ,w__767 ,w__2295);
  or g__2251(w__767 ,w__687 ,w__766);
  and g__2252(w__766 ,w__712 ,w__765);
  xnor g__2253(w__2280 ,w__764 ,w__714);
  or g__2254(w__765 ,w__653 ,w__764);
  and g__2255(w__764 ,w__717 ,w__763);
  or g__2256(w__763 ,w__718 ,w__762);
  and g__2257(w__762 ,w__715 ,w__761);
  or g__2258(w__761 ,w__725 ,w__760);
  and g__2259(w__760 ,w__722 ,w__759);
  or g__2260(w__759 ,w__724 ,w__758);
  and g__2261(w__758 ,w__727 ,w__757);
  or g__2262(w__757 ,w__720 ,w__756);
  and g__2263(w__756 ,w__719 ,w__755);
  xnor g__2264(w__2275 ,w__753 ,w__731);
  or g__2265(w__755 ,w__716 ,w__754);
  not g__2266(w__754 ,w__753);
  or g__2267(w__753 ,w__739 ,w__752);
  xor g__2268(w__2274 ,w__751 ,w__740);
  and g__2269(w__752 ,w__738 ,w__751);
  or g__2270(w__751 ,w__745 ,w__750);
  xnor g__2271(w__2273 ,w__749 ,w__746);
  and g__2272(w__750 ,w__744 ,w__749);
  xor g__2273(w__2272 ,w__741 ,w__747);
  or g__2274(w__749 ,w__743 ,w__748);
  and g__2275(w__748 ,w__742 ,w__741);
  xnor g__2276(w__747 ,w__698 ,w__644);
  xnor g__2277(w__746 ,w__730 ,w__645);
  xor g__2278(w__2271 ,w__721 ,w__652);
  and g__2279(w__745 ,w__730 ,w__645);
  or g__2280(w__744 ,w__730 ,w__645);
  nor g__2281(w__743 ,w__698 ,w__736);
  or g__2282(w__742 ,w__697 ,w__644);
  or g__2283(w__741 ,w__723 ,w__737);
  xnor g__2284(w__740 ,w__648 ,w__729);
  nor g__2285(w__739 ,w__648 ,w__728);
  or g__2286(w__738 ,w__713 ,w__729);
  and g__2287(w__737 ,w__721 ,w__726);
  not g__2288(w__736 ,w__644);
  xnor g__2289(w__735 ,w__646 ,w__695);
  xnor g__2290(w__734 ,w__650 ,w__704);
  xnor g__2291(w__733 ,w__643 ,w__693);
  xnor g__2292(w__732 ,w__647 ,w__694);
  xnor g__2293(w__731 ,w__649 ,w__696);
  not g__2294(w__728 ,w__729);
  or g__2295(w__727 ,w__694 ,w__647);
  or g__2296(w__726 ,w__664 ,w__708);
  and g__2297(w__725 ,w__704 ,w__650);
  and g__2298(w__724 ,w__695 ,w__646);
  nor g__2299(w__723 ,w__690 ,w__651);
  or g__2300(w__722 ,w__695 ,w__646);
  or g__2301(w__730 ,w__702 ,w__711);
  or g__2302(w__729 ,w__699 ,w__709);
  and g__2303(w__720 ,w__694 ,w__647);
  or g__2304(w__719 ,w__696 ,w__649);
  and g__2305(w__718 ,w__693 ,w__643);
  or g__2306(w__717 ,w__693 ,w__643);
  and g__2307(w__716 ,w__696 ,w__649);
  or g__2308(w__715 ,w__704 ,w__650);
  xnor g__2309(w__714 ,w__703 ,w__658);
  or g__2310(w__721 ,w__691 ,w__710);
  not g__2311(w__713 ,w__648);
  or g__2312(w__712 ,w__688 ,w__703);
  and g__2313(w__711 ,in23[2] ,w__692);
  and g__2314(w__710 ,in23[0] ,w__701);
  and g__2315(w__709 ,in23[3] ,w__700);
  not g__2316(w__708 ,w__651);
  xnor g__2317(w__707 ,w__672 ,in23[2]);
  xnor g__2318(w__706 ,w__669 ,in23[3]);
  xnor g__2319(w__705 ,w__656 ,in23[0]);
  and g__2320(w__702 ,w__671 ,w__660);
  or g__2321(w__701 ,w__666 ,w__655);
  or g__2322(w__700 ,w__668 ,w__662);
  and g__2323(w__699 ,w__669 ,w__662);
  or g__2324(w__704 ,w__678 ,w__684);
  or g__2325(w__703 ,w__682 ,w__676);
  not g__2326(w__697 ,w__698);
  or g__2327(w__692 ,w__672 ,w__660);
  and g__2328(w__691 ,w__666 ,w__656);
  or g__2329(w__698 ,w__675 ,w__689);
  or g__2330(w__696 ,w__677 ,w__674);
  or g__2331(w__695 ,w__683 ,w__679);
  or g__2332(w__694 ,w__681 ,w__685);
  or g__2333(w__693 ,w__686 ,w__680);
  not g__2334(w__690 ,w__664);
  not g__2335(w__689 ,in23[1]);
  not g__2336(w__688 ,w__658);
  not g__2337(w__682 ,w__673);
  not g__2338(w__672 ,w__670);
  not g__2339(w__671 ,w__670);
  not g__2340(w__670 ,w__2331);
  not g__2341(w__669 ,w__667);
  not g__2342(w__668 ,w__667);
  not g__2343(w__667 ,w__2332);
  not g__2344(w__666 ,w__665);
  not g__2345(w__665 ,w__2316);
  not g__2346(w__664 ,w__663);
  not g__2347(w__663 ,w__2284);
  not g__2348(w__675 ,w__2330);
  not g__2349(w__686 ,w__2337);
  not g__2350(w__681 ,w__2334);
  not g__2351(w__677 ,w__2333);
  not g__2352(w__683 ,w__2335);
  not g__2353(w__678 ,w__2336);
  not g__2354(w__662 ,w__661);
  not g__2355(w__661 ,w__2286);
  not g__2356(w__660 ,w__659);
  not g__2357(w__659 ,w__2285);
  not g__2358(w__685 ,w__2288);
  not g__2359(w__674 ,w__2287);
  not g__2360(w__658 ,w__657);
  not g__2361(w__657 ,w__2293);
  not g__2362(w__656 ,w__654);
  not g__2363(w__655 ,w__654);
  not g__2364(w__654 ,w__2283);
  not g__2365(w__687 ,w__2294);
  not g__2366(w__684 ,w__2290);
  not g__2367(w__680 ,w__2291);
  not g__2368(w__676 ,w__2292);
  not g__2369(w__679 ,w__2289);
  buf g__2370(w__673 ,w__2338);
  xor g__2371(w__2279 ,w__762 ,w__733);
  xor g__2372(w__2278 ,w__760 ,w__734);
  xor g__2373(w__2277 ,w__758 ,w__735);
  xor g__2374(w__2276 ,w__756 ,w__732);
  and g__2375(w__653 ,w__657 ,w__703);
  xor g__2376(w__2270 ,w__705 ,w__665);
  xor g__2377(w__652 ,w__651 ,w__663);
  xor g__2378(w__651 ,w__675 ,in23[1]);
  xnor g__2379(w__650 ,w__686 ,w__680);
  xnor g__2380(w__649 ,w__681 ,w__685);
  xnor g__2381(w__648 ,w__677 ,w__674);
  xnor g__2382(w__647 ,w__683 ,w__679);
  xnor g__2383(w__646 ,w__678 ,w__684);
  xor g__2384(w__645 ,w__706 ,w__661);
  xor g__2385(w__644 ,w__707 ,w__659);
  xor g__2386(w__2281 ,w__766 ,w__687);
  xor g__2387(w__643 ,w__673 ,w__676);
  xnor g__2388(w__2490 ,w__775 ,w__776);
  xnor g__2389(w__2491 ,w__778 ,w__777);
  xnor g__2390(w__2492 ,w__780 ,w__779);
  xnor g__2391(w__2493 ,w__774 ,w__773);
  or g__2392(w__2528 ,w__926 ,w__938);
  or g__2393(w__2532 ,w__905 ,w__937);
  or g__2394(w__2529 ,w__931 ,w__939);
  or g__2395(w__2530 ,w__928 ,w__936);
  or g__2396(w__2531 ,w__933 ,w__935);
  xnor g__2397(w__2485 ,w__923 ,w__800);
  xnor g__2398(w__2486 ,w__924 ,w__802);
  xnor g__2399(w__2487 ,w__922 ,w__804);
  xnor g__2400(w__2488 ,w__921 ,w__806);
  xnor g__2401(w__2494 ,w__934 ,w__907);
  xor g__2402(w__2489 ,w__913 ,w__781);
  and g__2403(w__939 ,w__930 ,w__778);
  and g__2404(w__938 ,w__932 ,w__775);
  nor g__2405(w__937 ,w__904 ,w__934);
  or g__2406(w__2527 ,w__916 ,w__927);
  and g__2407(w__936 ,w__929 ,w__780);
  and g__2408(w__935 ,w__925 ,w__774);
  xnor g__2409(w__2484 ,w__883 ,w__908);
  or g__2410(w__2524 ,w__890 ,w__914);
  and g__2411(w__933 ,w__823 ,w__911);
  or g__2412(w__932 ,w__831 ,w__919);
  or g__2413(w__2526 ,w__901 ,w__918);
  and g__2414(w__931 ,w__833 ,w__920);
  or g__2415(w__930 ,w__833 ,w__920);
  or g__2416(w__2523 ,w__900 ,w__910);
  or g__2417(w__929 ,w__837 ,w__912);
  or g__2418(w__2525 ,w__895 ,w__909);
  and g__2419(w__928 ,w__837 ,w__912);
  and g__2420(w__927 ,w__913 ,w__917);
  and g__2421(w__934 ,w__879 ,w__915);
  and g__2422(w__926 ,w__831 ,w__919);
  or g__2423(w__925 ,w__823 ,w__911);
  xor g__2424(w__2495 ,w__768 ,w__884);
  xnor g__2425(w__924 ,w__892 ,w__880);
  xnor g__2426(w__923 ,w__772 ,w__874);
  xnor g__2427(w__922 ,w__770 ,w__873);
  xnor g__2428(w__921 ,w__769 ,w__882);
  nor g__2429(w__918 ,w__898 ,w__769);
  or g__2430(w__917 ,w__843 ,w__891);
  nor g__2431(w__916 ,w__856 ,w__771);
  or g__2432(w__915 ,w__782 ,w__768);
  nor g__2433(w__914 ,w__899 ,w__892);
  or g__2434(w__920 ,w__867 ,w__897);
  or g__2435(w__919 ,w__878 ,w__903);
  nor g__2436(w__910 ,w__902 ,w__772);
  nor g__2437(w__909 ,w__893 ,w__770);
  xnor g__2438(w__908 ,w__866 ,w__2217);
  xnor g__2439(w__907 ,w__881 ,w__798);
  or g__2440(w__913 ,w__875 ,w__894);
  or g__2441(w__912 ,w__869 ,w__896);
  or g__2442(w__911 ,w__872 ,w__906);
  and g__2443(w__906 ,w__792 ,w__877);
  nor g__2444(w__905 ,w__865 ,w__881);
  and g__2445(w__904 ,w__865 ,w__881);
  and g__2446(w__903 ,w__794 ,w__870);
  and g__2447(w__902 ,w__860 ,w__874);
  nor g__2448(w__901 ,w__862 ,w__882);
  nor g__2449(w__900 ,w__860 ,w__874);
  and g__2450(w__899 ,w__857 ,w__880);
  and g__2451(w__898 ,w__862 ,w__882);
  and g__2452(w__897 ,w__790 ,w__876);
  and g__2453(w__896 ,w__786 ,w__868);
  nor g__2454(w__895 ,w__863 ,w__873);
  and g__2455(w__894 ,w__796 ,w__871);
  and g__2456(w__893 ,w__863 ,w__873);
  not g__2457(w__891 ,w__771);
  nor g__2458(w__890 ,w__857 ,w__880);
  xor g__2459(w__2496 ,w__784 ,w__788);
  xnor g__2460(w__889 ,w__812 ,w__794);
  xnor g__2461(w__888 ,w__821 ,w__786);
  xnor g__2462(w__887 ,w__815 ,w__790);
  xnor g__2463(w__886 ,w__818 ,w__792);
  xnor g__2464(w__885 ,w__809 ,w__796);
  xnor g__2465(w__884 ,w__825 ,w__845);
  xnor g__2466(w__883 ,w__2364 ,w__2351);
  xnor g__2467(w__892 ,w__2362 ,w__2349);
  or g__2468(w__879 ,w__864 ,w__861);
  and g__2469(w__878 ,w__835 ,w__811);
  or g__2470(w__877 ,w__841 ,w__817);
  or g__2471(w__876 ,w__839 ,w__814);
  and g__2472(w__875 ,w__829 ,w__808);
  and g__2473(w__2534 ,w__784 ,w__788);
  or g__2474(w__882 ,w__854 ,w__855);
  or g__2475(w__881 ,w__852 ,w__850);
  or g__2476(w__880 ,w__846 ,w__851);
  and g__2477(w__872 ,w__841 ,w__818);
  or g__2478(w__871 ,w__829 ,w__809);
  or g__2479(w__870 ,w__835 ,w__812);
  and g__2480(w__869 ,w__820 ,w__827);
  or g__2481(w__868 ,w__821 ,w__827);
  and g__2482(w__867 ,w__839 ,w__815);
  or g__2483(w__866 ,w__848 ,w__847);
  or g__2484(w__874 ,w__858 ,w__859);
  or g__2485(w__873 ,w__849 ,w__853);
  not g__2486(w__865 ,w__798);
  not g__2487(w__864 ,w__825);
  not g__2488(w__863 ,w__804);
  not g__2489(w__862 ,w__806);
  not g__2490(w__861 ,w__845);
  not g__2491(w__860 ,w__800);
  not g__2492(w__859 ,w__2349);
  not g__2493(w__858 ,w__2362);
  not g__2494(w__857 ,w__802);
  not g__2495(w__856 ,w__843);
  not g__2496(w__845 ,w__844);
  not g__2497(w__844 ,w__2206);
  not g__2498(w__843 ,w__842);
  not g__2499(w__842 ,w__2212);
  not g__2500(w__841 ,w__840);
  not g__2501(w__840 ,w__2354);
  not g__2502(w__839 ,w__838);
  not g__2503(w__838 ,w__2356);
  not g__2504(w__837 ,w__836);
  not g__2505(w__836 ,w__2209);
  not g__2506(w__835 ,w__834);
  not g__2507(w__834 ,w__2357);
  not g__2508(w__833 ,w__832);
  not g__2509(w__832 ,w__2210);
  not g__2510(w__831 ,w__830);
  not g__2511(w__830 ,w__2211);
  not g__2512(w__829 ,w__828);
  not g__2513(w__828 ,w__2358);
  not g__2514(w__827 ,w__826);
  not g__2515(w__826 ,w__2208);
  not g__2516(w__825 ,w__824);
  not g__2517(w__824 ,w__2353);
  not g__2518(w__823 ,w__822);
  not g__2519(w__822 ,w__2355);
  not g__2520(w__821 ,w__819);
  not g__2521(w__820 ,w__819);
  not g__2522(w__819 ,w__2342);
  not g__2523(w__818 ,w__816);
  not g__2524(w__817 ,w__816);
  not g__2525(w__816 ,w__2341);
  not g__2526(w__815 ,w__813);
  not g__2527(w__814 ,w__813);
  not g__2528(w__813 ,w__2343);
  not g__2529(w__812 ,w__810);
  not g__2530(w__811 ,w__810);
  not g__2531(w__810 ,w__2344);
  not g__2532(w__809 ,w__807);
  not g__2533(w__808 ,w__807);
  not g__2534(w__807 ,w__2345);
  not g__2535(w__806 ,w__805);
  not g__2536(w__805 ,w__2213);
  not g__2537(w__804 ,w__803);
  not g__2538(w__803 ,w__2214);
  not g__2539(w__802 ,w__801);
  not g__2540(w__801 ,w__2215);
  not g__2541(w__800 ,w__799);
  not g__2542(w__799 ,w__2216);
  not g__2543(w__798 ,w__797);
  not g__2544(w__797 ,w__2207);
  not g__2545(w__847 ,w__2350);
  not g__2546(w__796 ,w__795);
  not g__2547(w__795 ,w__2204);
  not g__2548(w__794 ,w__793);
  not g__2549(w__793 ,w__2203);
  not g__2550(w__792 ,w__791);
  not g__2551(w__791 ,w__2200);
  not g__2552(w__790 ,w__789);
  not g__2553(w__789 ,w__2202);
  not g__2554(w__848 ,w__2363);
  not g__2555(w__855 ,w__2346);
  not g__2556(w__851 ,w__2348);
  not g__2557(w__788 ,w__787);
  not g__2558(w__787 ,w__2198);
  not g__2559(w__786 ,w__785);
  not g__2560(w__785 ,w__2201);
  not g__2561(w__853 ,w__2347);
  not g__2562(w__850 ,w__2199);
  not g__2563(w__849 ,w__2360);
  not g__2564(w__854 ,w__2359);
  not g__2565(w__846 ,w__2361);
  not g__2566(w__852 ,w__2340);
  not g__2567(w__784 ,w__783);
  not g__2568(w__783 ,w__2352);
  buf g__2569(w__2535 ,w__2339);
  and g__2570(w__782 ,w__824 ,w__844);
  xor g__2571(w__781 ,w__771 ,w__842);
  xor g__2572(w__2533 ,w__886 ,w__840);
  xor g__2573(w__780 ,w__887 ,w__838);
  xor g__2574(w__779 ,w__912 ,w__836);
  xor g__2575(w__778 ,w__889 ,w__834);
  xor g__2576(w__777 ,w__920 ,w__832);
  xor g__2577(w__776 ,w__919 ,w__830);
  xor g__2578(w__775 ,w__885 ,w__828);
  xor g__2579(w__774 ,w__888 ,w__826);
  xor g__2580(w__773 ,w__911 ,w__822);
  xnor g__2581(w__772 ,w__848 ,w__847);
  xnor g__2582(w__771 ,w__854 ,w__855);
  xnor g__2583(w__770 ,w__846 ,w__851);
  xnor g__2584(w__769 ,w__849 ,w__853);
  xnor g__2585(w__768 ,w__852 ,w__850);
  xnor g__2586(w__2809 ,w__948 ,w__2112);
  xnor g__2587(w__2801 ,w__941 ,w__2120);
  xnor g__2588(w__2800 ,w__1011 ,w__2121);
  xnor g__2589(w__2810 ,w__949 ,w__2111);
  xnor g__2590(w__2802 ,w__942 ,w__2119);
  xnor g__2591(w__2803 ,w__940 ,w__2118);
  xnor g__2592(w__2804 ,w__943 ,w__2117);
  xnor g__2593(w__2805 ,w__946 ,w__2116);
  xnor g__2594(w__2806 ,w__945 ,w__2115);
  xnor g__2595(w__2807 ,w__947 ,w__2114);
  xnor g__2596(w__2808 ,w__944 ,w__2113);
  or g__2597(w__2839 ,w__1008 ,w__1017);
  or g__2598(w__2843 ,w__1009 ,w__1018);
  or g__2599(w__2841 ,w__993 ,w__1014);
  or g__2600(w__2844 ,w__1003 ,w__1021);
  or g__2601(w__2838 ,w__1002 ,w__1016);
  or g__2602(w__2842 ,w__995 ,w__1012);
  or g__2603(w__2845 ,w__1006 ,w__1015);
  or g__2604(w__2840 ,w__1000 ,w__1019);
  or g__2605(w__2847 ,w__1005 ,w__1020);
  and g__2606(w__1021 ,w__2114 ,w__996);
  and g__2607(w__1020 ,w__2111 ,w__1001);
  and g__2608(w__1019 ,w__2118 ,w__1007);
  and g__2609(w__1018 ,w__2115 ,w__1004);
  and g__2610(w__1017 ,w__2119 ,w__999);
  and g__2611(w__1016 ,w__2120 ,w__997);
  and g__2612(w__1015 ,w__2113 ,w__992);
  and g__2613(w__1014 ,w__2117 ,w__994);
  and g__2614(w__1013 ,w__2112 ,w__998);
  and g__2615(w__1012 ,w__2116 ,w__1010);
  xor g__2616(w__2811 ,w__2123 ,w__2110);
  xnor g__2617(w__1011 ,w__991 ,w__2134);
  or g__2618(w__1010 ,w__951 ,w__984);
  and g__2619(w__1009 ,w__954 ,w__982);
  and g__2620(w__1008 ,w__976 ,w__991);
  or g__2621(w__1007 ,w__972 ,w__991);
  and g__2622(w__1006 ,w__969 ,w__980);
  and g__2623(w__1005 ,w__963 ,w__990);
  or g__2624(w__1004 ,w__955 ,w__982);
  and g__2625(w__1003 ,w__960 ,w__986);
  and g__2626(w__1002 ,w__974 ,w__991);
  and g__2627(w__2848 ,w__2123 ,w__2110);
  or g__2628(w__1001 ,w__964 ,w__990);
  and g__2629(w__1000 ,w__972 ,w__991);
  or g__2630(w__999 ,w__976 ,w__991);
  or g__2631(w__998 ,w__957 ,w__988);
  or g__2632(w__997 ,w__974 ,w__991);
  or g__2633(w__996 ,w__961 ,w__986);
  and g__2634(w__995 ,w__952 ,w__984);
  or g__2635(w__994 ,w__966 ,w__978);
  and g__2636(w__993 ,w__967 ,w__978);
  or g__2637(w__992 ,w__970 ,w__980);
  not g__2638(w__990 ,w__989);
  not g__2639(w__989 ,w__2150);
  not g__2640(w__988 ,w__987);
  not g__2641(w__987 ,w__2151);
  not g__2642(w__986 ,w__985);
  not g__2643(w__985 ,w__2153);
  not g__2644(w__984 ,w__983);
  not g__2645(w__983 ,w__2155);
  not g__2646(w__982 ,w__981);
  not g__2647(w__981 ,w__2154);
  not g__2648(w__980 ,w__979);
  not g__2649(w__979 ,w__2152);
  not g__2650(w__978 ,w__977);
  not g__2651(w__977 ,w__2156);
  not g__2652(w__976 ,w__975);
  not g__2653(w__975 ,w__2132);
  not g__2654(w__974 ,w__973);
  not g__2655(w__973 ,w__2133);
  not g__2656(w__972 ,w__971);
  not g__2657(w__971 ,w__2131);
  not g__2658(w__970 ,w__968);
  not g__2659(w__969 ,w__968);
  not g__2660(w__968 ,w__2126);
  not g__2661(w__967 ,w__965);
  not g__2662(w__966 ,w__965);
  not g__2663(w__965 ,w__2130);
  not g__2664(w__964 ,w__962);
  not g__2665(w__963 ,w__962);
  not g__2666(w__962 ,w__2124);
  not g__2667(w__961 ,w__959);
  not g__2668(w__960 ,w__959);
  not g__2669(w__959 ,w__2127);
  not g__2670(w__958 ,w__956);
  not g__2671(w__957 ,w__956);
  not g__2672(w__956 ,w__2125);
  not g__2673(w__955 ,w__953);
  not g__2674(w__954 ,w__953);
  not g__2675(w__953 ,w__2128);
  not g__2676(w__952 ,w__950);
  not g__2677(w__951 ,w__950);
  not g__2678(w__950 ,w__2129);
  buf g__2679(w__2812 ,w__2148);
  buf g__2680(w__991 ,w__2157);
  xor g__2681(w__949 ,w__964 ,w__989);
  xor g__2682(w__948 ,w__958 ,w__987);
  xor g__2683(w__947 ,w__961 ,w__985);
  xor g__2684(w__946 ,w__952 ,w__983);
  xor g__2685(w__945 ,w__955 ,w__981);
  xor g__2686(w__944 ,w__970 ,w__979);
  xor g__2687(w__943 ,w__967 ,w__977);
  xor g__2688(w__942 ,w__991 ,w__975);
  xor g__2689(w__941 ,w__991 ,w__973);
  xor g__2690(w__940 ,w__991 ,w__971);
  xnor g__2691(w__2476 ,w__1151 ,w__1202);
  xnor g__2692(w__2477 ,w__1192 ,w__1201);
  xnor g__2693(w__2478 ,w__1190 ,w__1200);
  xnor g__2694(w__2480 ,w__1030 ,w__1029);
  xor g__2695(w__2479 ,w__1189 ,w__1199);
  or g__2696(w__2516 ,w__1197 ,w__1207);
  or g__2697(w__2519 ,w__1169 ,w__1208);
  or g__2698(w__2517 ,w__1194 ,w__1206);
  or g__2699(w__2514 ,w__1195 ,w__1205);
  or g__2700(w__2515 ,w__1187 ,w__1203);
  or g__2701(w__2518 ,w__1188 ,w__1204);
  xnor g__2702(w__2471 ,w__1129 ,w__1184);
  xnor g__2703(w__2481 ,w__1191 ,w__1171);
  xnor g__2704(w__2472 ,w__1154 ,w__1025);
  nor g__2705(w__1208 ,w__1167 ,w__1191);
  nor g__2706(w__1207 ,w__1196 ,w__1190);
  nor g__2707(w__1206 ,w__1193 ,w__1189);
  and g__2708(w__1205 ,w__1151 ,w__1185);
  and g__2709(w__1204 ,w__1186 ,w__1030);
  nor g__2710(w__1203 ,w__1198 ,w__1192);
  xnor g__2711(w__2474 ,w__1152 ,w__1022);
  xnor g__2712(w__2475 ,w__1153 ,w__1023);
  xnor g__2713(w__2473 ,w__1155 ,w__1024);
  xnor g__2714(w__1202 ,w__1183 ,w__1106);
  xnor g__2715(w__1201 ,w__1173 ,w__1098);
  xnor g__2716(w__1200 ,w__1178 ,w__1093);
  xnor g__2717(w__1199 ,w__1180 ,w__1103);
  and g__2718(w__1198 ,w__1098 ,w__1174);
  or g__2719(w__2510 ,w__1160 ,w__1177);
  nor g__2720(w__1197 ,w__1092 ,w__1179);
  or g__2721(w__2512 ,w__1170 ,w__1172);
  or g__2722(w__2513 ,w__1166 ,w__1175);
  and g__2723(w__1196 ,w__1093 ,w__1179);
  nor g__2724(w__1195 ,w__1105 ,w__1183);
  nor g__2725(w__1194 ,w__1102 ,w__1180);
  and g__2726(w__1193 ,w__1103 ,w__1180);
  or g__2727(w__2511 ,w__1158 ,w__1176);
  and g__2728(w__1188 ,w__1082 ,w__1181);
  nor g__2729(w__1187 ,w__1097 ,w__1174);
  or g__2730(w__1186 ,w__1082 ,w__1181);
  xnor g__2731(w__2482 ,w__1142 ,w__1146);
  or g__2732(w__1185 ,w__1125 ,w__1182);
  xnor g__2733(w__1184 ,w__1148 ,w__2217);
  xnor g__2734(w__1192 ,w__1149 ,w__1088);
  xnor g__2735(w__1191 ,w__1144 ,w__1100);
  xnor g__2736(w__1190 ,w__1143 ,w__1090);
  xnor g__2737(w__1189 ,w__1145 ,w__1095);
  not g__2738(w__1183 ,w__1182);
  not g__2739(w__1179 ,w__1178);
  and g__2740(w__1177 ,w__1168 ,w__1154);
  and g__2741(w__1176 ,w__1165 ,w__1155);
  and g__2742(w__1175 ,w__1157 ,w__1153);
  or g__2743(w__1182 ,w__1131 ,w__1161);
  or g__2744(w__1181 ,w__1130 ,w__1159);
  and g__2745(w__1180 ,w__1137 ,w__1162);
  or g__2746(w__1178 ,w__1136 ,w__1164);
  not g__2747(w__1174 ,w__1173);
  or g__2748(w__2520 ,w__1037 ,w__1150);
  and g__2749(w__1172 ,w__1156 ,w__1152);
  xnor g__2750(w__1171 ,w__1057 ,w__1138);
  or g__2751(w__1173 ,w__1132 ,w__1163);
  nor g__2752(w__1170 ,w__1069 ,w__1134);
  nor g__2753(w__1169 ,w__1058 ,w__1139);
  or g__2754(w__1168 ,w__1126 ,w__1119);
  and g__2755(w__1167 ,w__1057 ,w__1139);
  nor g__2756(w__1166 ,w__1060 ,w__1135);
  or g__2757(w__1165 ,w__1127 ,w__1120);
  nor g__2758(w__1164 ,w__1053 ,w__1033);
  nor g__2759(w__1163 ,w__1049 ,w__1032);
  or g__2760(w__1162 ,w__1043 ,w__1036);
  nor g__2761(w__1161 ,w__1047 ,w__1031);
  nor g__2762(w__1160 ,w__1063 ,w__1140);
  nor g__2763(w__1159 ,w__1055 ,w__1034);
  nor g__2764(w__1158 ,w__1066 ,w__1141);
  or g__2765(w__1157 ,w__1121 ,w__1118);
  or g__2766(w__1156 ,w__1122 ,w__1117);
  nor g__2767(w__1150 ,w__1035 ,w__1142);
  xnor g__2768(w__1149 ,w__1072 ,w__1047);
  xnor g__2769(w__1148 ,w__2364 ,w__2351);
  xnor g__2770(w__1147 ,w__1080 ,w__1043);
  xnor g__2771(w__1146 ,w__1086 ,w__1108);
  xnor g__2772(w__1145 ,w__1076 ,w__1053);
  xnor g__2773(w__1144 ,w__1078 ,w__1055);
  xnor g__2774(w__1143 ,w__1074 ,w__1049);
  or g__2775(w__1155 ,w__1133 ,w__1140);
  xnor g__2776(w__1154 ,w__1045 ,w__1051);
  or g__2777(w__1153 ,w__1028 ,w__1134);
  or g__2778(w__1152 ,w__1026 ,w__1141);
  or g__2779(w__1151 ,w__1027 ,w__1135);
  not g__2780(w__1139 ,w__1138);
  or g__2781(w__1137 ,w__1123 ,w__1084);
  and g__2782(w__1136 ,w__1095 ,w__1076);
  or g__2783(w__1142 ,w__1114 ,w__1041);
  and g__2784(w__1141 ,w__1109 ,w__1110);
  and g__2785(w__1140 ,w__1128 ,w__1124);
  or g__2786(w__1138 ,w__1115 ,w__1039);
  nor g__2787(w__1133 ,w__1128 ,w__1124);
  and g__2788(w__1132 ,w__1090 ,w__1074);
  and g__2789(w__1131 ,w__1088 ,w__1072);
  and g__2790(w__1130 ,w__1100 ,w__1078);
  nor g__2791(w__1129 ,w__1045 ,w__1051);
  and g__2792(w__1135 ,w__1113 ,w__1116);
  and g__2793(w__1134 ,w__1111 ,w__1112);
  not g__2794(w__2549 ,w__2205);
  not g__2795(w__1128 ,w__2362);
  not g__2796(w__1127 ,w__1067);
  not g__2797(w__1126 ,w__1064);
  not g__2798(w__1125 ,w__1106);
  not g__2799(w__1124 ,w__2349);
  not g__2800(w__1123 ,w__1080);
  not g__2801(w__1122 ,w__1070);
  not g__2802(w__1121 ,w__1061);
  not g__2803(w__1108 ,w__1107);
  not g__2804(w__1107 ,w__2206);
  not g__2805(w__1106 ,w__1104);
  not g__2806(w__1105 ,w__1104);
  not g__2807(w__1104 ,w__2212);
  not g__2808(w__1103 ,w__1101);
  not g__2809(w__1102 ,w__1101);
  not g__2810(w__1101 ,w__2209);
  not g__2811(w__1100 ,w__1099);
  not g__2812(w__1099 ,w__2354);
  not g__2813(w__1098 ,w__1096);
  not g__2814(w__1097 ,w__1096);
  not g__2815(w__1096 ,w__2211);
  not g__2816(w__1095 ,w__1094);
  not g__2817(w__1094 ,w__2356);
  not g__2818(w__1093 ,w__1091);
  not g__2819(w__1092 ,w__1091);
  not g__2820(w__1091 ,w__2210);
  not g__2821(w__1090 ,w__1089);
  not g__2822(w__1089 ,w__2357);
  not g__2823(w__1088 ,w__1087);
  not g__2824(w__1087 ,w__2358);
  not g__2825(w__1086 ,w__1085);
  not g__2826(w__1085 ,w__2353);
  not g__2827(w__1084 ,w__1083);
  not g__2828(w__1083 ,w__2208);
  not g__2829(w__1082 ,w__1081);
  not g__2830(w__1081 ,w__2355);
  not g__2831(w__1080 ,w__1079);
  not g__2832(w__1079 ,w__2342);
  not g__2833(w__1078 ,w__1077);
  not g__2834(w__1077 ,w__2341);
  not g__2835(w__1076 ,w__1075);
  not g__2836(w__1075 ,w__2343);
  not g__2837(w__1074 ,w__1073);
  not g__2838(w__1073 ,w__2344);
  not g__2839(w__1072 ,w__1071);
  not g__2840(w__1071 ,w__2345);
  not g__2841(w__1070 ,w__1068);
  not g__2842(w__1069 ,w__1068);
  not g__2843(w__1068 ,w__2214);
  not g__2844(w__1067 ,w__1065);
  not g__2845(w__1066 ,w__1065);
  not g__2846(w__1065 ,w__2215);
  not g__2847(w__1064 ,w__1062);
  not g__2848(w__1063 ,w__1062);
  not g__2849(w__1062 ,w__2216);
  not g__2850(w__1061 ,w__1059);
  not g__2851(w__1060 ,w__1059);
  not g__2852(w__1059 ,w__2213);
  not g__2853(w__1058 ,w__1056);
  not g__2854(w__1057 ,w__1056);
  not g__2855(w__1056 ,w__2207);
  not g__2856(w__1119 ,w__1140);
  not g__2857(w__1120 ,w__1141);
  not g__2858(w__1118 ,w__1135);
  not g__2859(w__1117 ,w__1134);
  not g__2860(w__1055 ,w__1054);
  not g__2861(w__1054 ,w__2200);
  not g__2862(w__1053 ,w__1052);
  not g__2863(w__1052 ,w__2202);
  not g__2864(w__1051 ,w__1050);
  not g__2865(w__1050 ,w__2350);
  not g__2866(w__1049 ,w__1048);
  not g__2867(w__1048 ,w__2203);
  not g__2868(w__1047 ,w__1046);
  not g__2869(w__1046 ,w__2204);
  not g__2870(w__1045 ,w__1044);
  not g__2871(w__1044 ,w__2363);
  not g__2872(w__1043 ,w__1042);
  not g__2873(w__1042 ,w__2201);
  not g__2874(w__1112 ,w__2347);
  not g__2875(w__1116 ,w__2346);
  not g__2876(w__1115 ,w__2199);
  not g__2877(w__1041 ,w__1040);
  not g__2878(w__1040 ,w__2198);
  not g__2879(w__1110 ,w__2348);
  not g__2880(w__1111 ,w__2360);
  not g__2881(w__1113 ,w__2359);
  not g__2882(w__1109 ,w__2361);
  not g__2883(w__1039 ,w__1038);
  not g__2884(w__1038 ,w__2340);
  not g__2885(w__1114 ,w__2352);
  buf g__2886(w__2522 ,w__2339);
  and g__2887(w__1037 ,w__1086 ,w__1107);
  and g__2888(w__1036 ,w__1084 ,w__1079);
  and g__2889(w__1035 ,w__1108 ,w__1085);
  and g__2890(w__1034 ,w__1099 ,w__1077);
  and g__2891(w__1033 ,w__1094 ,w__1075);
  and g__2892(w__1032 ,w__1089 ,w__1073);
  and g__2893(w__1031 ,w__1087 ,w__1071);
  xor g__2894(w__1030 ,w__1147 ,w__1083);
  xor g__2895(w__1029 ,w__1181 ,w__1081);
  nor g__2896(w__1028 ,w__1111 ,w__1112);
  nor g__2897(w__1027 ,w__1113 ,w__1116);
  xnor g__2898(w__2521 ,w__1115 ,w__1039);
  nor g__2899(w__1026 ,w__1109 ,w__1110);
  xor g__2900(w__2483 ,w__1114 ,w__1041);
  xor g__2901(w__1025 ,w__1119 ,w__1064);
  xor g__2902(w__1024 ,w__1120 ,w__1067);
  xor g__2903(w__1023 ,w__1118 ,w__1061);
  xor g__2904(w__1022 ,w__1117 ,w__1070);
  xor g__2905(w__2679 ,w__1270 ,w__2147);
  xor g__2906(w__2680 ,w__1275 ,w__2146);
  xor g__2907(w__2687 ,w__1272 ,w__1218);
  xor g__2908(w__2688 ,w__1271 ,w__2138);
  xor g__2909(w__2689 ,w__1276 ,w__2137);
  xor g__2910(w__2690 ,w__1269 ,w__2136);
  xor g__2911(w__2681 ,w__1274 ,w__2145);
  xor g__2912(w__2682 ,w__1273 ,w__1220);
  xor g__2913(w__2683 ,w__1268 ,w__1214);
  xor g__2914(w__2684 ,w__1267 ,w__2142);
  xor g__2915(w__2685 ,w__1266 ,w__1216);
  xor g__2916(w__2686 ,w__1265 ,w__2140);
  or g__2917(w__2827 ,w__1247 ,w__1287);
  or g__2918(w__2826 ,w__1254 ,w__1286);
  or g__2919(w__2836 ,w__1259 ,w__1285);
  or g__2920(w__2831 ,w__1210 ,w__1283);
  or g__2921(w__2829 ,w__1212 ,w__1279);
  or g__2922(w__2832 ,w__1256 ,w__1281);
  or g__2923(w__2828 ,w__1209 ,w__1284);
  or g__2924(w__2830 ,w__1250 ,w__1277);
  or g__2925(w__2833 ,w__1211 ,w__1280);
  or g__2926(w__2834 ,w__1260 ,w__1278);
  or g__2927(w__2835 ,w__1257 ,w__1282);
  nor g__2928(w__1287 ,w__2145 ,w__1249);
  nor g__2929(w__1286 ,w__2146 ,w__1251);
  nor g__2930(w__1285 ,w__2136 ,w__1255);
  and g__2931(w__1284 ,w__1242 ,w__1263);
  and g__2932(w__1283 ,w__1227 ,w__1262);
  nor g__2933(w__1282 ,w__2137 ,w__1258);
  nor g__2934(w__1281 ,w__2140 ,w__1253);
  and g__2935(w__1280 ,w__1229 ,w__1261);
  and g__2936(w__1279 ,w__1225 ,w__1264);
  nor g__2937(w__1278 ,w__2138 ,w__1248);
  nor g__2938(w__1277 ,w__2142 ,w__1252);
  xnor g__2939(w__1276 ,w__1234 ,w__2160);
  xnor g__2940(w__1275 ,w__1242 ,w__2169);
  xnor g__2941(w__1274 ,w__1242 ,w__2168);
  xnor g__2942(w__1273 ,w__1242 ,w__2167);
  xnor g__2943(w__1272 ,w__2162 ,w__1229);
  xnor g__2944(w__1271 ,w__1231 ,w__2161);
  xnor g__2945(w__1270 ,w__1242 ,w__2170);
  xnor g__2946(w__1269 ,w__1222 ,w__2159);
  xnor g__2947(w__1268 ,w__2166 ,w__1225);
  xnor g__2948(w__1267 ,w__1237 ,w__2165);
  xnor g__2949(w__1266 ,w__2164 ,w__1227);
  xnor g__2950(w__1265 ,w__1240 ,w__2163);
  or g__2951(w__1264 ,w__1244 ,w__2166);
  or g__2952(w__1263 ,w__1245 ,w__2167);
  or g__2953(w__1262 ,w__1246 ,w__2164);
  or g__2954(w__1261 ,w__1243 ,w__2162);
  and g__2955(w__1260 ,w__2161 ,w__1231);
  and g__2956(w__1259 ,w__2159 ,w__1222);
  nor g__2957(w__1258 ,w__2160 ,w__1235);
  and g__2958(w__1257 ,w__2160 ,w__1234);
  and g__2959(w__1256 ,w__2163 ,w__1240);
  nor g__2960(w__1255 ,w__2159 ,w__1223);
  and g__2961(w__1254 ,w__2169 ,w__1242);
  nor g__2962(w__1253 ,w__2163 ,w__1241);
  nor g__2963(w__1252 ,w__2165 ,w__1238);
  nor g__2964(w__1251 ,w__1242 ,w__2169);
  and g__2965(w__1250 ,w__2165 ,w__1237);
  nor g__2966(w__1249 ,w__1242 ,w__2168);
  nor g__2967(w__1248 ,w__2161 ,w__1232);
  and g__2968(w__1247 ,w__2168 ,w__1242);
  not g__2969(w__2691 ,w__2158);
  not g__2970(w__1246 ,w__1216);
  not g__2971(w__1245 ,w__1220);
  not g__2972(w__2862 ,w__2135);
  not g__2973(w__1244 ,w__1214);
  not g__2974(w__1243 ,w__1218);
  not g__2975(w__1241 ,w__1239);
  not g__2976(w__1240 ,w__1239);
  not g__2977(w__1239 ,w__2153);
  not g__2978(w__1238 ,w__1236);
  not g__2979(w__1237 ,w__1236);
  not g__2980(w__1236 ,w__2155);
  not g__2981(w__1235 ,w__1233);
  not g__2982(w__1234 ,w__1233);
  not g__2983(w__1233 ,w__2150);
  not g__2984(w__1232 ,w__1230);
  not g__2985(w__1231 ,w__1230);
  not g__2986(w__1230 ,w__2151);
  not g__2987(w__1229 ,w__1228);
  not g__2988(w__1228 ,w__2152);
  not g__2989(w__1227 ,w__1226);
  not g__2990(w__1226 ,w__2154);
  not g__2991(w__1225 ,w__1224);
  not g__2992(w__1224 ,w__2156);
  not g__2993(w__1223 ,w__1221);
  not g__2994(w__1222 ,w__1221);
  not g__2995(w__1221 ,w__2149);
  not g__2996(w__1220 ,w__1219);
  not g__2997(w__1219 ,w__2144);
  not g__2998(w__1218 ,w__1217);
  not g__2999(w__1217 ,w__2139);
  not g__3000(w__1216 ,w__1215);
  not g__3001(w__1215 ,w__2141);
  not g__3002(w__1214 ,w__1213);
  not g__3003(w__1213 ,w__2143);
  buf g__3004(w__2837 ,w__2148);
  buf g__3005(w__1242 ,w__2157);
  and g__3006(w__1212 ,w__2166 ,w__1213);
  and g__3007(w__1211 ,w__2162 ,w__1217);
  and g__3008(w__1210 ,w__2164 ,w__1215);
  and g__3009(w__1209 ,w__2167 ,w__1219);
  xnor g__3010(out1[12] ,w__1348 ,w__1317);
  or g__3011(w__1348 ,w__1301 ,w__1347);
  xnor g__3012(out1[11] ,w__1346 ,w__1320);
  and g__3013(w__1347 ,w__1306 ,w__1346);
  or g__3014(w__1346 ,w__1288 ,w__1345);
  xnor g__3015(out1[10] ,w__1344 ,w__1319);
  and g__3016(w__1345 ,w__1304 ,w__1344);
  or g__3017(w__1344 ,w__1300 ,w__1343);
  xnor g__3018(out1[9] ,w__1342 ,w__1312);
  and g__3019(w__1343 ,w__1299 ,w__1342);
  or g__3020(w__1342 ,w__1292 ,w__1341);
  xnor g__3021(out1[8] ,w__1340 ,w__1316);
  and g__3022(w__1341 ,w__1290 ,w__1340);
  or g__3023(w__1340 ,w__1311 ,w__1339);
  xnor g__3024(out1[7] ,w__1338 ,w__1315);
  and g__3025(w__1339 ,w__1310 ,w__1338);
  or g__3026(w__1338 ,w__1305 ,w__1337);
  xnor g__3027(out1[6] ,w__1336 ,w__1314);
  and g__3028(w__1337 ,w__1294 ,w__1336);
  or g__3029(w__1336 ,w__1298 ,w__1335);
  xnor g__3030(out1[5] ,w__1334 ,w__1313);
  and g__3031(w__1335 ,w__1303 ,w__1334);
  or g__3032(w__1334 ,w__1309 ,w__1333);
  xnor g__3033(out1[4] ,w__1332 ,w__1318);
  and g__3034(w__1333 ,w__1308 ,w__1332);
  or g__3035(w__1332 ,w__1291 ,w__1331);
  xnor g__3036(out1[3] ,w__1330 ,w__1324);
  and g__3037(w__1331 ,w__1307 ,w__1330);
  or g__3038(w__1330 ,w__1296 ,w__1329);
  xnor g__3039(out1[2] ,w__1328 ,w__1323);
  and g__3040(w__1329 ,w__1289 ,w__1328);
  or g__3041(w__1328 ,w__1295 ,w__1327);
  xnor g__3042(out1[1] ,w__1326 ,w__1322);
  and g__3043(w__1327 ,w__1297 ,w__1326);
  xnor g__3044(out1[0] ,w__1321 ,w__2171);
  or g__3045(w__1326 ,w__1293 ,w__1325);
  and g__3046(w__1325 ,w__2185 ,w__1302);
  xnor g__3047(w__1324 ,w__2188 ,w__2175);
  xnor g__3048(w__1323 ,w__2187 ,w__2174);
  xnor g__3049(w__1322 ,w__2186 ,w__2173);
  xnor g__3050(w__1321 ,w__2185 ,w__2172);
  xnor g__3051(w__1320 ,w__2196 ,w__2183);
  xnor g__3052(w__1319 ,w__2195 ,w__2182);
  xnor g__3053(w__1318 ,w__2189 ,w__2176);
  xnor g__3054(w__1317 ,w__2197 ,w__2184);
  xnor g__3055(w__1316 ,w__2193 ,w__2180);
  xnor g__3056(w__1315 ,w__2192 ,w__2179);
  xnor g__3057(w__1314 ,w__2191 ,w__2178);
  xnor g__3058(w__1313 ,w__2190 ,w__2177);
  xnor g__3059(w__1312 ,w__2194 ,w__2181);
  and g__3060(w__1311 ,w__2192 ,w__2179);
  or g__3061(w__1310 ,w__2192 ,w__2179);
  and g__3062(w__1309 ,w__2189 ,w__2176);
  or g__3063(w__1308 ,w__2189 ,w__2176);
  or g__3064(w__1307 ,w__2188 ,w__2175);
  or g__3065(w__1306 ,w__2196 ,w__2183);
  and g__3066(w__1305 ,w__2191 ,w__2178);
  or g__3067(w__1304 ,w__2195 ,w__2182);
  or g__3068(w__1303 ,w__2190 ,w__2177);
  or g__3069(w__1302 ,w__2172 ,w__2171);
  and g__3070(w__1301 ,w__2196 ,w__2183);
  and g__3071(w__1300 ,w__2194 ,w__2181);
  or g__3072(w__1299 ,w__2194 ,w__2181);
  and g__3073(w__1298 ,w__2190 ,w__2177);
  or g__3074(w__1297 ,w__2186 ,w__2173);
  and g__3075(w__1296 ,w__2187 ,w__2174);
  and g__3076(w__1295 ,w__2186 ,w__2173);
  or g__3077(w__1294 ,w__2191 ,w__2178);
  and g__3078(w__1293 ,w__2172 ,w__2171);
  and g__3079(w__1292 ,w__2193 ,w__2180);
  and g__3080(w__1291 ,w__2188 ,w__2175);
  or g__3081(w__1290 ,w__2193 ,w__2180);
  or g__3082(w__1289 ,w__2187 ,w__2174);
  and g__3083(w__1288 ,w__2195 ,w__2182);
  xnor g__3084(out2[12] ,w__1409 ,w__1378);
  or g__3085(w__1409 ,w__1362 ,w__1408);
  xnor g__3086(out2[11] ,w__1407 ,w__1381);
  and g__3087(w__1408 ,w__1367 ,w__1407);
  or g__3088(w__1407 ,w__1349 ,w__1406);
  xnor g__3089(out2[10] ,w__1405 ,w__1380);
  and g__3090(w__1406 ,w__1365 ,w__1405);
  or g__3091(w__1405 ,w__1361 ,w__1404);
  xnor g__3092(out2[9] ,w__1403 ,w__1373);
  and g__3093(w__1404 ,w__1360 ,w__1403);
  or g__3094(w__1403 ,w__1353 ,w__1402);
  xnor g__3095(out2[8] ,w__1401 ,w__1377);
  and g__3096(w__1402 ,w__1351 ,w__1401);
  or g__3097(w__1401 ,w__1372 ,w__1400);
  xnor g__3098(out2[7] ,w__1399 ,w__1376);
  and g__3099(w__1400 ,w__1371 ,w__1399);
  or g__3100(w__1399 ,w__1366 ,w__1398);
  xnor g__3101(out2[6] ,w__1397 ,w__1375);
  and g__3102(w__1398 ,w__1355 ,w__1397);
  or g__3103(w__1397 ,w__1359 ,w__1396);
  xnor g__3104(out2[5] ,w__1395 ,w__1374);
  and g__3105(w__1396 ,w__1364 ,w__1395);
  or g__3106(w__1395 ,w__1370 ,w__1394);
  xnor g__3107(out2[4] ,w__1393 ,w__1379);
  and g__3108(w__1394 ,w__1369 ,w__1393);
  or g__3109(w__1393 ,w__1352 ,w__1392);
  xnor g__3110(out2[3] ,w__1391 ,w__1385);
  and g__3111(w__1392 ,w__1368 ,w__1391);
  or g__3112(w__1391 ,w__1357 ,w__1390);
  xnor g__3113(out2[2] ,w__1389 ,w__1384);
  and g__3114(w__1390 ,w__1350 ,w__1389);
  or g__3115(w__1389 ,w__1356 ,w__1388);
  xnor g__3116(out2[1] ,w__1387 ,w__1383);
  and g__3117(w__1388 ,w__1358 ,w__1387);
  xnor g__3118(out2[0] ,w__1382 ,w__2082);
  or g__3119(w__1387 ,w__1354 ,w__1386);
  and g__3120(w__1386 ,w__2096 ,w__1363);
  xnor g__3121(w__1385 ,w__2099 ,w__2086);
  xnor g__3122(w__1384 ,w__2098 ,w__2085);
  xnor g__3123(w__1383 ,w__2097 ,w__2084);
  xnor g__3124(w__1382 ,w__2096 ,w__2083);
  xnor g__3125(w__1381 ,w__2107 ,w__2094);
  xnor g__3126(w__1380 ,w__2106 ,w__2093);
  xnor g__3127(w__1379 ,w__2100 ,w__2087);
  xnor g__3128(w__1378 ,w__2108 ,w__2095);
  xnor g__3129(w__1377 ,w__2104 ,w__2091);
  xnor g__3130(w__1376 ,w__2103 ,w__2090);
  xnor g__3131(w__1375 ,w__2102 ,w__2089);
  xnor g__3132(w__1374 ,w__2101 ,w__2088);
  xnor g__3133(w__1373 ,w__2105 ,w__2092);
  and g__3134(w__1372 ,w__2103 ,w__2090);
  or g__3135(w__1371 ,w__2103 ,w__2090);
  and g__3136(w__1370 ,w__2100 ,w__2087);
  or g__3137(w__1369 ,w__2100 ,w__2087);
  or g__3138(w__1368 ,w__2099 ,w__2086);
  or g__3139(w__1367 ,w__2107 ,w__2094);
  and g__3140(w__1366 ,w__2102 ,w__2089);
  or g__3141(w__1365 ,w__2106 ,w__2093);
  or g__3142(w__1364 ,w__2101 ,w__2088);
  or g__3143(w__1363 ,w__2083 ,w__2082);
  and g__3144(w__1362 ,w__2107 ,w__2094);
  and g__3145(w__1361 ,w__2105 ,w__2092);
  or g__3146(w__1360 ,w__2105 ,w__2092);
  and g__3147(w__1359 ,w__2101 ,w__2088);
  or g__3148(w__1358 ,w__2097 ,w__2084);
  and g__3149(w__1357 ,w__2098 ,w__2085);
  and g__3150(w__1356 ,w__2097 ,w__2084);
  or g__3151(w__1355 ,w__2102 ,w__2089);
  and g__3152(w__1354 ,w__2083 ,w__2082);
  and g__3153(w__1353 ,w__2104 ,w__2091);
  and g__3154(w__1352 ,w__2099 ,w__2086);
  or g__3155(w__1351 ,w__2104 ,w__2091);
  or g__3156(w__1350 ,w__2098 ,w__2085);
  and g__3157(w__1349 ,w__2106 ,w__2093);
  buf g__3158(w__2871 ,w__2924);
  buf g__3159(w__2888 ,w__2926);
  buf g__3160(w__2846 ,w__1013);
endmodule
